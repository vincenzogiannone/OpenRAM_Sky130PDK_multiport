magic
tech sky130A
magscale 1 2
timestamp 1644949024
<< checkpaint >>
rect -1260 -1286 3030 1410
<< scnmos >>
rect 60 0 90 94
rect 168 0 198 94
rect 276 0 306 94
rect 384 0 414 94
rect 492 0 522 94
rect 600 0 630 94
rect 708 0 738 94
rect 816 0 846 94
rect 924 0 954 94
rect 1032 0 1062 94
rect 1140 0 1170 94
rect 1248 0 1278 94
rect 1356 0 1386 94
rect 1464 0 1494 94
rect 1572 0 1602 94
rect 1680 0 1710 94
<< ndiff >>
rect 0 64 60 94
rect 0 30 8 64
rect 42 30 60 64
rect 0 0 60 30
rect 90 64 168 94
rect 90 30 112 64
rect 146 30 168 64
rect 90 0 168 30
rect 198 64 276 94
rect 198 30 220 64
rect 254 30 276 64
rect 198 0 276 30
rect 306 64 384 94
rect 306 30 328 64
rect 362 30 384 64
rect 306 0 384 30
rect 414 64 492 94
rect 414 30 436 64
rect 470 30 492 64
rect 414 0 492 30
rect 522 64 600 94
rect 522 30 544 64
rect 578 30 600 64
rect 522 0 600 30
rect 630 64 708 94
rect 630 30 652 64
rect 686 30 708 64
rect 630 0 708 30
rect 738 64 816 94
rect 738 30 760 64
rect 794 30 816 64
rect 738 0 816 30
rect 846 64 924 94
rect 846 30 868 64
rect 902 30 924 64
rect 846 0 924 30
rect 954 64 1032 94
rect 954 30 976 64
rect 1010 30 1032 64
rect 954 0 1032 30
rect 1062 64 1140 94
rect 1062 30 1084 64
rect 1118 30 1140 64
rect 1062 0 1140 30
rect 1170 64 1248 94
rect 1170 30 1192 64
rect 1226 30 1248 64
rect 1170 0 1248 30
rect 1278 64 1356 94
rect 1278 30 1300 64
rect 1334 30 1356 64
rect 1278 0 1356 30
rect 1386 64 1464 94
rect 1386 30 1408 64
rect 1442 30 1464 64
rect 1386 0 1464 30
rect 1494 64 1572 94
rect 1494 30 1516 64
rect 1550 30 1572 64
rect 1494 0 1572 30
rect 1602 64 1680 94
rect 1602 30 1624 64
rect 1658 30 1680 64
rect 1602 0 1680 30
rect 1710 64 1770 94
rect 1710 30 1728 64
rect 1762 30 1770 64
rect 1710 0 1770 30
<< ndiffc >>
rect 8 30 42 64
rect 112 30 146 64
rect 220 30 254 64
rect 328 30 362 64
rect 436 30 470 64
rect 544 30 578 64
rect 652 30 686 64
rect 760 30 794 64
rect 868 30 902 64
rect 976 30 1010 64
rect 1084 30 1118 64
rect 1192 30 1226 64
rect 1300 30 1334 64
rect 1408 30 1442 64
rect 1516 30 1550 64
rect 1624 30 1658 64
rect 1728 30 1762 64
<< poly >>
rect 60 120 1710 150
rect 60 94 90 120
rect 168 94 198 120
rect 276 94 306 120
rect 384 94 414 120
rect 492 94 522 120
rect 600 94 630 120
rect 708 94 738 120
rect 816 94 846 120
rect 924 94 954 120
rect 1032 94 1062 120
rect 1140 94 1170 120
rect 1248 94 1278 120
rect 1356 94 1386 120
rect 1464 94 1494 120
rect 1572 94 1602 120
rect 1680 94 1710 120
rect 60 -26 90 0
rect 168 -26 198 0
rect 276 -26 306 0
rect 384 -26 414 0
rect 492 -26 522 0
rect 600 -26 630 0
rect 708 -26 738 0
rect 816 -26 846 0
rect 924 -26 954 0
rect 1032 -26 1062 0
rect 1140 -26 1170 0
rect 1248 -26 1278 0
rect 1356 -26 1386 0
rect 1464 -26 1494 0
rect 1572 -26 1602 0
rect 1680 -26 1710 0
<< locali >>
rect 112 114 1658 148
rect 8 64 42 80
rect 8 14 42 30
rect 112 64 146 114
rect 112 14 146 30
rect 220 64 254 80
rect 220 14 254 30
rect 328 64 362 114
rect 328 14 362 30
rect 436 64 470 80
rect 436 14 470 30
rect 544 64 578 114
rect 544 14 578 30
rect 652 64 686 80
rect 652 14 686 30
rect 760 64 794 114
rect 760 14 794 30
rect 868 64 902 80
rect 868 14 902 30
rect 976 64 1010 114
rect 976 14 1010 30
rect 1084 64 1118 80
rect 1084 14 1118 30
rect 1192 64 1226 114
rect 1192 14 1226 30
rect 1300 64 1334 80
rect 1300 14 1334 30
rect 1408 64 1442 114
rect 1408 14 1442 30
rect 1516 64 1550 80
rect 1516 14 1550 30
rect 1624 64 1658 114
rect 1624 14 1658 30
rect 1728 64 1762 80
rect 1728 14 1762 30
use contact_8  contact_8_0
timestamp 1644949024
transform 1 0 1720 0 1 6
box 0 0 1 1
use contact_8  contact_8_1
timestamp 1644949024
transform 1 0 1616 0 1 6
box 0 0 1 1
use contact_8  contact_8_2
timestamp 1644949024
transform 1 0 1508 0 1 6
box 0 0 1 1
use contact_8  contact_8_3
timestamp 1644949024
transform 1 0 1400 0 1 6
box 0 0 1 1
use contact_8  contact_8_4
timestamp 1644949024
transform 1 0 1292 0 1 6
box 0 0 1 1
use contact_8  contact_8_5
timestamp 1644949024
transform 1 0 1184 0 1 6
box 0 0 1 1
use contact_8  contact_8_6
timestamp 1644949024
transform 1 0 1076 0 1 6
box 0 0 1 1
use contact_8  contact_8_7
timestamp 1644949024
transform 1 0 968 0 1 6
box 0 0 1 1
use contact_8  contact_8_8
timestamp 1644949024
transform 1 0 860 0 1 6
box 0 0 1 1
use contact_8  contact_8_9
timestamp 1644949024
transform 1 0 752 0 1 6
box 0 0 1 1
use contact_8  contact_8_10
timestamp 1644949024
transform 1 0 644 0 1 6
box 0 0 1 1
use contact_8  contact_8_11
timestamp 1644949024
transform 1 0 536 0 1 6
box 0 0 1 1
use contact_8  contact_8_12
timestamp 1644949024
transform 1 0 428 0 1 6
box 0 0 1 1
use contact_8  contact_8_13
timestamp 1644949024
transform 1 0 320 0 1 6
box 0 0 1 1
use contact_8  contact_8_14
timestamp 1644949024
transform 1 0 212 0 1 6
box 0 0 1 1
use contact_8  contact_8_15
timestamp 1644949024
transform 1 0 104 0 1 6
box 0 0 1 1
use contact_8  contact_8_16
timestamp 1644949024
transform 1 0 0 0 1 6
box 0 0 1 1
<< labels >>
rlabel mvvaractor s 885 135 885 135 4 G
rlabel locali s 1101 47 1101 47 4 S
rlabel locali s 237 47 237 47 4 S
rlabel locali s 885 47 885 47 4 S
rlabel locali s 1533 47 1533 47 4 S
rlabel locali s 1745 47 1745 47 4 S
rlabel locali s 25 47 25 47 4 S
rlabel locali s 669 47 669 47 4 S
rlabel locali s 1317 47 1317 47 4 S
rlabel locali s 453 47 453 47 4 S
rlabel locali s 885 131 885 131 4 D
<< properties >>
string FIXED_BBOX -25 -26 1795 150
string GDS_FILE sram_0rw2r1w_4_16_sky130A.gds
string GDS_END 484414
string GDS_START 480618
<< end >>
