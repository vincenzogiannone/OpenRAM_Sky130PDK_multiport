magic
tech sky130A
magscale 1 2
timestamp 1644949024
<< checkpaint >>
rect -1260 -1302 6520 25929
<< viali >>
rect 2422 23887 2456 23921
rect 2422 22263 2456 22297
rect 2422 20807 2456 20841
rect 2422 19183 2456 19217
rect 2422 14651 2456 14685
rect 2422 13027 2456 13061
rect 2422 11571 2456 11605
rect 2422 9947 2456 9981
rect 2422 5415 2456 5449
rect 2422 3791 2456 3825
rect 2422 2335 2456 2369
rect 2422 711 2456 745
<< metal1 >>
rect 5162 24582 5168 24634
rect 5220 24582 5226 24634
rect 3500 24200 3506 24252
rect 3558 24240 3564 24252
rect 3558 24212 4674 24240
rect 3558 24200 3564 24212
rect 3248 24114 3254 24166
rect 3306 24154 3312 24166
rect 3306 24126 4578 24154
rect 3306 24114 3312 24126
rect 2828 24028 2834 24080
rect 2886 24068 2892 24080
rect 2886 24040 4482 24068
rect 2886 24028 2892 24040
rect 4814 24000 5180 24028
rect 3500 23942 3506 23994
rect 3558 23982 3564 23994
rect 3558 23954 4278 23982
rect 3558 23942 3564 23954
rect 2407 23878 2413 23930
rect 2465 23878 2471 23930
rect 3248 23856 3254 23908
rect 3306 23896 3312 23908
rect 3306 23868 4182 23896
rect 4896 23878 5180 23906
rect 3306 23856 3312 23868
rect 2744 23770 2750 23822
rect 2802 23810 2808 23822
rect 2802 23782 4086 23810
rect 2802 23770 2808 23782
rect 3500 23684 3506 23736
rect 3558 23724 3564 23736
rect 5104 23732 5180 23760
rect 3558 23696 3990 23724
rect 3558 23684 3564 23696
rect 3248 23598 3254 23650
rect 3306 23638 3312 23650
rect 3306 23610 3894 23638
rect 3306 23598 3312 23610
rect 2660 23512 2666 23564
rect 2718 23552 2724 23564
rect 2718 23524 3798 23552
rect 2718 23512 2724 23524
rect 5162 23044 5168 23096
rect 5220 23044 5226 23096
rect 2744 22576 2750 22628
rect 2802 22616 2808 22628
rect 2802 22588 3798 22616
rect 2802 22576 2808 22588
rect 3164 22490 3170 22542
rect 3222 22530 3228 22542
rect 3222 22502 3894 22530
rect 3222 22490 3228 22502
rect 3500 22404 3506 22456
rect 3558 22444 3564 22456
rect 3558 22416 3990 22444
rect 3558 22404 3564 22416
rect 5104 22380 5180 22408
rect 2828 22318 2834 22370
rect 2886 22358 2892 22370
rect 2886 22330 4086 22358
rect 2886 22318 2892 22330
rect 2407 22254 2413 22306
rect 2465 22254 2471 22306
rect 3164 22232 3170 22284
rect 3222 22272 3228 22284
rect 3222 22244 4182 22272
rect 3222 22232 3228 22244
rect 4896 22234 5180 22262
rect 3500 22146 3506 22198
rect 3558 22186 3564 22198
rect 3558 22158 4278 22186
rect 3558 22146 3564 22158
rect 4814 22112 5180 22140
rect 2912 22060 2918 22112
rect 2970 22100 2976 22112
rect 2970 22072 4482 22100
rect 2970 22060 2976 22072
rect 3164 21974 3170 22026
rect 3222 22014 3228 22026
rect 3222 21986 4578 22014
rect 3222 21974 3228 21986
rect 3500 21888 3506 21940
rect 3558 21928 3564 21940
rect 3558 21900 4674 21928
rect 3558 21888 3564 21900
rect 5162 21506 5168 21558
rect 5220 21506 5226 21558
rect 3500 21124 3506 21176
rect 3558 21164 3564 21176
rect 3558 21136 4674 21164
rect 3558 21124 3564 21136
rect 3164 21038 3170 21090
rect 3222 21078 3228 21090
rect 3222 21050 4578 21078
rect 3222 21038 3228 21050
rect 2660 20952 2666 21004
rect 2718 20992 2724 21004
rect 2718 20964 4482 20992
rect 2718 20952 2724 20964
rect 4814 20924 5180 20952
rect 3500 20866 3506 20918
rect 3558 20906 3564 20918
rect 3558 20878 4278 20906
rect 3558 20866 3564 20878
rect 420 20798 426 20850
rect 478 20838 484 20850
rect 700 20838 706 20850
rect 478 20810 706 20838
rect 478 20798 484 20810
rect 700 20798 706 20810
rect 758 20798 764 20850
rect 2407 20798 2413 20850
rect 2465 20798 2471 20850
rect 3080 20780 3086 20832
rect 3138 20820 3144 20832
rect 3138 20792 4182 20820
rect 4896 20802 5180 20830
rect 3138 20780 3144 20792
rect 2912 20694 2918 20746
rect 2970 20734 2976 20746
rect 2970 20706 4086 20734
rect 2970 20694 2976 20706
rect 3500 20608 3506 20660
rect 3558 20648 3564 20660
rect 5104 20656 5180 20684
rect 3558 20620 3990 20648
rect 3558 20608 3564 20620
rect 3080 20522 3086 20574
rect 3138 20562 3144 20574
rect 3138 20534 3894 20562
rect 3138 20522 3144 20534
rect 2828 20436 2834 20488
rect 2886 20476 2892 20488
rect 2886 20448 3798 20476
rect 2886 20436 2892 20448
rect 5162 19968 5168 20020
rect 5220 19968 5226 20020
rect 2912 19500 2918 19552
rect 2970 19540 2976 19552
rect 2970 19512 3798 19540
rect 2970 19500 2976 19512
rect 2996 19414 3002 19466
rect 3054 19454 3060 19466
rect 3054 19426 3894 19454
rect 3054 19414 3060 19426
rect 3500 19328 3506 19380
rect 3558 19368 3564 19380
rect 3558 19340 3990 19368
rect 3558 19328 3564 19340
rect 5104 19304 5180 19332
rect 2660 19242 2666 19294
rect 2718 19282 2724 19294
rect 2718 19254 4086 19282
rect 2718 19242 2724 19254
rect 336 19174 342 19226
rect 394 19214 400 19226
rect 616 19214 622 19226
rect 394 19186 622 19214
rect 394 19174 400 19186
rect 616 19174 622 19186
rect 674 19174 680 19226
rect 2407 19174 2413 19226
rect 2465 19174 2471 19226
rect 3080 19156 3086 19208
rect 3138 19196 3144 19208
rect 3138 19168 4182 19196
rect 3138 19156 3144 19168
rect 4896 19158 5180 19186
rect 3500 19070 3506 19122
rect 3558 19110 3564 19122
rect 3558 19082 4278 19110
rect 3558 19070 3564 19082
rect 4814 19036 5180 19064
rect 2744 18984 2750 19036
rect 2802 19024 2808 19036
rect 2802 18996 4482 19024
rect 2802 18984 2808 18996
rect 3080 18898 3086 18950
rect 3138 18938 3144 18950
rect 3138 18910 4578 18938
rect 3138 18898 3144 18910
rect 3500 18812 3506 18864
rect 3558 18852 3564 18864
rect 3558 18824 4674 18852
rect 3558 18812 3564 18824
rect 5162 18430 5168 18482
rect 5220 18430 5226 18482
rect 3500 18048 3506 18100
rect 3558 18088 3564 18100
rect 3558 18060 4674 18088
rect 3558 18048 3564 18060
rect 2996 17962 3002 18014
rect 3054 18002 3060 18014
rect 3054 17974 4578 18002
rect 3054 17962 3060 17974
rect 2828 17876 2834 17928
rect 2886 17916 2892 17928
rect 2886 17888 4482 17916
rect 2886 17876 2892 17888
rect 4814 17848 5180 17876
rect 3500 17790 3506 17842
rect 3558 17830 3564 17842
rect 3558 17802 4278 17830
rect 3558 17790 3564 17802
rect 2996 17704 3002 17756
rect 3054 17744 3060 17756
rect 3054 17716 4182 17744
rect 4896 17726 5180 17754
rect 3054 17704 3060 17716
rect 2744 17618 2750 17670
rect 2802 17658 2808 17670
rect 2802 17630 4086 17658
rect 2802 17618 2808 17630
rect 3500 17532 3506 17584
rect 3558 17572 3564 17584
rect 5104 17580 5180 17608
rect 3558 17544 3990 17572
rect 3558 17532 3564 17544
rect 2996 17446 3002 17498
rect 3054 17486 3060 17498
rect 3054 17458 3894 17486
rect 3054 17446 3060 17458
rect 2660 17360 2666 17412
rect 2718 17400 2724 17412
rect 2718 17372 3798 17400
rect 2718 17360 2724 17372
rect 5162 16892 5168 16944
rect 5220 16892 5226 16944
rect 2744 16424 2750 16476
rect 2802 16464 2808 16476
rect 2802 16436 3798 16464
rect 2802 16424 2808 16436
rect 3248 16338 3254 16390
rect 3306 16378 3312 16390
rect 3306 16350 3894 16378
rect 3306 16338 3312 16350
rect 3416 16252 3422 16304
rect 3474 16292 3480 16304
rect 3474 16264 3990 16292
rect 3474 16252 3480 16264
rect 5104 16228 5180 16256
rect 2828 16166 2834 16218
rect 2886 16206 2892 16218
rect 2886 16178 4086 16206
rect 2886 16166 2892 16178
rect 3248 16080 3254 16132
rect 3306 16120 3312 16132
rect 3306 16092 4182 16120
rect 3306 16080 3312 16092
rect 4896 16082 5180 16110
rect 3416 15994 3422 16046
rect 3474 16034 3480 16046
rect 3474 16006 4278 16034
rect 3474 15994 3480 16006
rect 4814 15960 5180 15988
rect 2912 15908 2918 15960
rect 2970 15948 2976 15960
rect 2970 15920 4482 15948
rect 2970 15908 2976 15920
rect 3248 15822 3254 15874
rect 3306 15862 3312 15874
rect 3306 15834 4578 15862
rect 3306 15822 3312 15834
rect 3416 15736 3422 15788
rect 3474 15776 3480 15788
rect 3474 15748 4674 15776
rect 3474 15736 3480 15748
rect 5162 15354 5168 15406
rect 5220 15354 5226 15406
rect 3416 14972 3422 15024
rect 3474 15012 3480 15024
rect 3474 14984 4674 15012
rect 3474 14972 3480 14984
rect 3248 14886 3254 14938
rect 3306 14926 3312 14938
rect 3306 14898 4578 14926
rect 3306 14886 3312 14898
rect 2660 14800 2666 14852
rect 2718 14840 2724 14852
rect 2718 14812 4482 14840
rect 2718 14800 2724 14812
rect 4814 14772 5180 14800
rect 3416 14714 3422 14766
rect 3474 14754 3480 14766
rect 3474 14726 4278 14754
rect 3474 14714 3480 14726
rect 2407 14642 2413 14694
rect 2465 14642 2471 14694
rect 3164 14628 3170 14680
rect 3222 14668 3228 14680
rect 3222 14640 4182 14668
rect 4896 14650 5180 14678
rect 3222 14628 3228 14640
rect 2912 14542 2918 14594
rect 2970 14582 2976 14594
rect 2970 14554 4086 14582
rect 2970 14542 2976 14554
rect 3416 14456 3422 14508
rect 3474 14496 3480 14508
rect 5104 14504 5180 14532
rect 3474 14468 3990 14496
rect 3474 14456 3480 14468
rect 3164 14370 3170 14422
rect 3222 14410 3228 14422
rect 3222 14382 3894 14410
rect 3222 14370 3228 14382
rect 2828 14284 2834 14336
rect 2886 14324 2892 14336
rect 2886 14296 3798 14324
rect 2886 14284 2892 14296
rect 5162 13816 5168 13868
rect 5220 13816 5226 13868
rect 2912 13348 2918 13400
rect 2970 13388 2976 13400
rect 2970 13360 3798 13388
rect 2970 13348 2976 13360
rect 3080 13262 3086 13314
rect 3138 13302 3144 13314
rect 3138 13274 3894 13302
rect 3138 13262 3144 13274
rect 3416 13176 3422 13228
rect 3474 13216 3480 13228
rect 3474 13188 3990 13216
rect 3474 13176 3480 13188
rect 5104 13152 5180 13180
rect 2660 13090 2666 13142
rect 2718 13130 2724 13142
rect 2718 13102 4086 13130
rect 2718 13090 2724 13102
rect 2407 13018 2413 13070
rect 2465 13018 2471 13070
rect 3164 13004 3170 13056
rect 3222 13044 3228 13056
rect 3222 13016 4182 13044
rect 3222 13004 3228 13016
rect 4896 13006 5180 13034
rect 3416 12918 3422 12970
rect 3474 12958 3480 12970
rect 3474 12930 4278 12958
rect 3474 12918 3480 12930
rect 4814 12884 5180 12912
rect 2744 12832 2750 12884
rect 2802 12872 2808 12884
rect 2802 12844 4482 12872
rect 2802 12832 2808 12844
rect 3164 12746 3170 12798
rect 3222 12786 3228 12798
rect 3222 12758 4578 12786
rect 3222 12746 3228 12758
rect 3416 12660 3422 12712
rect 3474 12700 3480 12712
rect 3474 12672 4674 12700
rect 3474 12660 3480 12672
rect 5162 12278 5168 12330
rect 5220 12278 5226 12330
rect 3416 11896 3422 11948
rect 3474 11936 3480 11948
rect 3474 11908 4674 11936
rect 3474 11896 3480 11908
rect 3080 11810 3086 11862
rect 3138 11850 3144 11862
rect 3138 11822 4578 11850
rect 3138 11810 3144 11822
rect 2828 11724 2834 11776
rect 2886 11764 2892 11776
rect 2886 11736 4482 11764
rect 2886 11724 2892 11736
rect 4814 11696 5180 11724
rect 3416 11638 3422 11690
rect 3474 11678 3480 11690
rect 3474 11650 4278 11678
rect 3474 11638 3480 11650
rect 252 11562 258 11614
rect 310 11602 316 11614
rect 700 11602 706 11614
rect 310 11574 706 11602
rect 310 11562 316 11574
rect 700 11562 706 11574
rect 758 11562 764 11614
rect 2407 11562 2413 11614
rect 2465 11562 2471 11614
rect 3080 11552 3086 11604
rect 3138 11592 3144 11604
rect 3138 11564 4182 11592
rect 4896 11574 5180 11602
rect 3138 11552 3144 11564
rect 2744 11466 2750 11518
rect 2802 11506 2808 11518
rect 2802 11478 4086 11506
rect 2802 11466 2808 11478
rect 3416 11380 3422 11432
rect 3474 11420 3480 11432
rect 5104 11428 5180 11456
rect 3474 11392 3990 11420
rect 3474 11380 3480 11392
rect 3080 11294 3086 11346
rect 3138 11334 3144 11346
rect 3138 11306 3894 11334
rect 3138 11294 3144 11306
rect 2660 11208 2666 11260
rect 2718 11248 2724 11260
rect 2718 11220 3798 11248
rect 2718 11208 2724 11220
rect 5162 10740 5168 10792
rect 5220 10740 5226 10792
rect 2744 10272 2750 10324
rect 2802 10312 2808 10324
rect 2802 10284 3798 10312
rect 2802 10272 2808 10284
rect 2996 10186 3002 10238
rect 3054 10226 3060 10238
rect 3054 10198 3894 10226
rect 3054 10186 3060 10198
rect 3416 10100 3422 10152
rect 3474 10140 3480 10152
rect 3474 10112 3990 10140
rect 3474 10100 3480 10112
rect 5104 10076 5180 10104
rect 2828 10014 2834 10066
rect 2886 10054 2892 10066
rect 2886 10026 4086 10054
rect 2886 10014 2892 10026
rect 168 9938 174 9990
rect 226 9978 232 9990
rect 616 9978 622 9990
rect 226 9950 622 9978
rect 226 9938 232 9950
rect 616 9938 622 9950
rect 674 9938 680 9990
rect 2407 9938 2413 9990
rect 2465 9938 2471 9990
rect 2996 9928 3002 9980
rect 3054 9968 3060 9980
rect 3054 9940 4182 9968
rect 3054 9928 3060 9940
rect 4896 9930 5180 9958
rect 3416 9842 3422 9894
rect 3474 9882 3480 9894
rect 3474 9854 4278 9882
rect 3474 9842 3480 9854
rect 4814 9808 5180 9836
rect 2912 9756 2918 9808
rect 2970 9796 2976 9808
rect 2970 9768 4482 9796
rect 2970 9756 2976 9768
rect 2996 9670 3002 9722
rect 3054 9710 3060 9722
rect 3054 9682 4578 9710
rect 3054 9670 3060 9682
rect 3416 9584 3422 9636
rect 3474 9624 3480 9636
rect 3474 9596 4674 9624
rect 3474 9584 3480 9596
rect 5162 9202 5168 9254
rect 5220 9202 5226 9254
rect 3416 8820 3422 8872
rect 3474 8860 3480 8872
rect 3474 8832 4674 8860
rect 3474 8820 3480 8832
rect 2996 8734 3002 8786
rect 3054 8774 3060 8786
rect 3054 8746 4578 8774
rect 3054 8734 3060 8746
rect 2660 8648 2666 8700
rect 2718 8688 2724 8700
rect 2718 8660 4482 8688
rect 2718 8648 2724 8660
rect 4814 8620 5180 8648
rect 3332 8562 3338 8614
rect 3390 8602 3396 8614
rect 3390 8574 4278 8602
rect 3390 8562 3396 8574
rect 3248 8476 3254 8528
rect 3306 8516 3312 8528
rect 3306 8488 4182 8516
rect 4896 8498 5180 8526
rect 3306 8476 3312 8488
rect 2912 8390 2918 8442
rect 2970 8430 2976 8442
rect 2970 8402 4086 8430
rect 2970 8390 2976 8402
rect 3332 8304 3338 8356
rect 3390 8344 3396 8356
rect 5104 8352 5180 8380
rect 3390 8316 3990 8344
rect 3390 8304 3396 8316
rect 3248 8218 3254 8270
rect 3306 8258 3312 8270
rect 3306 8230 3894 8258
rect 3306 8218 3312 8230
rect 2828 8132 2834 8184
rect 2886 8172 2892 8184
rect 2886 8144 3798 8172
rect 2886 8132 2892 8144
rect 5162 7664 5168 7716
rect 5220 7664 5226 7716
rect 2912 7196 2918 7248
rect 2970 7236 2976 7248
rect 2970 7208 3798 7236
rect 2970 7196 2976 7208
rect 3164 7110 3170 7162
rect 3222 7150 3228 7162
rect 3222 7122 3894 7150
rect 3222 7110 3228 7122
rect 3332 7024 3338 7076
rect 3390 7064 3396 7076
rect 3390 7036 3990 7064
rect 3390 7024 3396 7036
rect 5104 7000 5180 7028
rect 2660 6938 2666 6990
rect 2718 6978 2724 6990
rect 2718 6950 4086 6978
rect 2718 6938 2724 6950
rect 3248 6852 3254 6904
rect 3306 6892 3312 6904
rect 3306 6864 4182 6892
rect 3306 6852 3312 6864
rect 4896 6854 5180 6882
rect 3332 6766 3338 6818
rect 3390 6806 3396 6818
rect 3390 6778 4278 6806
rect 3390 6766 3396 6778
rect 4814 6732 5180 6760
rect 2744 6680 2750 6732
rect 2802 6720 2808 6732
rect 2802 6692 4482 6720
rect 2802 6680 2808 6692
rect 3248 6594 3254 6646
rect 3306 6634 3312 6646
rect 3306 6606 4578 6634
rect 3306 6594 3312 6606
rect 3332 6508 3338 6560
rect 3390 6548 3396 6560
rect 3390 6520 4674 6548
rect 3390 6508 3396 6520
rect 5162 6126 5168 6178
rect 5220 6126 5226 6178
rect 3332 5744 3338 5796
rect 3390 5784 3396 5796
rect 3390 5756 4674 5784
rect 3390 5744 3396 5756
rect 3164 5658 3170 5710
rect 3222 5698 3228 5710
rect 3222 5670 4578 5698
rect 3222 5658 3228 5670
rect 2828 5572 2834 5624
rect 2886 5612 2892 5624
rect 2886 5584 4482 5612
rect 2886 5572 2892 5584
rect 4814 5544 5180 5572
rect 3332 5486 3338 5538
rect 3390 5526 3396 5538
rect 3390 5498 4278 5526
rect 3390 5486 3396 5498
rect 2407 5406 2413 5458
rect 2465 5406 2471 5458
rect 3164 5400 3170 5452
rect 3222 5440 3228 5452
rect 3222 5412 4182 5440
rect 4896 5422 5180 5450
rect 3222 5400 3228 5412
rect 2744 5314 2750 5366
rect 2802 5354 2808 5366
rect 2802 5326 4086 5354
rect 2802 5314 2808 5326
rect 3332 5228 3338 5280
rect 3390 5268 3396 5280
rect 5104 5276 5180 5304
rect 3390 5240 3990 5268
rect 3390 5228 3396 5240
rect 3164 5142 3170 5194
rect 3222 5182 3228 5194
rect 3222 5154 3894 5182
rect 3222 5142 3228 5154
rect 2660 5056 2666 5108
rect 2718 5096 2724 5108
rect 2718 5068 3798 5096
rect 2718 5056 2724 5068
rect 5162 4588 5168 4640
rect 5220 4588 5226 4640
rect 2744 4120 2750 4172
rect 2802 4160 2808 4172
rect 2802 4132 3798 4160
rect 2802 4120 2808 4132
rect 3080 4034 3086 4086
rect 3138 4074 3144 4086
rect 3138 4046 3894 4074
rect 3138 4034 3144 4046
rect 3332 3948 3338 4000
rect 3390 3988 3396 4000
rect 3390 3960 3990 3988
rect 3390 3948 3396 3960
rect 5104 3924 5180 3952
rect 2828 3862 2834 3914
rect 2886 3902 2892 3914
rect 2886 3874 4086 3902
rect 2886 3862 2892 3874
rect 2407 3782 2413 3834
rect 2465 3782 2471 3834
rect 3080 3776 3086 3828
rect 3138 3816 3144 3828
rect 3138 3788 4182 3816
rect 3138 3776 3144 3788
rect 4896 3778 5180 3806
rect 3332 3690 3338 3742
rect 3390 3730 3396 3742
rect 3390 3702 4278 3730
rect 3390 3690 3396 3702
rect 4814 3656 5180 3684
rect 2912 3604 2918 3656
rect 2970 3644 2976 3656
rect 2970 3616 4482 3644
rect 2970 3604 2976 3616
rect 3080 3518 3086 3570
rect 3138 3558 3144 3570
rect 3138 3530 4578 3558
rect 3138 3518 3144 3530
rect 3332 3432 3338 3484
rect 3390 3472 3396 3484
rect 3390 3444 4674 3472
rect 3390 3432 3396 3444
rect 5162 3050 5168 3102
rect 5220 3050 5226 3102
rect 3332 2668 3338 2720
rect 3390 2708 3396 2720
rect 3390 2680 4674 2708
rect 3390 2668 3396 2680
rect 3080 2582 3086 2634
rect 3138 2622 3144 2634
rect 3138 2594 4578 2622
rect 3138 2582 3144 2594
rect 2660 2496 2666 2548
rect 2718 2536 2724 2548
rect 2718 2508 4482 2536
rect 2718 2496 2724 2508
rect 4814 2468 5180 2496
rect 3332 2410 3338 2462
rect 3390 2450 3396 2462
rect 3390 2422 4278 2450
rect 3390 2410 3396 2422
rect 84 2326 90 2378
rect 142 2366 148 2378
rect 700 2366 706 2378
rect 142 2338 706 2366
rect 142 2326 148 2338
rect 700 2326 706 2338
rect 758 2326 764 2378
rect 2407 2326 2413 2378
rect 2465 2326 2471 2378
rect 2996 2324 3002 2376
rect 3054 2364 3060 2376
rect 3054 2336 4182 2364
rect 4896 2346 5180 2374
rect 3054 2324 3060 2336
rect 2912 2238 2918 2290
rect 2970 2278 2976 2290
rect 2970 2250 4086 2278
rect 2970 2238 2976 2250
rect 3332 2152 3338 2204
rect 3390 2192 3396 2204
rect 5104 2200 5180 2228
rect 3390 2164 3990 2192
rect 3390 2152 3396 2164
rect 2996 2066 3002 2118
rect 3054 2106 3060 2118
rect 3054 2078 3894 2106
rect 3054 2066 3060 2078
rect 2828 1980 2834 2032
rect 2886 2020 2892 2032
rect 2886 1992 3798 2020
rect 2886 1980 2892 1992
rect 5162 1512 5168 1564
rect 5220 1512 5226 1564
rect 5104 848 5180 876
rect 2660 786 2666 838
rect 2718 826 2724 838
rect 2718 798 4086 826
rect 2718 786 2724 798
rect 0 702 6 754
rect 58 742 64 754
rect 616 742 622 754
rect 58 714 622 742
rect 58 702 64 714
rect 616 702 622 714
rect 674 702 680 754
rect 2407 702 2413 754
rect 2465 702 2471 754
rect 2996 700 3002 752
rect 3054 740 3060 752
rect 3054 712 4182 740
rect 3054 700 3060 712
rect 4896 702 5180 730
rect 3332 614 3338 666
rect 3390 654 3396 666
rect 3390 626 4278 654
rect 3390 614 3396 626
rect 4814 580 5180 608
rect 2744 528 2750 580
rect 2802 568 2808 580
rect 2802 540 4482 568
rect 2802 528 2808 540
rect 2996 442 3002 494
rect 3054 482 3060 494
rect 3054 454 4578 482
rect 3054 442 3060 454
rect 3332 356 3338 408
rect 3390 396 3396 408
rect 3390 368 4674 396
rect 3390 356 3396 368
rect 5162 -26 5168 26
rect 5220 -26 5226 26
<< via1 >>
rect 5168 24582 5220 24634
rect 3506 24200 3558 24252
rect 3254 24114 3306 24166
rect 2834 24028 2886 24080
rect 3506 23942 3558 23994
rect 2413 23921 2465 23930
rect 2413 23887 2422 23921
rect 2422 23887 2456 23921
rect 2456 23887 2465 23921
rect 2413 23878 2465 23887
rect 3254 23856 3306 23908
rect 2750 23770 2802 23822
rect 3506 23684 3558 23736
rect 3254 23598 3306 23650
rect 2666 23512 2718 23564
rect 5168 23044 5220 23096
rect 2750 22576 2802 22628
rect 3170 22490 3222 22542
rect 3506 22404 3558 22456
rect 2834 22318 2886 22370
rect 2413 22297 2465 22306
rect 2413 22263 2422 22297
rect 2422 22263 2456 22297
rect 2456 22263 2465 22297
rect 2413 22254 2465 22263
rect 3170 22232 3222 22284
rect 3506 22146 3558 22198
rect 2918 22060 2970 22112
rect 3170 21974 3222 22026
rect 3506 21888 3558 21940
rect 5168 21506 5220 21558
rect 3506 21124 3558 21176
rect 3170 21038 3222 21090
rect 2666 20952 2718 21004
rect 3506 20866 3558 20918
rect 426 20798 478 20850
rect 706 20798 758 20850
rect 2413 20841 2465 20850
rect 2413 20807 2422 20841
rect 2422 20807 2456 20841
rect 2456 20807 2465 20841
rect 2413 20798 2465 20807
rect 3086 20780 3138 20832
rect 2918 20694 2970 20746
rect 3506 20608 3558 20660
rect 3086 20522 3138 20574
rect 2834 20436 2886 20488
rect 5168 19968 5220 20020
rect 2918 19500 2970 19552
rect 3002 19414 3054 19466
rect 3506 19328 3558 19380
rect 2666 19242 2718 19294
rect 342 19174 394 19226
rect 622 19174 674 19226
rect 2413 19217 2465 19226
rect 2413 19183 2422 19217
rect 2422 19183 2456 19217
rect 2456 19183 2465 19217
rect 2413 19174 2465 19183
rect 3086 19156 3138 19208
rect 3506 19070 3558 19122
rect 2750 18984 2802 19036
rect 3086 18898 3138 18950
rect 3506 18812 3558 18864
rect 5168 18430 5220 18482
rect 3506 18048 3558 18100
rect 3002 17962 3054 18014
rect 2834 17876 2886 17928
rect 3506 17790 3558 17842
rect 3002 17704 3054 17756
rect 2750 17618 2802 17670
rect 3506 17532 3558 17584
rect 3002 17446 3054 17498
rect 2666 17360 2718 17412
rect 5168 16892 5220 16944
rect 2750 16424 2802 16476
rect 3254 16338 3306 16390
rect 3422 16252 3474 16304
rect 2834 16166 2886 16218
rect 3254 16080 3306 16132
rect 3422 15994 3474 16046
rect 2918 15908 2970 15960
rect 3254 15822 3306 15874
rect 3422 15736 3474 15788
rect 5168 15354 5220 15406
rect 3422 14972 3474 15024
rect 3254 14886 3306 14938
rect 2666 14800 2718 14852
rect 3422 14714 3474 14766
rect 2413 14685 2465 14694
rect 2413 14651 2422 14685
rect 2422 14651 2456 14685
rect 2456 14651 2465 14685
rect 2413 14642 2465 14651
rect 3170 14628 3222 14680
rect 2918 14542 2970 14594
rect 3422 14456 3474 14508
rect 3170 14370 3222 14422
rect 2834 14284 2886 14336
rect 5168 13816 5220 13868
rect 2918 13348 2970 13400
rect 3086 13262 3138 13314
rect 3422 13176 3474 13228
rect 2666 13090 2718 13142
rect 2413 13061 2465 13070
rect 2413 13027 2422 13061
rect 2422 13027 2456 13061
rect 2456 13027 2465 13061
rect 2413 13018 2465 13027
rect 3170 13004 3222 13056
rect 3422 12918 3474 12970
rect 2750 12832 2802 12884
rect 3170 12746 3222 12798
rect 3422 12660 3474 12712
rect 5168 12278 5220 12330
rect 3422 11896 3474 11948
rect 3086 11810 3138 11862
rect 2834 11724 2886 11776
rect 3422 11638 3474 11690
rect 258 11562 310 11614
rect 706 11562 758 11614
rect 2413 11605 2465 11614
rect 2413 11571 2422 11605
rect 2422 11571 2456 11605
rect 2456 11571 2465 11605
rect 2413 11562 2465 11571
rect 3086 11552 3138 11604
rect 2750 11466 2802 11518
rect 3422 11380 3474 11432
rect 3086 11294 3138 11346
rect 2666 11208 2718 11260
rect 5168 10740 5220 10792
rect 2750 10272 2802 10324
rect 3002 10186 3054 10238
rect 3422 10100 3474 10152
rect 2834 10014 2886 10066
rect 174 9938 226 9990
rect 622 9938 674 9990
rect 2413 9981 2465 9990
rect 2413 9947 2422 9981
rect 2422 9947 2456 9981
rect 2456 9947 2465 9981
rect 2413 9938 2465 9947
rect 3002 9928 3054 9980
rect 3422 9842 3474 9894
rect 2918 9756 2970 9808
rect 3002 9670 3054 9722
rect 3422 9584 3474 9636
rect 5168 9202 5220 9254
rect 3422 8820 3474 8872
rect 3002 8734 3054 8786
rect 2666 8648 2718 8700
rect 3338 8562 3390 8614
rect 3254 8476 3306 8528
rect 2918 8390 2970 8442
rect 3338 8304 3390 8356
rect 3254 8218 3306 8270
rect 2834 8132 2886 8184
rect 5168 7664 5220 7716
rect 2918 7196 2970 7248
rect 3170 7110 3222 7162
rect 3338 7024 3390 7076
rect 2666 6938 2718 6990
rect 3254 6852 3306 6904
rect 3338 6766 3390 6818
rect 2750 6680 2802 6732
rect 3254 6594 3306 6646
rect 3338 6508 3390 6560
rect 5168 6126 5220 6178
rect 3338 5744 3390 5796
rect 3170 5658 3222 5710
rect 2834 5572 2886 5624
rect 3338 5486 3390 5538
rect 2413 5449 2465 5458
rect 2413 5415 2422 5449
rect 2422 5415 2456 5449
rect 2456 5415 2465 5449
rect 2413 5406 2465 5415
rect 3170 5400 3222 5452
rect 2750 5314 2802 5366
rect 3338 5228 3390 5280
rect 3170 5142 3222 5194
rect 2666 5056 2718 5108
rect 5168 4588 5220 4640
rect 2750 4120 2802 4172
rect 3086 4034 3138 4086
rect 3338 3948 3390 4000
rect 2834 3862 2886 3914
rect 2413 3825 2465 3834
rect 2413 3791 2422 3825
rect 2422 3791 2456 3825
rect 2456 3791 2465 3825
rect 2413 3782 2465 3791
rect 3086 3776 3138 3828
rect 3338 3690 3390 3742
rect 2918 3604 2970 3656
rect 3086 3518 3138 3570
rect 3338 3432 3390 3484
rect 5168 3050 5220 3102
rect 3338 2668 3390 2720
rect 3086 2582 3138 2634
rect 2666 2496 2718 2548
rect 3338 2410 3390 2462
rect 90 2326 142 2378
rect 706 2326 758 2378
rect 2413 2369 2465 2378
rect 2413 2335 2422 2369
rect 2422 2335 2456 2369
rect 2456 2335 2465 2369
rect 2413 2326 2465 2335
rect 3002 2324 3054 2376
rect 2918 2238 2970 2290
rect 3338 2152 3390 2204
rect 3002 2066 3054 2118
rect 2834 1980 2886 2032
rect 5168 1512 5220 1564
rect 2666 786 2718 838
rect 6 702 58 754
rect 622 702 674 754
rect 2413 745 2465 754
rect 2413 711 2422 745
rect 2422 711 2456 745
rect 2456 711 2465 745
rect 2413 702 2465 711
rect 3002 700 3054 752
rect 3338 614 3390 666
rect 2750 528 2802 580
rect 3002 442 3054 494
rect 3338 356 3390 408
rect 5168 -26 5220 26
<< metal2 >>
rect 18 760 46 24632
rect 102 2384 130 24632
rect 186 9996 214 24632
rect 270 11620 298 24632
rect 354 19232 382 24632
rect 438 20856 466 24632
rect 2411 23932 2467 23941
rect 2411 23867 2467 23876
rect 2678 23570 2706 24660
rect 2762 23828 2790 24660
rect 2846 24086 2874 24660
rect 2834 24080 2886 24086
rect 2834 24022 2886 24028
rect 2750 23822 2802 23828
rect 2750 23764 2802 23770
rect 2666 23564 2718 23570
rect 2666 23506 2718 23512
rect 2411 22308 2467 22317
rect 2411 22243 2467 22252
rect 2678 21010 2706 23506
rect 2762 22634 2790 23764
rect 2750 22628 2802 22634
rect 2750 22570 2802 22576
rect 2666 21004 2718 21010
rect 2666 20946 2718 20952
rect 426 20850 478 20856
rect 426 20792 478 20798
rect 706 20850 758 20856
rect 706 20792 758 20798
rect 2411 20852 2467 20861
rect 342 19226 394 19232
rect 342 19168 394 19174
rect 258 11614 310 11620
rect 258 11556 310 11562
rect 174 9990 226 9996
rect 174 9932 226 9938
rect 90 2378 142 2384
rect 90 2320 142 2326
rect 6 754 58 760
rect 6 696 58 702
rect 18 0 46 696
rect 102 0 130 2320
rect 186 0 214 9932
rect 270 0 298 11556
rect 354 0 382 19168
rect 438 0 466 20792
rect 2411 20787 2467 20796
rect 2678 19300 2706 20946
rect 2666 19294 2718 19300
rect 622 19226 674 19232
rect 622 19168 674 19174
rect 2411 19228 2467 19237
rect 2666 19236 2718 19242
rect 2411 19163 2467 19172
rect 2678 17418 2706 19236
rect 2762 19042 2790 22570
rect 2846 22376 2874 24022
rect 2834 22370 2886 22376
rect 2834 22312 2886 22318
rect 2846 20494 2874 22312
rect 2930 22118 2958 24660
rect 2918 22112 2970 22118
rect 2918 22054 2970 22060
rect 2930 20752 2958 22054
rect 2918 20746 2970 20752
rect 2918 20688 2970 20694
rect 2834 20488 2886 20494
rect 2834 20430 2886 20436
rect 2750 19036 2802 19042
rect 2750 18978 2802 18984
rect 2762 17676 2790 18978
rect 2846 17934 2874 20430
rect 2930 19558 2958 20688
rect 2918 19552 2970 19558
rect 2918 19494 2970 19500
rect 2834 17928 2886 17934
rect 2834 17870 2886 17876
rect 2750 17670 2802 17676
rect 2750 17612 2802 17618
rect 2666 17412 2718 17418
rect 2666 17354 2718 17360
rect 2678 14858 2706 17354
rect 2762 16482 2790 17612
rect 2750 16476 2802 16482
rect 2750 16418 2802 16424
rect 2666 14852 2718 14858
rect 2666 14794 2718 14800
rect 2411 14696 2467 14705
rect 2411 14631 2467 14640
rect 2678 13148 2706 14794
rect 2666 13142 2718 13148
rect 2666 13084 2718 13090
rect 2411 13072 2467 13081
rect 2411 13007 2467 13016
rect 706 11614 758 11620
rect 706 11556 758 11562
rect 2411 11616 2467 11625
rect 2411 11551 2467 11560
rect 2678 11266 2706 13084
rect 2762 12890 2790 16418
rect 2846 16224 2874 17870
rect 2834 16218 2886 16224
rect 2834 16160 2886 16166
rect 2846 14342 2874 16160
rect 2930 15966 2958 19494
rect 3014 19472 3042 24660
rect 3098 20838 3126 24660
rect 3182 22548 3210 24660
rect 3266 24172 3294 24660
rect 3254 24166 3306 24172
rect 3254 24108 3306 24114
rect 3266 23914 3294 24108
rect 3254 23908 3306 23914
rect 3254 23850 3306 23856
rect 3266 23656 3294 23850
rect 3254 23650 3306 23656
rect 3254 23592 3306 23598
rect 3170 22542 3222 22548
rect 3170 22484 3222 22490
rect 3182 22290 3210 22484
rect 3170 22284 3222 22290
rect 3170 22226 3222 22232
rect 3182 22032 3210 22226
rect 3170 22026 3222 22032
rect 3170 21968 3222 21974
rect 3182 21096 3210 21968
rect 3170 21090 3222 21096
rect 3170 21032 3222 21038
rect 3086 20832 3138 20838
rect 3086 20774 3138 20780
rect 3098 20580 3126 20774
rect 3086 20574 3138 20580
rect 3086 20516 3138 20522
rect 3002 19466 3054 19472
rect 3002 19408 3054 19414
rect 3014 18020 3042 19408
rect 3098 19214 3126 20516
rect 3086 19208 3138 19214
rect 3086 19150 3138 19156
rect 3098 18956 3126 19150
rect 3086 18950 3138 18956
rect 3086 18892 3138 18898
rect 3002 18014 3054 18020
rect 3002 17956 3054 17962
rect 3014 17762 3042 17956
rect 3002 17756 3054 17762
rect 3002 17698 3054 17704
rect 3014 17504 3042 17698
rect 3002 17498 3054 17504
rect 3002 17440 3054 17446
rect 2918 15960 2970 15966
rect 2918 15902 2970 15908
rect 2930 14600 2958 15902
rect 2918 14594 2970 14600
rect 2918 14536 2970 14542
rect 2834 14336 2886 14342
rect 2834 14278 2886 14284
rect 2750 12884 2802 12890
rect 2750 12826 2802 12832
rect 2762 11524 2790 12826
rect 2846 11782 2874 14278
rect 2930 13406 2958 14536
rect 2918 13400 2970 13406
rect 2918 13342 2970 13348
rect 2834 11776 2886 11782
rect 2834 11718 2886 11724
rect 2750 11518 2802 11524
rect 2750 11460 2802 11466
rect 2666 11260 2718 11266
rect 2666 11202 2718 11208
rect 622 9990 674 9996
rect 622 9932 674 9938
rect 2411 9992 2467 10001
rect 2411 9927 2467 9936
rect 2678 8706 2706 11202
rect 2762 10330 2790 11460
rect 2750 10324 2802 10330
rect 2750 10266 2802 10272
rect 2666 8700 2718 8706
rect 2666 8642 2718 8648
rect 2678 6996 2706 8642
rect 2666 6990 2718 6996
rect 2666 6932 2718 6938
rect 2411 5460 2467 5469
rect 2411 5395 2467 5404
rect 2678 5114 2706 6932
rect 2762 6738 2790 10266
rect 2846 10072 2874 11718
rect 2834 10066 2886 10072
rect 2834 10008 2886 10014
rect 2846 8190 2874 10008
rect 2930 9814 2958 13342
rect 3014 10244 3042 17440
rect 3098 13320 3126 18892
rect 3182 14686 3210 21032
rect 3266 16396 3294 23592
rect 3350 18509 3378 24660
rect 3434 20049 3462 24660
rect 3518 24258 3546 24660
rect 3506 24252 3558 24258
rect 3506 24194 3558 24200
rect 3518 24000 3546 24194
rect 3506 23994 3558 24000
rect 3506 23936 3558 23942
rect 3518 23742 3546 23936
rect 3506 23736 3558 23742
rect 3506 23678 3558 23684
rect 3518 22462 3546 23678
rect 3602 23129 3630 24660
rect 5166 24636 5222 24645
rect 5166 24571 5222 24580
rect 3588 23120 3644 23129
rect 3588 23055 3644 23064
rect 5166 23098 5222 23107
rect 3506 22456 3558 22462
rect 3506 22398 3558 22404
rect 3518 22204 3546 22398
rect 3506 22198 3558 22204
rect 3506 22140 3558 22146
rect 3518 21946 3546 22140
rect 3506 21940 3558 21946
rect 3506 21882 3558 21888
rect 3518 21589 3546 21882
rect 3504 21580 3560 21589
rect 3504 21515 3560 21524
rect 3518 21182 3546 21515
rect 3506 21176 3558 21182
rect 3506 21118 3558 21124
rect 3518 20924 3546 21118
rect 3506 20918 3558 20924
rect 3506 20860 3558 20866
rect 3518 20666 3546 20860
rect 3506 20660 3558 20666
rect 3506 20602 3558 20608
rect 3420 20040 3476 20049
rect 3420 19975 3476 19984
rect 3336 18500 3392 18509
rect 3336 18435 3392 18444
rect 3254 16390 3306 16396
rect 3254 16332 3306 16338
rect 3266 16138 3294 16332
rect 3254 16132 3306 16138
rect 3254 16074 3306 16080
rect 3266 15880 3294 16074
rect 3254 15874 3306 15880
rect 3254 15816 3306 15822
rect 3266 14944 3294 15816
rect 3254 14938 3306 14944
rect 3254 14880 3306 14886
rect 3170 14680 3222 14686
rect 3170 14622 3222 14628
rect 3182 14428 3210 14622
rect 3170 14422 3222 14428
rect 3170 14364 3222 14370
rect 3086 13314 3138 13320
rect 3086 13256 3138 13262
rect 3098 11868 3126 13256
rect 3182 13062 3210 14364
rect 3266 13893 3294 14880
rect 3252 13884 3308 13893
rect 3252 13819 3308 13828
rect 3170 13056 3222 13062
rect 3170 12998 3222 13004
rect 3182 12804 3210 12998
rect 3170 12798 3222 12804
rect 3170 12740 3222 12746
rect 3182 12353 3210 12740
rect 3168 12344 3224 12353
rect 3168 12279 3224 12288
rect 3086 11862 3138 11868
rect 3086 11804 3138 11810
rect 3098 11610 3126 11804
rect 3086 11604 3138 11610
rect 3086 11546 3138 11552
rect 3098 11352 3126 11546
rect 3086 11346 3138 11352
rect 3086 11288 3138 11294
rect 3098 10813 3126 11288
rect 3084 10804 3140 10813
rect 3084 10739 3140 10748
rect 3002 10238 3054 10244
rect 3002 10180 3054 10186
rect 3014 9986 3042 10180
rect 3002 9980 3054 9986
rect 3002 9922 3054 9928
rect 2918 9808 2970 9814
rect 2918 9750 2970 9756
rect 2930 8448 2958 9750
rect 3014 9728 3042 9922
rect 3002 9722 3054 9728
rect 3002 9664 3054 9670
rect 3014 9273 3042 9664
rect 3000 9264 3056 9273
rect 3000 9199 3056 9208
rect 3014 8792 3042 9199
rect 3002 8786 3054 8792
rect 3002 8728 3054 8734
rect 2918 8442 2970 8448
rect 2918 8384 2970 8390
rect 2834 8184 2886 8190
rect 2834 8126 2886 8132
rect 2750 6732 2802 6738
rect 2750 6674 2802 6680
rect 2762 5372 2790 6674
rect 2846 5630 2874 8126
rect 2930 7254 2958 8384
rect 2918 7248 2970 7254
rect 2918 7190 2970 7196
rect 2834 5624 2886 5630
rect 2834 5566 2886 5572
rect 2750 5366 2802 5372
rect 2750 5308 2802 5314
rect 2666 5108 2718 5114
rect 2666 5050 2718 5056
rect 2411 3836 2467 3845
rect 2411 3771 2467 3780
rect 2678 2554 2706 5050
rect 2762 4178 2790 5308
rect 2750 4172 2802 4178
rect 2750 4114 2802 4120
rect 2666 2548 2718 2554
rect 2666 2490 2718 2496
rect 706 2378 758 2384
rect 706 2320 758 2326
rect 2411 2380 2467 2389
rect 2411 2315 2467 2324
rect 2678 844 2706 2490
rect 2762 1577 2790 4114
rect 2846 3920 2874 5566
rect 2930 4657 2958 7190
rect 2916 4648 2972 4657
rect 2916 4583 2972 4592
rect 2834 3914 2886 3920
rect 2834 3856 2886 3862
rect 2846 3117 2874 3856
rect 2930 3662 2958 4583
rect 2918 3656 2970 3662
rect 2918 3598 2970 3604
rect 2832 3108 2888 3117
rect 2832 3043 2888 3052
rect 2846 2038 2874 3043
rect 2930 2296 2958 3598
rect 3014 2382 3042 8728
rect 3098 4092 3126 10739
rect 3182 7168 3210 12279
rect 3266 8534 3294 13819
rect 3350 8620 3378 18435
rect 3434 16310 3462 19975
rect 3518 19386 3546 20602
rect 3506 19380 3558 19386
rect 3506 19322 3558 19328
rect 3518 19128 3546 19322
rect 3506 19122 3558 19128
rect 3506 19064 3558 19070
rect 3518 18870 3546 19064
rect 3506 18864 3558 18870
rect 3506 18806 3558 18812
rect 3518 18106 3546 18806
rect 3506 18100 3558 18106
rect 3506 18042 3558 18048
rect 3518 17848 3546 18042
rect 3506 17842 3558 17848
rect 3506 17784 3558 17790
rect 3518 17590 3546 17784
rect 3506 17584 3558 17590
rect 3506 17526 3558 17532
rect 3422 16304 3474 16310
rect 3422 16246 3474 16252
rect 3434 16052 3462 16246
rect 3422 16046 3474 16052
rect 3422 15988 3474 15994
rect 3434 15794 3462 15988
rect 3422 15788 3474 15794
rect 3422 15730 3474 15736
rect 3434 15030 3462 15730
rect 3422 15024 3474 15030
rect 3422 14966 3474 14972
rect 3434 14772 3462 14966
rect 3422 14766 3474 14772
rect 3422 14708 3474 14714
rect 3434 14514 3462 14708
rect 3422 14508 3474 14514
rect 3422 14450 3474 14456
rect 3434 13234 3462 14450
rect 3422 13228 3474 13234
rect 3422 13170 3474 13176
rect 3434 12976 3462 13170
rect 3422 12970 3474 12976
rect 3422 12912 3474 12918
rect 3434 12718 3462 12912
rect 3422 12712 3474 12718
rect 3422 12654 3474 12660
rect 3434 11954 3462 12654
rect 3422 11948 3474 11954
rect 3422 11890 3474 11896
rect 3434 11696 3462 11890
rect 3422 11690 3474 11696
rect 3422 11632 3474 11638
rect 3434 11438 3462 11632
rect 3422 11432 3474 11438
rect 3422 11374 3474 11380
rect 3434 10158 3462 11374
rect 3422 10152 3474 10158
rect 3422 10094 3474 10100
rect 3434 9900 3462 10094
rect 3422 9894 3474 9900
rect 3422 9836 3474 9842
rect 3434 9642 3462 9836
rect 3422 9636 3474 9642
rect 3422 9578 3474 9584
rect 3434 8878 3462 9578
rect 3422 8872 3474 8878
rect 3422 8814 3474 8820
rect 3338 8614 3390 8620
rect 3338 8556 3390 8562
rect 3254 8528 3306 8534
rect 3254 8470 3306 8476
rect 3266 8276 3294 8470
rect 3350 8362 3378 8556
rect 3338 8356 3390 8362
rect 3338 8298 3390 8304
rect 3254 8270 3306 8276
rect 3254 8212 3306 8218
rect 3170 7162 3222 7168
rect 3170 7104 3222 7110
rect 3182 5716 3210 7104
rect 3266 6910 3294 8212
rect 3350 7082 3378 8298
rect 3338 7076 3390 7082
rect 3338 7018 3390 7024
rect 3254 6904 3306 6910
rect 3254 6846 3306 6852
rect 3266 6652 3294 6846
rect 3350 6824 3378 7018
rect 3338 6818 3390 6824
rect 3338 6760 3390 6766
rect 3254 6646 3306 6652
rect 3254 6588 3306 6594
rect 3170 5710 3222 5716
rect 3170 5652 3222 5658
rect 3182 5458 3210 5652
rect 3170 5452 3222 5458
rect 3170 5394 3222 5400
rect 3182 5200 3210 5394
rect 3170 5194 3222 5200
rect 3170 5136 3222 5142
rect 3086 4086 3138 4092
rect 3086 4028 3138 4034
rect 3098 3834 3126 4028
rect 3086 3828 3138 3834
rect 3086 3770 3138 3776
rect 3098 3576 3126 3770
rect 3086 3570 3138 3576
rect 3086 3512 3138 3518
rect 3098 2640 3126 3512
rect 3086 2634 3138 2640
rect 3086 2576 3138 2582
rect 3002 2376 3054 2382
rect 3002 2318 3054 2324
rect 2918 2290 2970 2296
rect 2918 2232 2970 2238
rect 2834 2032 2886 2038
rect 2834 1974 2886 1980
rect 2748 1568 2804 1577
rect 2748 1503 2804 1512
rect 2666 838 2718 844
rect 2666 780 2718 786
rect 622 754 674 760
rect 622 696 674 702
rect 2411 756 2467 765
rect 2411 691 2467 700
rect 2678 37 2706 780
rect 2762 586 2790 1503
rect 2750 580 2802 586
rect 2750 522 2802 528
rect 2664 28 2720 37
rect 2762 0 2790 522
rect 2846 0 2874 1974
rect 2930 0 2958 2232
rect 3014 2124 3042 2318
rect 3002 2118 3054 2124
rect 3002 2060 3054 2066
rect 3014 758 3042 2060
rect 3002 752 3054 758
rect 3002 694 3054 700
rect 3014 500 3042 694
rect 3002 494 3054 500
rect 3002 436 3054 442
rect 3014 0 3042 436
rect 3098 0 3126 2576
rect 3182 0 3210 5136
rect 3266 0 3294 6588
rect 3350 6566 3378 6760
rect 3338 6560 3390 6566
rect 3338 6502 3390 6508
rect 3350 5802 3378 6502
rect 3338 5796 3390 5802
rect 3338 5738 3390 5744
rect 3350 5544 3378 5738
rect 3338 5538 3390 5544
rect 3338 5480 3390 5486
rect 3350 5286 3378 5480
rect 3338 5280 3390 5286
rect 3338 5222 3390 5228
rect 3350 4006 3378 5222
rect 3338 4000 3390 4006
rect 3338 3942 3390 3948
rect 3350 3748 3378 3942
rect 3338 3742 3390 3748
rect 3338 3684 3390 3690
rect 3350 3490 3378 3684
rect 3338 3484 3390 3490
rect 3338 3426 3390 3432
rect 3350 2726 3378 3426
rect 3338 2720 3390 2726
rect 3338 2662 3390 2668
rect 3350 2468 3378 2662
rect 3338 2462 3390 2468
rect 3338 2404 3390 2410
rect 3350 2210 3378 2404
rect 3338 2204 3390 2210
rect 3338 2146 3390 2152
rect 3350 672 3378 2146
rect 3338 666 3390 672
rect 3338 608 3390 614
rect 3350 414 3378 608
rect 3338 408 3390 414
rect 3338 350 3390 356
rect 3350 0 3378 350
rect 3434 0 3462 8814
rect 3518 0 3546 17526
rect 3602 0 3630 23055
rect 5166 23033 5222 23042
rect 5166 21560 5222 21569
rect 5166 21495 5222 21504
rect 5166 20022 5222 20031
rect 5166 19957 5222 19966
rect 5166 18484 5222 18493
rect 5166 18419 5222 18428
rect 5166 16946 5222 16955
rect 5166 16881 5222 16890
rect 5166 15408 5222 15417
rect 5166 15343 5222 15352
rect 5166 13870 5222 13879
rect 5166 13805 5222 13814
rect 5166 12332 5222 12341
rect 5166 12267 5222 12276
rect 5166 10794 5222 10803
rect 5166 10729 5222 10738
rect 5166 9256 5222 9265
rect 5166 9191 5222 9200
rect 5166 7718 5222 7727
rect 5166 7653 5222 7662
rect 5166 6180 5222 6189
rect 5166 6115 5222 6124
rect 5166 4642 5222 4651
rect 5166 4577 5222 4586
rect 5166 3104 5222 3113
rect 5166 3039 5222 3048
rect 5166 1566 5222 1575
rect 5166 1501 5222 1510
rect 5166 28 5222 37
rect 2664 -37 2720 -28
rect 5166 -37 5222 -28
<< via2 >>
rect 2411 23930 2467 23932
rect 2411 23878 2413 23930
rect 2413 23878 2465 23930
rect 2465 23878 2467 23930
rect 2411 23876 2467 23878
rect 2411 22306 2467 22308
rect 2411 22254 2413 22306
rect 2413 22254 2465 22306
rect 2465 22254 2467 22306
rect 2411 22252 2467 22254
rect 2411 20850 2467 20852
rect 2411 20798 2413 20850
rect 2413 20798 2465 20850
rect 2465 20798 2467 20850
rect 2411 20796 2467 20798
rect 2411 19226 2467 19228
rect 2411 19174 2413 19226
rect 2413 19174 2465 19226
rect 2465 19174 2467 19226
rect 2411 19172 2467 19174
rect 2411 14694 2467 14696
rect 2411 14642 2413 14694
rect 2413 14642 2465 14694
rect 2465 14642 2467 14694
rect 2411 14640 2467 14642
rect 2411 13070 2467 13072
rect 2411 13018 2413 13070
rect 2413 13018 2465 13070
rect 2465 13018 2467 13070
rect 2411 13016 2467 13018
rect 2411 11614 2467 11616
rect 2411 11562 2413 11614
rect 2413 11562 2465 11614
rect 2465 11562 2467 11614
rect 2411 11560 2467 11562
rect 2411 9990 2467 9992
rect 2411 9938 2413 9990
rect 2413 9938 2465 9990
rect 2465 9938 2467 9990
rect 2411 9936 2467 9938
rect 2411 5458 2467 5460
rect 2411 5406 2413 5458
rect 2413 5406 2465 5458
rect 2465 5406 2467 5458
rect 2411 5404 2467 5406
rect 5166 24634 5222 24636
rect 5166 24582 5168 24634
rect 5168 24582 5220 24634
rect 5220 24582 5222 24634
rect 5166 24580 5222 24582
rect 3588 23064 3644 23120
rect 5166 23096 5222 23098
rect 3504 21524 3560 21580
rect 3420 19984 3476 20040
rect 3336 18444 3392 18500
rect 3252 13828 3308 13884
rect 3168 12288 3224 12344
rect 3084 10748 3140 10804
rect 3000 9208 3056 9264
rect 2411 3834 2467 3836
rect 2411 3782 2413 3834
rect 2413 3782 2465 3834
rect 2465 3782 2467 3834
rect 2411 3780 2467 3782
rect 2411 2378 2467 2380
rect 2411 2326 2413 2378
rect 2413 2326 2465 2378
rect 2465 2326 2467 2378
rect 2411 2324 2467 2326
rect 2916 4592 2972 4648
rect 2832 3052 2888 3108
rect 2748 1512 2804 1568
rect 2411 754 2467 756
rect 2411 702 2413 754
rect 2413 702 2465 754
rect 2465 702 2467 754
rect 2411 700 2467 702
rect 2664 -28 2720 28
rect 5166 23044 5168 23096
rect 5168 23044 5220 23096
rect 5220 23044 5222 23096
rect 5166 23042 5222 23044
rect 5166 21558 5222 21560
rect 5166 21506 5168 21558
rect 5168 21506 5220 21558
rect 5220 21506 5222 21558
rect 5166 21504 5222 21506
rect 5166 20020 5222 20022
rect 5166 19968 5168 20020
rect 5168 19968 5220 20020
rect 5220 19968 5222 20020
rect 5166 19966 5222 19968
rect 5166 18482 5222 18484
rect 5166 18430 5168 18482
rect 5168 18430 5220 18482
rect 5220 18430 5222 18482
rect 5166 18428 5222 18430
rect 5166 16944 5222 16946
rect 5166 16892 5168 16944
rect 5168 16892 5220 16944
rect 5220 16892 5222 16944
rect 5166 16890 5222 16892
rect 5166 15406 5222 15408
rect 5166 15354 5168 15406
rect 5168 15354 5220 15406
rect 5220 15354 5222 15406
rect 5166 15352 5222 15354
rect 5166 13868 5222 13870
rect 5166 13816 5168 13868
rect 5168 13816 5220 13868
rect 5220 13816 5222 13868
rect 5166 13814 5222 13816
rect 5166 12330 5222 12332
rect 5166 12278 5168 12330
rect 5168 12278 5220 12330
rect 5220 12278 5222 12330
rect 5166 12276 5222 12278
rect 5166 10792 5222 10794
rect 5166 10740 5168 10792
rect 5168 10740 5220 10792
rect 5220 10740 5222 10792
rect 5166 10738 5222 10740
rect 5166 9254 5222 9256
rect 5166 9202 5168 9254
rect 5168 9202 5220 9254
rect 5220 9202 5222 9254
rect 5166 9200 5222 9202
rect 5166 7716 5222 7718
rect 5166 7664 5168 7716
rect 5168 7664 5220 7716
rect 5220 7664 5222 7716
rect 5166 7662 5222 7664
rect 5166 6178 5222 6180
rect 5166 6126 5168 6178
rect 5168 6126 5220 6178
rect 5220 6126 5222 6178
rect 5166 6124 5222 6126
rect 5166 4640 5222 4642
rect 5166 4588 5168 4640
rect 5168 4588 5220 4640
rect 5220 4588 5222 4640
rect 5166 4586 5222 4588
rect 5166 3102 5222 3104
rect 5166 3050 5168 3102
rect 5168 3050 5220 3102
rect 5220 3050 5222 3102
rect 5166 3048 5222 3050
rect 5166 1564 5222 1566
rect 5166 1512 5168 1564
rect 5168 1512 5220 1564
rect 5220 1512 5222 1564
rect 5166 1510 5222 1512
rect 5166 26 5222 28
rect 5166 -26 5168 26
rect 5168 -26 5220 26
rect 5220 -26 5222 26
rect 5166 -28 5222 -26
<< metal3 >>
rect 792 24595 924 24669
rect 1664 24595 1796 24669
rect 5128 24636 5260 24645
rect 5128 24580 5166 24636
rect 5222 24580 5260 24636
rect 5128 24571 5260 24580
rect 2373 23932 2505 23937
rect 2373 23876 2411 23932
rect 2467 23876 2505 23932
rect 2373 23871 2505 23876
rect 792 23055 924 23129
rect 1664 23055 1796 23129
rect 2409 23122 2469 23871
rect 3550 23122 3682 23125
rect 2409 23120 3682 23122
rect 2409 23064 3588 23120
rect 3644 23064 3682 23120
rect 2409 23062 3682 23064
rect 3550 23059 3682 23062
rect 5128 23098 5260 23107
rect 5128 23042 5166 23098
rect 5222 23042 5260 23098
rect 5128 23033 5260 23042
rect 2373 22308 2505 22313
rect 2373 22252 2411 22308
rect 2467 22252 2505 22308
rect 2373 22247 2505 22252
rect 792 21515 924 21589
rect 1664 21515 1796 21589
rect 2409 21582 2469 22247
rect 3466 21582 3598 21585
rect 2409 21580 3598 21582
rect 2409 21524 3504 21580
rect 3560 21524 3598 21580
rect 2409 21522 3598 21524
rect 3466 21519 3598 21522
rect 5128 21560 5260 21569
rect 5128 21504 5166 21560
rect 5222 21504 5260 21560
rect 5128 21495 5260 21504
rect 2373 20852 2505 20857
rect 2373 20796 2411 20852
rect 2467 20796 2505 20852
rect 2373 20791 2505 20796
rect 792 19975 924 20049
rect 1664 19975 1796 20049
rect 2409 20042 2469 20791
rect 3382 20042 3514 20045
rect 2409 20040 3514 20042
rect 2409 19984 3420 20040
rect 3476 19984 3514 20040
rect 2409 19982 3514 19984
rect 3382 19979 3514 19982
rect 5128 20022 5260 20031
rect 5128 19966 5166 20022
rect 5222 19966 5260 20022
rect 5128 19957 5260 19966
rect 2373 19228 2505 19233
rect 2373 19172 2411 19228
rect 2467 19172 2505 19228
rect 2373 19167 2505 19172
rect 792 18435 924 18509
rect 1664 18435 1796 18509
rect 2409 18502 2469 19167
rect 3298 18502 3430 18505
rect 2409 18500 3430 18502
rect 2409 18444 3336 18500
rect 3392 18444 3430 18500
rect 2409 18442 3430 18444
rect 3298 18439 3430 18442
rect 5128 18484 5260 18493
rect 5128 18428 5166 18484
rect 5222 18428 5260 18484
rect 5128 18419 5260 18428
rect 5128 16946 5260 16955
rect 5128 16890 5166 16946
rect 5222 16890 5260 16946
rect 5128 16881 5260 16890
rect 792 15359 924 15433
rect 1664 15359 1796 15433
rect 5128 15408 5260 15417
rect 5128 15352 5166 15408
rect 5222 15352 5260 15408
rect 5128 15343 5260 15352
rect 2373 14696 2505 14701
rect 2373 14640 2411 14696
rect 2467 14640 2505 14696
rect 2373 14635 2505 14640
rect 792 13819 924 13893
rect 1664 13819 1796 13893
rect 2409 13886 2469 14635
rect 3214 13886 3346 13889
rect 2409 13884 3346 13886
rect 2409 13828 3252 13884
rect 3308 13828 3346 13884
rect 2409 13826 3346 13828
rect 3214 13823 3346 13826
rect 5128 13870 5260 13879
rect 5128 13814 5166 13870
rect 5222 13814 5260 13870
rect 5128 13805 5260 13814
rect 2373 13072 2505 13077
rect 2373 13016 2411 13072
rect 2467 13016 2505 13072
rect 2373 13011 2505 13016
rect 792 12279 924 12353
rect 1664 12279 1796 12353
rect 2409 12346 2469 13011
rect 3130 12346 3262 12349
rect 2409 12344 3262 12346
rect 2409 12288 3168 12344
rect 3224 12288 3262 12344
rect 2409 12286 3262 12288
rect 3130 12283 3262 12286
rect 5128 12332 5260 12341
rect 5128 12276 5166 12332
rect 5222 12276 5260 12332
rect 5128 12267 5260 12276
rect 2373 11616 2505 11621
rect 2373 11560 2411 11616
rect 2467 11560 2505 11616
rect 2373 11555 2505 11560
rect 792 10739 924 10813
rect 1664 10739 1796 10813
rect 2409 10806 2469 11555
rect 3046 10806 3178 10809
rect 2409 10804 3178 10806
rect 2409 10748 3084 10804
rect 3140 10748 3178 10804
rect 2409 10746 3178 10748
rect 3046 10743 3178 10746
rect 5128 10794 5260 10803
rect 5128 10738 5166 10794
rect 5222 10738 5260 10794
rect 5128 10729 5260 10738
rect 2373 9992 2505 9997
rect 2373 9936 2411 9992
rect 2467 9936 2505 9992
rect 2373 9931 2505 9936
rect 792 9199 924 9273
rect 1664 9199 1796 9273
rect 2409 9266 2469 9931
rect 2962 9266 3094 9269
rect 2409 9264 3094 9266
rect 2409 9208 3000 9264
rect 3056 9208 3094 9264
rect 2409 9206 3094 9208
rect 2962 9203 3094 9206
rect 5128 9256 5260 9265
rect 5128 9200 5166 9256
rect 5222 9200 5260 9256
rect 5128 9191 5260 9200
rect 5128 7718 5260 7727
rect 5128 7662 5166 7718
rect 5222 7662 5260 7718
rect 5128 7653 5260 7662
rect 792 6123 924 6197
rect 1664 6123 1796 6197
rect 5128 6180 5260 6189
rect 5128 6124 5166 6180
rect 5222 6124 5260 6180
rect 5128 6115 5260 6124
rect 2373 5460 2505 5465
rect 2373 5404 2411 5460
rect 2467 5404 2505 5460
rect 2373 5399 2505 5404
rect 792 4583 924 4657
rect 1664 4583 1796 4657
rect 2409 4650 2469 5399
rect 2878 4650 3010 4653
rect 2409 4648 3010 4650
rect 2409 4592 2916 4648
rect 2972 4592 3010 4648
rect 2409 4590 3010 4592
rect 2878 4587 3010 4590
rect 5128 4642 5260 4651
rect 5128 4586 5166 4642
rect 5222 4586 5260 4642
rect 5128 4577 5260 4586
rect 2373 3836 2505 3841
rect 2373 3780 2411 3836
rect 2467 3780 2505 3836
rect 2373 3775 2505 3780
rect 792 3043 924 3117
rect 1664 3043 1796 3117
rect 2409 3110 2469 3775
rect 2794 3110 2926 3113
rect 2409 3108 2926 3110
rect 2409 3052 2832 3108
rect 2888 3052 2926 3108
rect 2409 3050 2926 3052
rect 2794 3047 2926 3050
rect 5128 3104 5260 3113
rect 5128 3048 5166 3104
rect 5222 3048 5260 3104
rect 5128 3039 5260 3048
rect 2373 2380 2505 2385
rect 2373 2324 2411 2380
rect 2467 2324 2505 2380
rect 2373 2319 2505 2324
rect 792 1503 924 1577
rect 1664 1503 1796 1577
rect 2409 1570 2469 2319
rect 2710 1570 2842 1573
rect 2409 1568 2842 1570
rect 2409 1512 2748 1568
rect 2804 1512 2842 1568
rect 2409 1510 2842 1512
rect 2710 1507 2842 1510
rect 5128 1566 5260 1575
rect 5128 1510 5166 1566
rect 5222 1510 5260 1566
rect 5128 1501 5260 1510
rect 2373 756 2505 761
rect 2373 700 2411 756
rect 2467 700 2505 756
rect 2373 695 2505 700
rect 792 -37 924 37
rect 1664 -37 1796 37
rect 2409 30 2469 695
rect 2626 30 2758 33
rect 2409 28 2758 30
rect 2409 -28 2664 28
rect 2720 -28 2758 28
rect 2409 -30 2758 -28
rect 2626 -33 2758 -30
rect 5128 28 5260 37
rect 5128 -28 5166 28
rect 5222 -28 5260 28
rect 5128 -37 5260 -28
use contact_18  contact_18_0
timestamp 1644949024
transform 1 0 5128 0 1 24571
box 0 0 1 1
use contact_17  contact_17_0
timestamp 1644949024
transform 1 0 5162 0 1 24576
box 0 0 1 1
use contact_18  contact_18_1
timestamp 1644949024
transform 1 0 5128 0 1 23033
box 0 0 1 1
use contact_17  contact_17_1
timestamp 1644949024
transform 1 0 5162 0 1 23038
box 0 0 1 1
use contact_18  contact_18_2
timestamp 1644949024
transform 1 0 5128 0 1 21495
box 0 0 1 1
use contact_17  contact_17_2
timestamp 1644949024
transform 1 0 5162 0 1 21500
box 0 0 1 1
use contact_18  contact_18_3
timestamp 1644949024
transform 1 0 5128 0 1 23033
box 0 0 1 1
use contact_17  contact_17_3
timestamp 1644949024
transform 1 0 5162 0 1 23038
box 0 0 1 1
use contact_18  contact_18_4
timestamp 1644949024
transform 1 0 5128 0 1 21495
box 0 0 1 1
use contact_17  contact_17_4
timestamp 1644949024
transform 1 0 5162 0 1 21500
box 0 0 1 1
use contact_18  contact_18_5
timestamp 1644949024
transform 1 0 5128 0 1 19957
box 0 0 1 1
use contact_17  contact_17_5
timestamp 1644949024
transform 1 0 5162 0 1 19962
box 0 0 1 1
use contact_18  contact_18_6
timestamp 1644949024
transform 1 0 5128 0 1 18419
box 0 0 1 1
use contact_17  contact_17_6
timestamp 1644949024
transform 1 0 5162 0 1 18424
box 0 0 1 1
use contact_18  contact_18_7
timestamp 1644949024
transform 1 0 5128 0 1 19957
box 0 0 1 1
use contact_17  contact_17_7
timestamp 1644949024
transform 1 0 5162 0 1 19962
box 0 0 1 1
use contact_18  contact_18_8
timestamp 1644949024
transform 1 0 5128 0 1 18419
box 0 0 1 1
use contact_17  contact_17_8
timestamp 1644949024
transform 1 0 5162 0 1 18424
box 0 0 1 1
use contact_18  contact_18_9
timestamp 1644949024
transform 1 0 5128 0 1 16881
box 0 0 1 1
use contact_17  contact_17_9
timestamp 1644949024
transform 1 0 5162 0 1 16886
box 0 0 1 1
use contact_18  contact_18_10
timestamp 1644949024
transform 1 0 5128 0 1 15343
box 0 0 1 1
use contact_17  contact_17_10
timestamp 1644949024
transform 1 0 5162 0 1 15348
box 0 0 1 1
use contact_18  contact_18_11
timestamp 1644949024
transform 1 0 5128 0 1 16881
box 0 0 1 1
use contact_17  contact_17_11
timestamp 1644949024
transform 1 0 5162 0 1 16886
box 0 0 1 1
use contact_18  contact_18_12
timestamp 1644949024
transform 1 0 5128 0 1 15343
box 0 0 1 1
use contact_17  contact_17_12
timestamp 1644949024
transform 1 0 5162 0 1 15348
box 0 0 1 1
use contact_18  contact_18_13
timestamp 1644949024
transform 1 0 5128 0 1 13805
box 0 0 1 1
use contact_17  contact_17_13
timestamp 1644949024
transform 1 0 5162 0 1 13810
box 0 0 1 1
use contact_18  contact_18_14
timestamp 1644949024
transform 1 0 5128 0 1 12267
box 0 0 1 1
use contact_17  contact_17_14
timestamp 1644949024
transform 1 0 5162 0 1 12272
box 0 0 1 1
use contact_18  contact_18_15
timestamp 1644949024
transform 1 0 5128 0 1 13805
box 0 0 1 1
use contact_17  contact_17_15
timestamp 1644949024
transform 1 0 5162 0 1 13810
box 0 0 1 1
use contact_18  contact_18_16
timestamp 1644949024
transform 1 0 5128 0 1 12267
box 0 0 1 1
use contact_17  contact_17_16
timestamp 1644949024
transform 1 0 5162 0 1 12272
box 0 0 1 1
use contact_18  contact_18_17
timestamp 1644949024
transform 1 0 5128 0 1 10729
box 0 0 1 1
use contact_17  contact_17_17
timestamp 1644949024
transform 1 0 5162 0 1 10734
box 0 0 1 1
use contact_18  contact_18_18
timestamp 1644949024
transform 1 0 5128 0 1 9191
box 0 0 1 1
use contact_17  contact_17_18
timestamp 1644949024
transform 1 0 5162 0 1 9196
box 0 0 1 1
use contact_18  contact_18_19
timestamp 1644949024
transform 1 0 5128 0 1 10729
box 0 0 1 1
use contact_17  contact_17_19
timestamp 1644949024
transform 1 0 5162 0 1 10734
box 0 0 1 1
use contact_18  contact_18_20
timestamp 1644949024
transform 1 0 5128 0 1 9191
box 0 0 1 1
use contact_17  contact_17_20
timestamp 1644949024
transform 1 0 5162 0 1 9196
box 0 0 1 1
use contact_18  contact_18_21
timestamp 1644949024
transform 1 0 5128 0 1 7653
box 0 0 1 1
use contact_17  contact_17_21
timestamp 1644949024
transform 1 0 5162 0 1 7658
box 0 0 1 1
use contact_18  contact_18_22
timestamp 1644949024
transform 1 0 5128 0 1 6115
box 0 0 1 1
use contact_17  contact_17_22
timestamp 1644949024
transform 1 0 5162 0 1 6120
box 0 0 1 1
use contact_18  contact_18_23
timestamp 1644949024
transform 1 0 5128 0 1 7653
box 0 0 1 1
use contact_17  contact_17_23
timestamp 1644949024
transform 1 0 5162 0 1 7658
box 0 0 1 1
use contact_18  contact_18_24
timestamp 1644949024
transform 1 0 5128 0 1 6115
box 0 0 1 1
use contact_17  contact_17_24
timestamp 1644949024
transform 1 0 5162 0 1 6120
box 0 0 1 1
use contact_18  contact_18_25
timestamp 1644949024
transform 1 0 5128 0 1 4577
box 0 0 1 1
use contact_17  contact_17_25
timestamp 1644949024
transform 1 0 5162 0 1 4582
box 0 0 1 1
use contact_18  contact_18_26
timestamp 1644949024
transform 1 0 5128 0 1 3039
box 0 0 1 1
use contact_17  contact_17_26
timestamp 1644949024
transform 1 0 5162 0 1 3044
box 0 0 1 1
use contact_18  contact_18_27
timestamp 1644949024
transform 1 0 5128 0 1 4577
box 0 0 1 1
use contact_17  contact_17_27
timestamp 1644949024
transform 1 0 5162 0 1 4582
box 0 0 1 1
use contact_18  contact_18_28
timestamp 1644949024
transform 1 0 5128 0 1 3039
box 0 0 1 1
use contact_17  contact_17_28
timestamp 1644949024
transform 1 0 5162 0 1 3044
box 0 0 1 1
use contact_18  contact_18_29
timestamp 1644949024
transform 1 0 5128 0 1 1501
box 0 0 1 1
use contact_17  contact_17_29
timestamp 1644949024
transform 1 0 5162 0 1 1506
box 0 0 1 1
use contact_18  contact_18_30
timestamp 1644949024
transform 1 0 5128 0 1 -37
box 0 0 1 1
use contact_17  contact_17_30
timestamp 1644949024
transform 1 0 5162 0 1 -32
box 0 0 1 1
use contact_18  contact_18_31
timestamp 1644949024
transform 1 0 5128 0 1 1501
box 0 0 1 1
use contact_17  contact_17_31
timestamp 1644949024
transform 1 0 5162 0 1 1506
box 0 0 1 1
use contact_20  contact_20_0
timestamp 1644949024
transform 1 0 3550 0 1 23055
box 0 0 1 1
use contact_18  contact_18_32
timestamp 1644949024
transform 1 0 2373 0 1 23867
box 0 0 1 1
use contact_17  contact_17_32
timestamp 1644949024
transform 1 0 2407 0 1 23872
box 0 0 1 1
use contact_13  contact_13_0
timestamp 1644949024
transform 1 0 2410 0 1 23881
box 0 0 1 1
use contact_20  contact_20_1
timestamp 1644949024
transform 1 0 3466 0 1 21515
box 0 0 1 1
use contact_18  contact_18_33
timestamp 1644949024
transform 1 0 2373 0 1 22243
box 0 0 1 1
use contact_17  contact_17_33
timestamp 1644949024
transform 1 0 2407 0 1 22248
box 0 0 1 1
use contact_13  contact_13_1
timestamp 1644949024
transform 1 0 2410 0 1 22257
box 0 0 1 1
use contact_20  contact_20_2
timestamp 1644949024
transform 1 0 3382 0 1 19975
box 0 0 1 1
use contact_18  contact_18_34
timestamp 1644949024
transform 1 0 2373 0 1 20787
box 0 0 1 1
use contact_17  contact_17_34
timestamp 1644949024
transform 1 0 2407 0 1 20792
box 0 0 1 1
use contact_13  contact_13_2
timestamp 1644949024
transform 1 0 2410 0 1 20801
box 0 0 1 1
use contact_20  contact_20_3
timestamp 1644949024
transform 1 0 3298 0 1 18435
box 0 0 1 1
use contact_18  contact_18_35
timestamp 1644949024
transform 1 0 2373 0 1 19163
box 0 0 1 1
use contact_17  contact_17_35
timestamp 1644949024
transform 1 0 2407 0 1 19168
box 0 0 1 1
use contact_13  contact_13_3
timestamp 1644949024
transform 1 0 2410 0 1 19177
box 0 0 1 1
use contact_20  contact_20_4
timestamp 1644949024
transform 1 0 3214 0 1 13819
box 0 0 1 1
use contact_18  contact_18_36
timestamp 1644949024
transform 1 0 2373 0 1 14631
box 0 0 1 1
use contact_17  contact_17_36
timestamp 1644949024
transform 1 0 2407 0 1 14636
box 0 0 1 1
use contact_13  contact_13_4
timestamp 1644949024
transform 1 0 2410 0 1 14645
box 0 0 1 1
use contact_20  contact_20_5
timestamp 1644949024
transform 1 0 3130 0 1 12279
box 0 0 1 1
use contact_18  contact_18_37
timestamp 1644949024
transform 1 0 2373 0 1 13007
box 0 0 1 1
use contact_17  contact_17_37
timestamp 1644949024
transform 1 0 2407 0 1 13012
box 0 0 1 1
use contact_13  contact_13_5
timestamp 1644949024
transform 1 0 2410 0 1 13021
box 0 0 1 1
use contact_20  contact_20_6
timestamp 1644949024
transform 1 0 3046 0 1 10739
box 0 0 1 1
use contact_18  contact_18_38
timestamp 1644949024
transform 1 0 2373 0 1 11551
box 0 0 1 1
use contact_17  contact_17_38
timestamp 1644949024
transform 1 0 2407 0 1 11556
box 0 0 1 1
use contact_13  contact_13_6
timestamp 1644949024
transform 1 0 2410 0 1 11565
box 0 0 1 1
use contact_20  contact_20_7
timestamp 1644949024
transform 1 0 2962 0 1 9199
box 0 0 1 1
use contact_18  contact_18_39
timestamp 1644949024
transform 1 0 2373 0 1 9927
box 0 0 1 1
use contact_17  contact_17_39
timestamp 1644949024
transform 1 0 2407 0 1 9932
box 0 0 1 1
use contact_13  contact_13_7
timestamp 1644949024
transform 1 0 2410 0 1 9941
box 0 0 1 1
use contact_20  contact_20_8
timestamp 1644949024
transform 1 0 2878 0 1 4583
box 0 0 1 1
use contact_18  contact_18_40
timestamp 1644949024
transform 1 0 2373 0 1 5395
box 0 0 1 1
use contact_17  contact_17_40
timestamp 1644949024
transform 1 0 2407 0 1 5400
box 0 0 1 1
use contact_13  contact_13_8
timestamp 1644949024
transform 1 0 2410 0 1 5409
box 0 0 1 1
use contact_20  contact_20_9
timestamp 1644949024
transform 1 0 2794 0 1 3043
box 0 0 1 1
use contact_18  contact_18_41
timestamp 1644949024
transform 1 0 2373 0 1 3771
box 0 0 1 1
use contact_17  contact_17_41
timestamp 1644949024
transform 1 0 2407 0 1 3776
box 0 0 1 1
use contact_13  contact_13_9
timestamp 1644949024
transform 1 0 2410 0 1 3785
box 0 0 1 1
use contact_20  contact_20_10
timestamp 1644949024
transform 1 0 2710 0 1 1503
box 0 0 1 1
use contact_18  contact_18_42
timestamp 1644949024
transform 1 0 2373 0 1 2315
box 0 0 1 1
use contact_17  contact_17_42
timestamp 1644949024
transform 1 0 2407 0 1 2320
box 0 0 1 1
use contact_13  contact_13_10
timestamp 1644949024
transform 1 0 2410 0 1 2329
box 0 0 1 1
use contact_20  contact_20_11
timestamp 1644949024
transform 1 0 2626 0 1 -37
box 0 0 1 1
use contact_18  contact_18_43
timestamp 1644949024
transform 1 0 2373 0 1 691
box 0 0 1 1
use contact_17  contact_17_43
timestamp 1644949024
transform 1 0 2407 0 1 696
box 0 0 1 1
use contact_13  contact_13_11
timestamp 1644949024
transform 1 0 2410 0 1 705
box 0 0 1 1
use contact_14  contact_14_0
timestamp 1644949024
transform 1 0 3500 0 1 24194
box 0 0 1 1
use contact_14  contact_14_1
timestamp 1644949024
transform 1 0 3248 0 1 24108
box 0 0 1 1
use contact_14  contact_14_2
timestamp 1644949024
transform 1 0 2828 0 1 24022
box 0 0 1 1
use contact_14  contact_14_3
timestamp 1644949024
transform 1 0 3500 0 1 23936
box 0 0 1 1
use contact_14  contact_14_4
timestamp 1644949024
transform 1 0 3248 0 1 23850
box 0 0 1 1
use contact_14  contact_14_5
timestamp 1644949024
transform 1 0 2744 0 1 23764
box 0 0 1 1
use contact_14  contact_14_6
timestamp 1644949024
transform 1 0 3500 0 1 23678
box 0 0 1 1
use contact_14  contact_14_7
timestamp 1644949024
transform 1 0 3248 0 1 23592
box 0 0 1 1
use contact_14  contact_14_8
timestamp 1644949024
transform 1 0 2660 0 1 23506
box 0 0 1 1
use contact_14  contact_14_9
timestamp 1644949024
transform 1 0 3500 0 1 21882
box 0 0 1 1
use contact_14  contact_14_10
timestamp 1644949024
transform 1 0 3164 0 1 21968
box 0 0 1 1
use contact_14  contact_14_11
timestamp 1644949024
transform 1 0 2912 0 1 22054
box 0 0 1 1
use contact_14  contact_14_12
timestamp 1644949024
transform 1 0 3500 0 1 22140
box 0 0 1 1
use contact_14  contact_14_13
timestamp 1644949024
transform 1 0 3164 0 1 22226
box 0 0 1 1
use contact_14  contact_14_14
timestamp 1644949024
transform 1 0 2828 0 1 22312
box 0 0 1 1
use contact_14  contact_14_15
timestamp 1644949024
transform 1 0 3500 0 1 22398
box 0 0 1 1
use contact_14  contact_14_16
timestamp 1644949024
transform 1 0 3164 0 1 22484
box 0 0 1 1
use contact_14  contact_14_17
timestamp 1644949024
transform 1 0 2744 0 1 22570
box 0 0 1 1
use contact_14  contact_14_18
timestamp 1644949024
transform 1 0 3500 0 1 21118
box 0 0 1 1
use contact_14  contact_14_19
timestamp 1644949024
transform 1 0 3164 0 1 21032
box 0 0 1 1
use contact_14  contact_14_20
timestamp 1644949024
transform 1 0 2660 0 1 20946
box 0 0 1 1
use contact_14  contact_14_21
timestamp 1644949024
transform 1 0 3500 0 1 20860
box 0 0 1 1
use contact_14  contact_14_22
timestamp 1644949024
transform 1 0 3080 0 1 20774
box 0 0 1 1
use contact_14  contact_14_23
timestamp 1644949024
transform 1 0 2912 0 1 20688
box 0 0 1 1
use contact_14  contact_14_24
timestamp 1644949024
transform 1 0 3500 0 1 20602
box 0 0 1 1
use contact_14  contact_14_25
timestamp 1644949024
transform 1 0 3080 0 1 20516
box 0 0 1 1
use contact_14  contact_14_26
timestamp 1644949024
transform 1 0 2828 0 1 20430
box 0 0 1 1
use contact_14  contact_14_27
timestamp 1644949024
transform 1 0 3500 0 1 18806
box 0 0 1 1
use contact_14  contact_14_28
timestamp 1644949024
transform 1 0 3080 0 1 18892
box 0 0 1 1
use contact_14  contact_14_29
timestamp 1644949024
transform 1 0 2744 0 1 18978
box 0 0 1 1
use contact_14  contact_14_30
timestamp 1644949024
transform 1 0 3500 0 1 19064
box 0 0 1 1
use contact_14  contact_14_31
timestamp 1644949024
transform 1 0 3080 0 1 19150
box 0 0 1 1
use contact_14  contact_14_32
timestamp 1644949024
transform 1 0 2660 0 1 19236
box 0 0 1 1
use contact_14  contact_14_33
timestamp 1644949024
transform 1 0 3500 0 1 19322
box 0 0 1 1
use contact_14  contact_14_34
timestamp 1644949024
transform 1 0 2996 0 1 19408
box 0 0 1 1
use contact_14  contact_14_35
timestamp 1644949024
transform 1 0 2912 0 1 19494
box 0 0 1 1
use contact_14  contact_14_36
timestamp 1644949024
transform 1 0 3500 0 1 18042
box 0 0 1 1
use contact_14  contact_14_37
timestamp 1644949024
transform 1 0 2996 0 1 17956
box 0 0 1 1
use contact_14  contact_14_38
timestamp 1644949024
transform 1 0 2828 0 1 17870
box 0 0 1 1
use contact_14  contact_14_39
timestamp 1644949024
transform 1 0 3500 0 1 17784
box 0 0 1 1
use contact_14  contact_14_40
timestamp 1644949024
transform 1 0 2996 0 1 17698
box 0 0 1 1
use contact_14  contact_14_41
timestamp 1644949024
transform 1 0 2744 0 1 17612
box 0 0 1 1
use contact_14  contact_14_42
timestamp 1644949024
transform 1 0 3500 0 1 17526
box 0 0 1 1
use contact_14  contact_14_43
timestamp 1644949024
transform 1 0 2996 0 1 17440
box 0 0 1 1
use contact_14  contact_14_44
timestamp 1644949024
transform 1 0 2660 0 1 17354
box 0 0 1 1
use contact_14  contact_14_45
timestamp 1644949024
transform 1 0 3416 0 1 15730
box 0 0 1 1
use contact_14  contact_14_46
timestamp 1644949024
transform 1 0 3248 0 1 15816
box 0 0 1 1
use contact_14  contact_14_47
timestamp 1644949024
transform 1 0 2912 0 1 15902
box 0 0 1 1
use contact_14  contact_14_48
timestamp 1644949024
transform 1 0 3416 0 1 15988
box 0 0 1 1
use contact_14  contact_14_49
timestamp 1644949024
transform 1 0 3248 0 1 16074
box 0 0 1 1
use contact_14  contact_14_50
timestamp 1644949024
transform 1 0 2828 0 1 16160
box 0 0 1 1
use contact_14  contact_14_51
timestamp 1644949024
transform 1 0 3416 0 1 16246
box 0 0 1 1
use contact_14  contact_14_52
timestamp 1644949024
transform 1 0 3248 0 1 16332
box 0 0 1 1
use contact_14  contact_14_53
timestamp 1644949024
transform 1 0 2744 0 1 16418
box 0 0 1 1
use contact_14  contact_14_54
timestamp 1644949024
transform 1 0 3416 0 1 14966
box 0 0 1 1
use contact_14  contact_14_55
timestamp 1644949024
transform 1 0 3248 0 1 14880
box 0 0 1 1
use contact_14  contact_14_56
timestamp 1644949024
transform 1 0 2660 0 1 14794
box 0 0 1 1
use contact_14  contact_14_57
timestamp 1644949024
transform 1 0 3416 0 1 14708
box 0 0 1 1
use contact_14  contact_14_58
timestamp 1644949024
transform 1 0 3164 0 1 14622
box 0 0 1 1
use contact_14  contact_14_59
timestamp 1644949024
transform 1 0 2912 0 1 14536
box 0 0 1 1
use contact_14  contact_14_60
timestamp 1644949024
transform 1 0 3416 0 1 14450
box 0 0 1 1
use contact_14  contact_14_61
timestamp 1644949024
transform 1 0 3164 0 1 14364
box 0 0 1 1
use contact_14  contact_14_62
timestamp 1644949024
transform 1 0 2828 0 1 14278
box 0 0 1 1
use contact_14  contact_14_63
timestamp 1644949024
transform 1 0 3416 0 1 12654
box 0 0 1 1
use contact_14  contact_14_64
timestamp 1644949024
transform 1 0 3164 0 1 12740
box 0 0 1 1
use contact_14  contact_14_65
timestamp 1644949024
transform 1 0 2744 0 1 12826
box 0 0 1 1
use contact_14  contact_14_66
timestamp 1644949024
transform 1 0 3416 0 1 12912
box 0 0 1 1
use contact_14  contact_14_67
timestamp 1644949024
transform 1 0 3164 0 1 12998
box 0 0 1 1
use contact_14  contact_14_68
timestamp 1644949024
transform 1 0 2660 0 1 13084
box 0 0 1 1
use contact_14  contact_14_69
timestamp 1644949024
transform 1 0 3416 0 1 13170
box 0 0 1 1
use contact_14  contact_14_70
timestamp 1644949024
transform 1 0 3080 0 1 13256
box 0 0 1 1
use contact_14  contact_14_71
timestamp 1644949024
transform 1 0 2912 0 1 13342
box 0 0 1 1
use contact_14  contact_14_72
timestamp 1644949024
transform 1 0 3416 0 1 11890
box 0 0 1 1
use contact_14  contact_14_73
timestamp 1644949024
transform 1 0 3080 0 1 11804
box 0 0 1 1
use contact_14  contact_14_74
timestamp 1644949024
transform 1 0 2828 0 1 11718
box 0 0 1 1
use contact_14  contact_14_75
timestamp 1644949024
transform 1 0 3416 0 1 11632
box 0 0 1 1
use contact_14  contact_14_76
timestamp 1644949024
transform 1 0 3080 0 1 11546
box 0 0 1 1
use contact_14  contact_14_77
timestamp 1644949024
transform 1 0 2744 0 1 11460
box 0 0 1 1
use contact_14  contact_14_78
timestamp 1644949024
transform 1 0 3416 0 1 11374
box 0 0 1 1
use contact_14  contact_14_79
timestamp 1644949024
transform 1 0 3080 0 1 11288
box 0 0 1 1
use contact_14  contact_14_80
timestamp 1644949024
transform 1 0 2660 0 1 11202
box 0 0 1 1
use contact_14  contact_14_81
timestamp 1644949024
transform 1 0 3416 0 1 9578
box 0 0 1 1
use contact_14  contact_14_82
timestamp 1644949024
transform 1 0 2996 0 1 9664
box 0 0 1 1
use contact_14  contact_14_83
timestamp 1644949024
transform 1 0 2912 0 1 9750
box 0 0 1 1
use contact_14  contact_14_84
timestamp 1644949024
transform 1 0 3416 0 1 9836
box 0 0 1 1
use contact_14  contact_14_85
timestamp 1644949024
transform 1 0 2996 0 1 9922
box 0 0 1 1
use contact_14  contact_14_86
timestamp 1644949024
transform 1 0 2828 0 1 10008
box 0 0 1 1
use contact_14  contact_14_87
timestamp 1644949024
transform 1 0 3416 0 1 10094
box 0 0 1 1
use contact_14  contact_14_88
timestamp 1644949024
transform 1 0 2996 0 1 10180
box 0 0 1 1
use contact_14  contact_14_89
timestamp 1644949024
transform 1 0 2744 0 1 10266
box 0 0 1 1
use contact_14  contact_14_90
timestamp 1644949024
transform 1 0 3416 0 1 8814
box 0 0 1 1
use contact_14  contact_14_91
timestamp 1644949024
transform 1 0 2996 0 1 8728
box 0 0 1 1
use contact_14  contact_14_92
timestamp 1644949024
transform 1 0 2660 0 1 8642
box 0 0 1 1
use contact_14  contact_14_93
timestamp 1644949024
transform 1 0 3332 0 1 8556
box 0 0 1 1
use contact_14  contact_14_94
timestamp 1644949024
transform 1 0 3248 0 1 8470
box 0 0 1 1
use contact_14  contact_14_95
timestamp 1644949024
transform 1 0 2912 0 1 8384
box 0 0 1 1
use contact_14  contact_14_96
timestamp 1644949024
transform 1 0 3332 0 1 8298
box 0 0 1 1
use contact_14  contact_14_97
timestamp 1644949024
transform 1 0 3248 0 1 8212
box 0 0 1 1
use contact_14  contact_14_98
timestamp 1644949024
transform 1 0 2828 0 1 8126
box 0 0 1 1
use contact_14  contact_14_99
timestamp 1644949024
transform 1 0 3332 0 1 6502
box 0 0 1 1
use contact_14  contact_14_100
timestamp 1644949024
transform 1 0 3248 0 1 6588
box 0 0 1 1
use contact_14  contact_14_101
timestamp 1644949024
transform 1 0 2744 0 1 6674
box 0 0 1 1
use contact_14  contact_14_102
timestamp 1644949024
transform 1 0 3332 0 1 6760
box 0 0 1 1
use contact_14  contact_14_103
timestamp 1644949024
transform 1 0 3248 0 1 6846
box 0 0 1 1
use contact_14  contact_14_104
timestamp 1644949024
transform 1 0 2660 0 1 6932
box 0 0 1 1
use contact_14  contact_14_105
timestamp 1644949024
transform 1 0 3332 0 1 7018
box 0 0 1 1
use contact_14  contact_14_106
timestamp 1644949024
transform 1 0 3164 0 1 7104
box 0 0 1 1
use contact_14  contact_14_107
timestamp 1644949024
transform 1 0 2912 0 1 7190
box 0 0 1 1
use contact_14  contact_14_108
timestamp 1644949024
transform 1 0 3332 0 1 5738
box 0 0 1 1
use contact_14  contact_14_109
timestamp 1644949024
transform 1 0 3164 0 1 5652
box 0 0 1 1
use contact_14  contact_14_110
timestamp 1644949024
transform 1 0 2828 0 1 5566
box 0 0 1 1
use contact_14  contact_14_111
timestamp 1644949024
transform 1 0 3332 0 1 5480
box 0 0 1 1
use contact_14  contact_14_112
timestamp 1644949024
transform 1 0 3164 0 1 5394
box 0 0 1 1
use contact_14  contact_14_113
timestamp 1644949024
transform 1 0 2744 0 1 5308
box 0 0 1 1
use contact_14  contact_14_114
timestamp 1644949024
transform 1 0 3332 0 1 5222
box 0 0 1 1
use contact_14  contact_14_115
timestamp 1644949024
transform 1 0 3164 0 1 5136
box 0 0 1 1
use contact_14  contact_14_116
timestamp 1644949024
transform 1 0 2660 0 1 5050
box 0 0 1 1
use contact_14  contact_14_117
timestamp 1644949024
transform 1 0 3332 0 1 3426
box 0 0 1 1
use contact_14  contact_14_118
timestamp 1644949024
transform 1 0 3080 0 1 3512
box 0 0 1 1
use contact_14  contact_14_119
timestamp 1644949024
transform 1 0 2912 0 1 3598
box 0 0 1 1
use contact_14  contact_14_120
timestamp 1644949024
transform 1 0 3332 0 1 3684
box 0 0 1 1
use contact_14  contact_14_121
timestamp 1644949024
transform 1 0 3080 0 1 3770
box 0 0 1 1
use contact_14  contact_14_122
timestamp 1644949024
transform 1 0 2828 0 1 3856
box 0 0 1 1
use contact_14  contact_14_123
timestamp 1644949024
transform 1 0 3332 0 1 3942
box 0 0 1 1
use contact_14  contact_14_124
timestamp 1644949024
transform 1 0 3080 0 1 4028
box 0 0 1 1
use contact_14  contact_14_125
timestamp 1644949024
transform 1 0 2744 0 1 4114
box 0 0 1 1
use contact_14  contact_14_126
timestamp 1644949024
transform 1 0 3332 0 1 2662
box 0 0 1 1
use contact_14  contact_14_127
timestamp 1644949024
transform 1 0 3080 0 1 2576
box 0 0 1 1
use contact_14  contact_14_128
timestamp 1644949024
transform 1 0 2660 0 1 2490
box 0 0 1 1
use contact_14  contact_14_129
timestamp 1644949024
transform 1 0 3332 0 1 2404
box 0 0 1 1
use contact_14  contact_14_130
timestamp 1644949024
transform 1 0 2996 0 1 2318
box 0 0 1 1
use contact_14  contact_14_131
timestamp 1644949024
transform 1 0 2912 0 1 2232
box 0 0 1 1
use contact_14  contact_14_132
timestamp 1644949024
transform 1 0 3332 0 1 2146
box 0 0 1 1
use contact_14  contact_14_133
timestamp 1644949024
transform 1 0 2996 0 1 2060
box 0 0 1 1
use contact_14  contact_14_134
timestamp 1644949024
transform 1 0 2828 0 1 1974
box 0 0 1 1
use contact_14  contact_14_135
timestamp 1644949024
transform 1 0 3332 0 1 350
box 0 0 1 1
use contact_14  contact_14_136
timestamp 1644949024
transform 1 0 2996 0 1 436
box 0 0 1 1
use contact_14  contact_14_137
timestamp 1644949024
transform 1 0 2744 0 1 522
box 0 0 1 1
use contact_14  contact_14_138
timestamp 1644949024
transform 1 0 3332 0 1 608
box 0 0 1 1
use contact_14  contact_14_139
timestamp 1644949024
transform 1 0 2996 0 1 694
box 0 0 1 1
use contact_14  contact_14_140
timestamp 1644949024
transform 1 0 2660 0 1 780
box 0 0 1 1
use contact_14  contact_14_141
timestamp 1644949024
transform 1 0 420 0 1 20792
box 0 0 1 1
use contact_17  contact_17_44
timestamp 1644949024
transform 1 0 700 0 1 20792
box 0 0 1 1
use contact_14  contact_14_142
timestamp 1644949024
transform 1 0 336 0 1 19168
box 0 0 1 1
use contact_17  contact_17_45
timestamp 1644949024
transform 1 0 616 0 1 19168
box 0 0 1 1
use contact_14  contact_14_143
timestamp 1644949024
transform 1 0 252 0 1 11556
box 0 0 1 1
use contact_17  contact_17_46
timestamp 1644949024
transform 1 0 700 0 1 11556
box 0 0 1 1
use contact_14  contact_14_144
timestamp 1644949024
transform 1 0 168 0 1 9932
box 0 0 1 1
use contact_17  contact_17_47
timestamp 1644949024
transform 1 0 616 0 1 9932
box 0 0 1 1
use contact_14  contact_14_145
timestamp 1644949024
transform 1 0 84 0 1 2320
box 0 0 1 1
use contact_17  contact_17_48
timestamp 1644949024
transform 1 0 700 0 1 2320
box 0 0 1 1
use contact_14  contact_14_146
timestamp 1644949024
transform 1 0 0 0 1 696
box 0 0 1 1
use contact_17  contact_17_49
timestamp 1644949024
transform 1 0 616 0 1 696
box 0 0 1 1
use dec_cell3_2r1w  dec_cell3_2r1w_0
timestamp 1644949024
transform 1 0 3686 0 -1 24608
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_1
timestamp 1644949024
transform 1 0 3686 0 1 21532
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_2
timestamp 1644949024
transform 1 0 3686 0 -1 21532
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_3
timestamp 1644949024
transform 1 0 3686 0 1 18456
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_4
timestamp 1644949024
transform 1 0 3686 0 -1 18456
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_5
timestamp 1644949024
transform 1 0 3686 0 1 15380
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_6
timestamp 1644949024
transform 1 0 3686 0 -1 15380
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_7
timestamp 1644949024
transform 1 0 3686 0 1 12304
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_8
timestamp 1644949024
transform 1 0 3686 0 -1 12304
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_9
timestamp 1644949024
transform 1 0 3686 0 1 9228
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_10
timestamp 1644949024
transform 1 0 3686 0 -1 9228
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_11
timestamp 1644949024
transform 1 0 3686 0 1 6152
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_12
timestamp 1644949024
transform 1 0 3686 0 -1 6152
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_13
timestamp 1644949024
transform 1 0 3686 0 1 3076
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_14
timestamp 1644949024
transform 1 0 3686 0 -1 3076
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_15
timestamp 1644949024
transform 1 0 3686 0 1 0
box 0 -42 1494 1616
use hierarchical_predecode2x4  hierarchical_predecode2x4_0
timestamp 1644949024
transform 1 0 550 0 1 18472
box 0 -37 2080 6197
use hierarchical_predecode2x4  hierarchical_predecode2x4_1
timestamp 1644949024
transform 1 0 550 0 1 9236
box 0 -37 2080 6197
use hierarchical_predecode2x4  hierarchical_predecode2x4_2
timestamp 1644949024
transform 1 0 550 0 1 0
box 0 -37 2080 6197
<< labels >>
rlabel metal2 s 18 0 46 24632 4 addr_0
rlabel metal2 s 102 0 130 24632 4 addr_1
rlabel metal2 s 186 0 214 24632 4 addr_2
rlabel metal2 s 270 0 298 24632 4 addr_3
rlabel metal2 s 354 0 382 24632 4 addr_4
rlabel metal2 s 438 0 466 24632 4 addr_5
rlabel metal1 s 5104 848 5180 876 4 decode0_0
rlabel metal1 s 4896 702 5180 730 4 decode1_0
rlabel metal1 s 4814 580 5180 608 4 decode2_0
rlabel metal1 s 5104 2200 5180 2228 4 decode0_1
rlabel metal1 s 4896 2346 5180 2374 4 decode1_1
rlabel metal1 s 4814 2468 5180 2496 4 decode2_1
rlabel metal1 s 5104 3924 5180 3952 4 decode0_2
rlabel metal1 s 4896 3778 5180 3806 4 decode1_2
rlabel metal1 s 4814 3656 5180 3684 4 decode2_2
rlabel metal1 s 5104 5276 5180 5304 4 decode0_3
rlabel metal1 s 4896 5422 5180 5450 4 decode1_3
rlabel metal1 s 4814 5544 5180 5572 4 decode2_3
rlabel metal1 s 5104 7000 5180 7028 4 decode0_4
rlabel metal1 s 4896 6854 5180 6882 4 decode1_4
rlabel metal1 s 4814 6732 5180 6760 4 decode2_4
rlabel metal1 s 5104 8352 5180 8380 4 decode0_5
rlabel metal1 s 4896 8498 5180 8526 4 decode1_5
rlabel metal1 s 4814 8620 5180 8648 4 decode2_5
rlabel metal1 s 5104 10076 5180 10104 4 decode0_6
rlabel metal1 s 4896 9930 5180 9958 4 decode1_6
rlabel metal1 s 4814 9808 5180 9836 4 decode2_6
rlabel metal1 s 5104 11428 5180 11456 4 decode0_7
rlabel metal1 s 4896 11574 5180 11602 4 decode1_7
rlabel metal1 s 4814 11696 5180 11724 4 decode2_7
rlabel metal1 s 5104 13152 5180 13180 4 decode0_8
rlabel metal1 s 4896 13006 5180 13034 4 decode1_8
rlabel metal1 s 4814 12884 5180 12912 4 decode2_8
rlabel metal1 s 5104 14504 5180 14532 4 decode0_9
rlabel metal1 s 4896 14650 5180 14678 4 decode1_9
rlabel metal1 s 4814 14772 5180 14800 4 decode2_9
rlabel metal1 s 5104 16228 5180 16256 4 decode0_10
rlabel metal1 s 4896 16082 5180 16110 4 decode1_10
rlabel metal1 s 4814 15960 5180 15988 4 decode2_10
rlabel metal1 s 5104 17580 5180 17608 4 decode0_11
rlabel metal1 s 4896 17726 5180 17754 4 decode1_11
rlabel metal1 s 4814 17848 5180 17876 4 decode2_11
rlabel metal1 s 5104 19304 5180 19332 4 decode0_12
rlabel metal1 s 4896 19158 5180 19186 4 decode1_12
rlabel metal1 s 4814 19036 5180 19064 4 decode2_12
rlabel metal1 s 5104 20656 5180 20684 4 decode0_13
rlabel metal1 s 4896 20802 5180 20830 4 decode1_13
rlabel metal1 s 4814 20924 5180 20952 4 decode2_13
rlabel metal1 s 5104 22380 5180 22408 4 decode0_14
rlabel metal1 s 4896 22234 5180 22262 4 decode1_14
rlabel metal1 s 4814 22112 5180 22140 4 decode2_14
rlabel metal1 s 5104 23732 5180 23760 4 decode0_15
rlabel metal1 s 4896 23878 5180 23906 4 decode1_15
rlabel metal1 s 4814 24000 5180 24028 4 decode2_15
rlabel metal2 s 2678 0 2706 24660 4 predecode_0
rlabel metal2 s 2762 0 2790 24660 4 predecode_1
rlabel metal2 s 2846 0 2874 24660 4 predecode_2
rlabel metal2 s 2930 0 2958 24660 4 predecode_3
rlabel metal2 s 3014 0 3042 24660 4 predecode_4
rlabel metal2 s 3098 0 3126 24660 4 predecode_5
rlabel metal2 s 3182 0 3210 24660 4 predecode_6
rlabel metal2 s 3266 0 3294 24660 4 predecode_7
rlabel metal2 s 3350 0 3378 24660 4 predecode_8
rlabel metal2 s 3434 0 3462 24660 4 predecode_9
rlabel metal2 s 3518 0 3546 24660 4 predecode_10
rlabel metal2 s 3602 0 3630 24660 4 predecode_11
rlabel metal3 s 1664 19975 1796 20049 4 vdd
rlabel metal3 s 792 23055 924 23129 4 vdd
rlabel metal3 s 1664 1503 1796 1577 4 vdd
rlabel metal3 s 792 13819 924 13893 4 vdd
rlabel metal3 s 792 4583 924 4657 4 vdd
rlabel metal3 s 1664 23055 1796 23129 4 vdd
rlabel metal3 s 5128 7653 5260 7727 4 vdd
rlabel metal3 s 1664 4583 1796 4657 4 vdd
rlabel metal3 s 5128 1501 5260 1575 4 vdd
rlabel metal3 s 1664 13819 1796 13893 4 vdd
rlabel metal3 s 5194 1538 5194 1538 4 vdd
rlabel metal3 s 1664 10739 1796 10813 4 vdd
rlabel metal3 s 5128 4577 5260 4651 4 vdd
rlabel metal3 s 792 1503 924 1577 4 vdd
rlabel metal3 s 5128 13805 5260 13879 4 vdd
rlabel metal3 s 5128 10729 5260 10803 4 vdd
rlabel metal3 s 5194 10766 5194 10766 4 vdd
rlabel metal3 s 5128 16881 5260 16955 4 vdd
rlabel metal3 s 792 10739 924 10813 4 vdd
rlabel metal3 s 5128 19957 5260 20031 4 vdd
rlabel metal3 s 792 19975 924 20049 4 vdd
rlabel metal3 s 5128 23033 5260 23107 4 vdd
rlabel metal3 s 792 9199 924 9273 4 gnd
rlabel metal3 s 5128 18419 5260 18493 4 gnd
rlabel metal3 s 5128 15343 5260 15417 4 gnd
rlabel metal3 s 792 15359 924 15433 4 gnd
rlabel metal3 s 792 6123 924 6197 4 gnd
rlabel metal3 s 1664 21515 1796 21589 4 gnd
rlabel metal3 s 5128 -37 5260 37 4 gnd
rlabel metal3 s 792 24595 924 24669 4 gnd
rlabel metal3 s 5128 21495 5260 21569 4 gnd
rlabel metal3 s 792 18435 924 18509 4 gnd
rlabel metal3 s 1664 9199 1796 9273 4 gnd
rlabel metal3 s 5128 9191 5260 9265 4 gnd
rlabel metal3 s 5128 12267 5260 12341 4 gnd
rlabel metal3 s 792 21515 924 21589 4 gnd
rlabel metal3 s 1664 18435 1796 18509 4 gnd
rlabel metal3 s 1664 15359 1796 15433 4 gnd
rlabel metal3 s 1664 3043 1796 3117 4 gnd
rlabel metal3 s 5128 3039 5260 3113 4 gnd
rlabel metal3 s 792 12279 924 12353 4 gnd
rlabel metal3 s 1664 12279 1796 12353 4 gnd
rlabel metal3 s 792 3043 924 3117 4 gnd
rlabel metal3 s 1664 -37 1796 37 4 gnd
rlabel metal3 s 1664 6123 1796 6197 4 gnd
rlabel metal3 s 5128 24571 5260 24645 4 gnd
rlabel metal3 s 5128 6115 5260 6189 4 gnd
rlabel metal3 s 792 -37 924 37 4 gnd
rlabel metal3 s 1664 24595 1796 24669 4 gnd
<< properties >>
string FIXED_BBOX 5128 -37 5260 0
string GDS_FILE sram_0rw2r1w_4_16_sky130A.gds
string GDS_END 325804
string GDS_START 268094
<< end >>
