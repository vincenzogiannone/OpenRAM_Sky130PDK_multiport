magic
tech sky130A
magscale 1 2
timestamp 1644969367
<< checkpaint >>
rect -1296 -1277 1880 2155
<< nwell >>
rect -36 402 620 895
<< pwell >>
rect 474 51 524 133
<< psubdiff >>
rect 474 109 524 133
rect 474 75 482 109
rect 516 75 524 109
rect 474 51 524 75
<< nsubdiff >>
rect 474 763 524 787
rect 474 729 482 763
rect 516 729 524 763
rect 474 705 524 729
<< psubdiffcont >>
rect 482 75 516 109
<< nsubdiffcont >>
rect 482 729 516 763
<< poly >>
rect 114 410 144 479
rect 48 394 144 410
rect 48 360 64 394
rect 98 360 144 394
rect 48 344 144 360
rect 114 191 144 344
<< polycont >>
rect 64 360 98 394
<< locali >>
rect 0 821 584 855
rect 62 628 96 821
rect 274 628 308 821
rect 482 763 516 821
rect 482 713 516 729
rect 48 394 114 410
rect 48 360 64 394
rect 98 360 114 394
rect 48 344 114 360
rect 272 394 306 594
rect 272 360 323 394
rect 272 160 306 360
rect 482 109 516 125
rect 62 17 96 60
rect 274 17 308 60
rect 482 17 516 75
rect 0 -17 584 17
use contact_12  contact_12_0
timestamp 1644969367
transform 1 0 48 0 1 344
box 0 0 1 1
use contact_11  contact_11_0
timestamp 1644969367
transform 1 0 474 0 1 51
box 0 0 1 1
use contact_10  contact_10_0
timestamp 1644969367
transform 1 0 474 0 1 705
box 0 0 1 1
use nmos_m3_w0_420_sli_dli_da_p  nmos_m3_w0_420_sli_dli_da_p_0
timestamp 1644969367
transform 1 0 54 0 1 51
box 0 -26 366 143
use pmos_m3_w1_260_sli_dli_da_p  pmos_m3_w1_260_sli_dli_da_p_0
timestamp 1644969367
transform 1 0 54 0 1 535
box -59 -56 425 306
<< labels >>
rlabel locali s 81 377 81 377 4 A
rlabel locali s 306 377 306 377 4 Z
rlabel locali s 292 0 292 0 4 gnd
rlabel locali s 292 838 292 838 4 vdd
<< properties >>
string FIXED_BBOX 0 0 584 838
string GDS_FILE sram_0rw2r1w_32_128_sky130A.gds
string GDS_END 3308428
string GDS_START 3306808
<< end >>
