magic
tech sky130A
magscale 1 2
timestamp 1644951705
<< checkpaint >>
rect -1319 -1316 5681 1610
<< nwell >>
rect -54 232 4416 350
rect -59 64 4421 232
rect -54 -54 4416 64
<< scpmos >>
rect 60 0 90 296
rect 168 0 198 296
rect 276 0 306 296
rect 384 0 414 296
rect 492 0 522 296
rect 600 0 630 296
rect 708 0 738 296
rect 816 0 846 296
rect 924 0 954 296
rect 1032 0 1062 296
rect 1140 0 1170 296
rect 1248 0 1278 296
rect 1356 0 1386 296
rect 1464 0 1494 296
rect 1572 0 1602 296
rect 1680 0 1710 296
rect 1788 0 1818 296
rect 1896 0 1926 296
rect 2004 0 2034 296
rect 2112 0 2142 296
rect 2220 0 2250 296
rect 2328 0 2358 296
rect 2436 0 2466 296
rect 2544 0 2574 296
rect 2652 0 2682 296
rect 2760 0 2790 296
rect 2868 0 2898 296
rect 2976 0 3006 296
rect 3084 0 3114 296
rect 3192 0 3222 296
rect 3300 0 3330 296
rect 3408 0 3438 296
rect 3516 0 3546 296
rect 3624 0 3654 296
rect 3732 0 3762 296
rect 3840 0 3870 296
rect 3948 0 3978 296
rect 4056 0 4086 296
rect 4164 0 4194 296
rect 4272 0 4302 296
<< pdiff >>
rect 0 165 60 296
rect 0 131 8 165
rect 42 131 60 165
rect 0 0 60 131
rect 90 165 168 296
rect 90 131 112 165
rect 146 131 168 165
rect 90 0 168 131
rect 198 165 276 296
rect 198 131 220 165
rect 254 131 276 165
rect 198 0 276 131
rect 306 165 384 296
rect 306 131 328 165
rect 362 131 384 165
rect 306 0 384 131
rect 414 165 492 296
rect 414 131 436 165
rect 470 131 492 165
rect 414 0 492 131
rect 522 165 600 296
rect 522 131 544 165
rect 578 131 600 165
rect 522 0 600 131
rect 630 165 708 296
rect 630 131 652 165
rect 686 131 708 165
rect 630 0 708 131
rect 738 165 816 296
rect 738 131 760 165
rect 794 131 816 165
rect 738 0 816 131
rect 846 165 924 296
rect 846 131 868 165
rect 902 131 924 165
rect 846 0 924 131
rect 954 165 1032 296
rect 954 131 976 165
rect 1010 131 1032 165
rect 954 0 1032 131
rect 1062 165 1140 296
rect 1062 131 1084 165
rect 1118 131 1140 165
rect 1062 0 1140 131
rect 1170 165 1248 296
rect 1170 131 1192 165
rect 1226 131 1248 165
rect 1170 0 1248 131
rect 1278 165 1356 296
rect 1278 131 1300 165
rect 1334 131 1356 165
rect 1278 0 1356 131
rect 1386 165 1464 296
rect 1386 131 1408 165
rect 1442 131 1464 165
rect 1386 0 1464 131
rect 1494 165 1572 296
rect 1494 131 1516 165
rect 1550 131 1572 165
rect 1494 0 1572 131
rect 1602 165 1680 296
rect 1602 131 1624 165
rect 1658 131 1680 165
rect 1602 0 1680 131
rect 1710 165 1788 296
rect 1710 131 1732 165
rect 1766 131 1788 165
rect 1710 0 1788 131
rect 1818 165 1896 296
rect 1818 131 1840 165
rect 1874 131 1896 165
rect 1818 0 1896 131
rect 1926 165 2004 296
rect 1926 131 1948 165
rect 1982 131 2004 165
rect 1926 0 2004 131
rect 2034 165 2112 296
rect 2034 131 2056 165
rect 2090 131 2112 165
rect 2034 0 2112 131
rect 2142 165 2220 296
rect 2142 131 2164 165
rect 2198 131 2220 165
rect 2142 0 2220 131
rect 2250 165 2328 296
rect 2250 131 2272 165
rect 2306 131 2328 165
rect 2250 0 2328 131
rect 2358 165 2436 296
rect 2358 131 2380 165
rect 2414 131 2436 165
rect 2358 0 2436 131
rect 2466 165 2544 296
rect 2466 131 2488 165
rect 2522 131 2544 165
rect 2466 0 2544 131
rect 2574 165 2652 296
rect 2574 131 2596 165
rect 2630 131 2652 165
rect 2574 0 2652 131
rect 2682 165 2760 296
rect 2682 131 2704 165
rect 2738 131 2760 165
rect 2682 0 2760 131
rect 2790 165 2868 296
rect 2790 131 2812 165
rect 2846 131 2868 165
rect 2790 0 2868 131
rect 2898 165 2976 296
rect 2898 131 2920 165
rect 2954 131 2976 165
rect 2898 0 2976 131
rect 3006 165 3084 296
rect 3006 131 3028 165
rect 3062 131 3084 165
rect 3006 0 3084 131
rect 3114 165 3192 296
rect 3114 131 3136 165
rect 3170 131 3192 165
rect 3114 0 3192 131
rect 3222 165 3300 296
rect 3222 131 3244 165
rect 3278 131 3300 165
rect 3222 0 3300 131
rect 3330 165 3408 296
rect 3330 131 3352 165
rect 3386 131 3408 165
rect 3330 0 3408 131
rect 3438 165 3516 296
rect 3438 131 3460 165
rect 3494 131 3516 165
rect 3438 0 3516 131
rect 3546 165 3624 296
rect 3546 131 3568 165
rect 3602 131 3624 165
rect 3546 0 3624 131
rect 3654 165 3732 296
rect 3654 131 3676 165
rect 3710 131 3732 165
rect 3654 0 3732 131
rect 3762 165 3840 296
rect 3762 131 3784 165
rect 3818 131 3840 165
rect 3762 0 3840 131
rect 3870 165 3948 296
rect 3870 131 3892 165
rect 3926 131 3948 165
rect 3870 0 3948 131
rect 3978 165 4056 296
rect 3978 131 4000 165
rect 4034 131 4056 165
rect 3978 0 4056 131
rect 4086 165 4164 296
rect 4086 131 4108 165
rect 4142 131 4164 165
rect 4086 0 4164 131
rect 4194 165 4272 296
rect 4194 131 4216 165
rect 4250 131 4272 165
rect 4194 0 4272 131
rect 4302 165 4362 296
rect 4302 131 4320 165
rect 4354 131 4362 165
rect 4302 0 4362 131
<< pdiffc >>
rect 8 131 42 165
rect 112 131 146 165
rect 220 131 254 165
rect 328 131 362 165
rect 436 131 470 165
rect 544 131 578 165
rect 652 131 686 165
rect 760 131 794 165
rect 868 131 902 165
rect 976 131 1010 165
rect 1084 131 1118 165
rect 1192 131 1226 165
rect 1300 131 1334 165
rect 1408 131 1442 165
rect 1516 131 1550 165
rect 1624 131 1658 165
rect 1732 131 1766 165
rect 1840 131 1874 165
rect 1948 131 1982 165
rect 2056 131 2090 165
rect 2164 131 2198 165
rect 2272 131 2306 165
rect 2380 131 2414 165
rect 2488 131 2522 165
rect 2596 131 2630 165
rect 2704 131 2738 165
rect 2812 131 2846 165
rect 2920 131 2954 165
rect 3028 131 3062 165
rect 3136 131 3170 165
rect 3244 131 3278 165
rect 3352 131 3386 165
rect 3460 131 3494 165
rect 3568 131 3602 165
rect 3676 131 3710 165
rect 3784 131 3818 165
rect 3892 131 3926 165
rect 4000 131 4034 165
rect 4108 131 4142 165
rect 4216 131 4250 165
rect 4320 131 4354 165
<< poly >>
rect 60 296 90 322
rect 168 296 198 322
rect 276 296 306 322
rect 384 296 414 322
rect 492 296 522 322
rect 600 296 630 322
rect 708 296 738 322
rect 816 296 846 322
rect 924 296 954 322
rect 1032 296 1062 322
rect 1140 296 1170 322
rect 1248 296 1278 322
rect 1356 296 1386 322
rect 1464 296 1494 322
rect 1572 296 1602 322
rect 1680 296 1710 322
rect 1788 296 1818 322
rect 1896 296 1926 322
rect 2004 296 2034 322
rect 2112 296 2142 322
rect 2220 296 2250 322
rect 2328 296 2358 322
rect 2436 296 2466 322
rect 2544 296 2574 322
rect 2652 296 2682 322
rect 2760 296 2790 322
rect 2868 296 2898 322
rect 2976 296 3006 322
rect 3084 296 3114 322
rect 3192 296 3222 322
rect 3300 296 3330 322
rect 3408 296 3438 322
rect 3516 296 3546 322
rect 3624 296 3654 322
rect 3732 296 3762 322
rect 3840 296 3870 322
rect 3948 296 3978 322
rect 4056 296 4086 322
rect 4164 296 4194 322
rect 4272 296 4302 322
rect 60 -26 90 0
rect 168 -26 198 0
rect 276 -26 306 0
rect 384 -26 414 0
rect 492 -26 522 0
rect 600 -26 630 0
rect 708 -26 738 0
rect 816 -26 846 0
rect 924 -26 954 0
rect 1032 -26 1062 0
rect 1140 -26 1170 0
rect 1248 -26 1278 0
rect 1356 -26 1386 0
rect 1464 -26 1494 0
rect 1572 -26 1602 0
rect 1680 -26 1710 0
rect 1788 -26 1818 0
rect 1896 -26 1926 0
rect 2004 -26 2034 0
rect 2112 -26 2142 0
rect 2220 -26 2250 0
rect 2328 -26 2358 0
rect 2436 -26 2466 0
rect 2544 -26 2574 0
rect 2652 -26 2682 0
rect 2760 -26 2790 0
rect 2868 -26 2898 0
rect 2976 -26 3006 0
rect 3084 -26 3114 0
rect 3192 -26 3222 0
rect 3300 -26 3330 0
rect 3408 -26 3438 0
rect 3516 -26 3546 0
rect 3624 -26 3654 0
rect 3732 -26 3762 0
rect 3840 -26 3870 0
rect 3948 -26 3978 0
rect 4056 -26 4086 0
rect 4164 -26 4194 0
rect 4272 -26 4302 0
rect 60 -56 4302 -26
<< locali >>
rect 8 165 42 181
rect 8 115 42 131
rect 112 165 146 181
rect 112 81 146 131
rect 220 165 254 181
rect 220 115 254 131
rect 328 165 362 181
rect 328 81 362 131
rect 436 165 470 181
rect 436 115 470 131
rect 544 165 578 181
rect 544 81 578 131
rect 652 165 686 181
rect 652 115 686 131
rect 760 165 794 181
rect 760 81 794 131
rect 868 165 902 181
rect 868 115 902 131
rect 976 165 1010 181
rect 976 81 1010 131
rect 1084 165 1118 181
rect 1084 115 1118 131
rect 1192 165 1226 181
rect 1192 81 1226 131
rect 1300 165 1334 181
rect 1300 115 1334 131
rect 1408 165 1442 181
rect 1408 81 1442 131
rect 1516 165 1550 181
rect 1516 115 1550 131
rect 1624 165 1658 181
rect 1624 81 1658 131
rect 1732 165 1766 181
rect 1732 115 1766 131
rect 1840 165 1874 181
rect 1840 81 1874 131
rect 1948 165 1982 181
rect 1948 115 1982 131
rect 2056 165 2090 181
rect 2056 81 2090 131
rect 2164 165 2198 181
rect 2164 115 2198 131
rect 2272 165 2306 181
rect 2272 81 2306 131
rect 2380 165 2414 181
rect 2380 115 2414 131
rect 2488 165 2522 181
rect 2488 81 2522 131
rect 2596 165 2630 181
rect 2596 115 2630 131
rect 2704 165 2738 181
rect 2704 81 2738 131
rect 2812 165 2846 181
rect 2812 115 2846 131
rect 2920 165 2954 181
rect 2920 81 2954 131
rect 3028 165 3062 181
rect 3028 115 3062 131
rect 3136 165 3170 181
rect 3136 81 3170 131
rect 3244 165 3278 181
rect 3244 115 3278 131
rect 3352 165 3386 181
rect 3352 81 3386 131
rect 3460 165 3494 181
rect 3460 115 3494 131
rect 3568 165 3602 181
rect 3568 81 3602 131
rect 3676 165 3710 181
rect 3676 115 3710 131
rect 3784 165 3818 181
rect 3784 81 3818 131
rect 3892 165 3926 181
rect 3892 115 3926 131
rect 4000 165 4034 181
rect 4000 81 4034 131
rect 4108 165 4142 181
rect 4108 115 4142 131
rect 4216 165 4250 181
rect 4216 81 4250 131
rect 4320 165 4354 181
rect 4320 115 4354 131
rect 112 47 4250 81
use contact_9  contact_9_0
timestamp 1644951705
transform 1 0 4312 0 1 107
box 0 0 2 2
use contact_9  contact_9_1
timestamp 1644951705
transform 1 0 4208 0 1 107
box 0 0 2 2
use contact_9  contact_9_2
timestamp 1644951705
transform 1 0 4100 0 1 107
box 0 0 2 2
use contact_9  contact_9_3
timestamp 1644951705
transform 1 0 3992 0 1 107
box 0 0 2 2
use contact_9  contact_9_4
timestamp 1644951705
transform 1 0 3884 0 1 107
box 0 0 2 2
use contact_9  contact_9_5
timestamp 1644951705
transform 1 0 3776 0 1 107
box 0 0 2 2
use contact_9  contact_9_6
timestamp 1644951705
transform 1 0 3668 0 1 107
box 0 0 2 2
use contact_9  contact_9_7
timestamp 1644951705
transform 1 0 3560 0 1 107
box 0 0 2 2
use contact_9  contact_9_8
timestamp 1644951705
transform 1 0 3452 0 1 107
box 0 0 2 2
use contact_9  contact_9_9
timestamp 1644951705
transform 1 0 3344 0 1 107
box 0 0 2 2
use contact_9  contact_9_10
timestamp 1644951705
transform 1 0 3236 0 1 107
box 0 0 2 2
use contact_9  contact_9_11
timestamp 1644951705
transform 1 0 3128 0 1 107
box 0 0 2 2
use contact_9  contact_9_12
timestamp 1644951705
transform 1 0 3020 0 1 107
box 0 0 2 2
use contact_9  contact_9_13
timestamp 1644951705
transform 1 0 2912 0 1 107
box 0 0 2 2
use contact_9  contact_9_14
timestamp 1644951705
transform 1 0 2804 0 1 107
box 0 0 2 2
use contact_9  contact_9_15
timestamp 1644951705
transform 1 0 2696 0 1 107
box 0 0 2 2
use contact_9  contact_9_16
timestamp 1644951705
transform 1 0 2588 0 1 107
box 0 0 2 2
use contact_9  contact_9_17
timestamp 1644951705
transform 1 0 2480 0 1 107
box 0 0 2 2
use contact_9  contact_9_18
timestamp 1644951705
transform 1 0 2372 0 1 107
box 0 0 2 2
use contact_9  contact_9_19
timestamp 1644951705
transform 1 0 2264 0 1 107
box 0 0 2 2
use contact_9  contact_9_20
timestamp 1644951705
transform 1 0 2156 0 1 107
box 0 0 2 2
use contact_9  contact_9_21
timestamp 1644951705
transform 1 0 2048 0 1 107
box 0 0 2 2
use contact_9  contact_9_22
timestamp 1644951705
transform 1 0 1940 0 1 107
box 0 0 2 2
use contact_9  contact_9_23
timestamp 1644951705
transform 1 0 1832 0 1 107
box 0 0 2 2
use contact_9  contact_9_24
timestamp 1644951705
transform 1 0 1724 0 1 107
box 0 0 2 2
use contact_9  contact_9_25
timestamp 1644951705
transform 1 0 1616 0 1 107
box 0 0 2 2
use contact_9  contact_9_26
timestamp 1644951705
transform 1 0 1508 0 1 107
box 0 0 2 2
use contact_9  contact_9_27
timestamp 1644951705
transform 1 0 1400 0 1 107
box 0 0 2 2
use contact_9  contact_9_28
timestamp 1644951705
transform 1 0 1292 0 1 107
box 0 0 2 2
use contact_9  contact_9_29
timestamp 1644951705
transform 1 0 1184 0 1 107
box 0 0 2 2
use contact_9  contact_9_30
timestamp 1644951705
transform 1 0 1076 0 1 107
box 0 0 2 2
use contact_9  contact_9_31
timestamp 1644951705
transform 1 0 968 0 1 107
box 0 0 2 2
use contact_9  contact_9_32
timestamp 1644951705
transform 1 0 860 0 1 107
box 0 0 2 2
use contact_9  contact_9_33
timestamp 1644951705
transform 1 0 752 0 1 107
box 0 0 2 2
use contact_9  contact_9_34
timestamp 1644951705
transform 1 0 644 0 1 107
box 0 0 2 2
use contact_9  contact_9_35
timestamp 1644951705
transform 1 0 536 0 1 107
box 0 0 2 2
use contact_9  contact_9_36
timestamp 1644951705
transform 1 0 428 0 1 107
box 0 0 2 2
use contact_9  contact_9_37
timestamp 1644951705
transform 1 0 320 0 1 107
box 0 0 2 2
use contact_9  contact_9_38
timestamp 1644951705
transform 1 0 212 0 1 107
box 0 0 2 2
use contact_9  contact_9_39
timestamp 1644951705
transform 1 0 104 0 1 107
box 0 0 2 2
use contact_9  contact_9_40
timestamp 1644951705
transform 1 0 0 0 1 107
box 0 0 2 2
<< labels >>
rlabel mvvaractor s 2181 -41 2181 -41 4 G
rlabel locali s 3045 148 3045 148 4 S
rlabel locali s 2397 148 2397 148 4 S
rlabel locali s 1533 148 1533 148 4 S
rlabel locali s 2181 148 2181 148 4 S
rlabel locali s 2613 148 2613 148 4 S
rlabel locali s 3693 148 3693 148 4 S
rlabel locali s 1965 148 1965 148 4 S
rlabel locali s 3261 148 3261 148 4 S
rlabel locali s 669 148 669 148 4 S
rlabel locali s 1749 148 1749 148 4 S
rlabel locali s 3477 148 3477 148 4 S
rlabel locali s 4337 148 4337 148 4 S
rlabel locali s 2829 148 2829 148 4 S
rlabel locali s 237 148 237 148 4 S
rlabel locali s 1317 148 1317 148 4 S
rlabel locali s 885 148 885 148 4 S
rlabel locali s 3909 148 3909 148 4 S
rlabel locali s 1101 148 1101 148 4 S
rlabel locali s 453 148 453 148 4 S
rlabel locali s 25 148 25 148 4 S
rlabel locali s 4125 148 4125 148 4 S
rlabel locali s 2181 64 2181 64 4 D
<< properties >>
string FIXED_BBOX -54 -56 4416 64
string GDS_FILE sram_0rw2r1w_16_128_sky130A.gds
string GDS_END 2011208
string GDS_START 2002644
<< end >>
