magic
tech sky130A
magscale 1 2
timestamp 1644969367
<< checkpaint >>
rect -1260 -1286 7890 1415
<< scnmos >>
rect 60 0 90 99
rect 168 0 198 99
rect 276 0 306 99
rect 384 0 414 99
rect 492 0 522 99
rect 600 0 630 99
rect 708 0 738 99
rect 816 0 846 99
rect 924 0 954 99
rect 1032 0 1062 99
rect 1140 0 1170 99
rect 1248 0 1278 99
rect 1356 0 1386 99
rect 1464 0 1494 99
rect 1572 0 1602 99
rect 1680 0 1710 99
rect 1788 0 1818 99
rect 1896 0 1926 99
rect 2004 0 2034 99
rect 2112 0 2142 99
rect 2220 0 2250 99
rect 2328 0 2358 99
rect 2436 0 2466 99
rect 2544 0 2574 99
rect 2652 0 2682 99
rect 2760 0 2790 99
rect 2868 0 2898 99
rect 2976 0 3006 99
rect 3084 0 3114 99
rect 3192 0 3222 99
rect 3300 0 3330 99
rect 3408 0 3438 99
rect 3516 0 3546 99
rect 3624 0 3654 99
rect 3732 0 3762 99
rect 3840 0 3870 99
rect 3948 0 3978 99
rect 4056 0 4086 99
rect 4164 0 4194 99
rect 4272 0 4302 99
rect 4380 0 4410 99
rect 4488 0 4518 99
rect 4596 0 4626 99
rect 4704 0 4734 99
rect 4812 0 4842 99
rect 4920 0 4950 99
rect 5028 0 5058 99
rect 5136 0 5166 99
rect 5244 0 5274 99
rect 5352 0 5382 99
rect 5460 0 5490 99
rect 5568 0 5598 99
rect 5676 0 5706 99
rect 5784 0 5814 99
rect 5892 0 5922 99
rect 6000 0 6030 99
rect 6108 0 6138 99
rect 6216 0 6246 99
rect 6324 0 6354 99
rect 6432 0 6462 99
rect 6540 0 6570 99
<< ndiff >>
rect 0 66 60 99
rect 0 32 8 66
rect 42 32 60 66
rect 0 0 60 32
rect 90 66 168 99
rect 90 32 112 66
rect 146 32 168 66
rect 90 0 168 32
rect 198 66 276 99
rect 198 32 220 66
rect 254 32 276 66
rect 198 0 276 32
rect 306 66 384 99
rect 306 32 328 66
rect 362 32 384 66
rect 306 0 384 32
rect 414 66 492 99
rect 414 32 436 66
rect 470 32 492 66
rect 414 0 492 32
rect 522 66 600 99
rect 522 32 544 66
rect 578 32 600 66
rect 522 0 600 32
rect 630 66 708 99
rect 630 32 652 66
rect 686 32 708 66
rect 630 0 708 32
rect 738 66 816 99
rect 738 32 760 66
rect 794 32 816 66
rect 738 0 816 32
rect 846 66 924 99
rect 846 32 868 66
rect 902 32 924 66
rect 846 0 924 32
rect 954 66 1032 99
rect 954 32 976 66
rect 1010 32 1032 66
rect 954 0 1032 32
rect 1062 66 1140 99
rect 1062 32 1084 66
rect 1118 32 1140 66
rect 1062 0 1140 32
rect 1170 66 1248 99
rect 1170 32 1192 66
rect 1226 32 1248 66
rect 1170 0 1248 32
rect 1278 66 1356 99
rect 1278 32 1300 66
rect 1334 32 1356 66
rect 1278 0 1356 32
rect 1386 66 1464 99
rect 1386 32 1408 66
rect 1442 32 1464 66
rect 1386 0 1464 32
rect 1494 66 1572 99
rect 1494 32 1516 66
rect 1550 32 1572 66
rect 1494 0 1572 32
rect 1602 66 1680 99
rect 1602 32 1624 66
rect 1658 32 1680 66
rect 1602 0 1680 32
rect 1710 66 1788 99
rect 1710 32 1732 66
rect 1766 32 1788 66
rect 1710 0 1788 32
rect 1818 66 1896 99
rect 1818 32 1840 66
rect 1874 32 1896 66
rect 1818 0 1896 32
rect 1926 66 2004 99
rect 1926 32 1948 66
rect 1982 32 2004 66
rect 1926 0 2004 32
rect 2034 66 2112 99
rect 2034 32 2056 66
rect 2090 32 2112 66
rect 2034 0 2112 32
rect 2142 66 2220 99
rect 2142 32 2164 66
rect 2198 32 2220 66
rect 2142 0 2220 32
rect 2250 66 2328 99
rect 2250 32 2272 66
rect 2306 32 2328 66
rect 2250 0 2328 32
rect 2358 66 2436 99
rect 2358 32 2380 66
rect 2414 32 2436 66
rect 2358 0 2436 32
rect 2466 66 2544 99
rect 2466 32 2488 66
rect 2522 32 2544 66
rect 2466 0 2544 32
rect 2574 66 2652 99
rect 2574 32 2596 66
rect 2630 32 2652 66
rect 2574 0 2652 32
rect 2682 66 2760 99
rect 2682 32 2704 66
rect 2738 32 2760 66
rect 2682 0 2760 32
rect 2790 66 2868 99
rect 2790 32 2812 66
rect 2846 32 2868 66
rect 2790 0 2868 32
rect 2898 66 2976 99
rect 2898 32 2920 66
rect 2954 32 2976 66
rect 2898 0 2976 32
rect 3006 66 3084 99
rect 3006 32 3028 66
rect 3062 32 3084 66
rect 3006 0 3084 32
rect 3114 66 3192 99
rect 3114 32 3136 66
rect 3170 32 3192 66
rect 3114 0 3192 32
rect 3222 66 3300 99
rect 3222 32 3244 66
rect 3278 32 3300 66
rect 3222 0 3300 32
rect 3330 66 3408 99
rect 3330 32 3352 66
rect 3386 32 3408 66
rect 3330 0 3408 32
rect 3438 66 3516 99
rect 3438 32 3460 66
rect 3494 32 3516 66
rect 3438 0 3516 32
rect 3546 66 3624 99
rect 3546 32 3568 66
rect 3602 32 3624 66
rect 3546 0 3624 32
rect 3654 66 3732 99
rect 3654 32 3676 66
rect 3710 32 3732 66
rect 3654 0 3732 32
rect 3762 66 3840 99
rect 3762 32 3784 66
rect 3818 32 3840 66
rect 3762 0 3840 32
rect 3870 66 3948 99
rect 3870 32 3892 66
rect 3926 32 3948 66
rect 3870 0 3948 32
rect 3978 66 4056 99
rect 3978 32 4000 66
rect 4034 32 4056 66
rect 3978 0 4056 32
rect 4086 66 4164 99
rect 4086 32 4108 66
rect 4142 32 4164 66
rect 4086 0 4164 32
rect 4194 66 4272 99
rect 4194 32 4216 66
rect 4250 32 4272 66
rect 4194 0 4272 32
rect 4302 66 4380 99
rect 4302 32 4324 66
rect 4358 32 4380 66
rect 4302 0 4380 32
rect 4410 66 4488 99
rect 4410 32 4432 66
rect 4466 32 4488 66
rect 4410 0 4488 32
rect 4518 66 4596 99
rect 4518 32 4540 66
rect 4574 32 4596 66
rect 4518 0 4596 32
rect 4626 66 4704 99
rect 4626 32 4648 66
rect 4682 32 4704 66
rect 4626 0 4704 32
rect 4734 66 4812 99
rect 4734 32 4756 66
rect 4790 32 4812 66
rect 4734 0 4812 32
rect 4842 66 4920 99
rect 4842 32 4864 66
rect 4898 32 4920 66
rect 4842 0 4920 32
rect 4950 66 5028 99
rect 4950 32 4972 66
rect 5006 32 5028 66
rect 4950 0 5028 32
rect 5058 66 5136 99
rect 5058 32 5080 66
rect 5114 32 5136 66
rect 5058 0 5136 32
rect 5166 66 5244 99
rect 5166 32 5188 66
rect 5222 32 5244 66
rect 5166 0 5244 32
rect 5274 66 5352 99
rect 5274 32 5296 66
rect 5330 32 5352 66
rect 5274 0 5352 32
rect 5382 66 5460 99
rect 5382 32 5404 66
rect 5438 32 5460 66
rect 5382 0 5460 32
rect 5490 66 5568 99
rect 5490 32 5512 66
rect 5546 32 5568 66
rect 5490 0 5568 32
rect 5598 66 5676 99
rect 5598 32 5620 66
rect 5654 32 5676 66
rect 5598 0 5676 32
rect 5706 66 5784 99
rect 5706 32 5728 66
rect 5762 32 5784 66
rect 5706 0 5784 32
rect 5814 66 5892 99
rect 5814 32 5836 66
rect 5870 32 5892 66
rect 5814 0 5892 32
rect 5922 66 6000 99
rect 5922 32 5944 66
rect 5978 32 6000 66
rect 5922 0 6000 32
rect 6030 66 6108 99
rect 6030 32 6052 66
rect 6086 32 6108 66
rect 6030 0 6108 32
rect 6138 66 6216 99
rect 6138 32 6160 66
rect 6194 32 6216 66
rect 6138 0 6216 32
rect 6246 66 6324 99
rect 6246 32 6268 66
rect 6302 32 6324 66
rect 6246 0 6324 32
rect 6354 66 6432 99
rect 6354 32 6376 66
rect 6410 32 6432 66
rect 6354 0 6432 32
rect 6462 66 6540 99
rect 6462 32 6484 66
rect 6518 32 6540 66
rect 6462 0 6540 32
rect 6570 66 6630 99
rect 6570 32 6588 66
rect 6622 32 6630 66
rect 6570 0 6630 32
<< ndiffc >>
rect 8 32 42 66
rect 112 32 146 66
rect 220 32 254 66
rect 328 32 362 66
rect 436 32 470 66
rect 544 32 578 66
rect 652 32 686 66
rect 760 32 794 66
rect 868 32 902 66
rect 976 32 1010 66
rect 1084 32 1118 66
rect 1192 32 1226 66
rect 1300 32 1334 66
rect 1408 32 1442 66
rect 1516 32 1550 66
rect 1624 32 1658 66
rect 1732 32 1766 66
rect 1840 32 1874 66
rect 1948 32 1982 66
rect 2056 32 2090 66
rect 2164 32 2198 66
rect 2272 32 2306 66
rect 2380 32 2414 66
rect 2488 32 2522 66
rect 2596 32 2630 66
rect 2704 32 2738 66
rect 2812 32 2846 66
rect 2920 32 2954 66
rect 3028 32 3062 66
rect 3136 32 3170 66
rect 3244 32 3278 66
rect 3352 32 3386 66
rect 3460 32 3494 66
rect 3568 32 3602 66
rect 3676 32 3710 66
rect 3784 32 3818 66
rect 3892 32 3926 66
rect 4000 32 4034 66
rect 4108 32 4142 66
rect 4216 32 4250 66
rect 4324 32 4358 66
rect 4432 32 4466 66
rect 4540 32 4574 66
rect 4648 32 4682 66
rect 4756 32 4790 66
rect 4864 32 4898 66
rect 4972 32 5006 66
rect 5080 32 5114 66
rect 5188 32 5222 66
rect 5296 32 5330 66
rect 5404 32 5438 66
rect 5512 32 5546 66
rect 5620 32 5654 66
rect 5728 32 5762 66
rect 5836 32 5870 66
rect 5944 32 5978 66
rect 6052 32 6086 66
rect 6160 32 6194 66
rect 6268 32 6302 66
rect 6376 32 6410 66
rect 6484 32 6518 66
rect 6588 32 6622 66
<< poly >>
rect 60 125 6570 155
rect 60 99 90 125
rect 168 99 198 125
rect 276 99 306 125
rect 384 99 414 125
rect 492 99 522 125
rect 600 99 630 125
rect 708 99 738 125
rect 816 99 846 125
rect 924 99 954 125
rect 1032 99 1062 125
rect 1140 99 1170 125
rect 1248 99 1278 125
rect 1356 99 1386 125
rect 1464 99 1494 125
rect 1572 99 1602 125
rect 1680 99 1710 125
rect 1788 99 1818 125
rect 1896 99 1926 125
rect 2004 99 2034 125
rect 2112 99 2142 125
rect 2220 99 2250 125
rect 2328 99 2358 125
rect 2436 99 2466 125
rect 2544 99 2574 125
rect 2652 99 2682 125
rect 2760 99 2790 125
rect 2868 99 2898 125
rect 2976 99 3006 125
rect 3084 99 3114 125
rect 3192 99 3222 125
rect 3300 99 3330 125
rect 3408 99 3438 125
rect 3516 99 3546 125
rect 3624 99 3654 125
rect 3732 99 3762 125
rect 3840 99 3870 125
rect 3948 99 3978 125
rect 4056 99 4086 125
rect 4164 99 4194 125
rect 4272 99 4302 125
rect 4380 99 4410 125
rect 4488 99 4518 125
rect 4596 99 4626 125
rect 4704 99 4734 125
rect 4812 99 4842 125
rect 4920 99 4950 125
rect 5028 99 5058 125
rect 5136 99 5166 125
rect 5244 99 5274 125
rect 5352 99 5382 125
rect 5460 99 5490 125
rect 5568 99 5598 125
rect 5676 99 5706 125
rect 5784 99 5814 125
rect 5892 99 5922 125
rect 6000 99 6030 125
rect 6108 99 6138 125
rect 6216 99 6246 125
rect 6324 99 6354 125
rect 6432 99 6462 125
rect 6540 99 6570 125
rect 60 -26 90 0
rect 168 -26 198 0
rect 276 -26 306 0
rect 384 -26 414 0
rect 492 -26 522 0
rect 600 -26 630 0
rect 708 -26 738 0
rect 816 -26 846 0
rect 924 -26 954 0
rect 1032 -26 1062 0
rect 1140 -26 1170 0
rect 1248 -26 1278 0
rect 1356 -26 1386 0
rect 1464 -26 1494 0
rect 1572 -26 1602 0
rect 1680 -26 1710 0
rect 1788 -26 1818 0
rect 1896 -26 1926 0
rect 2004 -26 2034 0
rect 2112 -26 2142 0
rect 2220 -26 2250 0
rect 2328 -26 2358 0
rect 2436 -26 2466 0
rect 2544 -26 2574 0
rect 2652 -26 2682 0
rect 2760 -26 2790 0
rect 2868 -26 2898 0
rect 2976 -26 3006 0
rect 3084 -26 3114 0
rect 3192 -26 3222 0
rect 3300 -26 3330 0
rect 3408 -26 3438 0
rect 3516 -26 3546 0
rect 3624 -26 3654 0
rect 3732 -26 3762 0
rect 3840 -26 3870 0
rect 3948 -26 3978 0
rect 4056 -26 4086 0
rect 4164 -26 4194 0
rect 4272 -26 4302 0
rect 4380 -26 4410 0
rect 4488 -26 4518 0
rect 4596 -26 4626 0
rect 4704 -26 4734 0
rect 4812 -26 4842 0
rect 4920 -26 4950 0
rect 5028 -26 5058 0
rect 5136 -26 5166 0
rect 5244 -26 5274 0
rect 5352 -26 5382 0
rect 5460 -26 5490 0
rect 5568 -26 5598 0
rect 5676 -26 5706 0
rect 5784 -26 5814 0
rect 5892 -26 5922 0
rect 6000 -26 6030 0
rect 6108 -26 6138 0
rect 6216 -26 6246 0
rect 6324 -26 6354 0
rect 6432 -26 6462 0
rect 6540 -26 6570 0
<< locali >>
rect 112 116 6622 150
rect 8 66 42 82
rect 8 16 42 32
rect 112 66 146 116
rect 112 16 146 32
rect 220 66 254 82
rect 220 16 254 32
rect 328 66 362 116
rect 328 16 362 32
rect 436 66 470 82
rect 436 16 470 32
rect 544 66 578 116
rect 544 16 578 32
rect 652 66 686 82
rect 652 16 686 32
rect 760 66 794 116
rect 760 16 794 32
rect 868 66 902 82
rect 868 16 902 32
rect 976 66 1010 116
rect 976 16 1010 32
rect 1084 66 1118 82
rect 1084 16 1118 32
rect 1192 66 1226 116
rect 1192 16 1226 32
rect 1300 66 1334 82
rect 1300 16 1334 32
rect 1408 66 1442 116
rect 1408 16 1442 32
rect 1516 66 1550 82
rect 1516 16 1550 32
rect 1624 66 1658 116
rect 1624 16 1658 32
rect 1732 66 1766 82
rect 1732 16 1766 32
rect 1840 66 1874 116
rect 1840 16 1874 32
rect 1948 66 1982 82
rect 1948 16 1982 32
rect 2056 66 2090 116
rect 2056 16 2090 32
rect 2164 66 2198 82
rect 2164 16 2198 32
rect 2272 66 2306 116
rect 2272 16 2306 32
rect 2380 66 2414 82
rect 2380 16 2414 32
rect 2488 66 2522 116
rect 2488 16 2522 32
rect 2596 66 2630 82
rect 2596 16 2630 32
rect 2704 66 2738 116
rect 2704 16 2738 32
rect 2812 66 2846 82
rect 2812 16 2846 32
rect 2920 66 2954 116
rect 2920 16 2954 32
rect 3028 66 3062 82
rect 3028 16 3062 32
rect 3136 66 3170 116
rect 3136 16 3170 32
rect 3244 66 3278 82
rect 3244 16 3278 32
rect 3352 66 3386 116
rect 3352 16 3386 32
rect 3460 66 3494 82
rect 3460 16 3494 32
rect 3568 66 3602 116
rect 3568 16 3602 32
rect 3676 66 3710 82
rect 3676 16 3710 32
rect 3784 66 3818 116
rect 3784 16 3818 32
rect 3892 66 3926 82
rect 3892 16 3926 32
rect 4000 66 4034 116
rect 4000 16 4034 32
rect 4108 66 4142 82
rect 4108 16 4142 32
rect 4216 66 4250 116
rect 4216 16 4250 32
rect 4324 66 4358 82
rect 4324 16 4358 32
rect 4432 66 4466 116
rect 4432 16 4466 32
rect 4540 66 4574 82
rect 4540 16 4574 32
rect 4648 66 4682 116
rect 4648 16 4682 32
rect 4756 66 4790 82
rect 4756 16 4790 32
rect 4864 66 4898 116
rect 4864 16 4898 32
rect 4972 66 5006 82
rect 4972 16 5006 32
rect 5080 66 5114 116
rect 5080 16 5114 32
rect 5188 66 5222 82
rect 5188 16 5222 32
rect 5296 66 5330 116
rect 5296 16 5330 32
rect 5404 66 5438 82
rect 5404 16 5438 32
rect 5512 66 5546 116
rect 5512 16 5546 32
rect 5620 66 5654 82
rect 5620 16 5654 32
rect 5728 66 5762 116
rect 5728 16 5762 32
rect 5836 66 5870 82
rect 5836 16 5870 32
rect 5944 66 5978 116
rect 5944 16 5978 32
rect 6052 66 6086 82
rect 6052 16 6086 32
rect 6160 66 6194 116
rect 6160 16 6194 32
rect 6268 66 6302 82
rect 6268 16 6302 32
rect 6376 66 6410 116
rect 6376 16 6410 32
rect 6484 66 6518 82
rect 6484 16 6518 32
rect 6588 66 6622 116
rect 6588 16 6622 32
use contact_8  contact_8_0
timestamp 1644969367
transform 1 0 6580 0 1 8
box 0 0 1 1
use contact_8  contact_8_1
timestamp 1644969367
transform 1 0 6476 0 1 8
box 0 0 1 1
use contact_8  contact_8_2
timestamp 1644969367
transform 1 0 6368 0 1 8
box 0 0 1 1
use contact_8  contact_8_3
timestamp 1644969367
transform 1 0 6260 0 1 8
box 0 0 1 1
use contact_8  contact_8_4
timestamp 1644969367
transform 1 0 6152 0 1 8
box 0 0 1 1
use contact_8  contact_8_5
timestamp 1644969367
transform 1 0 6044 0 1 8
box 0 0 1 1
use contact_8  contact_8_6
timestamp 1644969367
transform 1 0 5936 0 1 8
box 0 0 1 1
use contact_8  contact_8_7
timestamp 1644969367
transform 1 0 5828 0 1 8
box 0 0 1 1
use contact_8  contact_8_8
timestamp 1644969367
transform 1 0 5720 0 1 8
box 0 0 1 1
use contact_8  contact_8_9
timestamp 1644969367
transform 1 0 5612 0 1 8
box 0 0 1 1
use contact_8  contact_8_10
timestamp 1644969367
transform 1 0 5504 0 1 8
box 0 0 1 1
use contact_8  contact_8_11
timestamp 1644969367
transform 1 0 5396 0 1 8
box 0 0 1 1
use contact_8  contact_8_12
timestamp 1644969367
transform 1 0 5288 0 1 8
box 0 0 1 1
use contact_8  contact_8_13
timestamp 1644969367
transform 1 0 5180 0 1 8
box 0 0 1 1
use contact_8  contact_8_14
timestamp 1644969367
transform 1 0 5072 0 1 8
box 0 0 1 1
use contact_8  contact_8_15
timestamp 1644969367
transform 1 0 4964 0 1 8
box 0 0 1 1
use contact_8  contact_8_16
timestamp 1644969367
transform 1 0 4856 0 1 8
box 0 0 1 1
use contact_8  contact_8_17
timestamp 1644969367
transform 1 0 4748 0 1 8
box 0 0 1 1
use contact_8  contact_8_18
timestamp 1644969367
transform 1 0 4640 0 1 8
box 0 0 1 1
use contact_8  contact_8_19
timestamp 1644969367
transform 1 0 4532 0 1 8
box 0 0 1 1
use contact_8  contact_8_20
timestamp 1644969367
transform 1 0 4424 0 1 8
box 0 0 1 1
use contact_8  contact_8_21
timestamp 1644969367
transform 1 0 4316 0 1 8
box 0 0 1 1
use contact_8  contact_8_22
timestamp 1644969367
transform 1 0 4208 0 1 8
box 0 0 1 1
use contact_8  contact_8_23
timestamp 1644969367
transform 1 0 4100 0 1 8
box 0 0 1 1
use contact_8  contact_8_24
timestamp 1644969367
transform 1 0 3992 0 1 8
box 0 0 1 1
use contact_8  contact_8_25
timestamp 1644969367
transform 1 0 3884 0 1 8
box 0 0 1 1
use contact_8  contact_8_26
timestamp 1644969367
transform 1 0 3776 0 1 8
box 0 0 1 1
use contact_8  contact_8_27
timestamp 1644969367
transform 1 0 3668 0 1 8
box 0 0 1 1
use contact_8  contact_8_28
timestamp 1644969367
transform 1 0 3560 0 1 8
box 0 0 1 1
use contact_8  contact_8_29
timestamp 1644969367
transform 1 0 3452 0 1 8
box 0 0 1 1
use contact_8  contact_8_30
timestamp 1644969367
transform 1 0 3344 0 1 8
box 0 0 1 1
use contact_8  contact_8_31
timestamp 1644969367
transform 1 0 3236 0 1 8
box 0 0 1 1
use contact_8  contact_8_32
timestamp 1644969367
transform 1 0 3128 0 1 8
box 0 0 1 1
use contact_8  contact_8_33
timestamp 1644969367
transform 1 0 3020 0 1 8
box 0 0 1 1
use contact_8  contact_8_34
timestamp 1644969367
transform 1 0 2912 0 1 8
box 0 0 1 1
use contact_8  contact_8_35
timestamp 1644969367
transform 1 0 2804 0 1 8
box 0 0 1 1
use contact_8  contact_8_36
timestamp 1644969367
transform 1 0 2696 0 1 8
box 0 0 1 1
use contact_8  contact_8_37
timestamp 1644969367
transform 1 0 2588 0 1 8
box 0 0 1 1
use contact_8  contact_8_38
timestamp 1644969367
transform 1 0 2480 0 1 8
box 0 0 1 1
use contact_8  contact_8_39
timestamp 1644969367
transform 1 0 2372 0 1 8
box 0 0 1 1
use contact_8  contact_8_40
timestamp 1644969367
transform 1 0 2264 0 1 8
box 0 0 1 1
use contact_8  contact_8_41
timestamp 1644969367
transform 1 0 2156 0 1 8
box 0 0 1 1
use contact_8  contact_8_42
timestamp 1644969367
transform 1 0 2048 0 1 8
box 0 0 1 1
use contact_8  contact_8_43
timestamp 1644969367
transform 1 0 1940 0 1 8
box 0 0 1 1
use contact_8  contact_8_44
timestamp 1644969367
transform 1 0 1832 0 1 8
box 0 0 1 1
use contact_8  contact_8_45
timestamp 1644969367
transform 1 0 1724 0 1 8
box 0 0 1 1
use contact_8  contact_8_46
timestamp 1644969367
transform 1 0 1616 0 1 8
box 0 0 1 1
use contact_8  contact_8_47
timestamp 1644969367
transform 1 0 1508 0 1 8
box 0 0 1 1
use contact_8  contact_8_48
timestamp 1644969367
transform 1 0 1400 0 1 8
box 0 0 1 1
use contact_8  contact_8_49
timestamp 1644969367
transform 1 0 1292 0 1 8
box 0 0 1 1
use contact_8  contact_8_50
timestamp 1644969367
transform 1 0 1184 0 1 8
box 0 0 1 1
use contact_8  contact_8_51
timestamp 1644969367
transform 1 0 1076 0 1 8
box 0 0 1 1
use contact_8  contact_8_52
timestamp 1644969367
transform 1 0 968 0 1 8
box 0 0 1 1
use contact_8  contact_8_53
timestamp 1644969367
transform 1 0 860 0 1 8
box 0 0 1 1
use contact_8  contact_8_54
timestamp 1644969367
transform 1 0 752 0 1 8
box 0 0 1 1
use contact_8  contact_8_55
timestamp 1644969367
transform 1 0 644 0 1 8
box 0 0 1 1
use contact_8  contact_8_56
timestamp 1644969367
transform 1 0 536 0 1 8
box 0 0 1 1
use contact_8  contact_8_57
timestamp 1644969367
transform 1 0 428 0 1 8
box 0 0 1 1
use contact_8  contact_8_58
timestamp 1644969367
transform 1 0 320 0 1 8
box 0 0 1 1
use contact_8  contact_8_59
timestamp 1644969367
transform 1 0 212 0 1 8
box 0 0 1 1
use contact_8  contact_8_60
timestamp 1644969367
transform 1 0 104 0 1 8
box 0 0 1 1
use contact_8  contact_8_61
timestamp 1644969367
transform 1 0 0 0 1 8
box 0 0 1 1
<< labels >>
rlabel mvvaractor s 3315 140 3315 140 4 G
rlabel locali s 1533 49 1533 49 4 S
rlabel locali s 3045 49 3045 49 4 S
rlabel locali s 4125 49 4125 49 4 S
rlabel locali s 1101 49 1101 49 4 S
rlabel locali s 2613 49 2613 49 4 S
rlabel locali s 6501 49 6501 49 4 S
rlabel locali s 2829 49 2829 49 4 S
rlabel locali s 3909 49 3909 49 4 S
rlabel locali s 4773 49 4773 49 4 S
rlabel locali s 5637 49 5637 49 4 S
rlabel locali s 2397 49 2397 49 4 S
rlabel locali s 1749 49 1749 49 4 S
rlabel locali s 4989 49 4989 49 4 S
rlabel locali s 1965 49 1965 49 4 S
rlabel locali s 6285 49 6285 49 4 S
rlabel locali s 4557 49 4557 49 4 S
rlabel locali s 3261 49 3261 49 4 S
rlabel locali s 5205 49 5205 49 4 S
rlabel locali s 2181 49 2181 49 4 S
rlabel locali s 1317 49 1317 49 4 S
rlabel locali s 237 49 237 49 4 S
rlabel locali s 669 49 669 49 4 S
rlabel locali s 3693 49 3693 49 4 S
rlabel locali s 25 49 25 49 4 S
rlabel locali s 5421 49 5421 49 4 S
rlabel locali s 6069 49 6069 49 4 S
rlabel locali s 4341 49 4341 49 4 S
rlabel locali s 885 49 885 49 4 S
rlabel locali s 3477 49 3477 49 4 S
rlabel locali s 453 49 453 49 4 S
rlabel locali s 5853 49 5853 49 4 S
rlabel locali s 3367 133 3367 133 4 D
<< properties >>
string FIXED_BBOX -25 -26 6655 155
string GDS_FILE sram_0rw2r1w_32_128_sky130A.gds
string GDS_END 3360380
string GDS_START 3347792
<< end >>
