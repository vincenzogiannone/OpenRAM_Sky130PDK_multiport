VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO sram_0rw2r1w_16_32_sky130A
   CLASS BLOCK ;
   SIZE 376.5 BY 187.5 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  84.6 0.0 84.9 0.9 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  91.2 0.0 91.5 0.9 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  98.4 0.0 98.7 0.9 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  106.8 0.0 107.1 0.9 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  114.0 0.0 114.3 0.9 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  121.8 0.0 122.1 0.9 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  129.0 0.0 129.3 0.9 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  136.2 0.0 136.5 0.9 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  144.0 0.0 144.3 0.9 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  151.2 0.0 151.5 0.9 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  158.4 0.0 158.7 0.9 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  165.6 0.0 165.9 0.9 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  172.8 0.0 173.1 0.9 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  180.0 0.0 180.3 0.9 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  188.4 0.0 188.7 0.9 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  195.6 0.0 195.9 0.9 ;
      END
   END din0[15]
   PIN addr[0]
      DIRECTION INPUT ;
      PORT
      END
   END addr[0]
   PIN addr[1]
      DIRECTION INPUT ;
      PORT
      END
   END addr[1]
   PIN addr[2]
      DIRECTION INPUT ;
      PORT
      END
   END addr[2]
   PIN addr[3]
      DIRECTION INPUT ;
      PORT
      END
   END addr[3]
   PIN addr[4]
      DIRECTION INPUT ;
      PORT
      END
   END addr[4]
   PIN addr[5]
      DIRECTION INPUT ;
      PORT
      END
   END addr[5]
   PIN addr[6]
      DIRECTION INPUT ;
      PORT
      END
   END addr[6]
   PIN csb
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  13.175 30.19 13.475 30.49 ;
      END
   END csb
   PIN web
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  13.175 24.27 13.475 24.57 ;
      END
   END web
   PIN clk
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  30.0 0.0 30.3 0.9 ;
      END
   END clk
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  124.2 0.0 124.5 0.9 ;
      END
   END dout0[0]
   PIN dout1[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  123.6 46.25 123.9 46.55 ;
      END
   END dout1[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  131.4 0.0 131.7 0.9 ;
      END
   END dout0[1]
   PIN dout1[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  131.38 46.25 131.68 46.55 ;
      END
   END dout1[1]
   PIN dout0[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  139.2 0.0 139.5 0.9 ;
      END
   END dout0[2]
   PIN dout1[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  139.16 46.25 139.46 46.55 ;
      END
   END dout1[2]
   PIN dout0[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  147.0 0.0 147.3 0.9 ;
      END
   END dout0[3]
   PIN dout1[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  146.94 46.25 147.24 46.55 ;
      END
   END dout1[3]
   PIN dout0[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  154.8 0.0 155.1 0.9 ;
      END
   END dout0[4]
   PIN dout1[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  154.72 46.25 155.02 46.55 ;
      END
   END dout1[4]
   PIN dout0[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  162.6 0.0 162.9 0.9 ;
      END
   END dout0[5]
   PIN dout1[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  162.5 46.25 162.8 46.55 ;
      END
   END dout1[5]
   PIN dout0[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  170.4 0.0 170.7 0.9 ;
      END
   END dout0[6]
   PIN dout1[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  170.28 46.25 170.58 46.55 ;
      END
   END dout1[6]
   PIN dout0[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  178.2 0.0 178.5 0.9 ;
      END
   END dout0[7]
   PIN dout1[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  178.06 46.25 178.36 46.55 ;
      END
   END dout1[7]
   PIN dout0[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  186.0 0.0 186.3 0.9 ;
      END
   END dout0[8]
   PIN dout1[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  185.84 46.25 186.14 46.55 ;
      END
   END dout1[8]
   PIN dout0[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  193.8 0.0 194.1 0.9 ;
      END
   END dout0[9]
   PIN dout1[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  193.62 46.25 193.92 46.55 ;
      END
   END dout1[9]
   PIN dout0[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  201.6 0.0 201.9 0.9 ;
      END
   END dout0[10]
   PIN dout1[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  201.4 46.25 201.7 46.55 ;
      END
   END dout1[10]
   PIN dout0[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  209.4 0.0 209.7 0.9 ;
      END
   END dout0[11]
   PIN dout1[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  209.18 46.25 209.48 46.55 ;
      END
   END dout1[11]
   PIN dout0[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  217.2 0.0 217.5 0.9 ;
      END
   END dout0[12]
   PIN dout1[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  216.96 46.25 217.26 46.55 ;
      END
   END dout1[12]
   PIN dout0[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  225.0 0.0 225.3 0.9 ;
      END
   END dout0[13]
   PIN dout1[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  224.74 46.25 225.04 46.55 ;
      END
   END dout1[13]
   PIN dout0[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  232.8 0.0 233.1 0.9 ;
      END
   END dout0[14]
   PIN dout1[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  232.52 46.25 232.82 46.55 ;
      END
   END dout1[14]
   PIN dout0[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  240.6 0.0 240.9 0.9 ;
      END
   END dout0[15]
   PIN dout1[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  240.3 46.25 240.6 46.55 ;
      END
   END dout1[15]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met4 ;
         RECT  372.0 4.2 373.5 184.5 ;
         LAYER met3 ;
         RECT  4.2 4.2 373.5 5.7 ;
         LAYER met4 ;
         RECT  4.2 4.2 5.7 184.5 ;
         LAYER met3 ;
         RECT  4.2 183.0 373.5 184.5 ;
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met4 ;
         RECT  1.2 1.2 2.7 187.5 ;
         LAYER met4 ;
         RECT  375.0 1.2 376.5 187.5 ;
         LAYER met3 ;
         RECT  1.2 186.0 376.5 187.5 ;
         LAYER met3 ;
         RECT  1.2 1.2 376.5 2.7 ;
      END
   END gnd
   OBS
   LAYER  met1 ;
      RECT  0.6 0.6 375.9 186.9 ;
   LAYER  met2 ;
      RECT  0.6 0.6 375.9 186.9 ;
   LAYER  met3 ;
      RECT  0.6 29.59 12.575 31.09 ;
      RECT  14.075 29.59 375.9 31.09 ;
      RECT  12.575 25.17 14.075 29.59 ;
      RECT  14.075 31.09 123.0 45.65 ;
      RECT  14.075 45.65 123.0 47.15 ;
      RECT  123.0 31.09 124.5 45.65 ;
      RECT  124.5 31.09 375.9 45.65 ;
      RECT  124.5 45.65 130.78 47.15 ;
      RECT  132.28 45.65 138.56 47.15 ;
      RECT  140.06 45.65 146.34 47.15 ;
      RECT  147.84 45.65 154.12 47.15 ;
      RECT  155.62 45.65 161.9 47.15 ;
      RECT  163.4 45.65 169.68 47.15 ;
      RECT  171.18 45.65 177.46 47.15 ;
      RECT  178.96 45.65 185.24 47.15 ;
      RECT  186.74 45.65 193.02 47.15 ;
      RECT  194.52 45.65 200.8 47.15 ;
      RECT  202.3 45.65 208.58 47.15 ;
      RECT  210.08 45.65 216.36 47.15 ;
      RECT  217.86 45.65 224.14 47.15 ;
      RECT  225.64 45.65 231.92 47.15 ;
      RECT  233.42 45.65 239.7 47.15 ;
      RECT  241.2 45.65 375.9 47.15 ;
      RECT  0.6 3.6 3.6 6.3 ;
      RECT  0.6 6.3 3.6 29.59 ;
      RECT  3.6 6.3 12.575 29.59 ;
      RECT  14.075 6.3 374.1 29.59 ;
      RECT  374.1 3.6 375.9 6.3 ;
      RECT  374.1 6.3 375.9 29.59 ;
      RECT  12.575 6.3 14.075 23.67 ;
      RECT  0.6 31.09 3.6 182.4 ;
      RECT  0.6 182.4 3.6 185.1 ;
      RECT  3.6 31.09 12.575 182.4 ;
      RECT  12.575 31.09 14.075 182.4 ;
      RECT  14.075 47.15 123.0 182.4 ;
      RECT  123.0 47.15 124.5 182.4 ;
      RECT  124.5 47.15 374.1 182.4 ;
      RECT  374.1 47.15 375.9 182.4 ;
      RECT  374.1 182.4 375.9 185.1 ;
      RECT  0.6 185.1 3.6 185.4 ;
      RECT  3.6 185.1 12.575 185.4 ;
      RECT  12.575 185.1 14.075 185.4 ;
      RECT  14.075 185.1 123.0 185.4 ;
      RECT  123.0 185.1 124.5 185.4 ;
      RECT  124.5 185.1 374.1 185.4 ;
      RECT  374.1 185.1 375.9 185.4 ;
      RECT  0.6 3.3 3.6 3.6 ;
      RECT  3.6 3.3 12.575 3.6 ;
      RECT  14.075 3.3 374.1 3.6 ;
      RECT  374.1 3.3 375.9 3.6 ;
      RECT  12.575 3.3 14.075 3.6 ;
   LAYER  met4 ;
      RECT  84.0 1.5 85.5 186.9 ;
      RECT  85.5 0.6 90.6 1.5 ;
      RECT  92.1 0.6 97.8 1.5 ;
      RECT  99.3 0.6 106.2 1.5 ;
      RECT  107.7 0.6 113.4 1.5 ;
      RECT  114.9 0.6 121.2 1.5 ;
      RECT  30.9 0.6 84.0 1.5 ;
      RECT  122.7 0.6 123.6 1.5 ;
      RECT  125.1 0.6 128.4 1.5 ;
      RECT  129.9 0.6 130.8 1.5 ;
      RECT  132.3 0.6 135.6 1.5 ;
      RECT  137.1 0.6 138.6 1.5 ;
      RECT  140.1 0.6 143.4 1.5 ;
      RECT  144.9 0.6 146.4 1.5 ;
      RECT  147.9 0.6 150.6 1.5 ;
      RECT  152.1 0.6 154.2 1.5 ;
      RECT  155.7 0.6 157.8 1.5 ;
      RECT  159.3 0.6 162.0 1.5 ;
      RECT  163.5 0.6 165.0 1.5 ;
      RECT  166.5 0.6 169.8 1.5 ;
      RECT  171.3 0.6 172.2 1.5 ;
      RECT  173.7 0.6 177.6 1.5 ;
      RECT  179.1 0.6 179.4 1.5 ;
      RECT  180.9 0.6 185.4 1.5 ;
      RECT  186.9 0.6 187.8 1.5 ;
      RECT  189.3 0.6 193.2 1.5 ;
      RECT  194.7 0.6 195.0 1.5 ;
      RECT  196.5 0.6 201.0 1.5 ;
      RECT  202.5 0.6 208.8 1.5 ;
      RECT  210.3 0.6 216.6 1.5 ;
      RECT  218.1 0.6 224.4 1.5 ;
      RECT  225.9 0.6 232.2 1.5 ;
      RECT  233.7 0.6 240.0 1.5 ;
      RECT  85.5 1.5 371.4 3.6 ;
      RECT  85.5 3.6 371.4 185.1 ;
      RECT  85.5 185.1 371.4 186.9 ;
      RECT  371.4 1.5 374.1 3.6 ;
      RECT  371.4 185.1 374.1 186.9 ;
      RECT  3.6 1.5 6.3 3.6 ;
      RECT  3.6 185.1 6.3 186.9 ;
      RECT  6.3 1.5 84.0 3.6 ;
      RECT  6.3 3.6 84.0 185.1 ;
      RECT  6.3 185.1 84.0 186.9 ;
      RECT  3.3 0.6 29.4 1.5 ;
      RECT  3.3 1.5 3.6 3.6 ;
      RECT  3.3 3.6 3.6 185.1 ;
      RECT  3.3 185.1 3.6 186.9 ;
      RECT  241.5 0.6 374.4 1.5 ;
      RECT  374.1 1.5 374.4 3.6 ;
      RECT  374.1 3.6 374.4 185.1 ;
      RECT  374.1 185.1 374.4 186.9 ;
   END
END    sram_0rw2r1w_16_32_sky130A
END    LIBRARY
