magic
tech sky130A
timestamp 1644949024
<< checkpaint >>
rect -630 -651 2186 12971
<< metal1 >>
rect 0 12305 1556 12336
rect 0 11984 1556 11998
rect 0 11921 1556 11935
rect 0 11808 1556 11822
rect 0 11534 1556 11566
rect 0 11278 1556 11292
rect 0 11165 1556 11179
rect 0 11102 1556 11116
rect 0 10764 1556 10796
rect 0 10444 1556 10458
rect 0 10381 1556 10395
rect 0 10268 1556 10282
rect 0 9994 1556 10026
rect 0 9738 1556 9752
rect 0 9625 1556 9639
rect 0 9562 1556 9576
rect 0 9224 1556 9256
rect 0 8904 1556 8918
rect 0 8841 1556 8855
rect 0 8728 1556 8742
rect 0 8454 1556 8486
rect 0 8198 1556 8212
rect 0 8085 1556 8099
rect 0 8022 1556 8036
rect 0 7684 1556 7716
rect 0 7364 1556 7378
rect 0 7301 1556 7315
rect 0 7188 1556 7202
rect 0 6914 1556 6946
rect 0 6658 1556 6672
rect 0 6545 1556 6559
rect 0 6482 1556 6496
rect 0 6144 1556 6176
rect 0 5824 1556 5838
rect 0 5761 1556 5775
rect 0 5648 1556 5662
rect 0 5374 1556 5406
rect 0 5118 1556 5132
rect 0 5005 1556 5019
rect 0 4942 1556 4956
rect 0 4604 1556 4636
rect 0 4284 1556 4298
rect 0 4221 1556 4235
rect 0 4108 1556 4122
rect 0 3834 1556 3866
rect 0 3578 1556 3592
rect 0 3465 1556 3479
rect 0 3402 1556 3416
rect 0 3064 1556 3096
rect 0 2744 1556 2758
rect 0 2681 1556 2695
rect 0 2568 1556 2582
rect 0 2294 1556 2326
rect 0 2038 1556 2052
rect 0 1925 1556 1939
rect 0 1862 1556 1876
rect 0 1524 1556 1556
rect 0 1204 1556 1218
rect 0 1141 1556 1155
rect 0 1028 1556 1042
rect 0 754 1556 786
rect 0 498 1556 512
rect 0 385 1556 399
rect 0 322 1556 336
rect 0 -16 1556 15
<< metal2 >>
rect 96 0 110 12320
rect 222 0 236 12320
rect 313 0 327 12320
rect 485 0 499 12320
rect 611 0 625 12320
rect 702 0 716 12320
rect 874 0 888 12320
rect 1000 0 1014 12320
rect 1091 0 1105 12320
rect 1263 0 1277 12320
rect 1389 0 1403 12320
rect 1480 0 1494 12320
use cell_2r1w  cell_2r1w_0
timestamp 1644949024
transform 1 0 1167 0 -1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1
timestamp 1644949024
transform 1 0 1167 0 1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_2
timestamp 1644949024
transform 1 0 1167 0 -1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_3
timestamp 1644949024
transform 1 0 1167 0 1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_4
timestamp 1644949024
transform 1 0 1167 0 -1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_5
timestamp 1644949024
transform 1 0 1167 0 1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_6
timestamp 1644949024
transform 1 0 1167 0 -1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_7
timestamp 1644949024
transform 1 0 1167 0 1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_8
timestamp 1644949024
transform 1 0 1167 0 -1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_9
timestamp 1644949024
transform 1 0 1167 0 1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_10
timestamp 1644949024
transform 1 0 1167 0 -1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_11
timestamp 1644949024
transform 1 0 1167 0 1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_12
timestamp 1644949024
transform 1 0 1167 0 -1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_13
timestamp 1644949024
transform 1 0 1167 0 1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_14
timestamp 1644949024
transform 1 0 1167 0 -1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_15
timestamp 1644949024
transform 1 0 1167 0 1 0
box 0 -21 389 808
use cell_2r1w  cell_2r1w_16
timestamp 1644949024
transform 1 0 778 0 -1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_17
timestamp 1644949024
transform 1 0 778 0 1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_18
timestamp 1644949024
transform 1 0 778 0 -1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_19
timestamp 1644949024
transform 1 0 778 0 1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_20
timestamp 1644949024
transform 1 0 778 0 -1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_21
timestamp 1644949024
transform 1 0 778 0 1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_22
timestamp 1644949024
transform 1 0 778 0 -1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_23
timestamp 1644949024
transform 1 0 778 0 1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_24
timestamp 1644949024
transform 1 0 778 0 -1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_25
timestamp 1644949024
transform 1 0 778 0 1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_26
timestamp 1644949024
transform 1 0 778 0 -1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_27
timestamp 1644949024
transform 1 0 778 0 1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_28
timestamp 1644949024
transform 1 0 778 0 -1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_29
timestamp 1644949024
transform 1 0 778 0 1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_30
timestamp 1644949024
transform 1 0 778 0 -1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_31
timestamp 1644949024
transform 1 0 778 0 1 0
box 0 -21 389 808
use cell_2r1w  cell_2r1w_32
timestamp 1644949024
transform 1 0 389 0 -1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_33
timestamp 1644949024
transform 1 0 389 0 1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_34
timestamp 1644949024
transform 1 0 389 0 -1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_35
timestamp 1644949024
transform 1 0 389 0 1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_36
timestamp 1644949024
transform 1 0 389 0 -1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_37
timestamp 1644949024
transform 1 0 389 0 1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_38
timestamp 1644949024
transform 1 0 389 0 -1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_39
timestamp 1644949024
transform 1 0 389 0 1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_40
timestamp 1644949024
transform 1 0 389 0 -1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_41
timestamp 1644949024
transform 1 0 389 0 1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_42
timestamp 1644949024
transform 1 0 389 0 -1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_43
timestamp 1644949024
transform 1 0 389 0 1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_44
timestamp 1644949024
transform 1 0 389 0 -1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_45
timestamp 1644949024
transform 1 0 389 0 1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_46
timestamp 1644949024
transform 1 0 389 0 -1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_47
timestamp 1644949024
transform 1 0 389 0 1 0
box 0 -21 389 808
use cell_2r1w  cell_2r1w_48
timestamp 1644949024
transform 1 0 0 0 -1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_49
timestamp 1644949024
transform 1 0 0 0 1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_50
timestamp 1644949024
transform 1 0 0 0 -1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_51
timestamp 1644949024
transform 1 0 0 0 1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_52
timestamp 1644949024
transform 1 0 0 0 -1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_53
timestamp 1644949024
transform 1 0 0 0 1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_54
timestamp 1644949024
transform 1 0 0 0 -1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_55
timestamp 1644949024
transform 1 0 0 0 1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_56
timestamp 1644949024
transform 1 0 0 0 -1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_57
timestamp 1644949024
transform 1 0 0 0 1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_58
timestamp 1644949024
transform 1 0 0 0 -1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_59
timestamp 1644949024
transform 1 0 0 0 1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_60
timestamp 1644949024
transform 1 0 0 0 -1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_61
timestamp 1644949024
transform 1 0 0 0 1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_62
timestamp 1644949024
transform 1 0 0 0 -1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_63
timestamp 1644949024
transform 1 0 0 0 1 0
box 0 -21 389 808
<< labels >>
rlabel metal2 s 96 0 110 12320 4 read_bl_0_0
rlabel metal2 s 222 0 236 12320 4 read_bl_1_0
rlabel metal2 s 313 0 327 12320 4 write_bl_0_0
rlabel metal2 s 485 0 499 12320 4 read_bl_0_1
rlabel metal2 s 611 0 625 12320 4 read_bl_1_1
rlabel metal2 s 702 0 716 12320 4 write_bl_0_1
rlabel metal2 s 874 0 888 12320 4 read_bl_0_2
rlabel metal2 s 1000 0 1014 12320 4 read_bl_1_2
rlabel metal2 s 1091 0 1105 12320 4 write_bl_0_2
rlabel metal2 s 1263 0 1277 12320 4 read_bl_0_3
rlabel metal2 s 1389 0 1403 12320 4 read_bl_1_3
rlabel metal2 s 1480 0 1494 12320 4 write_bl_0_3
rlabel metal1 s 0 385 1556 399 4 rwl_0_0
rlabel metal1 s 0 498 1556 512 4 rwl_1_0
rlabel metal1 s 0 322 1556 336 4 wwl_0_0
rlabel metal1 s 0 1141 1556 1155 4 rwl_0_1
rlabel metal1 s 0 1028 1556 1042 4 rwl_1_1
rlabel metal1 s 0 1204 1556 1218 4 wwl_0_1
rlabel metal1 s 0 1925 1556 1939 4 rwl_0_2
rlabel metal1 s 0 2038 1556 2052 4 rwl_1_2
rlabel metal1 s 0 1862 1556 1876 4 wwl_0_2
rlabel metal1 s 0 2681 1556 2695 4 rwl_0_3
rlabel metal1 s 0 2568 1556 2582 4 rwl_1_3
rlabel metal1 s 0 2744 1556 2758 4 wwl_0_3
rlabel metal1 s 0 3465 1556 3479 4 rwl_0_4
rlabel metal1 s 0 3578 1556 3592 4 rwl_1_4
rlabel metal1 s 0 3402 1556 3416 4 wwl_0_4
rlabel metal1 s 0 4221 1556 4235 4 rwl_0_5
rlabel metal1 s 0 4108 1556 4122 4 rwl_1_5
rlabel metal1 s 0 4284 1556 4298 4 wwl_0_5
rlabel metal1 s 0 5005 1556 5019 4 rwl_0_6
rlabel metal1 s 0 5118 1556 5132 4 rwl_1_6
rlabel metal1 s 0 4942 1556 4956 4 wwl_0_6
rlabel metal1 s 0 5761 1556 5775 4 rwl_0_7
rlabel metal1 s 0 5648 1556 5662 4 rwl_1_7
rlabel metal1 s 0 5824 1556 5838 4 wwl_0_7
rlabel metal1 s 0 6545 1556 6559 4 rwl_0_8
rlabel metal1 s 0 6658 1556 6672 4 rwl_1_8
rlabel metal1 s 0 6482 1556 6496 4 wwl_0_8
rlabel metal1 s 0 7301 1556 7315 4 rwl_0_9
rlabel metal1 s 0 7188 1556 7202 4 rwl_1_9
rlabel metal1 s 0 7364 1556 7378 4 wwl_0_9
rlabel metal1 s 0 8085 1556 8099 4 rwl_0_10
rlabel metal1 s 0 8198 1556 8212 4 rwl_1_10
rlabel metal1 s 0 8022 1556 8036 4 wwl_0_10
rlabel metal1 s 0 8841 1556 8855 4 rwl_0_11
rlabel metal1 s 0 8728 1556 8742 4 rwl_1_11
rlabel metal1 s 0 8904 1556 8918 4 wwl_0_11
rlabel metal1 s 0 9625 1556 9639 4 rwl_0_12
rlabel metal1 s 0 9738 1556 9752 4 rwl_1_12
rlabel metal1 s 0 9562 1556 9576 4 wwl_0_12
rlabel metal1 s 0 10381 1556 10395 4 rwl_0_13
rlabel metal1 s 0 10268 1556 10282 4 rwl_1_13
rlabel metal1 s 0 10444 1556 10458 4 wwl_0_13
rlabel metal1 s 0 11165 1556 11179 4 rwl_0_14
rlabel metal1 s 0 11278 1556 11292 4 rwl_1_14
rlabel metal1 s 0 11102 1556 11116 4 wwl_0_14
rlabel metal1 s 0 11921 1556 11935 4 rwl_0_15
rlabel metal1 s 0 11808 1556 11822 4 rwl_1_15
rlabel metal1 s 0 11984 1556 11998 4 wwl_0_15
rlabel metal1 s 389 5375 778 5406 4 vdd
rlabel metal1 s 389 5374 778 5405 4 vdd
rlabel metal1 s 389 9995 778 10026 4 vdd
rlabel metal1 s 778 9994 1167 10025 4 vdd
rlabel metal1 s 0 9994 389 10025 4 vdd
rlabel metal1 s 0 754 389 785 4 vdd
rlabel metal1 s 778 8455 1167 8486 4 vdd
rlabel metal1 s 778 2294 1167 2325 4 vdd
rlabel metal1 s 778 2295 1167 2326 4 vdd
rlabel metal1 s 0 2294 389 2325 4 vdd
rlabel metal1 s 778 6914 1167 6945 4 vdd
rlabel metal1 s 389 8454 778 8485 4 vdd
rlabel metal1 s 1167 11534 1556 11565 4 vdd
rlabel metal1 s 0 3835 389 3866 4 vdd
rlabel metal1 s 778 3835 1167 3866 4 vdd
rlabel metal1 s 778 8454 1167 8485 4 vdd
rlabel metal1 s 0 8455 389 8486 4 vdd
rlabel metal1 s 1167 9995 1556 10026 4 vdd
rlabel metal1 s 389 8455 778 8486 4 vdd
rlabel metal1 s 389 755 778 786 4 vdd
rlabel metal1 s 1167 8455 1556 8486 4 vdd
rlabel metal1 s 1167 2294 1556 2325 4 vdd
rlabel metal1 s 778 11535 1167 11566 4 vdd
rlabel metal1 s 389 3835 778 3866 4 vdd
rlabel metal1 s 778 9995 1167 10026 4 vdd
rlabel metal1 s 1167 6914 1556 6945 4 vdd
rlabel metal1 s 0 6915 389 6946 4 vdd
rlabel metal1 s 1167 755 1556 786 4 vdd
rlabel metal1 s 0 3834 389 3865 4 vdd
rlabel metal1 s 778 5374 1167 5405 4 vdd
rlabel metal1 s 0 6914 389 6945 4 vdd
rlabel metal1 s 1167 5375 1556 5406 4 vdd
rlabel metal1 s 0 9995 389 10026 4 vdd
rlabel metal1 s 0 11535 389 11566 4 vdd
rlabel metal1 s 389 3834 778 3865 4 vdd
rlabel metal1 s 0 5374 389 5405 4 vdd
rlabel metal1 s 1167 11535 1556 11566 4 vdd
rlabel metal1 s 1167 2295 1556 2326 4 vdd
rlabel metal1 s 0 11534 389 11565 4 vdd
rlabel metal1 s 389 2294 778 2325 4 vdd
rlabel metal1 s 1167 3834 1556 3865 4 vdd
rlabel metal1 s 389 6915 778 6946 4 vdd
rlabel metal1 s 778 3834 1167 3865 4 vdd
rlabel metal1 s 1167 9994 1556 10025 4 vdd
rlabel metal1 s 389 6914 778 6945 4 vdd
rlabel metal1 s 1167 3835 1556 3866 4 vdd
rlabel metal1 s 0 755 389 786 4 vdd
rlabel metal1 s 1167 754 1556 785 4 vdd
rlabel metal1 s 778 6915 1167 6946 4 vdd
rlabel metal1 s 389 11534 778 11565 4 vdd
rlabel metal1 s 778 5375 1167 5406 4 vdd
rlabel metal1 s 389 754 778 785 4 vdd
rlabel metal1 s 389 9994 778 10025 4 vdd
rlabel metal1 s 389 2295 778 2326 4 vdd
rlabel metal1 s 0 2295 389 2326 4 vdd
rlabel metal1 s 1167 5374 1556 5405 4 vdd
rlabel metal1 s 0 8454 389 8485 4 vdd
rlabel metal1 s 0 5375 389 5406 4 vdd
rlabel metal1 s 1167 6915 1556 6946 4 vdd
rlabel metal1 s 1167 8454 1556 8485 4 vdd
rlabel metal1 s 389 11535 778 11566 4 vdd
rlabel metal1 s 778 11534 1167 11565 4 vdd
rlabel metal1 s 778 754 1167 785 4 vdd
rlabel metal1 s 778 755 1167 786 4 vdd
rlabel metal1 s 0 3064 389 3095 4 gnd
rlabel metal1 s 1167 1524 1556 1555 4 gnd
rlabel metal1 s 778 3065 1167 3096 4 gnd
rlabel metal1 s 389 1525 778 1556 4 gnd
rlabel metal1 s 0 9225 389 9256 4 gnd
rlabel metal1 s 1167 9224 1556 9255 4 gnd
rlabel metal1 s 389 1524 778 1555 4 gnd
rlabel metal1 s 389 7685 778 7716 4 gnd
rlabel metal1 s 1167 9225 1556 9256 4 gnd
rlabel metal1 s 778 7685 1167 7716 4 gnd
rlabel metal1 s 389 4605 778 4636 4 gnd
rlabel metal1 s 0 4604 389 4635 4 gnd
rlabel metal1 s 0 12305 389 12336 4 gnd
rlabel metal1 s 1167 1525 1556 1556 4 gnd
rlabel metal1 s 778 10764 1167 10795 4 gnd
rlabel metal1 s 778 3064 1167 3095 4 gnd
rlabel metal1 s 389 7684 778 7715 4 gnd
rlabel metal1 s 389 6144 778 6175 4 gnd
rlabel metal1 s 389 9225 778 9256 4 gnd
rlabel metal1 s 778 4604 1167 4635 4 gnd
rlabel metal1 s 389 9224 778 9255 4 gnd
rlabel metal1 s 778 6145 1167 6176 4 gnd
rlabel metal1 s 0 3065 389 3096 4 gnd
rlabel metal1 s 778 12305 1167 12336 4 gnd
rlabel metal1 s 778 1525 1167 1556 4 gnd
rlabel metal1 s 389 10765 778 10796 4 gnd
rlabel metal1 s 1167 12305 1556 12336 4 gnd
rlabel metal1 s 0 1524 389 1555 4 gnd
rlabel metal1 s 389 10764 778 10795 4 gnd
rlabel metal1 s 1167 6144 1556 6175 4 gnd
rlabel metal1 s 389 3064 778 3095 4 gnd
rlabel metal1 s 778 6144 1167 6175 4 gnd
rlabel metal1 s 0 -16 389 15 4 gnd
rlabel metal1 s 1167 7684 1556 7715 4 gnd
rlabel metal1 s 0 6145 389 6176 4 gnd
rlabel metal1 s 389 -16 778 15 4 gnd
rlabel metal1 s 778 9224 1167 9255 4 gnd
rlabel metal1 s 778 1524 1167 1555 4 gnd
rlabel metal1 s 0 10764 389 10795 4 gnd
rlabel metal1 s 0 7685 389 7716 4 gnd
rlabel metal1 s 0 6144 389 6175 4 gnd
rlabel metal1 s 389 4604 778 4635 4 gnd
rlabel metal1 s 778 10765 1167 10796 4 gnd
rlabel metal1 s 0 7684 389 7715 4 gnd
rlabel metal1 s 778 -16 1167 15 4 gnd
rlabel metal1 s 0 4605 389 4636 4 gnd
rlabel metal1 s 389 6145 778 6176 4 gnd
rlabel metal1 s 778 4605 1167 4636 4 gnd
rlabel metal1 s 1167 10764 1556 10795 4 gnd
rlabel metal1 s 389 12305 778 12336 4 gnd
rlabel metal1 s 0 9224 389 9255 4 gnd
rlabel metal1 s 0 10765 389 10796 4 gnd
rlabel metal1 s 1167 4605 1556 4636 4 gnd
rlabel metal1 s 1167 7685 1556 7716 4 gnd
rlabel metal1 s 1167 10765 1556 10796 4 gnd
rlabel metal1 s 0 1525 389 1556 4 gnd
rlabel metal1 s 1167 4604 1556 4635 4 gnd
rlabel metal1 s 1167 -16 1556 15 4 gnd
rlabel metal1 s 1167 3065 1556 3096 4 gnd
rlabel metal1 s 778 7684 1167 7715 4 gnd
rlabel metal1 s 1167 6145 1556 6176 4 gnd
rlabel metal1 s 1167 3064 1556 3095 4 gnd
rlabel metal1 s 389 3065 778 3096 4 gnd
rlabel metal1 s 778 9225 1167 9256 4 gnd
<< properties >>
string FIXED_BBOX 0 0 3112 24640
string GDS_FILE sram_0rw2r1w_4_16_sky130A.gds
string GDS_END 159408
string GDS_START 121460
<< end >>
