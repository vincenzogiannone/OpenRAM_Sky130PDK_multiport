magic
tech sky130A
magscale 1 2
timestamp 1643678851
<< checkpaint >>
rect -1326 -1302 13144 7182
<< locali >>
rect 3833 4734 4035 4768
rect 4001 4550 4035 4734
rect 3807 2207 3983 2241
rect 3807 2154 3841 2207
rect 3682 2120 3841 2154
<< viali >>
rect 3550 5472 3584 5506
rect 5478 5476 5512 5510
rect 6685 4543 6719 4577
rect 3598 4463 3632 4497
rect 3598 3883 3632 3917
rect 5125 3802 5159 3836
rect 3698 3635 3732 3669
rect 3698 3035 3732 3069
rect 4585 2870 4619 2904
rect 3598 2787 3632 2821
rect 3550 2120 3584 2154
rect 4936 2124 4970 2158
rect 4049 1959 4083 1993
rect 3550 1198 3584 1232
rect 9420 1190 9454 1224
<< metal1 >>
rect 3538 5506 3596 5512
rect 5466 5508 5469 5516
rect 3538 5503 3550 5506
rect 2982 5475 3550 5503
rect 3538 5472 3550 5475
rect 3584 5472 3596 5506
rect 5440 5478 5469 5508
rect 3538 5466 3596 5472
rect 5466 5470 5469 5478
rect 5521 5508 5524 5516
rect 5521 5478 5551 5508
rect 5521 5470 5524 5478
rect 6673 4575 6676 4583
rect 6647 4545 6676 4575
rect 6673 4537 6676 4545
rect 6728 4575 6731 4583
rect 6728 4545 6758 4575
rect 6728 4537 6731 4545
rect 3586 4497 3644 4503
rect 3586 4494 3598 4497
rect 3050 4466 3598 4494
rect 3586 4463 3598 4466
rect 3632 4463 3644 4497
rect 3586 4457 3644 4463
rect 3586 3917 3644 3923
rect 3586 3914 3598 3917
rect 3118 3886 3598 3914
rect 3586 3883 3598 3886
rect 3632 3883 3644 3917
rect 3586 3877 3644 3883
rect 5113 3834 5116 3842
rect 5087 3804 5116 3834
rect 5113 3796 5116 3804
rect 5168 3834 5171 3842
rect 5168 3804 5198 3834
rect 5168 3796 5171 3804
rect 3686 3669 3744 3675
rect 3686 3666 3698 3669
rect 2982 3638 3698 3666
rect 3686 3635 3698 3638
rect 3732 3635 3744 3669
rect 3686 3629 3744 3635
rect 40 3280 3202 3308
rect 3686 3069 3744 3075
rect 3686 3066 3698 3069
rect 3322 3038 3698 3066
rect 3686 3035 3698 3038
rect 3732 3035 3744 3069
rect 3686 3029 3744 3035
rect 4573 2902 4576 2910
rect 4547 2872 4576 2902
rect 4573 2864 4576 2872
rect 4628 2902 4631 2910
rect 4628 2872 4658 2902
rect 4628 2864 4631 2872
rect 3586 2821 3644 2827
rect 3586 2818 3598 2821
rect 3254 2790 3598 2818
rect 3586 2787 3598 2790
rect 3632 2787 3644 2821
rect 3586 2781 3644 2787
rect 3538 2154 3596 2160
rect 4924 2156 4927 2164
rect 3538 2151 3550 2154
rect 3254 2123 3550 2151
rect 3538 2120 3550 2123
rect 3584 2120 3596 2154
rect 4898 2126 4927 2156
rect 3538 2114 3596 2120
rect 4924 2118 4927 2126
rect 4979 2156 4982 2164
rect 4979 2126 5009 2156
rect 4979 2118 4982 2126
rect 4037 1991 4040 1999
rect 4011 1961 4040 1991
rect 4037 1953 4040 1961
rect 4092 1991 4095 1999
rect 4092 1961 4122 1991
rect 4092 1953 4095 1961
rect 3538 1230 3541 1238
rect 3512 1200 3541 1230
rect 3538 1192 3541 1200
rect 3593 1230 3596 1238
rect 3593 1200 3623 1230
rect 9408 1222 9411 1230
rect 3593 1192 3596 1200
rect 9382 1192 9411 1222
rect 9408 1184 9411 1192
rect 9463 1222 9466 1230
rect 9463 1192 9493 1222
rect 9463 1184 9466 1192
<< via1 >>
rect 2930 5463 2982 5515
rect 5469 5510 5521 5519
rect 5469 5476 5478 5510
rect 5478 5476 5512 5510
rect 5512 5476 5521 5510
rect 5469 5467 5521 5476
rect 6676 4577 6728 4586
rect 6676 4543 6685 4577
rect 6685 4543 6719 4577
rect 6719 4543 6728 4577
rect 6676 4534 6728 4543
rect 2998 4454 3050 4506
rect 3066 3874 3118 3926
rect 5116 3836 5168 3845
rect 5116 3802 5125 3836
rect 5125 3802 5159 3836
rect 5159 3802 5168 3836
rect 5116 3793 5168 3802
rect 2930 3626 2982 3678
rect -12 3268 40 3320
rect 3202 3268 3254 3320
rect 3270 3026 3322 3078
rect 4576 2904 4628 2913
rect 4576 2870 4585 2904
rect 4585 2870 4619 2904
rect 4619 2870 4628 2904
rect 4576 2861 4628 2870
rect 3202 2778 3254 2830
rect 3202 2111 3254 2163
rect 4927 2158 4979 2167
rect 4927 2124 4936 2158
rect 4936 2124 4970 2158
rect 4970 2124 4979 2158
rect 4927 2115 4979 2124
rect 4040 1993 4092 2002
rect 4040 1959 4049 1993
rect 4049 1959 4083 1993
rect 4083 1959 4092 1993
rect 4040 1950 4092 1959
rect 3541 1232 3593 1241
rect 3541 1198 3550 1232
rect 3550 1198 3584 1232
rect 3584 1198 3593 1232
rect 9411 1224 9463 1233
rect 3541 1189 3593 1198
rect 9411 1190 9420 1224
rect 9420 1190 9454 1224
rect 9454 1190 9463 1224
rect 9411 1181 9463 1190
<< metal2 >>
rect 2942 5515 2970 5922
rect 2942 3678 2970 5463
rect 3010 4506 3038 5922
rect 0 1676 28 3268
rect 2942 1834 2970 3626
rect 3010 2915 3038 4454
rect 3078 3926 3106 5922
rect 180 1416 234 1444
rect 180 232 234 260
rect 2942 0 2970 1778
rect 3010 0 3038 2859
rect 3078 541 3106 3874
rect 3078 0 3106 485
rect 3146 269 3174 5922
rect 3214 3320 3242 5922
rect 3214 2830 3242 3268
rect 3282 3078 3310 5922
rect 3214 2163 3242 2778
rect 3214 900 3242 2111
rect 3282 2004 3310 3026
rect 3282 1191 3310 1948
rect 3350 1463 3378 5922
rect 5521 5479 11884 5507
rect 6728 4546 11884 4574
rect 5168 3805 11884 3833
rect 4582 2915 4622 2921
rect 4582 2853 4622 2859
rect 4046 2004 4086 2010
rect 4046 1942 4086 1948
rect 4939 1834 4967 2115
rect 3146 0 3174 213
rect 3214 0 3242 844
rect 3282 0 3310 1135
rect 3350 0 3378 1407
rect 9463 1193 11884 1221
rect 9423 900 9451 1181
<< via2 >>
rect 2996 2859 3052 2915
rect 2928 1778 2984 1834
rect 2615 1407 2671 1463
rect 2150 1135 2206 1191
rect 2150 485 2206 541
rect 2615 213 2671 269
rect 3064 485 3120 541
rect 3268 1948 3324 2004
rect 4574 2913 4630 2915
rect 4574 2861 4576 2913
rect 4576 2861 4628 2913
rect 4628 2861 4630 2913
rect 4574 2859 4630 2861
rect 4038 2002 4094 2004
rect 4038 1950 4040 2002
rect 4040 1950 4092 2002
rect 4092 1950 4094 2002
rect 4038 1948 4094 1950
rect 4925 1778 4981 1834
rect 3336 1407 3392 1463
rect 3268 1135 3324 1191
rect 3200 844 3256 900
rect 3132 213 3188 269
rect 9409 844 9465 900
<< metal3 >>
rect 2958 2917 3090 2920
rect 4536 2917 4668 2920
rect 2958 2915 4668 2917
rect 2958 2859 2996 2915
rect 3052 2859 4574 2915
rect 4630 2859 4668 2915
rect 2958 2857 4668 2859
rect 2958 2854 3090 2857
rect 4536 2854 4668 2857
rect 3230 2006 3362 2009
rect 4000 2006 4132 2009
rect 3230 2004 4132 2006
rect 3230 1948 3268 2004
rect 3324 1948 4038 2004
rect 4094 1948 4132 2004
rect 3230 1946 4132 1948
rect 3230 1943 3362 1946
rect 4000 1943 4132 1946
rect 2890 1836 3022 1839
rect 4887 1836 5019 1839
rect 2890 1834 5019 1836
rect 2890 1778 2928 1834
rect 2984 1778 4925 1834
rect 4981 1778 5019 1834
rect 2890 1776 5019 1778
rect 2890 1773 3022 1776
rect 4887 1773 5019 1776
rect -66 1643 66 1709
rect 2577 1465 2709 1468
rect 3298 1465 3430 1468
rect 2577 1463 3430 1465
rect 2577 1407 2615 1463
rect 2671 1407 3336 1463
rect 3392 1407 3430 1463
rect 2577 1405 3430 1407
rect 2577 1402 2709 1405
rect 3298 1402 3430 1405
rect 2112 1193 2244 1196
rect 3230 1193 3362 1196
rect 2112 1191 3362 1193
rect 2112 1135 2150 1191
rect 2206 1135 3268 1191
rect 3324 1135 3362 1191
rect 2112 1133 3362 1135
rect 2112 1130 2244 1133
rect 3230 1130 3362 1133
rect 3162 902 3294 905
rect 9371 902 9503 905
rect 3162 900 9503 902
rect -66 805 66 871
rect 3162 844 3200 900
rect 3256 844 9409 900
rect 9465 844 9503 900
rect 3162 842 9503 844
rect 3162 839 3294 842
rect 9371 839 9503 842
rect 2112 543 2244 546
rect 3026 543 3158 546
rect 2112 541 3158 543
rect 2112 485 2150 541
rect 2206 485 3064 541
rect 3120 485 3158 541
rect 2112 483 3158 485
rect 2112 480 2244 483
rect 3026 480 3158 483
rect 2577 271 2709 274
rect 3094 271 3226 274
rect 2577 269 3226 271
rect 2577 213 2615 269
rect 2671 213 3132 269
rect 3188 213 3226 269
rect 2577 211 3226 213
rect 2577 208 2709 211
rect 3094 208 3226 211
rect -66 -33 66 33
use contact_17  contact_17_0
timestamp 1643678851
transform 1 0 4587 0 1 2872
box 0 0 1 1
use contact_13  contact_13_0
timestamp 1643678851
transform 1 0 4573 0 1 2864
box 0 0 1 1
use contact_18  contact_18_0
timestamp 1643678851
transform 1 0 4536 0 1 2854
box 0 0 1 1
use contact_17  contact_17_1
timestamp 1643678851
transform 1 0 4587 0 1 2872
box 0 0 1 1
use contact_13  contact_13_1
timestamp 1643678851
transform 1 0 4573 0 1 2864
box 0 0 1 1
use contact_29  contact_29_0
timestamp 1643678851
transform 1 0 2958 0 1 2854
box 0 0 1 1
use contact_13  contact_13_2
timestamp 1643678851
transform 1 0 3686 0 1 3029
box 0 0 1 1
use contact_17  contact_17_2
timestamp 1643678851
transform 1 0 3281 0 1 3037
box 0 0 1 1
use contact_13  contact_13_3
timestamp 1643678851
transform 1 0 3586 0 1 2781
box 0 0 1 1
use contact_17  contact_17_3
timestamp 1643678851
transform 1 0 3213 0 1 2789
box 0 0 1 1
use contact_17  contact_17_4
timestamp 1643678851
transform 1 0 4938 0 1 2126
box 0 0 1 1
use contact_13  contact_13_4
timestamp 1643678851
transform 1 0 4924 0 1 2118
box 0 0 1 1
use contact_29  contact_29_1
timestamp 1643678851
transform 1 0 2890 0 1 1773
box 0 0 1 1
use contact_29  contact_29_2
timestamp 1643678851
transform 1 0 4887 0 1 1773
box 0 0 1 1
use contact_18  contact_18_1
timestamp 1643678851
transform 1 0 4000 0 1 1943
box 0 0 1 1
use contact_17  contact_17_5
timestamp 1643678851
transform 1 0 4051 0 1 1961
box 0 0 1 1
use contact_13  contact_13_5
timestamp 1643678851
transform 1 0 4037 0 1 1953
box 0 0 1 1
use contact_18  contact_18_2
timestamp 1643678851
transform 1 0 4000 0 1 1943
box 0 0 1 1
use contact_17  contact_17_6
timestamp 1643678851
transform 1 0 4051 0 1 1961
box 0 0 1 1
use contact_13  contact_13_6
timestamp 1643678851
transform 1 0 4037 0 1 1953
box 0 0 1 1
use contact_29  contact_29_3
timestamp 1643678851
transform 1 0 3230 0 1 1943
box 0 0 1 1
use contact_13  contact_13_7
timestamp 1643678851
transform 1 0 3538 0 1 2114
box 0 0 1 1
use contact_17  contact_17_7
timestamp 1643678851
transform 1 0 3213 0 1 2122
box 0 0 1 1
use contact_17  contact_17_8
timestamp 1643678851
transform 1 0 9422 0 1 1192
box 0 0 1 1
use contact_13  contact_13_8
timestamp 1643678851
transform 1 0 9408 0 1 1184
box 0 0 1 1
use contact_17  contact_17_9
timestamp 1643678851
transform 1 0 9422 0 1 1192
box 0 0 1 1
use contact_13  contact_13_9
timestamp 1643678851
transform 1 0 9408 0 1 1184
box 0 0 1 1
use contact_29  contact_29_4
timestamp 1643678851
transform 1 0 3162 0 1 839
box 0 0 1 1
use contact_29  contact_29_5
timestamp 1643678851
transform 1 0 9371 0 1 839
box 0 0 1 1
use contact_17  contact_17_10
timestamp 1643678851
transform 1 0 3552 0 1 1200
box 0 0 1 1
use contact_13  contact_13_10
timestamp 1643678851
transform 1 0 3538 0 1 1192
box 0 0 1 1
use contact_17  contact_17_11
timestamp 1643678851
transform 1 0 6687 0 1 4545
box 0 0 1 1
use contact_13  contact_13_11
timestamp 1643678851
transform 1 0 6673 0 1 4537
box 0 0 1 1
use contact_13  contact_13_12
timestamp 1643678851
transform 1 0 3586 0 1 4457
box 0 0 1 1
use contact_17  contact_17_12
timestamp 1643678851
transform 1 0 3009 0 1 4465
box 0 0 1 1
use contact_17  contact_17_13
timestamp 1643678851
transform 1 0 5127 0 1 3804
box 0 0 1 1
use contact_13  contact_13_13
timestamp 1643678851
transform 1 0 5113 0 1 3796
box 0 0 1 1
use contact_13  contact_13_14
timestamp 1643678851
transform 1 0 3686 0 1 3629
box 0 0 1 1
use contact_17  contact_17_14
timestamp 1643678851
transform 1 0 2941 0 1 3637
box 0 0 1 1
use contact_13  contact_13_15
timestamp 1643678851
transform 1 0 3586 0 1 3877
box 0 0 1 1
use contact_17  contact_17_15
timestamp 1643678851
transform 1 0 3077 0 1 3885
box 0 0 1 1
use contact_17  contact_17_16
timestamp 1643678851
transform 1 0 5480 0 1 5478
box 0 0 1 1
use contact_13  contact_13_16
timestamp 1643678851
transform 1 0 5466 0 1 5470
box 0 0 1 1
use contact_13  contact_13_17
timestamp 1643678851
transform 1 0 3538 0 1 5466
box 0 0 1 1
use contact_17  contact_17_17
timestamp 1643678851
transform 1 0 2941 0 1 5474
box 0 0 1 1
use contact_17  contact_17_18
timestamp 1643678851
transform 1 0 3213 0 1 3279
box 0 0 1 1
use contact_17  contact_17_19
timestamp 1643678851
transform 1 0 -1 0 1 3279
box 0 0 1 1
use contact_18  contact_18_3
timestamp 1643678851
transform 1 0 2577 0 1 1402
box 0 0 1 1
use contact_29  contact_29_6
timestamp 1643678851
transform 1 0 3298 0 1 1402
box 0 0 1 1
use contact_18  contact_18_4
timestamp 1643678851
transform 1 0 2112 0 1 1130
box 0 0 1 1
use contact_29  contact_29_7
timestamp 1643678851
transform 1 0 3230 0 1 1130
box 0 0 1 1
use contact_18  contact_18_5
timestamp 1643678851
transform 1 0 2577 0 1 208
box 0 0 1 1
use contact_29  contact_29_8
timestamp 1643678851
transform 1 0 3094 0 1 208
box 0 0 1 1
use contact_18  contact_18_6
timestamp 1643678851
transform 1 0 2112 0 1 480
box 0 0 1 1
use contact_29  contact_29_9
timestamp 1643678851
transform 1 0 3026 0 1 480
box 0 0 1 1
use pdriver_4  pdriver_4_0
timestamp 1643678851
transform 1 0 3937 0 1 4190
box -36 -17 3924 895
use pnand2_1  pnand2_1_0
timestamp 1643678851
transform 1 0 3486 0 1 4190
box -36 -17 487 895
use pand2_1  pand2_1_0
timestamp 1643678851
transform 1 0 3486 0 -1 4190
box -36 -17 2925 895
use pdriver_2  pdriver_2_0
timestamp 1643678851
transform 1 0 3486 0 -1 5866
box -36 -17 2736 895
use pand2_0  pand2_0_0
timestamp 1643678851
transform 1 0 3486 0 1 2514
box -36 -17 1845 895
use pand2_0  pand2_0_1
timestamp 1643678851
transform 1 0 3837 0 -1 2514
box -36 -17 1845 895
use pinv_1  pinv_1_0
timestamp 1643678851
transform 1 0 3486 0 -1 2514
box -36 -17 387 895
use pdriver_1  pdriver_1_0
timestamp 1643678851
transform 1 0 3486 0 1 838
box -36 -17 8298 895
use dff_buf_array  dff_buf_array_0
timestamp 1643678851
transform 1 0 0 0 1 0
box -66 -42 2978 1718
<< labels >>
rlabel metal2 s 180 1416 234 1444 4 csb
rlabel metal2 s 180 232 234 260 4 web
rlabel metal2 s 5495 5479 11884 5507 4 wl_en
rlabel metal2 s 5142 3805 11884 3833 4 w_en
rlabel metal2 s 6702 4546 11884 4574 4 p_en_bar
rlabel metal2 s 3553 1201 3581 1229 4 clk
rlabel metal2 s 9437 1193 11884 1221 4 clk_buf
rlabel metal3 s -66 1643 66 1709 4 gnd
rlabel metal3 s -66 -33 66 33 4 gnd
rlabel metal3 s -66 805 66 871 4 vdd
<< properties >>
string FIXED_BBOX 0 0 11884 116
string GDS_FILE sram_0rw2r1w_16_128_sky130A.gds
string GDS_END 2009958
string GDS_START 2001244
<< end >>
