magic
tech sky130A
magscale 1 2
timestamp 1643671299
<< checkpaint >>
rect -1271 -1302 7156 25926
<< metal1 >>
rect 4799 23998 5212 24026
rect 4799 23906 4827 23998
rect 5838 23928 5866 23956
rect 4708 23878 4910 23906
rect 4708 23760 4736 23878
rect 4655 23732 4736 23760
rect 4655 23644 4683 23732
rect 4708 23644 4736 23732
rect 4799 23644 4827 23878
rect 5838 23802 5866 23830
rect 4634 23616 4827 23644
rect 4655 23522 4683 23616
rect 4634 23494 4683 23522
rect 4708 23376 4736 23616
rect 5838 23576 5866 23604
rect 4634 23348 4736 23376
rect 5838 22536 5866 22564
rect 4655 22380 4732 22408
rect 4655 22072 4683 22380
rect 5838 22310 5866 22338
rect 4708 22234 4910 22262
rect 4708 22072 4736 22234
rect 5838 22184 5866 22212
rect 4634 22044 4736 22072
rect 4799 22114 5212 22142
rect 4655 21926 4683 22044
rect 4634 21898 4683 21926
rect 4799 21804 4827 22114
rect 4634 21776 4827 21804
rect 4799 20922 5212 20950
rect 4799 20830 4827 20922
rect 5838 20852 5866 20880
rect 4708 20802 4910 20830
rect 4708 20684 4736 20802
rect 4655 20656 4736 20684
rect 4655 20616 4683 20656
rect 4708 20616 4736 20656
rect 4799 20616 4827 20802
rect 5838 20726 5866 20754
rect 4634 20588 4827 20616
rect 4655 20494 4683 20588
rect 4634 20466 4683 20494
rect 4708 20348 4736 20588
rect 5838 20500 5866 20528
rect 4634 20320 4736 20348
rect 5838 19460 5866 19488
rect 4655 19304 4732 19332
rect 4655 19044 4683 19304
rect 5838 19234 5866 19262
rect 4708 19158 4910 19186
rect 4708 19044 4736 19158
rect 5838 19108 5866 19136
rect 4634 19016 4736 19044
rect 4799 19038 5212 19066
rect 4655 18898 4683 19016
rect 4634 18870 4683 18898
rect 4799 18776 4827 19038
rect 4634 18748 4827 18776
rect 4799 17846 5212 17874
rect 4799 17754 4827 17846
rect 5838 17776 5866 17804
rect 4708 17726 4910 17754
rect 4708 17608 4736 17726
rect 4655 17588 4736 17608
rect 4799 17588 4827 17726
rect 5838 17650 5866 17678
rect 4634 17560 4827 17588
rect 4655 17466 4683 17560
rect 4634 17438 4683 17466
rect 4708 17320 4736 17560
rect 5838 17424 5866 17452
rect 4634 17292 4736 17320
rect 5838 16384 5866 16412
rect 4655 16228 4732 16256
rect 4655 16016 4683 16228
rect 5838 16158 5866 16186
rect 4708 16082 4910 16110
rect 4708 16016 4736 16082
rect 5838 16032 5866 16060
rect 4634 15988 4736 16016
rect 4655 15870 4683 15988
rect 4634 15842 4683 15870
rect 4799 15962 5212 15990
rect 4799 15748 4827 15962
rect 4634 15720 4827 15748
rect 4799 14770 5212 14798
rect 4799 14678 4827 14770
rect 5838 14700 5866 14728
rect 4708 14650 4910 14678
rect 4708 14560 4736 14650
rect 4799 14560 4827 14650
rect 5838 14574 5866 14602
rect 4634 14532 4827 14560
rect 4655 14504 4736 14532
rect 4655 14438 4683 14504
rect 4634 14410 4683 14438
rect 4708 14292 4736 14504
rect 5838 14348 5866 14376
rect 4634 14264 4736 14292
rect 5838 13308 5866 13336
rect 4655 13152 4732 13180
rect 4655 12988 4683 13152
rect 5838 13082 5866 13110
rect 4708 13006 4910 13034
rect 4708 12988 4736 13006
rect 4634 12960 4736 12988
rect 4655 12842 4683 12960
rect 5838 12956 5866 12984
rect 4634 12814 4683 12842
rect 4799 12886 5212 12914
rect 4799 12720 4827 12886
rect 4634 12692 4827 12720
rect 4799 11694 5212 11722
rect 4799 11602 4827 11694
rect 5838 11624 5866 11652
rect 4708 11574 4910 11602
rect 4708 11532 4736 11574
rect 4799 11532 4827 11574
rect 4634 11504 4827 11532
rect 4708 11456 4736 11504
rect 5838 11498 5866 11526
rect 4655 11428 4736 11456
rect 4655 11410 4683 11428
rect 4634 11382 4683 11410
rect 4708 11264 4736 11428
rect 5838 11272 5866 11300
rect 4634 11236 4736 11264
rect 5838 10232 5866 10260
rect 4655 10076 4732 10104
rect 4655 9960 4683 10076
rect 5838 10006 5866 10034
rect 4634 9958 4736 9960
rect 4634 9932 4910 9958
rect 4655 9814 4683 9932
rect 4708 9930 4910 9932
rect 5838 9880 5866 9908
rect 4634 9786 4683 9814
rect 4799 9810 5212 9838
rect 4799 9692 4827 9810
rect 4634 9664 4827 9692
rect 4799 8618 5212 8646
rect 4799 8526 4827 8618
rect 5838 8548 5866 8576
rect 4708 8504 4910 8526
rect 4634 8498 4910 8504
rect 4634 8476 4827 8498
rect 4634 8380 4683 8382
rect 4708 8380 4736 8476
rect 5838 8422 5866 8450
rect 4634 8354 4736 8380
rect 4655 8352 4736 8354
rect 4708 8236 4736 8352
rect 4634 8208 4736 8236
rect 5838 8196 5866 8224
rect 5838 7156 5866 7184
rect 4655 7000 4732 7028
rect 4655 6932 4683 7000
rect 4634 6904 4736 6932
rect 5838 6930 5866 6958
rect 4655 6786 4683 6904
rect 4708 6882 4736 6904
rect 4708 6854 4910 6882
rect 5838 6804 5866 6832
rect 4634 6758 4683 6786
rect 4799 6734 5212 6762
rect 4799 6664 4827 6734
rect 4634 6636 4827 6664
rect 4799 5542 5212 5570
rect 4799 5476 4827 5542
rect 4634 5450 4827 5476
rect 5838 5472 5866 5500
rect 4634 5448 4910 5450
rect 4708 5422 4910 5448
rect 4634 5326 4683 5354
rect 4655 5304 4683 5326
rect 4708 5304 4736 5422
rect 5838 5346 5866 5374
rect 4655 5276 4736 5304
rect 4708 5208 4736 5276
rect 4634 5180 4736 5208
rect 5838 5120 5866 5148
rect 5838 4080 5866 4108
rect 4655 3924 4732 3952
rect 4655 3904 4683 3924
rect 4634 3876 4736 3904
rect 4655 3758 4683 3876
rect 4708 3806 4736 3876
rect 5838 3854 5866 3882
rect 4708 3778 4910 3806
rect 4634 3730 4683 3758
rect 5838 3728 5866 3756
rect 4799 3658 5212 3686
rect 4799 3636 4827 3658
rect 4634 3608 4827 3636
rect 4799 2466 5212 2494
rect 4799 2448 4827 2466
rect 4634 2420 4827 2448
rect 5838 2396 5866 2424
rect 4708 2346 4910 2374
rect 4634 2298 4683 2326
rect 4655 2228 4683 2298
rect 4708 2228 4736 2346
rect 5838 2270 5866 2298
rect 4655 2200 4736 2228
rect 4708 2180 4736 2200
rect 4634 2152 4736 2180
rect 5838 2044 5866 2072
rect 5838 1004 5866 1032
rect 4634 848 4736 876
rect 4655 730 4683 848
rect 4634 702 4683 730
rect 4708 730 4736 848
rect 5838 778 5866 806
rect 4708 702 4910 730
rect 5838 652 5866 680
rect 4799 608 5212 610
rect 4634 582 5212 608
rect 4634 580 4827 582
<< metal2 >>
rect 1 0 29 24632
rect 69 0 97 24632
rect 137 0 165 24632
rect 205 0 233 24632
rect 273 0 301 24632
rect 341 0 369 24632
rect 4476 24594 4690 24622
<< metal3 >>
rect 651 24602 711 24662
rect 1410 24602 1470 24662
rect 5836 24578 5896 24638
rect 4632 24194 4692 24254
rect 651 23062 711 23122
rect 1410 23062 1470 23122
rect 5836 23040 5896 23100
rect 4632 22680 4692 22740
rect 651 21522 711 21582
rect 1410 21522 1470 21582
rect 5836 21502 5896 21562
rect 4632 21166 4692 21226
rect 651 19982 711 20042
rect 1410 19982 1470 20042
rect 5836 19964 5896 20024
rect 4632 19652 4692 19712
rect 651 18442 711 18502
rect 1410 18442 1470 18502
rect 5836 18426 5896 18486
rect 4632 18138 4692 18198
rect 5836 16888 5896 16948
rect 4632 16624 4692 16684
rect 651 15366 711 15426
rect 1410 15366 1470 15426
rect 5836 15350 5896 15410
rect 4632 15110 4692 15170
rect 651 13826 711 13886
rect 1410 13826 1470 13886
rect 5836 13812 5896 13872
rect 4632 13596 4692 13656
rect 651 12286 711 12346
rect 1410 12286 1470 12346
rect 5836 12274 5896 12334
rect 4632 12082 4692 12142
rect 651 10746 711 10806
rect 1410 10746 1470 10806
rect 5836 10736 5896 10796
rect 4632 10568 4692 10628
rect 651 9206 711 9266
rect 1410 9206 1470 9266
rect 5836 9198 5896 9258
rect 4632 9054 4692 9114
rect 5836 7660 5896 7720
rect 4632 7540 4692 7600
rect 651 6130 711 6190
rect 1410 6130 1470 6190
rect 5836 6122 5896 6182
rect 4632 6026 4692 6086
rect 651 4590 711 4650
rect 1410 4590 1470 4650
rect 5836 4584 5896 4644
rect 4632 4512 4692 4572
rect 651 3050 711 3110
rect 1410 3050 1470 3110
rect 4632 2998 4692 3058
rect 5836 3046 5896 3106
rect 651 1510 711 1570
rect 1410 1510 1470 1570
rect 4632 1484 4692 1544
rect 5836 1508 5896 1568
rect 651 -30 711 30
rect 1410 -30 1470 30
rect 4632 -30 4692 30
rect 5836 -30 5896 30
use wordline_driver_array  wordline_driver_array_0
timestamp 1643671299
transform 1 0 4662 0 1 0
box 0 -42 1234 24650
use hierarchical_decoder  hierarchical_decoder_0
timestamp 1643671299
transform 1 0 0 0 1 0
box -11 -42 4692 24666
<< labels >>
rlabel metal2 s 1 0 29 24632 4 addr0
rlabel metal2 s 69 0 97 24632 4 addr1
rlabel metal2 s 137 0 165 24632 4 addr2
rlabel metal2 s 205 0 233 24632 4 addr3
rlabel metal2 s 273 0 301 24632 4 addr4
rlabel metal2 s 341 0 369 24632 4 addr5
rlabel metal1 s 5838 778 5866 806 4 rwl0_0
rlabel metal1 s 5838 1004 5866 1032 4 rwl1_0
rlabel metal1 s 5838 652 5866 680 4 wwl0_0
rlabel metal1 s 5838 2270 5866 2298 4 rwl0_1
rlabel metal1 s 5838 2044 5866 2072 4 rwl1_1
rlabel metal1 s 5838 2396 5866 2424 4 wwl0_1
rlabel metal1 s 5838 3854 5866 3882 4 rwl0_2
rlabel metal1 s 5838 4080 5866 4108 4 rwl1_2
rlabel metal1 s 5838 3728 5866 3756 4 wwl0_2
rlabel metal1 s 5838 5346 5866 5374 4 rwl0_3
rlabel metal1 s 5838 5120 5866 5148 4 rwl1_3
rlabel metal1 s 5838 5472 5866 5500 4 wwl0_3
rlabel metal1 s 5838 6930 5866 6958 4 rwl0_4
rlabel metal1 s 5838 7156 5866 7184 4 rwl1_4
rlabel metal1 s 5838 6804 5866 6832 4 wwl0_4
rlabel metal1 s 5838 8422 5866 8450 4 rwl0_5
rlabel metal1 s 5838 8196 5866 8224 4 rwl1_5
rlabel metal1 s 5838 8548 5866 8576 4 wwl0_5
rlabel metal1 s 5838 10006 5866 10034 4 rwl0_6
rlabel metal1 s 5838 10232 5866 10260 4 rwl1_6
rlabel metal1 s 5838 9880 5866 9908 4 wwl0_6
rlabel metal1 s 5838 11498 5866 11526 4 rwl0_7
rlabel metal1 s 5838 11272 5866 11300 4 rwl1_7
rlabel metal1 s 5838 11624 5866 11652 4 wwl0_7
rlabel metal1 s 5838 13082 5866 13110 4 rwl0_8
rlabel metal1 s 5838 13308 5866 13336 4 rwl1_8
rlabel metal1 s 5838 12956 5866 12984 4 wwl0_8
rlabel metal1 s 5838 14574 5866 14602 4 rwl0_9
rlabel metal1 s 5838 14348 5866 14376 4 rwl1_9
rlabel metal1 s 5838 14700 5866 14728 4 wwl0_9
rlabel metal1 s 5838 16158 5866 16186 4 rwl0_10
rlabel metal1 s 5838 16384 5866 16412 4 rwl1_10
rlabel metal1 s 5838 16032 5866 16060 4 wwl0_10
rlabel metal1 s 5838 17650 5866 17678 4 rwl0_11
rlabel metal1 s 5838 17424 5866 17452 4 rwl1_11
rlabel metal1 s 5838 17776 5866 17804 4 wwl0_11
rlabel metal1 s 5838 19234 5866 19262 4 rwl0_12
rlabel metal1 s 5838 19460 5866 19488 4 rwl1_12
rlabel metal1 s 5838 19108 5866 19136 4 wwl0_12
rlabel metal1 s 5838 20726 5866 20754 4 rwl0_13
rlabel metal1 s 5838 20500 5866 20528 4 rwl1_13
rlabel metal1 s 5838 20852 5866 20880 4 wwl0_13
rlabel metal1 s 5838 22310 5866 22338 4 rwl0_14
rlabel metal1 s 5838 22536 5866 22564 4 rwl1_14
rlabel metal1 s 5838 22184 5866 22212 4 wwl0_14
rlabel metal1 s 5838 23802 5866 23830 4 rwl0_15
rlabel metal1 s 5838 23576 5866 23604 4 rwl1_15
rlabel metal1 s 5838 23928 5866 23956 4 wwl0_15
rlabel metal2 s 4662 24594 4690 24622 4 wl_en
rlabel metal3 s 651 13826 711 13886 4 vdd
rlabel metal3 s 4632 22680 4692 22740 4 vdd
rlabel metal3 s 5836 4584 5896 4644 4 vdd
rlabel metal3 s 1410 10746 1470 10806 4 vdd
rlabel metal3 s 5836 19964 5896 20024 4 vdd
rlabel metal3 s 1410 23062 1470 23122 4 vdd
rlabel metal3 s 5836 10736 5896 10796 4 vdd
rlabel metal3 s 4632 1484 4692 1544 4 vdd
rlabel metal3 s 4632 19652 4692 19712 4 vdd
rlabel metal3 s 651 23062 711 23122 4 vdd
rlabel metal3 s 651 4590 711 4650 4 vdd
rlabel metal3 s 4632 4512 4692 4572 4 vdd
rlabel metal3 s 5836 16888 5896 16948 4 vdd
rlabel metal3 s 4632 7540 4692 7600 4 vdd
rlabel metal3 s 1410 13826 1470 13886 4 vdd
rlabel metal3 s 4632 16624 4692 16684 4 vdd
rlabel metal3 s 4632 13596 4692 13656 4 vdd
rlabel metal3 s 651 10746 711 10806 4 vdd
rlabel metal3 s 5836 23040 5896 23100 4 vdd
rlabel metal3 s 1410 4590 1470 4650 4 vdd
rlabel metal3 s 1410 19982 1470 20042 4 vdd
rlabel metal3 s 4632 10568 4692 10628 4 vdd
rlabel metal3 s 1410 1510 1470 1570 4 vdd
rlabel metal3 s 651 1510 711 1570 4 vdd
rlabel metal3 s 5836 7660 5896 7720 4 vdd
rlabel metal3 s 5836 1508 5896 1568 4 vdd
rlabel metal3 s 5836 13812 5896 13872 4 vdd
rlabel metal3 s 651 19982 711 20042 4 vdd
rlabel metal3 s 1410 18442 1470 18502 4 gnd
rlabel metal3 s 4632 2998 4692 3058 4 gnd
rlabel metal3 s 4632 21166 4692 21226 4 gnd
rlabel metal3 s 1410 9206 1470 9266 4 gnd
rlabel metal3 s 4632 15110 4692 15170 4 gnd
rlabel metal3 s 1410 12286 1470 12346 4 gnd
rlabel metal3 s 651 -30 711 30 4 gnd
rlabel metal3 s 5836 9198 5896 9258 4 gnd
rlabel metal3 s 5836 -30 5896 30 4 gnd
rlabel metal3 s 1410 21522 1470 21582 4 gnd
rlabel metal3 s 651 3050 711 3110 4 gnd
rlabel metal3 s 4632 18138 4692 18198 4 gnd
rlabel metal3 s 4632 12082 4692 12142 4 gnd
rlabel metal3 s 651 15366 711 15426 4 gnd
rlabel metal3 s 1410 -30 1470 30 4 gnd
rlabel metal3 s 4632 24194 4692 24254 4 gnd
rlabel metal3 s 651 6130 711 6190 4 gnd
rlabel metal3 s 4632 6026 4692 6086 4 gnd
rlabel metal3 s 1410 15366 1470 15426 4 gnd
rlabel metal3 s 1410 3050 1470 3110 4 gnd
rlabel metal3 s 1410 6130 1470 6190 4 gnd
rlabel metal3 s 5836 12274 5896 12334 4 gnd
rlabel metal3 s 5836 24578 5896 24638 4 gnd
rlabel metal3 s 1410 24602 1470 24662 4 gnd
rlabel metal3 s 5836 21502 5896 21562 4 gnd
rlabel metal3 s 651 21522 711 21582 4 gnd
rlabel metal3 s 4632 -30 4692 30 4 gnd
rlabel metal3 s 651 9206 711 9266 4 gnd
rlabel metal3 s 651 18442 711 18502 4 gnd
rlabel metal3 s 5836 3046 5896 3106 4 gnd
rlabel metal3 s 5836 18426 5896 18486 4 gnd
rlabel metal3 s 651 24602 711 24662 4 gnd
rlabel metal3 s 5836 15350 5896 15410 4 gnd
rlabel metal3 s 5836 6122 5896 6182 4 gnd
rlabel metal3 s 4632 9054 4692 9114 4 gnd
rlabel metal3 s 651 12286 711 12346 4 gnd
<< properties >>
string FIXED_BBOX 0 0 5902 24660
string GDS_FILE sram_0rw2r1w_16_32_sky130A.gds
string GDS_END 935618
string GDS_START 891536
<< end >>
