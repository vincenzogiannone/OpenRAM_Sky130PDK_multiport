magic
tech sky130A
magscale 1 2
timestamp 1643671299
<< checkpaint >>
rect -1260 -1260 1261 1261
<< properties >>
string GDS_FILE sram_0rw2r1w_16_32_sky130A.gds
string GDS_END 819958
string GDS_START 819634
<< end >>
