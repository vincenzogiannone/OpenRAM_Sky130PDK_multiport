magic
tech sky130A
magscale 1 2
timestamp 1643671299
<< checkpaint >>
rect -1263 -1302 24972 2176
<< via1 >>
rect 715 812 767 864
rect 2197 812 2249 864
rect 3679 812 3731 864
rect 5161 812 5213 864
rect 6643 812 6695 864
rect 8125 812 8177 864
rect 9607 812 9659 864
rect 11089 812 11141 864
rect 12571 812 12623 864
rect 14053 812 14105 864
rect 15535 812 15587 864
rect 17017 812 17069 864
rect 18499 812 18551 864
rect 19981 812 20033 864
rect 21463 812 21515 864
rect 22945 812 22997 864
rect 715 -26 767 26
rect 2197 -26 2249 26
rect 3679 -26 3731 26
rect 5161 -26 5213 26
rect 6643 -26 6695 26
rect 8125 -26 8177 26
rect 9607 -26 9659 26
rect 11089 -26 11141 26
rect 12571 -26 12623 26
rect 14053 -26 14105 26
rect 15535 -26 15587 26
rect 17017 -26 17069 26
rect 18499 -26 18551 26
rect 19981 -26 20033 26
rect 21463 -26 21515 26
rect 22945 -26 22997 26
<< metal2 >>
rect 721 866 761 872
rect 2203 866 2243 872
rect 3685 866 3725 872
rect 5167 866 5207 872
rect 6649 866 6689 872
rect 8131 866 8171 872
rect 9613 866 9653 872
rect 11095 866 11135 872
rect 12577 866 12617 872
rect 14059 866 14099 872
rect 15541 866 15581 872
rect 17023 866 17063 872
rect 18505 866 18545 872
rect 19987 866 20027 872
rect 21469 866 21509 872
rect 22951 866 22991 872
rect 0 328 28 838
rect 721 804 761 810
rect 1482 328 1510 838
rect 2203 804 2243 810
rect 2964 328 2992 838
rect 3685 804 3725 810
rect 4446 328 4474 838
rect 5167 804 5207 810
rect 5928 328 5956 838
rect 6649 804 6689 810
rect 7410 328 7438 838
rect 8131 804 8171 810
rect 8892 328 8920 838
rect 9613 804 9653 810
rect 10374 328 10402 838
rect 11095 804 11135 810
rect 11856 328 11884 838
rect 12577 804 12617 810
rect 13338 328 13366 838
rect 14059 804 14099 810
rect 14820 328 14848 838
rect 15541 804 15581 810
rect 16302 328 16330 838
rect 17023 804 17063 810
rect 17784 328 17812 838
rect 18505 804 18545 810
rect 19266 328 19294 838
rect 19987 804 20027 810
rect 20748 328 20776 838
rect 21469 804 21509 810
rect 22230 328 22258 838
rect 22951 804 22991 810
rect 0 0 28 272
rect 180 232 234 260
rect 1260 228 1314 256
rect 721 28 761 34
rect 1482 0 1510 272
rect 1662 232 1716 260
rect 2742 228 2796 256
rect 2203 28 2243 34
rect 2964 0 2992 272
rect 3144 232 3198 260
rect 4224 228 4278 256
rect 3685 28 3725 34
rect 4446 0 4474 272
rect 4626 232 4680 260
rect 5706 228 5760 256
rect 5167 28 5207 34
rect 5928 0 5956 272
rect 6108 232 6162 260
rect 7188 228 7242 256
rect 6649 28 6689 34
rect 7410 0 7438 272
rect 7590 232 7644 260
rect 8670 228 8724 256
rect 8131 28 8171 34
rect 8892 0 8920 272
rect 9072 232 9126 260
rect 10152 228 10206 256
rect 9613 28 9653 34
rect 10374 0 10402 272
rect 10554 232 10608 260
rect 11634 228 11688 256
rect 11095 28 11135 34
rect 11856 0 11884 272
rect 12036 232 12090 260
rect 13116 228 13170 256
rect 12577 28 12617 34
rect 13338 0 13366 272
rect 13518 232 13572 260
rect 14598 228 14652 256
rect 14059 28 14099 34
rect 14820 0 14848 272
rect 15000 232 15054 260
rect 16080 228 16134 256
rect 15541 28 15581 34
rect 16302 0 16330 272
rect 16482 232 16536 260
rect 17562 228 17616 256
rect 17023 28 17063 34
rect 17784 0 17812 272
rect 17964 232 18018 260
rect 19044 228 19098 256
rect 18505 28 18545 34
rect 19266 0 19294 272
rect 19446 232 19500 260
rect 20526 228 20580 256
rect 19987 28 20027 34
rect 20748 0 20776 272
rect 20928 232 20982 260
rect 22008 228 22062 256
rect 21469 28 21509 34
rect 22230 0 22258 272
rect 22410 232 22464 260
rect 23490 228 23544 256
rect 22951 28 22991 34
rect 721 -34 761 -28
rect 2203 -34 2243 -28
rect 3685 -34 3725 -28
rect 5167 -34 5207 -28
rect 6649 -34 6689 -28
rect 8131 -34 8171 -28
rect 9613 -34 9653 -28
rect 11095 -34 11135 -28
rect 12577 -34 12617 -28
rect 14059 -34 14099 -28
rect 15541 -34 15581 -28
rect 17023 -34 17063 -28
rect 18505 -34 18545 -28
rect 19987 -34 20027 -28
rect 21469 -34 21509 -28
rect 22951 -34 22991 -28
<< via2 >>
rect 713 864 769 866
rect 713 812 715 864
rect 715 812 767 864
rect 767 812 769 864
rect 2195 864 2251 866
rect 713 810 769 812
rect 2195 812 2197 864
rect 2197 812 2249 864
rect 2249 812 2251 864
rect 3677 864 3733 866
rect 2195 810 2251 812
rect 3677 812 3679 864
rect 3679 812 3731 864
rect 3731 812 3733 864
rect 5159 864 5215 866
rect 3677 810 3733 812
rect 5159 812 5161 864
rect 5161 812 5213 864
rect 5213 812 5215 864
rect 6641 864 6697 866
rect 5159 810 5215 812
rect 6641 812 6643 864
rect 6643 812 6695 864
rect 6695 812 6697 864
rect 8123 864 8179 866
rect 6641 810 6697 812
rect 8123 812 8125 864
rect 8125 812 8177 864
rect 8177 812 8179 864
rect 9605 864 9661 866
rect 8123 810 8179 812
rect 9605 812 9607 864
rect 9607 812 9659 864
rect 9659 812 9661 864
rect 11087 864 11143 866
rect 9605 810 9661 812
rect 11087 812 11089 864
rect 11089 812 11141 864
rect 11141 812 11143 864
rect 12569 864 12625 866
rect 11087 810 11143 812
rect 12569 812 12571 864
rect 12571 812 12623 864
rect 12623 812 12625 864
rect 14051 864 14107 866
rect 12569 810 12625 812
rect 14051 812 14053 864
rect 14053 812 14105 864
rect 14105 812 14107 864
rect 15533 864 15589 866
rect 14051 810 14107 812
rect 15533 812 15535 864
rect 15535 812 15587 864
rect 15587 812 15589 864
rect 17015 864 17071 866
rect 15533 810 15589 812
rect 17015 812 17017 864
rect 17017 812 17069 864
rect 17069 812 17071 864
rect 18497 864 18553 866
rect 17015 810 17071 812
rect 18497 812 18499 864
rect 18499 812 18551 864
rect 18551 812 18553 864
rect 19979 864 20035 866
rect 18497 810 18553 812
rect 19979 812 19981 864
rect 19981 812 20033 864
rect 20033 812 20035 864
rect 21461 864 21517 866
rect 19979 810 20035 812
rect 21461 812 21463 864
rect 21463 812 21515 864
rect 21515 812 21517 864
rect 22943 864 22999 866
rect 21461 810 21517 812
rect 22943 812 22945 864
rect 22945 812 22997 864
rect 22997 812 22999 864
rect 22943 810 22999 812
rect -1 272 55 328
rect 1481 272 1537 328
rect 2963 272 3019 328
rect 4445 272 4501 328
rect 5927 272 5983 328
rect 7409 272 7465 328
rect 8891 272 8947 328
rect 10373 272 10429 328
rect 11855 272 11911 328
rect 13337 272 13393 328
rect 14819 272 14875 328
rect 16301 272 16357 328
rect 17783 272 17839 328
rect 19265 272 19321 328
rect 20747 272 20803 328
rect 22229 272 22285 328
rect 713 26 769 28
rect 713 -26 715 26
rect 715 -26 767 26
rect 767 -26 769 26
rect 2195 26 2251 28
rect 713 -28 769 -26
rect 2195 -26 2197 26
rect 2197 -26 2249 26
rect 2249 -26 2251 26
rect 3677 26 3733 28
rect 2195 -28 2251 -26
rect 3677 -26 3679 26
rect 3679 -26 3731 26
rect 3731 -26 3733 26
rect 5159 26 5215 28
rect 3677 -28 3733 -26
rect 5159 -26 5161 26
rect 5161 -26 5213 26
rect 5213 -26 5215 26
rect 6641 26 6697 28
rect 5159 -28 5215 -26
rect 6641 -26 6643 26
rect 6643 -26 6695 26
rect 6695 -26 6697 26
rect 8123 26 8179 28
rect 6641 -28 6697 -26
rect 8123 -26 8125 26
rect 8125 -26 8177 26
rect 8177 -26 8179 26
rect 9605 26 9661 28
rect 8123 -28 8179 -26
rect 9605 -26 9607 26
rect 9607 -26 9659 26
rect 9659 -26 9661 26
rect 11087 26 11143 28
rect 9605 -28 9661 -26
rect 11087 -26 11089 26
rect 11089 -26 11141 26
rect 11141 -26 11143 26
rect 12569 26 12625 28
rect 11087 -28 11143 -26
rect 12569 -26 12571 26
rect 12571 -26 12623 26
rect 12623 -26 12625 26
rect 14051 26 14107 28
rect 12569 -28 12625 -26
rect 14051 -26 14053 26
rect 14053 -26 14105 26
rect 14105 -26 14107 26
rect 15533 26 15589 28
rect 14051 -28 14107 -26
rect 15533 -26 15535 26
rect 15535 -26 15587 26
rect 15587 -26 15589 26
rect 17015 26 17071 28
rect 15533 -28 15589 -26
rect 17015 -26 17017 26
rect 17017 -26 17069 26
rect 17069 -26 17071 26
rect 18497 26 18553 28
rect 17015 -28 17071 -26
rect 18497 -26 18499 26
rect 18499 -26 18551 26
rect 18551 -26 18553 26
rect 19979 26 20035 28
rect 18497 -28 18553 -26
rect 19979 -26 19981 26
rect 19981 -26 20033 26
rect 20033 -26 20035 26
rect 21461 26 21517 28
rect 19979 -28 20035 -26
rect 21461 -26 21463 26
rect 21463 -26 21515 26
rect 21515 -26 21517 26
rect 22943 26 22999 28
rect 21461 -28 21517 -26
rect 22943 -26 22945 26
rect 22945 -26 22997 26
rect 22997 -26 22999 26
rect 22943 -28 22999 -26
<< metal3 >>
rect 711 866 771 868
rect 711 810 713 866
rect 769 810 771 866
rect 711 808 771 810
rect 2193 866 2253 868
rect 2193 810 2195 866
rect 2251 810 2253 866
rect 2193 808 2253 810
rect 3675 866 3735 868
rect 3675 810 3677 866
rect 3733 810 3735 866
rect 3675 808 3735 810
rect 5157 866 5217 868
rect 5157 810 5159 866
rect 5215 810 5217 866
rect 5157 808 5217 810
rect 6639 866 6699 868
rect 6639 810 6641 866
rect 6697 810 6699 866
rect 6639 808 6699 810
rect 8121 866 8181 868
rect 8121 810 8123 866
rect 8179 810 8181 866
rect 8121 808 8181 810
rect 9603 866 9663 868
rect 9603 810 9605 866
rect 9661 810 9663 866
rect 9603 808 9663 810
rect 11085 866 11145 868
rect 11085 810 11087 866
rect 11143 810 11145 866
rect 11085 808 11145 810
rect 12567 866 12627 868
rect 12567 810 12569 866
rect 12625 810 12627 866
rect 12567 808 12627 810
rect 14049 866 14109 868
rect 14049 810 14051 866
rect 14107 810 14109 866
rect 14049 808 14109 810
rect 15531 866 15591 868
rect 15531 810 15533 866
rect 15589 810 15591 866
rect 15531 808 15591 810
rect 17013 866 17073 868
rect 17013 810 17015 866
rect 17071 810 17073 866
rect 17013 808 17073 810
rect 18495 866 18555 868
rect 18495 810 18497 866
rect 18553 810 18555 866
rect 18495 808 18555 810
rect 19977 866 20037 868
rect 19977 810 19979 866
rect 20035 810 20037 866
rect 19977 808 20037 810
rect 21459 866 21519 868
rect 21459 810 21461 866
rect 21517 810 21519 866
rect 21459 808 21519 810
rect 22941 866 23001 868
rect 22941 810 22943 866
rect 22999 810 23001 866
rect 22941 808 23001 810
rect -3 328 23712 330
rect -3 272 -1 328
rect 55 272 1481 328
rect 1537 272 2963 328
rect 3019 272 4445 328
rect 4501 272 5927 328
rect 5983 272 7409 328
rect 7465 272 8891 328
rect 8947 272 10373 328
rect 10429 272 11855 328
rect 11911 272 13337 328
rect 13393 272 14819 328
rect 14875 272 16301 328
rect 16357 272 17783 328
rect 17839 272 19265 328
rect 19321 272 20747 328
rect 20803 272 22229 328
rect 22285 272 23712 328
rect -3 270 23712 272
rect 711 28 771 30
rect 711 -28 713 28
rect 769 -28 771 28
rect 711 -30 771 -28
rect 2193 28 2253 30
rect 2193 -28 2195 28
rect 2251 -28 2253 28
rect 2193 -30 2253 -28
rect 3675 28 3735 30
rect 3675 -28 3677 28
rect 3733 -28 3735 28
rect 3675 -30 3735 -28
rect 5157 28 5217 30
rect 5157 -28 5159 28
rect 5215 -28 5217 28
rect 5157 -30 5217 -28
rect 6639 28 6699 30
rect 6639 -28 6641 28
rect 6697 -28 6699 28
rect 6639 -30 6699 -28
rect 8121 28 8181 30
rect 8121 -28 8123 28
rect 8179 -28 8181 28
rect 8121 -30 8181 -28
rect 9603 28 9663 30
rect 9603 -28 9605 28
rect 9661 -28 9663 28
rect 9603 -30 9663 -28
rect 11085 28 11145 30
rect 11085 -28 11087 28
rect 11143 -28 11145 28
rect 11085 -30 11145 -28
rect 12567 28 12627 30
rect 12567 -28 12569 28
rect 12625 -28 12627 28
rect 12567 -30 12627 -28
rect 14049 28 14109 30
rect 14049 -28 14051 28
rect 14107 -28 14109 28
rect 14049 -30 14109 -28
rect 15531 28 15591 30
rect 15531 -28 15533 28
rect 15589 -28 15591 28
rect 15531 -30 15591 -28
rect 17013 28 17073 30
rect 17013 -28 17015 28
rect 17071 -28 17073 28
rect 17013 -30 17073 -28
rect 18495 28 18555 30
rect 18495 -28 18497 28
rect 18553 -28 18555 28
rect 18495 -30 18555 -28
rect 19977 28 20037 30
rect 19977 -28 19979 28
rect 20035 -28 20037 28
rect 19977 -30 20037 -28
rect 21459 28 21519 30
rect 21459 -28 21461 28
rect 21517 -28 21519 28
rect 21459 -30 21519 -28
rect 22941 28 23001 30
rect 22941 -28 22943 28
rect 22999 -28 23001 28
rect 22941 -30 23001 -28
use contact_18  contact_18_0
timestamp 1643671299
transform 1 0 22227 0 1 270
box 0 0 1 1
use contact_18  contact_18_1
timestamp 1643671299
transform 1 0 20745 0 1 270
box 0 0 1 1
use contact_18  contact_18_2
timestamp 1643671299
transform 1 0 19263 0 1 270
box 0 0 1 1
use contact_18  contact_18_3
timestamp 1643671299
transform 1 0 17781 0 1 270
box 0 0 1 1
use contact_18  contact_18_4
timestamp 1643671299
transform 1 0 16299 0 1 270
box 0 0 1 1
use contact_18  contact_18_5
timestamp 1643671299
transform 1 0 14817 0 1 270
box 0 0 1 1
use contact_18  contact_18_6
timestamp 1643671299
transform 1 0 13335 0 1 270
box 0 0 1 1
use contact_18  contact_18_7
timestamp 1643671299
transform 1 0 11853 0 1 270
box 0 0 1 1
use contact_18  contact_18_8
timestamp 1643671299
transform 1 0 10371 0 1 270
box 0 0 1 1
use contact_18  contact_18_9
timestamp 1643671299
transform 1 0 8889 0 1 270
box 0 0 1 1
use contact_18  contact_18_10
timestamp 1643671299
transform 1 0 7407 0 1 270
box 0 0 1 1
use contact_18  contact_18_11
timestamp 1643671299
transform 1 0 5925 0 1 270
box 0 0 1 1
use contact_18  contact_18_12
timestamp 1643671299
transform 1 0 4443 0 1 270
box 0 0 1 1
use contact_18  contact_18_13
timestamp 1643671299
transform 1 0 2961 0 1 270
box 0 0 1 1
use contact_18  contact_18_14
timestamp 1643671299
transform 1 0 1479 0 1 270
box 0 0 1 1
use contact_18  contact_18_15
timestamp 1643671299
transform 1 0 -3 0 1 270
box 0 0 1 1
use contact_18  contact_18_16
timestamp 1643671299
transform 1 0 22941 0 1 -30
box 0 0 1 1
use contact_17  contact_17_0
timestamp 1643671299
transform 1 0 22956 0 1 -15
box 0 0 1 1
use contact_18  contact_18_17
timestamp 1643671299
transform 1 0 22941 0 1 808
box 0 0 1 1
use contact_17  contact_17_1
timestamp 1643671299
transform 1 0 22956 0 1 823
box 0 0 1 1
use contact_18  contact_18_18
timestamp 1643671299
transform 1 0 21459 0 1 -30
box 0 0 1 1
use contact_17  contact_17_2
timestamp 1643671299
transform 1 0 21474 0 1 -15
box 0 0 1 1
use contact_18  contact_18_19
timestamp 1643671299
transform 1 0 21459 0 1 808
box 0 0 1 1
use contact_17  contact_17_3
timestamp 1643671299
transform 1 0 21474 0 1 823
box 0 0 1 1
use contact_18  contact_18_20
timestamp 1643671299
transform 1 0 19977 0 1 -30
box 0 0 1 1
use contact_17  contact_17_4
timestamp 1643671299
transform 1 0 19992 0 1 -15
box 0 0 1 1
use contact_18  contact_18_21
timestamp 1643671299
transform 1 0 19977 0 1 808
box 0 0 1 1
use contact_17  contact_17_5
timestamp 1643671299
transform 1 0 19992 0 1 823
box 0 0 1 1
use contact_18  contact_18_22
timestamp 1643671299
transform 1 0 18495 0 1 -30
box 0 0 1 1
use contact_17  contact_17_6
timestamp 1643671299
transform 1 0 18510 0 1 -15
box 0 0 1 1
use contact_18  contact_18_23
timestamp 1643671299
transform 1 0 18495 0 1 808
box 0 0 1 1
use contact_17  contact_17_7
timestamp 1643671299
transform 1 0 18510 0 1 823
box 0 0 1 1
use contact_18  contact_18_24
timestamp 1643671299
transform 1 0 17013 0 1 -30
box 0 0 1 1
use contact_17  contact_17_8
timestamp 1643671299
transform 1 0 17028 0 1 -15
box 0 0 1 1
use contact_18  contact_18_25
timestamp 1643671299
transform 1 0 17013 0 1 808
box 0 0 1 1
use contact_17  contact_17_9
timestamp 1643671299
transform 1 0 17028 0 1 823
box 0 0 1 1
use contact_18  contact_18_26
timestamp 1643671299
transform 1 0 15531 0 1 -30
box 0 0 1 1
use contact_17  contact_17_10
timestamp 1643671299
transform 1 0 15546 0 1 -15
box 0 0 1 1
use contact_18  contact_18_27
timestamp 1643671299
transform 1 0 15531 0 1 808
box 0 0 1 1
use contact_17  contact_17_11
timestamp 1643671299
transform 1 0 15546 0 1 823
box 0 0 1 1
use contact_18  contact_18_28
timestamp 1643671299
transform 1 0 14049 0 1 -30
box 0 0 1 1
use contact_17  contact_17_12
timestamp 1643671299
transform 1 0 14064 0 1 -15
box 0 0 1 1
use contact_18  contact_18_29
timestamp 1643671299
transform 1 0 14049 0 1 808
box 0 0 1 1
use contact_17  contact_17_13
timestamp 1643671299
transform 1 0 14064 0 1 823
box 0 0 1 1
use contact_18  contact_18_30
timestamp 1643671299
transform 1 0 12567 0 1 -30
box 0 0 1 1
use contact_17  contact_17_14
timestamp 1643671299
transform 1 0 12582 0 1 -15
box 0 0 1 1
use contact_18  contact_18_31
timestamp 1643671299
transform 1 0 12567 0 1 808
box 0 0 1 1
use contact_17  contact_17_15
timestamp 1643671299
transform 1 0 12582 0 1 823
box 0 0 1 1
use contact_18  contact_18_32
timestamp 1643671299
transform 1 0 11085 0 1 -30
box 0 0 1 1
use contact_17  contact_17_16
timestamp 1643671299
transform 1 0 11100 0 1 -15
box 0 0 1 1
use contact_18  contact_18_33
timestamp 1643671299
transform 1 0 11085 0 1 808
box 0 0 1 1
use contact_17  contact_17_17
timestamp 1643671299
transform 1 0 11100 0 1 823
box 0 0 1 1
use contact_18  contact_18_34
timestamp 1643671299
transform 1 0 9603 0 1 -30
box 0 0 1 1
use contact_17  contact_17_18
timestamp 1643671299
transform 1 0 9618 0 1 -15
box 0 0 1 1
use contact_18  contact_18_35
timestamp 1643671299
transform 1 0 9603 0 1 808
box 0 0 1 1
use contact_17  contact_17_19
timestamp 1643671299
transform 1 0 9618 0 1 823
box 0 0 1 1
use contact_18  contact_18_36
timestamp 1643671299
transform 1 0 8121 0 1 -30
box 0 0 1 1
use contact_17  contact_17_20
timestamp 1643671299
transform 1 0 8136 0 1 -15
box 0 0 1 1
use contact_18  contact_18_37
timestamp 1643671299
transform 1 0 8121 0 1 808
box 0 0 1 1
use contact_17  contact_17_21
timestamp 1643671299
transform 1 0 8136 0 1 823
box 0 0 1 1
use contact_18  contact_18_38
timestamp 1643671299
transform 1 0 6639 0 1 -30
box 0 0 1 1
use contact_17  contact_17_22
timestamp 1643671299
transform 1 0 6654 0 1 -15
box 0 0 1 1
use contact_18  contact_18_39
timestamp 1643671299
transform 1 0 6639 0 1 808
box 0 0 1 1
use contact_17  contact_17_23
timestamp 1643671299
transform 1 0 6654 0 1 823
box 0 0 1 1
use contact_18  contact_18_40
timestamp 1643671299
transform 1 0 5157 0 1 -30
box 0 0 1 1
use contact_17  contact_17_24
timestamp 1643671299
transform 1 0 5172 0 1 -15
box 0 0 1 1
use contact_18  contact_18_41
timestamp 1643671299
transform 1 0 5157 0 1 808
box 0 0 1 1
use contact_17  contact_17_25
timestamp 1643671299
transform 1 0 5172 0 1 823
box 0 0 1 1
use contact_18  contact_18_42
timestamp 1643671299
transform 1 0 3675 0 1 -30
box 0 0 1 1
use contact_17  contact_17_26
timestamp 1643671299
transform 1 0 3690 0 1 -15
box 0 0 1 1
use contact_18  contact_18_43
timestamp 1643671299
transform 1 0 3675 0 1 808
box 0 0 1 1
use contact_17  contact_17_27
timestamp 1643671299
transform 1 0 3690 0 1 823
box 0 0 1 1
use contact_18  contact_18_44
timestamp 1643671299
transform 1 0 2193 0 1 -30
box 0 0 1 1
use contact_17  contact_17_28
timestamp 1643671299
transform 1 0 2208 0 1 -15
box 0 0 1 1
use contact_18  contact_18_45
timestamp 1643671299
transform 1 0 2193 0 1 808
box 0 0 1 1
use contact_17  contact_17_29
timestamp 1643671299
transform 1 0 2208 0 1 823
box 0 0 1 1
use contact_18  contact_18_46
timestamp 1643671299
transform 1 0 711 0 1 -30
box 0 0 1 1
use contact_17  contact_17_30
timestamp 1643671299
transform 1 0 726 0 1 -15
box 0 0 1 1
use contact_18  contact_18_47
timestamp 1643671299
transform 1 0 711 0 1 808
box 0 0 1 1
use contact_17  contact_17_31
timestamp 1643671299
transform 1 0 726 0 1 823
box 0 0 1 1
use dff  dff_0
timestamp 1643671299
transform 1 0 22230 0 1 0
box 0 -42 1482 916
use dff  dff_1
timestamp 1643671299
transform 1 0 20748 0 1 0
box 0 -42 1482 916
use dff  dff_2
timestamp 1643671299
transform 1 0 19266 0 1 0
box 0 -42 1482 916
use dff  dff_3
timestamp 1643671299
transform 1 0 17784 0 1 0
box 0 -42 1482 916
use dff  dff_4
timestamp 1643671299
transform 1 0 16302 0 1 0
box 0 -42 1482 916
use dff  dff_5
timestamp 1643671299
transform 1 0 14820 0 1 0
box 0 -42 1482 916
use dff  dff_6
timestamp 1643671299
transform 1 0 13338 0 1 0
box 0 -42 1482 916
use dff  dff_7
timestamp 1643671299
transform 1 0 11856 0 1 0
box 0 -42 1482 916
use dff  dff_8
timestamp 1643671299
transform 1 0 10374 0 1 0
box 0 -42 1482 916
use dff  dff_9
timestamp 1643671299
transform 1 0 8892 0 1 0
box 0 -42 1482 916
use dff  dff_10
timestamp 1643671299
transform 1 0 7410 0 1 0
box 0 -42 1482 916
use dff  dff_11
timestamp 1643671299
transform 1 0 5928 0 1 0
box 0 -42 1482 916
use dff  dff_12
timestamp 1643671299
transform 1 0 4446 0 1 0
box 0 -42 1482 916
use dff  dff_13
timestamp 1643671299
transform 1 0 2964 0 1 0
box 0 -42 1482 916
use dff  dff_14
timestamp 1643671299
transform 1 0 1482 0 1 0
box 0 -42 1482 916
use dff  dff_15
timestamp 1643671299
transform 1 0 0 0 1 0
box 0 -42 1482 916
<< labels >>
rlabel metal3 s 8121 808 8181 868 4 vdd
rlabel metal3 s 6639 808 6699 868 4 vdd
rlabel metal3 s 21459 808 21519 868 4 vdd
rlabel metal3 s 2193 808 2253 868 4 vdd
rlabel metal3 s 11085 808 11145 868 4 vdd
rlabel metal3 s 18495 808 18555 868 4 vdd
rlabel metal3 s 14049 808 14109 868 4 vdd
rlabel metal3 s 3675 808 3735 868 4 vdd
rlabel metal3 s 5157 808 5217 868 4 vdd
rlabel metal3 s 12567 808 12627 868 4 vdd
rlabel metal3 s 15531 808 15591 868 4 vdd
rlabel metal3 s 19977 808 20037 868 4 vdd
rlabel metal3 s 17013 808 17073 868 4 vdd
rlabel metal3 s 22941 808 23001 868 4 vdd
rlabel metal3 s 711 808 771 868 4 vdd
rlabel metal3 s 9603 808 9663 868 4 vdd
rlabel metal3 s 3675 -30 3735 30 4 gnd
rlabel metal3 s 5157 -30 5217 30 4 gnd
rlabel metal3 s 8121 -30 8181 30 4 gnd
rlabel metal3 s 11085 -30 11145 30 4 gnd
rlabel metal3 s 15531 -30 15591 30 4 gnd
rlabel metal3 s 6639 -30 6699 30 4 gnd
rlabel metal3 s 711 -30 771 30 4 gnd
rlabel metal3 s 19977 -30 20037 30 4 gnd
rlabel metal3 s 9603 -30 9663 30 4 gnd
rlabel metal3 s 14049 -30 14109 30 4 gnd
rlabel metal3 s 22941 -30 23001 30 4 gnd
rlabel metal3 s 17013 -30 17073 30 4 gnd
rlabel metal3 s 18495 -30 18555 30 4 gnd
rlabel metal3 s 21459 -30 21519 30 4 gnd
rlabel metal3 s 2193 -30 2253 30 4 gnd
rlabel metal3 s 12567 -30 12627 30 4 gnd
rlabel metal2 s 180 232 234 260 4 din_0
rlabel metal2 s 1260 228 1314 256 4 dout_0
rlabel metal2 s 1662 232 1716 260 4 din_1
rlabel metal2 s 2742 228 2796 256 4 dout_1
rlabel metal2 s 3144 232 3198 260 4 din_2
rlabel metal2 s 4224 228 4278 256 4 dout_2
rlabel metal2 s 4626 232 4680 260 4 din_3
rlabel metal2 s 5706 228 5760 256 4 dout_3
rlabel metal2 s 6108 232 6162 260 4 din_4
rlabel metal2 s 7188 228 7242 256 4 dout_4
rlabel metal2 s 7590 232 7644 260 4 din_5
rlabel metal2 s 8670 228 8724 256 4 dout_5
rlabel metal2 s 9072 232 9126 260 4 din_6
rlabel metal2 s 10152 228 10206 256 4 dout_6
rlabel metal2 s 10554 232 10608 260 4 din_7
rlabel metal2 s 11634 228 11688 256 4 dout_7
rlabel metal2 s 12036 232 12090 260 4 din_8
rlabel metal2 s 13116 228 13170 256 4 dout_8
rlabel metal2 s 13518 232 13572 260 4 din_9
rlabel metal2 s 14598 228 14652 256 4 dout_9
rlabel metal2 s 15000 232 15054 260 4 din_10
rlabel metal2 s 16080 228 16134 256 4 dout_10
rlabel metal2 s 16482 232 16536 260 4 din_11
rlabel metal2 s 17562 228 17616 256 4 dout_11
rlabel metal2 s 17964 232 18018 260 4 din_12
rlabel metal2 s 19044 228 19098 256 4 dout_12
rlabel metal2 s 19446 232 19500 260 4 din_13
rlabel metal2 s 20526 228 20580 256 4 dout_13
rlabel metal2 s 20928 232 20982 260 4 din_14
rlabel metal2 s 22008 228 22062 256 4 dout_14
rlabel metal2 s 22410 232 22464 260 4 din_15
rlabel metal2 s 23490 228 23544 256 4 dout_15
rlabel metal3 s 0 270 23712 330 4 clk
<< properties >>
string FIXED_BBOX 22941 -30 23001 0
string GDS_FILE sram_0rw2r1w_16_32_sky130A.gds
string GDS_END 1252726
string GDS_START 1233612
<< end >>
