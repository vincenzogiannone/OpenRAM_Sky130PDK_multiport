magic
tech sky130A
magscale 1 2
timestamp 1644969367
<< checkpaint >>
rect -1260 -1260 1958 2212
<< nwell >>
rect 0 472 698 952
<< pwell >>
rect 122 0 194 84
rect 314 0 386 84
rect 506 0 578 84
<< nmos >>
rect 108 138 138 222
rect 220 138 250 222
rect 448 138 478 222
rect 560 138 590 222
<< pmos >>
rect 108 508 138 778
rect 220 508 250 778
rect 448 508 478 778
rect 560 508 590 778
<< ndiff >>
rect 36 196 108 222
rect 36 162 50 196
rect 84 162 108 196
rect 36 138 108 162
rect 138 196 220 222
rect 138 162 162 196
rect 196 162 220 196
rect 138 138 220 162
rect 250 196 322 222
rect 250 162 274 196
rect 308 162 322 196
rect 250 138 322 162
rect 376 196 448 222
rect 376 162 390 196
rect 424 162 448 196
rect 376 138 448 162
rect 478 138 560 222
rect 590 196 662 222
rect 590 162 614 196
rect 648 162 662 196
rect 590 138 662 162
<< pdiff >>
rect 36 736 108 778
rect 36 702 50 736
rect 84 702 108 736
rect 36 660 108 702
rect 36 626 50 660
rect 84 626 108 660
rect 36 584 108 626
rect 36 550 50 584
rect 84 550 108 584
rect 36 508 108 550
rect 138 736 220 778
rect 138 702 162 736
rect 196 702 220 736
rect 138 660 220 702
rect 138 626 162 660
rect 196 626 220 660
rect 138 584 220 626
rect 138 550 162 584
rect 196 550 220 584
rect 138 508 220 550
rect 250 736 322 778
rect 250 702 274 736
rect 308 702 322 736
rect 250 660 322 702
rect 250 626 274 660
rect 308 626 322 660
rect 250 584 322 626
rect 250 550 274 584
rect 308 550 322 584
rect 250 508 322 550
rect 376 736 448 778
rect 376 702 390 736
rect 424 702 448 736
rect 376 660 448 702
rect 376 626 390 660
rect 424 626 448 660
rect 376 584 448 626
rect 376 550 390 584
rect 424 550 448 584
rect 376 508 448 550
rect 478 508 560 778
rect 590 736 662 778
rect 590 702 614 736
rect 648 702 662 736
rect 590 660 662 702
rect 590 626 614 660
rect 648 626 662 660
rect 590 584 662 626
rect 590 550 614 584
rect 648 550 662 584
rect 590 508 662 550
<< ndiffc >>
rect 50 162 84 196
rect 162 162 196 196
rect 274 162 308 196
rect 390 162 424 196
rect 614 162 648 196
<< pdiffc >>
rect 50 702 84 736
rect 50 626 84 660
rect 50 550 84 584
rect 162 702 196 736
rect 162 626 196 660
rect 162 550 196 584
rect 274 702 308 736
rect 274 626 308 660
rect 274 550 308 584
rect 390 702 424 736
rect 390 626 424 660
rect 390 550 424 584
rect 614 702 648 736
rect 614 626 648 660
rect 614 550 648 584
<< psubdiff >>
rect 122 59 194 84
rect 122 25 141 59
rect 175 25 194 59
rect 122 0 194 25
rect 314 59 386 84
rect 314 25 333 59
rect 367 25 386 59
rect 314 0 386 25
rect 506 59 578 84
rect 506 25 525 59
rect 559 25 578 59
rect 506 0 578 25
<< nsubdiff >>
rect 122 891 194 916
rect 122 857 141 891
rect 175 857 194 891
rect 122 832 194 857
rect 314 891 386 916
rect 314 857 333 891
rect 367 857 386 891
rect 314 832 386 857
rect 506 891 578 916
rect 506 857 525 891
rect 559 857 578 891
rect 506 832 578 857
<< psubdiffcont >>
rect 141 25 175 59
rect 333 25 367 59
rect 525 25 559 59
<< nsubdiffcont >>
rect 141 857 175 891
rect 333 857 367 891
rect 525 857 559 891
<< poly >>
rect 108 778 138 804
rect 220 778 250 804
rect 448 778 478 804
rect 560 778 590 804
rect 108 406 138 508
rect 8 390 138 406
rect 8 356 18 390
rect 52 376 138 390
rect 52 356 62 376
rect 8 340 62 356
rect 108 222 138 376
rect 220 322 250 508
rect 448 474 478 508
rect 560 474 590 508
rect 424 458 478 474
rect 424 424 434 458
rect 468 424 478 458
rect 424 408 478 424
rect 536 458 590 474
rect 536 424 546 458
rect 580 424 590 458
rect 536 408 590 424
rect 196 306 250 322
rect 196 272 206 306
rect 240 272 250 306
rect 196 256 250 272
rect 220 222 250 256
rect 448 222 478 408
rect 536 306 590 322
rect 536 272 546 306
rect 580 272 590 306
rect 536 256 590 272
rect 560 222 590 256
rect 108 112 138 138
rect 220 112 250 138
rect 448 112 478 138
rect 560 112 590 138
<< polycont >>
rect 18 356 52 390
rect 434 424 468 458
rect 546 424 580 458
rect 206 272 240 306
rect 546 272 580 306
<< locali >>
rect 140 891 182 908
rect 140 857 141 891
rect 175 857 182 891
rect 140 840 182 857
rect 332 891 368 908
rect 332 857 333 891
rect 367 874 368 891
rect 524 891 560 908
rect 367 857 410 874
rect 332 840 410 857
rect 524 857 525 891
rect 559 857 560 891
rect 524 840 560 857
rect 148 778 182 840
rect 376 778 410 840
rect 36 736 98 778
rect 36 702 50 736
rect 84 702 98 736
rect 36 660 98 702
rect 36 626 50 660
rect 84 626 98 660
rect 36 584 98 626
rect 36 550 50 584
rect 84 550 98 584
rect 36 508 98 550
rect 148 736 210 778
rect 148 702 162 736
rect 196 702 210 736
rect 148 660 210 702
rect 148 626 162 660
rect 196 626 210 660
rect 148 584 210 626
rect 148 550 162 584
rect 196 550 210 584
rect 148 508 210 550
rect 260 736 322 778
rect 260 702 274 736
rect 308 702 322 736
rect 260 660 322 702
rect 260 626 274 660
rect 308 626 322 660
rect 260 584 322 626
rect 260 550 274 584
rect 308 550 322 584
rect 260 508 322 550
rect 376 736 438 778
rect 376 702 390 736
rect 424 702 438 736
rect 376 660 438 702
rect 376 626 390 660
rect 424 626 438 660
rect 376 584 438 626
rect 376 550 390 584
rect 424 550 438 584
rect 376 508 438 550
rect 600 736 662 778
rect 600 702 614 736
rect 648 702 662 736
rect 600 660 662 702
rect 600 626 614 660
rect 648 626 662 660
rect 600 584 662 626
rect 600 550 614 584
rect 648 550 662 584
rect 600 508 662 550
rect 64 474 98 508
rect 64 440 138 474
rect 18 390 52 406
rect 18 340 52 356
rect 104 294 138 440
rect 288 460 322 508
rect 434 460 468 474
rect 288 458 468 460
rect 288 424 434 458
rect 64 258 138 294
rect 206 306 240 322
rect 64 222 98 258
rect 206 256 240 272
rect 288 222 322 424
rect 434 408 468 424
rect 546 458 580 474
rect 546 408 580 424
rect 546 306 580 322
rect 546 256 580 272
rect 628 306 662 508
rect 628 222 662 272
rect 36 196 98 222
rect 36 162 50 196
rect 84 162 98 196
rect 36 138 98 162
rect 148 196 210 222
rect 148 162 162 196
rect 196 162 210 196
rect 148 138 210 162
rect 260 196 322 222
rect 260 162 274 196
rect 308 162 322 196
rect 260 138 322 162
rect 376 196 438 222
rect 376 162 390 196
rect 424 162 438 196
rect 376 138 438 162
rect 600 196 662 222
rect 600 162 614 196
rect 648 162 662 196
rect 600 138 662 162
rect 148 76 182 138
rect 376 76 410 138
rect 140 59 182 76
rect 140 25 141 59
rect 175 25 182 59
rect 140 8 182 25
rect 332 59 410 76
rect 332 25 333 59
rect 367 42 410 59
rect 524 59 560 76
rect 367 25 368 42
rect 332 8 368 25
rect 524 25 525 59
rect 559 25 560 59
rect 524 8 560 25
<< viali >>
rect 141 857 175 891
rect 333 857 367 891
rect 525 857 559 891
rect 50 550 84 584
rect 18 356 52 390
rect 206 272 240 306
rect 546 424 580 458
rect 546 272 580 306
rect 628 272 662 306
rect 141 25 175 59
rect 333 25 367 59
rect 525 25 559 59
<< metal1 >>
rect 0 891 698 904
rect 0 857 141 891
rect 175 857 333 891
rect 367 857 525 891
rect 559 857 698 891
rect 0 844 698 857
rect 44 584 90 596
rect 44 550 50 584
rect 84 566 90 584
rect 84 550 568 566
rect 44 538 568 550
rect 540 470 568 538
rect 540 458 586 470
rect 540 424 546 458
rect 580 424 586 458
rect 540 412 586 424
rect 10 390 62 404
rect 10 384 18 390
rect 8 356 18 384
rect 52 384 62 390
rect 52 356 402 384
rect 10 340 62 356
rect 196 314 250 320
rect 196 262 198 314
rect 374 318 402 356
rect 374 306 586 318
rect 374 290 546 306
rect 196 256 250 262
rect 540 272 546 290
rect 580 272 586 306
rect 540 260 586 272
rect 618 316 670 322
rect 618 258 670 264
rect 0 59 698 72
rect 0 25 141 59
rect 175 25 333 59
rect 367 25 525 59
rect 559 25 698 59
rect 0 12 698 25
<< via1 >>
rect 198 306 250 314
rect 198 272 206 306
rect 206 272 240 306
rect 240 272 250 306
rect 198 262 250 272
rect 618 306 670 316
rect 618 272 628 306
rect 628 272 662 306
rect 662 272 670 306
rect 618 264 670 272
<< metal2 >>
rect 630 322 658 952
rect 198 314 250 320
rect 196 272 198 300
rect 198 256 250 262
rect 618 316 670 322
rect 618 258 670 264
rect 630 0 658 258
<< labels >>
rlabel locali s 76 270 76 270 4 enb
rlabel locali s 306 316 306 316 4 net1
rlabel mvpsubdiff s 520 664 520 664 4 net2
rlabel mvpsubdiff s 516 174 516 174 4 net3
rlabel metal2 s 196 272 250 300 4 din
port 1 nsew
rlabel metal1 s 0 844 698 904 4 vdd
port 2 nsew
rlabel metal1 s 0 12 698 72 4 gnd
port 3 nsew
rlabel metal1 s 8 356 402 384 4 en
port 4 nsew
rlabel metal2 s 630 322 658 952 4 wbl
port 5 nsew
rlabel metal2 s 223 286 223 286 4 din
rlabel metal1 s 205 370 205 370 4 en
rlabel metal2 s 644 637 644 637 4 wbl
rlabel metal1 s 349 874 349 874 4 vdd
rlabel metal1 s 349 42 349 42 4 gnd
<< properties >>
string FIXED_BBOX 0 0 698 952
string GDS_FILE sram_0rw2r1w_32_128_sky130A.gds
string GDS_END 2648184
string GDS_START 2638028
<< end >>
