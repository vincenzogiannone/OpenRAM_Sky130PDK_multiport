magic
tech sky130A
magscale 1 2
timestamp 1644969367
<< checkpaint >>
rect -1260 -1284 50583 2212
<< metal1 >>
rect 712 900 764 906
rect 712 842 764 848
rect 2268 900 2320 906
rect 2268 842 2320 848
rect 3824 900 3876 906
rect 3824 842 3876 848
rect 5380 900 5432 906
rect 5380 842 5432 848
rect 6936 900 6988 906
rect 6936 842 6988 848
rect 8492 900 8544 906
rect 8492 842 8544 848
rect 10048 900 10100 906
rect 10048 842 10100 848
rect 11604 900 11656 906
rect 11604 842 11656 848
rect 13160 900 13212 906
rect 13160 842 13212 848
rect 14716 900 14768 906
rect 14716 842 14768 848
rect 16272 900 16324 906
rect 16272 842 16324 848
rect 17828 900 17880 906
rect 17828 842 17880 848
rect 19384 900 19436 906
rect 19384 842 19436 848
rect 20940 900 20992 906
rect 20940 842 20992 848
rect 22496 900 22548 906
rect 22496 842 22548 848
rect 24052 900 24104 906
rect 24052 842 24104 848
rect 25608 900 25660 906
rect 25608 842 25660 848
rect 27164 900 27216 906
rect 27164 842 27216 848
rect 28720 900 28772 906
rect 28720 842 28772 848
rect 30276 900 30328 906
rect 30276 842 30328 848
rect 31832 900 31884 906
rect 31832 842 31884 848
rect 33388 900 33440 906
rect 33388 842 33440 848
rect 34944 900 34996 906
rect 34944 842 34996 848
rect 36500 900 36552 906
rect 36500 842 36552 848
rect 38056 900 38108 906
rect 38056 842 38108 848
rect 39612 900 39664 906
rect 39612 842 39664 848
rect 41168 900 41220 906
rect 41168 842 41220 848
rect 42724 900 42776 906
rect 42724 842 42776 848
rect 44280 900 44332 906
rect 44280 842 44332 848
rect 45836 900 45888 906
rect 45836 842 45888 848
rect 47392 900 47444 906
rect 47392 842 47444 848
rect 48948 900 49000 906
rect 48948 842 49000 848
rect 0 356 49323 384
rect 712 68 764 74
rect 712 10 764 16
rect 2268 68 2320 74
rect 2268 10 2320 16
rect 3824 68 3876 74
rect 3824 10 3876 16
rect 5380 68 5432 74
rect 5380 10 5432 16
rect 6936 68 6988 74
rect 6936 10 6988 16
rect 8492 68 8544 74
rect 8492 10 8544 16
rect 10048 68 10100 74
rect 10048 10 10100 16
rect 11604 68 11656 74
rect 11604 10 11656 16
rect 13160 68 13212 74
rect 13160 10 13212 16
rect 14716 68 14768 74
rect 14716 10 14768 16
rect 16272 68 16324 74
rect 16272 10 16324 16
rect 17828 68 17880 74
rect 17828 10 17880 16
rect 19384 68 19436 74
rect 19384 10 19436 16
rect 20940 68 20992 74
rect 20940 10 20992 16
rect 22496 68 22548 74
rect 22496 10 22548 16
rect 24052 68 24104 74
rect 24052 10 24104 16
rect 25608 68 25660 74
rect 25608 10 25660 16
rect 27164 68 27216 74
rect 27164 10 27216 16
rect 28720 68 28772 74
rect 28720 10 28772 16
rect 30276 68 30328 74
rect 30276 10 30328 16
rect 31832 68 31884 74
rect 31832 10 31884 16
rect 33388 68 33440 74
rect 33388 10 33440 16
rect 34944 68 34996 74
rect 34944 10 34996 16
rect 36500 68 36552 74
rect 36500 10 36552 16
rect 38056 68 38108 74
rect 38056 10 38108 16
rect 39612 68 39664 74
rect 39612 10 39664 16
rect 41168 68 41220 74
rect 41168 10 41220 16
rect 42724 68 42776 74
rect 42724 10 42776 16
rect 44280 68 44332 74
rect 44280 10 44332 16
rect 45836 68 45888 74
rect 45836 10 45888 16
rect 47392 68 47444 74
rect 47392 10 47444 16
rect 48948 68 49000 74
rect 48948 10 49000 16
<< via1 >>
rect 712 848 764 900
rect 2268 848 2320 900
rect 3824 848 3876 900
rect 5380 848 5432 900
rect 6936 848 6988 900
rect 8492 848 8544 900
rect 10048 848 10100 900
rect 11604 848 11656 900
rect 13160 848 13212 900
rect 14716 848 14768 900
rect 16272 848 16324 900
rect 17828 848 17880 900
rect 19384 848 19436 900
rect 20940 848 20992 900
rect 22496 848 22548 900
rect 24052 848 24104 900
rect 25608 848 25660 900
rect 27164 848 27216 900
rect 28720 848 28772 900
rect 30276 848 30328 900
rect 31832 848 31884 900
rect 33388 848 33440 900
rect 34944 848 34996 900
rect 36500 848 36552 900
rect 38056 848 38108 900
rect 39612 848 39664 900
rect 41168 848 41220 900
rect 42724 848 42776 900
rect 44280 848 44332 900
rect 45836 848 45888 900
rect 47392 848 47444 900
rect 48948 848 49000 900
rect 712 16 764 68
rect 2268 16 2320 68
rect 3824 16 3876 68
rect 5380 16 5432 68
rect 6936 16 6988 68
rect 8492 16 8544 68
rect 10048 16 10100 68
rect 11604 16 11656 68
rect 13160 16 13212 68
rect 14716 16 14768 68
rect 16272 16 16324 68
rect 17828 16 17880 68
rect 19384 16 19436 68
rect 20940 16 20992 68
rect 22496 16 22548 68
rect 24052 16 24104 68
rect 25608 16 25660 68
rect 27164 16 27216 68
rect 28720 16 28772 68
rect 30276 16 30328 68
rect 31832 16 31884 68
rect 33388 16 33440 68
rect 34944 16 34996 68
rect 36500 16 36552 68
rect 38056 16 38108 68
rect 39612 16 39664 68
rect 41168 16 41220 68
rect 42724 16 42776 68
rect 44280 16 44332 68
rect 45836 16 45888 68
rect 47392 16 47444 68
rect 48948 16 49000 68
<< metal2 >>
rect 710 902 766 911
rect 710 837 766 846
rect 1019 322 1047 952
rect 2266 902 2322 911
rect 2266 837 2322 846
rect 2575 322 2603 952
rect 3822 902 3878 911
rect 3822 837 3878 846
rect 4131 322 4159 952
rect 5378 902 5434 911
rect 5378 837 5434 846
rect 5687 322 5715 952
rect 6934 902 6990 911
rect 6934 837 6990 846
rect 7243 322 7271 952
rect 8490 902 8546 911
rect 8490 837 8546 846
rect 8799 322 8827 952
rect 10046 902 10102 911
rect 10046 837 10102 846
rect 10355 322 10383 952
rect 11602 902 11658 911
rect 11602 837 11658 846
rect 11911 322 11939 952
rect 13158 902 13214 911
rect 13158 837 13214 846
rect 13467 322 13495 952
rect 14714 902 14770 911
rect 14714 837 14770 846
rect 15023 322 15051 952
rect 16270 902 16326 911
rect 16270 837 16326 846
rect 16579 322 16607 952
rect 17826 902 17882 911
rect 17826 837 17882 846
rect 18135 322 18163 952
rect 19382 902 19438 911
rect 19382 837 19438 846
rect 19691 322 19719 952
rect 20938 902 20994 911
rect 20938 837 20994 846
rect 21247 322 21275 952
rect 22494 902 22550 911
rect 22494 837 22550 846
rect 22803 322 22831 952
rect 24050 902 24106 911
rect 24050 837 24106 846
rect 24359 322 24387 952
rect 25606 902 25662 911
rect 25606 837 25662 846
rect 25915 322 25943 952
rect 27162 902 27218 911
rect 27162 837 27218 846
rect 27471 322 27499 952
rect 28718 902 28774 911
rect 28718 837 28774 846
rect 29027 322 29055 952
rect 30274 902 30330 911
rect 30274 837 30330 846
rect 30583 322 30611 952
rect 31830 902 31886 911
rect 31830 837 31886 846
rect 32139 322 32167 952
rect 33386 902 33442 911
rect 33386 837 33442 846
rect 33695 322 33723 952
rect 34942 902 34998 911
rect 34942 837 34998 846
rect 35251 322 35279 952
rect 36498 902 36554 911
rect 36498 837 36554 846
rect 36807 322 36835 952
rect 38054 902 38110 911
rect 38054 837 38110 846
rect 38363 322 38391 952
rect 39610 902 39666 911
rect 39610 837 39666 846
rect 39919 322 39947 952
rect 41166 902 41222 911
rect 41166 837 41222 846
rect 41475 322 41503 952
rect 42722 902 42778 911
rect 42722 837 42778 846
rect 43031 322 43059 952
rect 44278 902 44334 911
rect 44278 837 44334 846
rect 44587 322 44615 952
rect 45834 902 45890 911
rect 45834 837 45890 846
rect 46143 322 46171 952
rect 47390 902 47446 911
rect 47390 837 47446 846
rect 47699 322 47727 952
rect 48946 902 49002 911
rect 48946 837 49002 846
rect 49255 322 49283 952
rect 585 272 639 300
rect 2141 272 2195 300
rect 3697 272 3751 300
rect 5253 272 5307 300
rect 6809 272 6863 300
rect 8365 272 8419 300
rect 9921 272 9975 300
rect 11477 272 11531 300
rect 13033 272 13087 300
rect 14589 272 14643 300
rect 16145 272 16199 300
rect 17701 272 17755 300
rect 19257 272 19311 300
rect 20813 272 20867 300
rect 22369 272 22423 300
rect 23925 272 23979 300
rect 25481 272 25535 300
rect 27037 272 27091 300
rect 28593 272 28647 300
rect 30149 272 30203 300
rect 31705 272 31759 300
rect 33261 272 33315 300
rect 34817 272 34871 300
rect 36373 272 36427 300
rect 37929 272 37983 300
rect 39485 272 39539 300
rect 41041 272 41095 300
rect 42597 272 42651 300
rect 44153 272 44207 300
rect 45709 272 45763 300
rect 47265 272 47319 300
rect 48821 272 48875 300
rect 710 70 766 79
rect 710 5 766 14
rect 2266 70 2322 79
rect 2266 5 2322 14
rect 3822 70 3878 79
rect 3822 5 3878 14
rect 5378 70 5434 79
rect 5378 5 5434 14
rect 6934 70 6990 79
rect 6934 5 6990 14
rect 8490 70 8546 79
rect 8490 5 8546 14
rect 10046 70 10102 79
rect 10046 5 10102 14
rect 11602 70 11658 79
rect 11602 5 11658 14
rect 13158 70 13214 79
rect 13158 5 13214 14
rect 14714 70 14770 79
rect 14714 5 14770 14
rect 16270 70 16326 79
rect 16270 5 16326 14
rect 17826 70 17882 79
rect 17826 5 17882 14
rect 19382 70 19438 79
rect 19382 5 19438 14
rect 20938 70 20994 79
rect 20938 5 20994 14
rect 22494 70 22550 79
rect 22494 5 22550 14
rect 24050 70 24106 79
rect 24050 5 24106 14
rect 25606 70 25662 79
rect 25606 5 25662 14
rect 27162 70 27218 79
rect 27162 5 27218 14
rect 28718 70 28774 79
rect 28718 5 28774 14
rect 30274 70 30330 79
rect 30274 5 30330 14
rect 31830 70 31886 79
rect 31830 5 31886 14
rect 33386 70 33442 79
rect 33386 5 33442 14
rect 34942 70 34998 79
rect 34942 5 34998 14
rect 36498 70 36554 79
rect 36498 5 36554 14
rect 38054 70 38110 79
rect 38054 5 38110 14
rect 39610 70 39666 79
rect 39610 5 39666 14
rect 41166 70 41222 79
rect 41166 5 41222 14
rect 42722 70 42778 79
rect 42722 5 42778 14
rect 44278 70 44334 79
rect 44278 5 44334 14
rect 45834 70 45890 79
rect 45834 5 45890 14
rect 47390 70 47446 79
rect 47390 5 47446 14
rect 48946 70 49002 79
rect 48946 5 49002 14
<< via2 >>
rect 710 900 766 902
rect 710 848 712 900
rect 712 848 764 900
rect 764 848 766 900
rect 710 846 766 848
rect 2266 900 2322 902
rect 2266 848 2268 900
rect 2268 848 2320 900
rect 2320 848 2322 900
rect 2266 846 2322 848
rect 3822 900 3878 902
rect 3822 848 3824 900
rect 3824 848 3876 900
rect 3876 848 3878 900
rect 3822 846 3878 848
rect 5378 900 5434 902
rect 5378 848 5380 900
rect 5380 848 5432 900
rect 5432 848 5434 900
rect 5378 846 5434 848
rect 6934 900 6990 902
rect 6934 848 6936 900
rect 6936 848 6988 900
rect 6988 848 6990 900
rect 6934 846 6990 848
rect 8490 900 8546 902
rect 8490 848 8492 900
rect 8492 848 8544 900
rect 8544 848 8546 900
rect 8490 846 8546 848
rect 10046 900 10102 902
rect 10046 848 10048 900
rect 10048 848 10100 900
rect 10100 848 10102 900
rect 10046 846 10102 848
rect 11602 900 11658 902
rect 11602 848 11604 900
rect 11604 848 11656 900
rect 11656 848 11658 900
rect 11602 846 11658 848
rect 13158 900 13214 902
rect 13158 848 13160 900
rect 13160 848 13212 900
rect 13212 848 13214 900
rect 13158 846 13214 848
rect 14714 900 14770 902
rect 14714 848 14716 900
rect 14716 848 14768 900
rect 14768 848 14770 900
rect 14714 846 14770 848
rect 16270 900 16326 902
rect 16270 848 16272 900
rect 16272 848 16324 900
rect 16324 848 16326 900
rect 16270 846 16326 848
rect 17826 900 17882 902
rect 17826 848 17828 900
rect 17828 848 17880 900
rect 17880 848 17882 900
rect 17826 846 17882 848
rect 19382 900 19438 902
rect 19382 848 19384 900
rect 19384 848 19436 900
rect 19436 848 19438 900
rect 19382 846 19438 848
rect 20938 900 20994 902
rect 20938 848 20940 900
rect 20940 848 20992 900
rect 20992 848 20994 900
rect 20938 846 20994 848
rect 22494 900 22550 902
rect 22494 848 22496 900
rect 22496 848 22548 900
rect 22548 848 22550 900
rect 22494 846 22550 848
rect 24050 900 24106 902
rect 24050 848 24052 900
rect 24052 848 24104 900
rect 24104 848 24106 900
rect 24050 846 24106 848
rect 25606 900 25662 902
rect 25606 848 25608 900
rect 25608 848 25660 900
rect 25660 848 25662 900
rect 25606 846 25662 848
rect 27162 900 27218 902
rect 27162 848 27164 900
rect 27164 848 27216 900
rect 27216 848 27218 900
rect 27162 846 27218 848
rect 28718 900 28774 902
rect 28718 848 28720 900
rect 28720 848 28772 900
rect 28772 848 28774 900
rect 28718 846 28774 848
rect 30274 900 30330 902
rect 30274 848 30276 900
rect 30276 848 30328 900
rect 30328 848 30330 900
rect 30274 846 30330 848
rect 31830 900 31886 902
rect 31830 848 31832 900
rect 31832 848 31884 900
rect 31884 848 31886 900
rect 31830 846 31886 848
rect 33386 900 33442 902
rect 33386 848 33388 900
rect 33388 848 33440 900
rect 33440 848 33442 900
rect 33386 846 33442 848
rect 34942 900 34998 902
rect 34942 848 34944 900
rect 34944 848 34996 900
rect 34996 848 34998 900
rect 34942 846 34998 848
rect 36498 900 36554 902
rect 36498 848 36500 900
rect 36500 848 36552 900
rect 36552 848 36554 900
rect 36498 846 36554 848
rect 38054 900 38110 902
rect 38054 848 38056 900
rect 38056 848 38108 900
rect 38108 848 38110 900
rect 38054 846 38110 848
rect 39610 900 39666 902
rect 39610 848 39612 900
rect 39612 848 39664 900
rect 39664 848 39666 900
rect 39610 846 39666 848
rect 41166 900 41222 902
rect 41166 848 41168 900
rect 41168 848 41220 900
rect 41220 848 41222 900
rect 41166 846 41222 848
rect 42722 900 42778 902
rect 42722 848 42724 900
rect 42724 848 42776 900
rect 42776 848 42778 900
rect 42722 846 42778 848
rect 44278 900 44334 902
rect 44278 848 44280 900
rect 44280 848 44332 900
rect 44332 848 44334 900
rect 44278 846 44334 848
rect 45834 900 45890 902
rect 45834 848 45836 900
rect 45836 848 45888 900
rect 45888 848 45890 900
rect 45834 846 45890 848
rect 47390 900 47446 902
rect 47390 848 47392 900
rect 47392 848 47444 900
rect 47444 848 47446 900
rect 47390 846 47446 848
rect 48946 900 49002 902
rect 48946 848 48948 900
rect 48948 848 49000 900
rect 49000 848 49002 900
rect 48946 846 49002 848
rect 710 68 766 70
rect 710 16 712 68
rect 712 16 764 68
rect 764 16 766 68
rect 710 14 766 16
rect 2266 68 2322 70
rect 2266 16 2268 68
rect 2268 16 2320 68
rect 2320 16 2322 68
rect 2266 14 2322 16
rect 3822 68 3878 70
rect 3822 16 3824 68
rect 3824 16 3876 68
rect 3876 16 3878 68
rect 3822 14 3878 16
rect 5378 68 5434 70
rect 5378 16 5380 68
rect 5380 16 5432 68
rect 5432 16 5434 68
rect 5378 14 5434 16
rect 6934 68 6990 70
rect 6934 16 6936 68
rect 6936 16 6988 68
rect 6988 16 6990 68
rect 6934 14 6990 16
rect 8490 68 8546 70
rect 8490 16 8492 68
rect 8492 16 8544 68
rect 8544 16 8546 68
rect 8490 14 8546 16
rect 10046 68 10102 70
rect 10046 16 10048 68
rect 10048 16 10100 68
rect 10100 16 10102 68
rect 10046 14 10102 16
rect 11602 68 11658 70
rect 11602 16 11604 68
rect 11604 16 11656 68
rect 11656 16 11658 68
rect 11602 14 11658 16
rect 13158 68 13214 70
rect 13158 16 13160 68
rect 13160 16 13212 68
rect 13212 16 13214 68
rect 13158 14 13214 16
rect 14714 68 14770 70
rect 14714 16 14716 68
rect 14716 16 14768 68
rect 14768 16 14770 68
rect 14714 14 14770 16
rect 16270 68 16326 70
rect 16270 16 16272 68
rect 16272 16 16324 68
rect 16324 16 16326 68
rect 16270 14 16326 16
rect 17826 68 17882 70
rect 17826 16 17828 68
rect 17828 16 17880 68
rect 17880 16 17882 68
rect 17826 14 17882 16
rect 19382 68 19438 70
rect 19382 16 19384 68
rect 19384 16 19436 68
rect 19436 16 19438 68
rect 19382 14 19438 16
rect 20938 68 20994 70
rect 20938 16 20940 68
rect 20940 16 20992 68
rect 20992 16 20994 68
rect 20938 14 20994 16
rect 22494 68 22550 70
rect 22494 16 22496 68
rect 22496 16 22548 68
rect 22548 16 22550 68
rect 22494 14 22550 16
rect 24050 68 24106 70
rect 24050 16 24052 68
rect 24052 16 24104 68
rect 24104 16 24106 68
rect 24050 14 24106 16
rect 25606 68 25662 70
rect 25606 16 25608 68
rect 25608 16 25660 68
rect 25660 16 25662 68
rect 25606 14 25662 16
rect 27162 68 27218 70
rect 27162 16 27164 68
rect 27164 16 27216 68
rect 27216 16 27218 68
rect 27162 14 27218 16
rect 28718 68 28774 70
rect 28718 16 28720 68
rect 28720 16 28772 68
rect 28772 16 28774 68
rect 28718 14 28774 16
rect 30274 68 30330 70
rect 30274 16 30276 68
rect 30276 16 30328 68
rect 30328 16 30330 68
rect 30274 14 30330 16
rect 31830 68 31886 70
rect 31830 16 31832 68
rect 31832 16 31884 68
rect 31884 16 31886 68
rect 31830 14 31886 16
rect 33386 68 33442 70
rect 33386 16 33388 68
rect 33388 16 33440 68
rect 33440 16 33442 68
rect 33386 14 33442 16
rect 34942 68 34998 70
rect 34942 16 34944 68
rect 34944 16 34996 68
rect 34996 16 34998 68
rect 34942 14 34998 16
rect 36498 68 36554 70
rect 36498 16 36500 68
rect 36500 16 36552 68
rect 36552 16 36554 68
rect 36498 14 36554 16
rect 38054 68 38110 70
rect 38054 16 38056 68
rect 38056 16 38108 68
rect 38108 16 38110 68
rect 38054 14 38110 16
rect 39610 68 39666 70
rect 39610 16 39612 68
rect 39612 16 39664 68
rect 39664 16 39666 68
rect 39610 14 39666 16
rect 41166 68 41222 70
rect 41166 16 41168 68
rect 41168 16 41220 68
rect 41220 16 41222 68
rect 41166 14 41222 16
rect 42722 68 42778 70
rect 42722 16 42724 68
rect 42724 16 42776 68
rect 42776 16 42778 68
rect 42722 14 42778 16
rect 44278 68 44334 70
rect 44278 16 44280 68
rect 44280 16 44332 68
rect 44332 16 44334 68
rect 44278 14 44334 16
rect 45834 68 45890 70
rect 45834 16 45836 68
rect 45836 16 45888 68
rect 45888 16 45890 68
rect 45834 14 45890 16
rect 47390 68 47446 70
rect 47390 16 47392 68
rect 47392 16 47444 68
rect 47444 16 47446 68
rect 47390 14 47446 16
rect 48946 68 49002 70
rect 48946 16 48948 68
rect 48948 16 49000 68
rect 49000 16 49002 68
rect 48946 14 49002 16
<< metal3 >>
rect 705 902 771 940
rect 705 846 710 902
rect 766 846 771 902
rect 705 808 771 846
rect 2261 902 2327 940
rect 2261 846 2266 902
rect 2322 846 2327 902
rect 2261 808 2327 846
rect 3817 902 3883 940
rect 3817 846 3822 902
rect 3878 846 3883 902
rect 3817 808 3883 846
rect 5373 902 5439 940
rect 5373 846 5378 902
rect 5434 846 5439 902
rect 5373 808 5439 846
rect 6929 902 6995 940
rect 6929 846 6934 902
rect 6990 846 6995 902
rect 6929 808 6995 846
rect 8485 902 8551 940
rect 8485 846 8490 902
rect 8546 846 8551 902
rect 8485 808 8551 846
rect 10041 902 10107 940
rect 10041 846 10046 902
rect 10102 846 10107 902
rect 10041 808 10107 846
rect 11597 902 11663 940
rect 11597 846 11602 902
rect 11658 846 11663 902
rect 11597 808 11663 846
rect 13153 902 13219 940
rect 13153 846 13158 902
rect 13214 846 13219 902
rect 13153 808 13219 846
rect 14709 902 14775 940
rect 14709 846 14714 902
rect 14770 846 14775 902
rect 14709 808 14775 846
rect 16265 902 16331 940
rect 16265 846 16270 902
rect 16326 846 16331 902
rect 16265 808 16331 846
rect 17821 902 17887 940
rect 17821 846 17826 902
rect 17882 846 17887 902
rect 17821 808 17887 846
rect 19377 902 19443 940
rect 19377 846 19382 902
rect 19438 846 19443 902
rect 19377 808 19443 846
rect 20933 902 20999 940
rect 20933 846 20938 902
rect 20994 846 20999 902
rect 20933 808 20999 846
rect 22489 902 22555 940
rect 22489 846 22494 902
rect 22550 846 22555 902
rect 22489 808 22555 846
rect 24045 902 24111 940
rect 24045 846 24050 902
rect 24106 846 24111 902
rect 24045 808 24111 846
rect 25601 902 25667 940
rect 25601 846 25606 902
rect 25662 846 25667 902
rect 25601 808 25667 846
rect 27157 902 27223 940
rect 27157 846 27162 902
rect 27218 846 27223 902
rect 27157 808 27223 846
rect 28713 902 28779 940
rect 28713 846 28718 902
rect 28774 846 28779 902
rect 28713 808 28779 846
rect 30269 902 30335 940
rect 30269 846 30274 902
rect 30330 846 30335 902
rect 30269 808 30335 846
rect 31825 902 31891 940
rect 31825 846 31830 902
rect 31886 846 31891 902
rect 31825 808 31891 846
rect 33381 902 33447 940
rect 33381 846 33386 902
rect 33442 846 33447 902
rect 33381 808 33447 846
rect 34937 902 35003 940
rect 34937 846 34942 902
rect 34998 846 35003 902
rect 34937 808 35003 846
rect 36493 902 36559 940
rect 36493 846 36498 902
rect 36554 846 36559 902
rect 36493 808 36559 846
rect 38049 902 38115 940
rect 38049 846 38054 902
rect 38110 846 38115 902
rect 38049 808 38115 846
rect 39605 902 39671 940
rect 39605 846 39610 902
rect 39666 846 39671 902
rect 39605 808 39671 846
rect 41161 902 41227 940
rect 41161 846 41166 902
rect 41222 846 41227 902
rect 41161 808 41227 846
rect 42717 902 42783 940
rect 42717 846 42722 902
rect 42778 846 42783 902
rect 42717 808 42783 846
rect 44273 902 44339 940
rect 44273 846 44278 902
rect 44334 846 44339 902
rect 44273 808 44339 846
rect 45829 902 45895 940
rect 45829 846 45834 902
rect 45890 846 45895 902
rect 45829 808 45895 846
rect 47385 902 47451 940
rect 47385 846 47390 902
rect 47446 846 47451 902
rect 47385 808 47451 846
rect 48941 902 49007 940
rect 48941 846 48946 902
rect 49002 846 49007 902
rect 48941 808 49007 846
rect 705 70 771 108
rect 705 14 710 70
rect 766 14 771 70
rect 705 -24 771 14
rect 2261 70 2327 108
rect 2261 14 2266 70
rect 2322 14 2327 70
rect 2261 -24 2327 14
rect 3817 70 3883 108
rect 3817 14 3822 70
rect 3878 14 3883 70
rect 3817 -24 3883 14
rect 5373 70 5439 108
rect 5373 14 5378 70
rect 5434 14 5439 70
rect 5373 -24 5439 14
rect 6929 70 6995 108
rect 6929 14 6934 70
rect 6990 14 6995 70
rect 6929 -24 6995 14
rect 8485 70 8551 108
rect 8485 14 8490 70
rect 8546 14 8551 70
rect 8485 -24 8551 14
rect 10041 70 10107 108
rect 10041 14 10046 70
rect 10102 14 10107 70
rect 10041 -24 10107 14
rect 11597 70 11663 108
rect 11597 14 11602 70
rect 11658 14 11663 70
rect 11597 -24 11663 14
rect 13153 70 13219 108
rect 13153 14 13158 70
rect 13214 14 13219 70
rect 13153 -24 13219 14
rect 14709 70 14775 108
rect 14709 14 14714 70
rect 14770 14 14775 70
rect 14709 -24 14775 14
rect 16265 70 16331 108
rect 16265 14 16270 70
rect 16326 14 16331 70
rect 16265 -24 16331 14
rect 17821 70 17887 108
rect 17821 14 17826 70
rect 17882 14 17887 70
rect 17821 -24 17887 14
rect 19377 70 19443 108
rect 19377 14 19382 70
rect 19438 14 19443 70
rect 19377 -24 19443 14
rect 20933 70 20999 108
rect 20933 14 20938 70
rect 20994 14 20999 70
rect 20933 -24 20999 14
rect 22489 70 22555 108
rect 22489 14 22494 70
rect 22550 14 22555 70
rect 22489 -24 22555 14
rect 24045 70 24111 108
rect 24045 14 24050 70
rect 24106 14 24111 70
rect 24045 -24 24111 14
rect 25601 70 25667 108
rect 25601 14 25606 70
rect 25662 14 25667 70
rect 25601 -24 25667 14
rect 27157 70 27223 108
rect 27157 14 27162 70
rect 27218 14 27223 70
rect 27157 -24 27223 14
rect 28713 70 28779 108
rect 28713 14 28718 70
rect 28774 14 28779 70
rect 28713 -24 28779 14
rect 30269 70 30335 108
rect 30269 14 30274 70
rect 30330 14 30335 70
rect 30269 -24 30335 14
rect 31825 70 31891 108
rect 31825 14 31830 70
rect 31886 14 31891 70
rect 31825 -24 31891 14
rect 33381 70 33447 108
rect 33381 14 33386 70
rect 33442 14 33447 70
rect 33381 -24 33447 14
rect 34937 70 35003 108
rect 34937 14 34942 70
rect 34998 14 35003 70
rect 34937 -24 35003 14
rect 36493 70 36559 108
rect 36493 14 36498 70
rect 36554 14 36559 70
rect 36493 -24 36559 14
rect 38049 70 38115 108
rect 38049 14 38054 70
rect 38110 14 38115 70
rect 38049 -24 38115 14
rect 39605 70 39671 108
rect 39605 14 39610 70
rect 39666 14 39671 70
rect 39605 -24 39671 14
rect 41161 70 41227 108
rect 41161 14 41166 70
rect 41222 14 41227 70
rect 41161 -24 41227 14
rect 42717 70 42783 108
rect 42717 14 42722 70
rect 42778 14 42783 70
rect 42717 -24 42783 14
rect 44273 70 44339 108
rect 44273 14 44278 70
rect 44334 14 44339 70
rect 44273 -24 44339 14
rect 45829 70 45895 108
rect 45829 14 45834 70
rect 45890 14 45895 70
rect 45829 -24 45895 14
rect 47385 70 47451 108
rect 47385 14 47390 70
rect 47446 14 47451 70
rect 47385 -24 47451 14
rect 48941 70 49007 108
rect 48941 14 48946 70
rect 49002 14 49007 70
rect 48941 -24 49007 14
use contact_23  contact_23_0
timestamp 1644969367
transform 1 0 48941 0 1 -24
box 0 0 1 1
use contact_22  contact_22_0
timestamp 1644969367
transform 1 0 48948 0 1 10
box 0 0 1 1
use contact_23  contact_23_1
timestamp 1644969367
transform 1 0 48941 0 1 808
box 0 0 1 1
use contact_22  contact_22_1
timestamp 1644969367
transform 1 0 48948 0 1 842
box 0 0 1 1
use contact_23  contact_23_2
timestamp 1644969367
transform 1 0 47385 0 1 -24
box 0 0 1 1
use contact_22  contact_22_2
timestamp 1644969367
transform 1 0 47392 0 1 10
box 0 0 1 1
use contact_23  contact_23_3
timestamp 1644969367
transform 1 0 47385 0 1 808
box 0 0 1 1
use contact_22  contact_22_3
timestamp 1644969367
transform 1 0 47392 0 1 842
box 0 0 1 1
use contact_23  contact_23_4
timestamp 1644969367
transform 1 0 45829 0 1 -24
box 0 0 1 1
use contact_22  contact_22_4
timestamp 1644969367
transform 1 0 45836 0 1 10
box 0 0 1 1
use contact_23  contact_23_5
timestamp 1644969367
transform 1 0 45829 0 1 808
box 0 0 1 1
use contact_22  contact_22_5
timestamp 1644969367
transform 1 0 45836 0 1 842
box 0 0 1 1
use contact_23  contact_23_6
timestamp 1644969367
transform 1 0 44273 0 1 -24
box 0 0 1 1
use contact_22  contact_22_6
timestamp 1644969367
transform 1 0 44280 0 1 10
box 0 0 1 1
use contact_23  contact_23_7
timestamp 1644969367
transform 1 0 44273 0 1 808
box 0 0 1 1
use contact_22  contact_22_7
timestamp 1644969367
transform 1 0 44280 0 1 842
box 0 0 1 1
use contact_23  contact_23_8
timestamp 1644969367
transform 1 0 42717 0 1 -24
box 0 0 1 1
use contact_22  contact_22_8
timestamp 1644969367
transform 1 0 42724 0 1 10
box 0 0 1 1
use contact_23  contact_23_9
timestamp 1644969367
transform 1 0 42717 0 1 808
box 0 0 1 1
use contact_22  contact_22_9
timestamp 1644969367
transform 1 0 42724 0 1 842
box 0 0 1 1
use contact_23  contact_23_10
timestamp 1644969367
transform 1 0 41161 0 1 -24
box 0 0 1 1
use contact_22  contact_22_10
timestamp 1644969367
transform 1 0 41168 0 1 10
box 0 0 1 1
use contact_23  contact_23_11
timestamp 1644969367
transform 1 0 41161 0 1 808
box 0 0 1 1
use contact_22  contact_22_11
timestamp 1644969367
transform 1 0 41168 0 1 842
box 0 0 1 1
use contact_23  contact_23_12
timestamp 1644969367
transform 1 0 39605 0 1 -24
box 0 0 1 1
use contact_22  contact_22_12
timestamp 1644969367
transform 1 0 39612 0 1 10
box 0 0 1 1
use contact_23  contact_23_13
timestamp 1644969367
transform 1 0 39605 0 1 808
box 0 0 1 1
use contact_22  contact_22_13
timestamp 1644969367
transform 1 0 39612 0 1 842
box 0 0 1 1
use contact_23  contact_23_14
timestamp 1644969367
transform 1 0 38049 0 1 -24
box 0 0 1 1
use contact_22  contact_22_14
timestamp 1644969367
transform 1 0 38056 0 1 10
box 0 0 1 1
use contact_23  contact_23_15
timestamp 1644969367
transform 1 0 38049 0 1 808
box 0 0 1 1
use contact_22  contact_22_15
timestamp 1644969367
transform 1 0 38056 0 1 842
box 0 0 1 1
use contact_23  contact_23_16
timestamp 1644969367
transform 1 0 36493 0 1 -24
box 0 0 1 1
use contact_22  contact_22_16
timestamp 1644969367
transform 1 0 36500 0 1 10
box 0 0 1 1
use contact_23  contact_23_17
timestamp 1644969367
transform 1 0 36493 0 1 808
box 0 0 1 1
use contact_22  contact_22_17
timestamp 1644969367
transform 1 0 36500 0 1 842
box 0 0 1 1
use contact_23  contact_23_18
timestamp 1644969367
transform 1 0 34937 0 1 -24
box 0 0 1 1
use contact_22  contact_22_18
timestamp 1644969367
transform 1 0 34944 0 1 10
box 0 0 1 1
use contact_23  contact_23_19
timestamp 1644969367
transform 1 0 34937 0 1 808
box 0 0 1 1
use contact_22  contact_22_19
timestamp 1644969367
transform 1 0 34944 0 1 842
box 0 0 1 1
use contact_23  contact_23_20
timestamp 1644969367
transform 1 0 33381 0 1 -24
box 0 0 1 1
use contact_22  contact_22_20
timestamp 1644969367
transform 1 0 33388 0 1 10
box 0 0 1 1
use contact_23  contact_23_21
timestamp 1644969367
transform 1 0 33381 0 1 808
box 0 0 1 1
use contact_22  contact_22_21
timestamp 1644969367
transform 1 0 33388 0 1 842
box 0 0 1 1
use contact_23  contact_23_22
timestamp 1644969367
transform 1 0 31825 0 1 -24
box 0 0 1 1
use contact_22  contact_22_22
timestamp 1644969367
transform 1 0 31832 0 1 10
box 0 0 1 1
use contact_23  contact_23_23
timestamp 1644969367
transform 1 0 31825 0 1 808
box 0 0 1 1
use contact_22  contact_22_23
timestamp 1644969367
transform 1 0 31832 0 1 842
box 0 0 1 1
use contact_23  contact_23_24
timestamp 1644969367
transform 1 0 30269 0 1 -24
box 0 0 1 1
use contact_22  contact_22_24
timestamp 1644969367
transform 1 0 30276 0 1 10
box 0 0 1 1
use contact_23  contact_23_25
timestamp 1644969367
transform 1 0 30269 0 1 808
box 0 0 1 1
use contact_22  contact_22_25
timestamp 1644969367
transform 1 0 30276 0 1 842
box 0 0 1 1
use contact_23  contact_23_26
timestamp 1644969367
transform 1 0 28713 0 1 -24
box 0 0 1 1
use contact_22  contact_22_26
timestamp 1644969367
transform 1 0 28720 0 1 10
box 0 0 1 1
use contact_23  contact_23_27
timestamp 1644969367
transform 1 0 28713 0 1 808
box 0 0 1 1
use contact_22  contact_22_27
timestamp 1644969367
transform 1 0 28720 0 1 842
box 0 0 1 1
use contact_23  contact_23_28
timestamp 1644969367
transform 1 0 27157 0 1 -24
box 0 0 1 1
use contact_22  contact_22_28
timestamp 1644969367
transform 1 0 27164 0 1 10
box 0 0 1 1
use contact_23  contact_23_29
timestamp 1644969367
transform 1 0 27157 0 1 808
box 0 0 1 1
use contact_22  contact_22_29
timestamp 1644969367
transform 1 0 27164 0 1 842
box 0 0 1 1
use contact_23  contact_23_30
timestamp 1644969367
transform 1 0 25601 0 1 -24
box 0 0 1 1
use contact_22  contact_22_30
timestamp 1644969367
transform 1 0 25608 0 1 10
box 0 0 1 1
use contact_23  contact_23_31
timestamp 1644969367
transform 1 0 25601 0 1 808
box 0 0 1 1
use contact_22  contact_22_31
timestamp 1644969367
transform 1 0 25608 0 1 842
box 0 0 1 1
use contact_23  contact_23_32
timestamp 1644969367
transform 1 0 24045 0 1 -24
box 0 0 1 1
use contact_22  contact_22_32
timestamp 1644969367
transform 1 0 24052 0 1 10
box 0 0 1 1
use contact_23  contact_23_33
timestamp 1644969367
transform 1 0 24045 0 1 808
box 0 0 1 1
use contact_22  contact_22_33
timestamp 1644969367
transform 1 0 24052 0 1 842
box 0 0 1 1
use contact_23  contact_23_34
timestamp 1644969367
transform 1 0 22489 0 1 -24
box 0 0 1 1
use contact_22  contact_22_34
timestamp 1644969367
transform 1 0 22496 0 1 10
box 0 0 1 1
use contact_23  contact_23_35
timestamp 1644969367
transform 1 0 22489 0 1 808
box 0 0 1 1
use contact_22  contact_22_35
timestamp 1644969367
transform 1 0 22496 0 1 842
box 0 0 1 1
use contact_23  contact_23_36
timestamp 1644969367
transform 1 0 20933 0 1 -24
box 0 0 1 1
use contact_22  contact_22_36
timestamp 1644969367
transform 1 0 20940 0 1 10
box 0 0 1 1
use contact_23  contact_23_37
timestamp 1644969367
transform 1 0 20933 0 1 808
box 0 0 1 1
use contact_22  contact_22_37
timestamp 1644969367
transform 1 0 20940 0 1 842
box 0 0 1 1
use contact_23  contact_23_38
timestamp 1644969367
transform 1 0 19377 0 1 -24
box 0 0 1 1
use contact_22  contact_22_38
timestamp 1644969367
transform 1 0 19384 0 1 10
box 0 0 1 1
use contact_23  contact_23_39
timestamp 1644969367
transform 1 0 19377 0 1 808
box 0 0 1 1
use contact_22  contact_22_39
timestamp 1644969367
transform 1 0 19384 0 1 842
box 0 0 1 1
use contact_23  contact_23_40
timestamp 1644969367
transform 1 0 17821 0 1 -24
box 0 0 1 1
use contact_22  contact_22_40
timestamp 1644969367
transform 1 0 17828 0 1 10
box 0 0 1 1
use contact_23  contact_23_41
timestamp 1644969367
transform 1 0 17821 0 1 808
box 0 0 1 1
use contact_22  contact_22_41
timestamp 1644969367
transform 1 0 17828 0 1 842
box 0 0 1 1
use contact_23  contact_23_42
timestamp 1644969367
transform 1 0 16265 0 1 -24
box 0 0 1 1
use contact_22  contact_22_42
timestamp 1644969367
transform 1 0 16272 0 1 10
box 0 0 1 1
use contact_23  contact_23_43
timestamp 1644969367
transform 1 0 16265 0 1 808
box 0 0 1 1
use contact_22  contact_22_43
timestamp 1644969367
transform 1 0 16272 0 1 842
box 0 0 1 1
use contact_23  contact_23_44
timestamp 1644969367
transform 1 0 14709 0 1 -24
box 0 0 1 1
use contact_22  contact_22_44
timestamp 1644969367
transform 1 0 14716 0 1 10
box 0 0 1 1
use contact_23  contact_23_45
timestamp 1644969367
transform 1 0 14709 0 1 808
box 0 0 1 1
use contact_22  contact_22_45
timestamp 1644969367
transform 1 0 14716 0 1 842
box 0 0 1 1
use contact_23  contact_23_46
timestamp 1644969367
transform 1 0 13153 0 1 -24
box 0 0 1 1
use contact_22  contact_22_46
timestamp 1644969367
transform 1 0 13160 0 1 10
box 0 0 1 1
use contact_23  contact_23_47
timestamp 1644969367
transform 1 0 13153 0 1 808
box 0 0 1 1
use contact_22  contact_22_47
timestamp 1644969367
transform 1 0 13160 0 1 842
box 0 0 1 1
use contact_23  contact_23_48
timestamp 1644969367
transform 1 0 11597 0 1 -24
box 0 0 1 1
use contact_22  contact_22_48
timestamp 1644969367
transform 1 0 11604 0 1 10
box 0 0 1 1
use contact_23  contact_23_49
timestamp 1644969367
transform 1 0 11597 0 1 808
box 0 0 1 1
use contact_22  contact_22_49
timestamp 1644969367
transform 1 0 11604 0 1 842
box 0 0 1 1
use contact_23  contact_23_50
timestamp 1644969367
transform 1 0 10041 0 1 -24
box 0 0 1 1
use contact_22  contact_22_50
timestamp 1644969367
transform 1 0 10048 0 1 10
box 0 0 1 1
use contact_23  contact_23_51
timestamp 1644969367
transform 1 0 10041 0 1 808
box 0 0 1 1
use contact_22  contact_22_51
timestamp 1644969367
transform 1 0 10048 0 1 842
box 0 0 1 1
use contact_23  contact_23_52
timestamp 1644969367
transform 1 0 8485 0 1 -24
box 0 0 1 1
use contact_22  contact_22_52
timestamp 1644969367
transform 1 0 8492 0 1 10
box 0 0 1 1
use contact_23  contact_23_53
timestamp 1644969367
transform 1 0 8485 0 1 808
box 0 0 1 1
use contact_22  contact_22_53
timestamp 1644969367
transform 1 0 8492 0 1 842
box 0 0 1 1
use contact_23  contact_23_54
timestamp 1644969367
transform 1 0 6929 0 1 -24
box 0 0 1 1
use contact_22  contact_22_54
timestamp 1644969367
transform 1 0 6936 0 1 10
box 0 0 1 1
use contact_23  contact_23_55
timestamp 1644969367
transform 1 0 6929 0 1 808
box 0 0 1 1
use contact_22  contact_22_55
timestamp 1644969367
transform 1 0 6936 0 1 842
box 0 0 1 1
use contact_23  contact_23_56
timestamp 1644969367
transform 1 0 5373 0 1 -24
box 0 0 1 1
use contact_22  contact_22_56
timestamp 1644969367
transform 1 0 5380 0 1 10
box 0 0 1 1
use contact_23  contact_23_57
timestamp 1644969367
transform 1 0 5373 0 1 808
box 0 0 1 1
use contact_22  contact_22_57
timestamp 1644969367
transform 1 0 5380 0 1 842
box 0 0 1 1
use contact_23  contact_23_58
timestamp 1644969367
transform 1 0 3817 0 1 -24
box 0 0 1 1
use contact_22  contact_22_58
timestamp 1644969367
transform 1 0 3824 0 1 10
box 0 0 1 1
use contact_23  contact_23_59
timestamp 1644969367
transform 1 0 3817 0 1 808
box 0 0 1 1
use contact_22  contact_22_59
timestamp 1644969367
transform 1 0 3824 0 1 842
box 0 0 1 1
use contact_23  contact_23_60
timestamp 1644969367
transform 1 0 2261 0 1 -24
box 0 0 1 1
use contact_22  contact_22_60
timestamp 1644969367
transform 1 0 2268 0 1 10
box 0 0 1 1
use contact_23  contact_23_61
timestamp 1644969367
transform 1 0 2261 0 1 808
box 0 0 1 1
use contact_22  contact_22_61
timestamp 1644969367
transform 1 0 2268 0 1 842
box 0 0 1 1
use contact_23  contact_23_62
timestamp 1644969367
transform 1 0 705 0 1 -24
box 0 0 1 1
use contact_22  contact_22_62
timestamp 1644969367
transform 1 0 712 0 1 10
box 0 0 1 1
use contact_23  contact_23_63
timestamp 1644969367
transform 1 0 705 0 1 808
box 0 0 1 1
use contact_22  contact_22_63
timestamp 1644969367
transform 1 0 712 0 1 842
box 0 0 1 1
use write_driver_multiport  write_driver_multiport_0
timestamp 1644969367
transform 1 0 48625 0 1 0
box 0 0 698 952
use write_driver_multiport  write_driver_multiport_1
timestamp 1644969367
transform 1 0 47069 0 1 0
box 0 0 698 952
use write_driver_multiport  write_driver_multiport_2
timestamp 1644969367
transform 1 0 45513 0 1 0
box 0 0 698 952
use write_driver_multiport  write_driver_multiport_3
timestamp 1644969367
transform 1 0 43957 0 1 0
box 0 0 698 952
use write_driver_multiport  write_driver_multiport_4
timestamp 1644969367
transform 1 0 42401 0 1 0
box 0 0 698 952
use write_driver_multiport  write_driver_multiport_5
timestamp 1644969367
transform 1 0 40845 0 1 0
box 0 0 698 952
use write_driver_multiport  write_driver_multiport_6
timestamp 1644969367
transform 1 0 39289 0 1 0
box 0 0 698 952
use write_driver_multiport  write_driver_multiport_7
timestamp 1644969367
transform 1 0 37733 0 1 0
box 0 0 698 952
use write_driver_multiport  write_driver_multiport_8
timestamp 1644969367
transform 1 0 36177 0 1 0
box 0 0 698 952
use write_driver_multiport  write_driver_multiport_9
timestamp 1644969367
transform 1 0 34621 0 1 0
box 0 0 698 952
use write_driver_multiport  write_driver_multiport_10
timestamp 1644969367
transform 1 0 33065 0 1 0
box 0 0 698 952
use write_driver_multiport  write_driver_multiport_11
timestamp 1644969367
transform 1 0 31509 0 1 0
box 0 0 698 952
use write_driver_multiport  write_driver_multiport_12
timestamp 1644969367
transform 1 0 29953 0 1 0
box 0 0 698 952
use write_driver_multiport  write_driver_multiport_13
timestamp 1644969367
transform 1 0 28397 0 1 0
box 0 0 698 952
use write_driver_multiport  write_driver_multiport_14
timestamp 1644969367
transform 1 0 26841 0 1 0
box 0 0 698 952
use write_driver_multiport  write_driver_multiport_15
timestamp 1644969367
transform 1 0 25285 0 1 0
box 0 0 698 952
use write_driver_multiport  write_driver_multiport_16
timestamp 1644969367
transform 1 0 23729 0 1 0
box 0 0 698 952
use write_driver_multiport  write_driver_multiport_17
timestamp 1644969367
transform 1 0 22173 0 1 0
box 0 0 698 952
use write_driver_multiport  write_driver_multiport_18
timestamp 1644969367
transform 1 0 20617 0 1 0
box 0 0 698 952
use write_driver_multiport  write_driver_multiport_19
timestamp 1644969367
transform 1 0 19061 0 1 0
box 0 0 698 952
use write_driver_multiport  write_driver_multiport_20
timestamp 1644969367
transform 1 0 17505 0 1 0
box 0 0 698 952
use write_driver_multiport  write_driver_multiport_21
timestamp 1644969367
transform 1 0 15949 0 1 0
box 0 0 698 952
use write_driver_multiport  write_driver_multiport_22
timestamp 1644969367
transform 1 0 14393 0 1 0
box 0 0 698 952
use write_driver_multiport  write_driver_multiport_23
timestamp 1644969367
transform 1 0 12837 0 1 0
box 0 0 698 952
use write_driver_multiport  write_driver_multiport_24
timestamp 1644969367
transform 1 0 11281 0 1 0
box 0 0 698 952
use write_driver_multiport  write_driver_multiport_25
timestamp 1644969367
transform 1 0 9725 0 1 0
box 0 0 698 952
use write_driver_multiport  write_driver_multiport_26
timestamp 1644969367
transform 1 0 8169 0 1 0
box 0 0 698 952
use write_driver_multiport  write_driver_multiport_27
timestamp 1644969367
transform 1 0 6613 0 1 0
box 0 0 698 952
use write_driver_multiport  write_driver_multiport_28
timestamp 1644969367
transform 1 0 5057 0 1 0
box 0 0 698 952
use write_driver_multiport  write_driver_multiport_29
timestamp 1644969367
transform 1 0 3501 0 1 0
box 0 0 698 952
use write_driver_multiport  write_driver_multiport_30
timestamp 1644969367
transform 1 0 1945 0 1 0
box 0 0 698 952
use write_driver_multiport  write_driver_multiport_31
timestamp 1644969367
transform 1 0 389 0 1 0
box 0 0 698 952
<< labels >>
rlabel metal2 s 585 272 639 300 4 din_0
rlabel metal2 s 1019 322 1047 952 4 wbl0_0
rlabel metal3 s 17821 808 17887 940 4 vdd
rlabel metal3 s 25601 808 25667 940 4 vdd
rlabel metal3 s 30269 808 30335 940 4 vdd
rlabel metal3 s 16265 808 16331 940 4 vdd
rlabel metal3 s 705 808 771 940 4 vdd
rlabel metal3 s 47385 808 47451 940 4 vdd
rlabel metal3 s 38049 808 38115 940 4 vdd
rlabel metal3 s 28713 808 28779 940 4 vdd
rlabel metal3 s 13153 808 13219 940 4 vdd
rlabel metal3 s 45829 808 45895 940 4 vdd
rlabel metal3 s 3817 808 3883 940 4 vdd
rlabel metal3 s 11597 808 11663 940 4 vdd
rlabel metal3 s 36493 808 36559 940 4 vdd
rlabel metal3 s 44273 808 44339 940 4 vdd
rlabel metal3 s 19377 808 19443 940 4 vdd
rlabel metal3 s 10041 808 10107 940 4 vdd
rlabel metal3 s 14709 808 14775 940 4 vdd
rlabel metal3 s 33381 808 33447 940 4 vdd
rlabel metal3 s 6929 808 6995 940 4 vdd
rlabel metal3 s 39605 808 39671 940 4 vdd
rlabel metal3 s 5373 808 5439 940 4 vdd
rlabel metal3 s 20933 808 20999 940 4 vdd
rlabel metal3 s 24045 808 24111 940 4 vdd
rlabel metal3 s 34937 808 35003 940 4 vdd
rlabel metal3 s 31825 808 31891 940 4 vdd
rlabel metal3 s 42717 808 42783 940 4 vdd
rlabel metal3 s 48941 808 49007 940 4 vdd
rlabel metal3 s 8485 808 8551 940 4 vdd
rlabel metal3 s 27157 808 27223 940 4 vdd
rlabel metal3 s 22489 808 22555 940 4 vdd
rlabel metal3 s 41161 808 41227 940 4 vdd
rlabel metal3 s 2261 808 2327 940 4 vdd
rlabel metal3 s 38049 -24 38115 108 4 gnd
rlabel metal3 s 8485 -24 8551 108 4 gnd
rlabel metal3 s 42717 -24 42783 108 4 gnd
rlabel metal3 s 24045 -24 24111 108 4 gnd
rlabel metal3 s 11597 -24 11663 108 4 gnd
rlabel metal3 s 10041 -24 10107 108 4 gnd
rlabel metal3 s 33381 -24 33447 108 4 gnd
rlabel metal3 s 39605 -24 39671 108 4 gnd
rlabel metal3 s 5373 -24 5439 108 4 gnd
rlabel metal3 s 25601 -24 25667 108 4 gnd
rlabel metal3 s 6929 -24 6995 108 4 gnd
rlabel metal3 s 20933 -24 20999 108 4 gnd
rlabel metal3 s 3817 -24 3883 108 4 gnd
rlabel metal3 s 27157 -24 27223 108 4 gnd
rlabel metal3 s 34937 -24 35003 108 4 gnd
rlabel metal3 s 13153 -24 13219 108 4 gnd
rlabel metal3 s 14709 -24 14775 108 4 gnd
rlabel metal3 s 22489 -24 22555 108 4 gnd
rlabel metal3 s 16265 -24 16331 108 4 gnd
rlabel metal3 s 28713 -24 28779 108 4 gnd
rlabel metal3 s 705 -24 771 108 4 gnd
rlabel metal3 s 45829 -24 45895 108 4 gnd
rlabel metal3 s 31825 -24 31891 108 4 gnd
rlabel metal3 s 2261 -24 2327 108 4 gnd
rlabel metal3 s 48941 -24 49007 108 4 gnd
rlabel metal3 s 44273 -24 44339 108 4 gnd
rlabel metal3 s 36493 -24 36559 108 4 gnd
rlabel metal3 s 47385 -24 47451 108 4 gnd
rlabel metal3 s 30269 -24 30335 108 4 gnd
rlabel metal3 s 17821 -24 17887 108 4 gnd
rlabel metal3 s 19377 -24 19443 108 4 gnd
rlabel metal3 s 41161 -24 41227 108 4 gnd
rlabel metal2 s 2141 272 2195 300 4 din_1
rlabel metal2 s 2575 322 2603 952 4 wbl0_1
rlabel metal2 s 3697 272 3751 300 4 din_2
rlabel metal2 s 4131 322 4159 952 4 wbl0_2
rlabel metal2 s 5253 272 5307 300 4 din_3
rlabel metal2 s 5687 322 5715 952 4 wbl0_3
rlabel metal2 s 6809 272 6863 300 4 din_4
rlabel metal2 s 7243 322 7271 952 4 wbl0_4
rlabel metal2 s 8365 272 8419 300 4 din_5
rlabel metal2 s 8799 322 8827 952 4 wbl0_5
rlabel metal2 s 9921 272 9975 300 4 din_6
rlabel metal2 s 10355 322 10383 952 4 wbl0_6
rlabel metal2 s 11477 272 11531 300 4 din_7
rlabel metal2 s 11911 322 11939 952 4 wbl0_7
rlabel metal2 s 13033 272 13087 300 4 din_8
rlabel metal2 s 13467 322 13495 952 4 wbl0_8
rlabel metal2 s 14589 272 14643 300 4 din_9
rlabel metal2 s 15023 322 15051 952 4 wbl0_9
rlabel metal2 s 16145 272 16199 300 4 din_10
rlabel metal2 s 16579 322 16607 952 4 wbl0_10
rlabel metal2 s 17701 272 17755 300 4 din_11
rlabel metal2 s 18135 322 18163 952 4 wbl0_11
rlabel metal2 s 19257 272 19311 300 4 din_12
rlabel metal2 s 19691 322 19719 952 4 wbl0_12
rlabel metal2 s 20813 272 20867 300 4 din_13
rlabel metal2 s 21247 322 21275 952 4 wbl0_13
rlabel metal2 s 22369 272 22423 300 4 din_14
rlabel metal2 s 22803 322 22831 952 4 wbl0_14
rlabel metal2 s 23925 272 23979 300 4 din_15
rlabel metal2 s 24359 322 24387 952 4 wbl0_15
rlabel metal2 s 25481 272 25535 300 4 din_16
rlabel metal2 s 25915 322 25943 952 4 wbl0_16
rlabel metal2 s 27037 272 27091 300 4 din_17
rlabel metal2 s 27471 322 27499 952 4 wbl0_17
rlabel metal2 s 28593 272 28647 300 4 din_18
rlabel metal2 s 29027 322 29055 952 4 wbl0_18
rlabel metal2 s 30149 272 30203 300 4 din_19
rlabel metal2 s 30583 322 30611 952 4 wbl0_19
rlabel metal2 s 31705 272 31759 300 4 din_20
rlabel metal2 s 32139 322 32167 952 4 wbl0_20
rlabel metal2 s 33261 272 33315 300 4 din_21
rlabel metal2 s 33695 322 33723 952 4 wbl0_21
rlabel metal2 s 34817 272 34871 300 4 din_22
rlabel metal2 s 35251 322 35279 952 4 wbl0_22
rlabel metal2 s 36373 272 36427 300 4 din_23
rlabel metal2 s 36807 322 36835 952 4 wbl0_23
rlabel metal2 s 37929 272 37983 300 4 din_24
rlabel metal2 s 38363 322 38391 952 4 wbl0_24
rlabel metal2 s 39485 272 39539 300 4 din_25
rlabel metal2 s 39919 322 39947 952 4 wbl0_25
rlabel metal2 s 41041 272 41095 300 4 din_26
rlabel metal2 s 41475 322 41503 952 4 wbl0_26
rlabel metal2 s 42597 272 42651 300 4 din_27
rlabel metal2 s 43031 322 43059 952 4 wbl0_27
rlabel metal2 s 44153 272 44207 300 4 din_28
rlabel metal2 s 44587 322 44615 952 4 wbl0_28
rlabel metal2 s 45709 272 45763 300 4 din_29
rlabel metal2 s 46143 322 46171 952 4 wbl0_29
rlabel metal2 s 47265 272 47319 300 4 din_30
rlabel metal2 s 47699 322 47727 952 4 wbl0_30
rlabel metal2 s 48821 272 48875 300 4 din_31
rlabel metal2 s 49255 322 49283 952 4 wbl0_31
rlabel metal1 s 0 356 49323 384 4 en
<< properties >>
string FIXED_BBOX 48941 -24 49007 0
string GDS_FILE sram_0rw2r1w_32_128_sky130A.gds
string GDS_END 2637974
string GDS_START 2602798
<< end >>
