magic
tech sky130A
magscale 1 2
timestamp 1643678851
<< checkpaint >>
rect -1227 -1260 2104 2768
<< pwell >>
rect 753 718 803 800
<< psubdiff >>
rect 753 776 803 800
rect 753 742 761 776
rect 795 742 803 776
rect 753 718 803 742
<< psubdiffcont >>
rect 761 742 795 776
<< poly >>
rect 374 726 404 780
rect 374 28 404 54
<< locali >>
rect 99 1435 456 1469
rect 422 1116 456 1435
rect 761 776 795 792
rect 761 726 795 742
rect 322 73 356 390
rect 322 39 707 73
<< viali >>
rect 65 1435 99 1469
rect 322 1099 356 1133
rect 761 742 795 776
rect 422 373 456 407
rect 707 39 741 73
<< metal1 >>
rect 53 1469 56 1475
rect 108 1469 111 1475
rect 33 1435 56 1469
rect 108 1435 131 1469
rect 53 1429 56 1435
rect 108 1429 111 1435
rect 310 1133 368 1139
rect 310 1099 322 1133
rect 356 1099 368 1133
rect 310 1093 368 1099
rect 325 470 353 1093
rect 710 952 738 1452
rect 68 442 353 470
rect 425 924 738 952
rect 68 56 96 442
rect 425 413 453 924
rect 749 736 752 782
rect 804 736 807 782
rect 410 407 468 413
rect 410 373 422 407
rect 456 373 468 407
rect 410 367 468 373
rect 695 73 698 79
rect 750 73 753 79
rect 675 39 698 73
rect 750 39 773 73
rect 695 33 698 39
rect 750 33 753 39
<< via1 >>
rect 56 1469 108 1478
rect 56 1435 65 1469
rect 65 1435 99 1469
rect 99 1435 108 1469
rect 56 1426 108 1435
rect 752 776 804 785
rect 752 742 761 776
rect 761 742 795 776
rect 795 742 804 776
rect 752 733 804 742
rect 698 73 750 82
rect 698 39 707 73
rect 707 39 741 73
rect 741 39 750 73
rect 698 30 750 39
<< metal2 >>
rect 68 1478 96 1508
rect 710 1452 738 1508
rect 758 787 798 793
rect 758 725 798 731
rect 68 0 96 56
rect 710 0 738 30
<< via2 >>
rect 750 785 806 787
rect 750 733 752 785
rect 752 733 804 785
rect 804 733 806 785
rect 750 731 806 733
<< metal3 >>
rect 712 787 844 792
rect 712 731 750 787
rect 806 731 844 787
rect 712 726 844 731
use contact_18  contact_18_0
timestamp 1643678851
transform 1 0 712 0 1 726
box 0 0 1 1
use contact_17  contact_17_0
timestamp 1643678851
transform 1 0 763 0 1 744
box 0 0 1 1
use contact_13  contact_13_0
timestamp 1643678851
transform 1 0 749 0 1 736
box 0 0 1 1
use contact_25  contact_25_0
timestamp 1643678851
transform 1 0 753 0 1 718
box 0 0 1 1
use contact_13  contact_13_1
timestamp 1643678851
transform 1 0 410 0 1 367
box 0 0 1 1
use contact_13  contact_13_2
timestamp 1643678851
transform 1 0 310 0 1 1093
box 0 0 1 1
use contact_13  contact_13_3
timestamp 1643678851
transform 1 0 695 0 1 33
box 0 0 1 1
use contact_17  contact_17_1
timestamp 1643678851
transform 1 0 709 0 1 41
box 0 0 1 1
use contact_13  contact_13_4
timestamp 1643678851
transform 1 0 53 0 1 1429
box 0 0 1 1
use contact_17  contact_17_2
timestamp 1643678851
transform 1 0 67 0 1 1437
box 0 0 1 1
use nmos_m1_w3_360_sli_dli  nmos_m1_w3_360_sli_dli_0
timestamp 1643678851
transform 1 0 314 0 1 780
box 0 -26 150 698
use nmos_m1_w3_360_sli_dli  nmos_m1_w3_360_sli_dli_1
timestamp 1643678851
transform 1 0 314 0 1 54
box 0 -26 150 698
<< labels >>
rlabel mvvaractor s 389 41 389 41 4 sel
rlabel metal2 s 68 1452 96 1508 4 rbl0
rlabel metal2 s 710 1452 738 1508 4 rbl1
rlabel metal2 s 68 0 96 56 4 rbl0_out
rlabel metal2 s 710 0 738 56 4 rbl1_out
rlabel metal3 s 712 726 844 792 4 gnd
<< properties >>
string FIXED_BBOX 0 0 778 693
string GDS_FILE sram_0rw2r1w_16_128_sky130A.gds
string GDS_END 1625874
string GDS_START 1622898
<< end >>
