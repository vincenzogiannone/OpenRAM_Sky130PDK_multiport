magic
tech sky130A
magscale 1 2
timestamp 1644949024
<< checkpaint >>
rect -1296 -1277 5036 2155
<< nwell >>
rect -36 402 3776 895
<< locali >>
rect 0 821 3740 855
rect 48 344 114 410
rect 196 360 449 394
rect 568 360 925 394
rect 1243 354 1833 388
rect 2691 354 2725 388
rect 0 -17 3740 17
use pinv_8  pinv_8_0
timestamp 1644949024
transform 1 0 1752 0 1 0
box -36 -17 2024 895
use pinv_7  pinv_7_0
timestamp 1644949024
transform 1 0 844 0 1 0
box -36 -17 944 895
use pinv_6  pinv_6_0
timestamp 1644949024
transform 1 0 368 0 1 0
box -36 -17 512 895
use pinv_5  pinv_5_0
timestamp 1644949024
transform 1 0 0 0 1 0
box -36 -17 404 895
<< labels >>
rlabel locali s 2708 371 2708 371 4 Z
rlabel locali s 81 377 81 377 4 A
rlabel locali s 1870 0 1870 0 4 gnd
rlabel locali s 1870 838 1870 838 4 vdd
<< properties >>
string FIXED_BBOX 0 0 3740 838
string GDS_FILE sram_0rw2r1w_4_16_sky130A.gds
string GDS_END 465126
string GDS_START 463854
<< end >>
