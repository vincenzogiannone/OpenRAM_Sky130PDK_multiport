magic
tech sky130A
magscale 1 2
timestamp 1644949024
<< checkpaint >>
rect -1260 -1286 1734 1403
<< scnmos >>
rect 60 0 90 84
rect 168 0 198 84
rect 276 0 306 84
rect 384 0 414 84
<< ndiff >>
rect 0 59 60 84
rect 0 25 8 59
rect 42 25 60 59
rect 0 0 60 25
rect 90 59 168 84
rect 90 25 112 59
rect 146 25 168 59
rect 90 0 168 25
rect 198 59 276 84
rect 198 25 220 59
rect 254 25 276 59
rect 198 0 276 25
rect 306 59 384 84
rect 306 25 328 59
rect 362 25 384 59
rect 306 0 384 25
rect 414 59 474 84
rect 414 25 432 59
rect 466 25 474 59
rect 414 0 474 25
<< ndiffc >>
rect 8 25 42 59
rect 112 25 146 59
rect 220 25 254 59
rect 328 25 362 59
rect 432 25 466 59
<< poly >>
rect 60 110 414 140
rect 60 84 90 110
rect 168 84 198 110
rect 276 84 306 110
rect 384 84 414 110
rect 60 -26 90 0
rect 168 -26 198 0
rect 276 -26 306 0
rect 384 -26 414 0
<< locali >>
rect 112 109 362 143
rect 8 59 42 75
rect 8 9 42 25
rect 112 59 146 109
rect 112 9 146 25
rect 220 59 254 75
rect 220 9 254 25
rect 328 59 362 109
rect 328 9 362 25
rect 432 59 466 75
rect 432 9 466 25
use contact_8  contact_8_0
timestamp 1644949024
transform 1 0 424 0 1 1
box 0 0 1 1
use contact_8  contact_8_1
timestamp 1644949024
transform 1 0 320 0 1 1
box 0 0 1 1
use contact_8  contact_8_2
timestamp 1644949024
transform 1 0 212 0 1 1
box 0 0 1 1
use contact_8  contact_8_3
timestamp 1644949024
transform 1 0 104 0 1 1
box 0 0 1 1
use contact_8  contact_8_4
timestamp 1644949024
transform 1 0 0 0 1 1
box 0 0 1 1
<< labels >>
rlabel mvvaractor s 237 125 237 125 4 G
rlabel locali s 449 42 449 42 4 S
rlabel locali s 237 42 237 42 4 S
rlabel locali s 25 42 25 42 4 S
rlabel locali s 237 126 237 126 4 D
<< properties >>
string FIXED_BBOX -25 -26 499 143
string GDS_FILE sram_0rw2r1w_4_16_sky130A.gds
string GDS_END 463812
string GDS_START 462368
<< end >>
