magic
tech sky130A
magscale 1 2
timestamp 1644969367
<< checkpaint >>
rect -1319 -1316 3305 1608
<< nwell >>
rect -54 231 2040 348
rect -59 63 2045 231
rect -54 -54 2040 63
<< scpmos >>
rect 60 0 90 294
rect 168 0 198 294
rect 276 0 306 294
rect 384 0 414 294
rect 492 0 522 294
rect 600 0 630 294
rect 708 0 738 294
rect 816 0 846 294
rect 924 0 954 294
rect 1032 0 1062 294
rect 1140 0 1170 294
rect 1248 0 1278 294
rect 1356 0 1386 294
rect 1464 0 1494 294
rect 1572 0 1602 294
rect 1680 0 1710 294
rect 1788 0 1818 294
rect 1896 0 1926 294
<< pdiff >>
rect 0 164 60 294
rect 0 130 8 164
rect 42 130 60 164
rect 0 0 60 130
rect 90 164 168 294
rect 90 130 112 164
rect 146 130 168 164
rect 90 0 168 130
rect 198 164 276 294
rect 198 130 220 164
rect 254 130 276 164
rect 198 0 276 130
rect 306 164 384 294
rect 306 130 328 164
rect 362 130 384 164
rect 306 0 384 130
rect 414 164 492 294
rect 414 130 436 164
rect 470 130 492 164
rect 414 0 492 130
rect 522 164 600 294
rect 522 130 544 164
rect 578 130 600 164
rect 522 0 600 130
rect 630 164 708 294
rect 630 130 652 164
rect 686 130 708 164
rect 630 0 708 130
rect 738 164 816 294
rect 738 130 760 164
rect 794 130 816 164
rect 738 0 816 130
rect 846 164 924 294
rect 846 130 868 164
rect 902 130 924 164
rect 846 0 924 130
rect 954 164 1032 294
rect 954 130 976 164
rect 1010 130 1032 164
rect 954 0 1032 130
rect 1062 164 1140 294
rect 1062 130 1084 164
rect 1118 130 1140 164
rect 1062 0 1140 130
rect 1170 164 1248 294
rect 1170 130 1192 164
rect 1226 130 1248 164
rect 1170 0 1248 130
rect 1278 164 1356 294
rect 1278 130 1300 164
rect 1334 130 1356 164
rect 1278 0 1356 130
rect 1386 164 1464 294
rect 1386 130 1408 164
rect 1442 130 1464 164
rect 1386 0 1464 130
rect 1494 164 1572 294
rect 1494 130 1516 164
rect 1550 130 1572 164
rect 1494 0 1572 130
rect 1602 164 1680 294
rect 1602 130 1624 164
rect 1658 130 1680 164
rect 1602 0 1680 130
rect 1710 164 1788 294
rect 1710 130 1732 164
rect 1766 130 1788 164
rect 1710 0 1788 130
rect 1818 164 1896 294
rect 1818 130 1840 164
rect 1874 130 1896 164
rect 1818 0 1896 130
rect 1926 164 1986 294
rect 1926 130 1944 164
rect 1978 130 1986 164
rect 1926 0 1986 130
<< pdiffc >>
rect 8 130 42 164
rect 112 130 146 164
rect 220 130 254 164
rect 328 130 362 164
rect 436 130 470 164
rect 544 130 578 164
rect 652 130 686 164
rect 760 130 794 164
rect 868 130 902 164
rect 976 130 1010 164
rect 1084 130 1118 164
rect 1192 130 1226 164
rect 1300 130 1334 164
rect 1408 130 1442 164
rect 1516 130 1550 164
rect 1624 130 1658 164
rect 1732 130 1766 164
rect 1840 130 1874 164
rect 1944 130 1978 164
<< poly >>
rect 60 294 90 320
rect 168 294 198 320
rect 276 294 306 320
rect 384 294 414 320
rect 492 294 522 320
rect 600 294 630 320
rect 708 294 738 320
rect 816 294 846 320
rect 924 294 954 320
rect 1032 294 1062 320
rect 1140 294 1170 320
rect 1248 294 1278 320
rect 1356 294 1386 320
rect 1464 294 1494 320
rect 1572 294 1602 320
rect 1680 294 1710 320
rect 1788 294 1818 320
rect 1896 294 1926 320
rect 60 -26 90 0
rect 168 -26 198 0
rect 276 -26 306 0
rect 384 -26 414 0
rect 492 -26 522 0
rect 600 -26 630 0
rect 708 -26 738 0
rect 816 -26 846 0
rect 924 -26 954 0
rect 1032 -26 1062 0
rect 1140 -26 1170 0
rect 1248 -26 1278 0
rect 1356 -26 1386 0
rect 1464 -26 1494 0
rect 1572 -26 1602 0
rect 1680 -26 1710 0
rect 1788 -26 1818 0
rect 1896 -26 1926 0
rect 60 -56 1926 -26
<< locali >>
rect 8 164 42 180
rect 8 114 42 130
rect 112 164 146 180
rect 112 80 146 130
rect 220 164 254 180
rect 220 114 254 130
rect 328 164 362 180
rect 328 80 362 130
rect 436 164 470 180
rect 436 114 470 130
rect 544 164 578 180
rect 544 80 578 130
rect 652 164 686 180
rect 652 114 686 130
rect 760 164 794 180
rect 760 80 794 130
rect 868 164 902 180
rect 868 114 902 130
rect 976 164 1010 180
rect 976 80 1010 130
rect 1084 164 1118 180
rect 1084 114 1118 130
rect 1192 164 1226 180
rect 1192 80 1226 130
rect 1300 164 1334 180
rect 1300 114 1334 130
rect 1408 164 1442 180
rect 1408 80 1442 130
rect 1516 164 1550 180
rect 1516 114 1550 130
rect 1624 164 1658 180
rect 1624 80 1658 130
rect 1732 164 1766 180
rect 1732 114 1766 130
rect 1840 164 1874 180
rect 1840 80 1874 130
rect 1944 164 1978 180
rect 1944 114 1978 130
rect 112 46 1874 80
use contact_9  contact_9_0
timestamp 1644969367
transform 1 0 1936 0 1 106
box 0 0 2 2
use contact_9  contact_9_1
timestamp 1644969367
transform 1 0 1832 0 1 106
box 0 0 2 2
use contact_9  contact_9_2
timestamp 1644969367
transform 1 0 1724 0 1 106
box 0 0 2 2
use contact_9  contact_9_3
timestamp 1644969367
transform 1 0 1616 0 1 106
box 0 0 2 2
use contact_9  contact_9_4
timestamp 1644969367
transform 1 0 1508 0 1 106
box 0 0 2 2
use contact_9  contact_9_5
timestamp 1644969367
transform 1 0 1400 0 1 106
box 0 0 2 2
use contact_9  contact_9_6
timestamp 1644969367
transform 1 0 1292 0 1 106
box 0 0 2 2
use contact_9  contact_9_7
timestamp 1644969367
transform 1 0 1184 0 1 106
box 0 0 2 2
use contact_9  contact_9_8
timestamp 1644969367
transform 1 0 1076 0 1 106
box 0 0 2 2
use contact_9  contact_9_9
timestamp 1644969367
transform 1 0 968 0 1 106
box 0 0 2 2
use contact_9  contact_9_10
timestamp 1644969367
transform 1 0 860 0 1 106
box 0 0 2 2
use contact_9  contact_9_11
timestamp 1644969367
transform 1 0 752 0 1 106
box 0 0 2 2
use contact_9  contact_9_12
timestamp 1644969367
transform 1 0 644 0 1 106
box 0 0 2 2
use contact_9  contact_9_13
timestamp 1644969367
transform 1 0 536 0 1 106
box 0 0 2 2
use contact_9  contact_9_14
timestamp 1644969367
transform 1 0 428 0 1 106
box 0 0 2 2
use contact_9  contact_9_15
timestamp 1644969367
transform 1 0 320 0 1 106
box 0 0 2 2
use contact_9  contact_9_16
timestamp 1644969367
transform 1 0 212 0 1 106
box 0 0 2 2
use contact_9  contact_9_17
timestamp 1644969367
transform 1 0 104 0 1 106
box 0 0 2 2
use contact_9  contact_9_18
timestamp 1644969367
transform 1 0 0 0 1 106
box 0 0 2 2
<< labels >>
rlabel mvvaractor s 993 -41 993 -41 4 G
rlabel locali s 885 147 885 147 4 S
rlabel locali s 25 147 25 147 4 S
rlabel locali s 1533 147 1533 147 4 S
rlabel locali s 1317 147 1317 147 4 S
rlabel locali s 1749 147 1749 147 4 S
rlabel locali s 669 147 669 147 4 S
rlabel locali s 237 147 237 147 4 S
rlabel locali s 1101 147 1101 147 4 S
rlabel locali s 1961 147 1961 147 4 S
rlabel locali s 453 147 453 147 4 S
rlabel locali s 993 63 993 63 4 D
<< properties >>
string FIXED_BBOX -54 -56 2040 63
string GDS_FILE sram_0rw2r1w_32_128_sky130A.gds
string GDS_END 3388336
string GDS_START 3384084
<< end >>
