magic
tech sky130A
magscale 1 2
timestamp 1644949024
<< checkpaint >>
rect -1260 -1260 12174 30220
<< metal1 >>
rect 6883 28184 7024 28212
rect 6883 28172 6911 28184
rect 6734 28144 6911 28172
rect 6883 28058 7024 28086
rect 6883 28046 6911 28058
rect 6734 28018 6911 28046
rect 6883 27832 7024 27860
rect 6883 27820 6911 27832
rect 6734 27792 6911 27820
rect 6883 26780 7024 26800
rect 6734 26772 7024 26780
rect 6734 26752 6911 26772
rect 6883 26554 7024 26574
rect 6734 26546 7024 26554
rect 6734 26526 6911 26546
rect 6883 26428 7024 26448
rect 6734 26420 7024 26428
rect 6734 26400 6911 26420
rect 6883 25104 7024 25132
rect 6883 25096 6911 25104
rect 6734 25068 6911 25096
rect 6883 24978 7024 25006
rect 6883 24970 6911 24978
rect 6734 24942 6911 24970
rect 6883 24752 7024 24780
rect 6883 24744 6911 24752
rect 6734 24716 6911 24744
rect 6883 23704 7024 23720
rect 6734 23692 7024 23704
rect 6734 23676 6911 23692
rect 6883 23478 7024 23494
rect 6734 23466 7024 23478
rect 6734 23450 6911 23466
rect 6883 23352 7024 23368
rect 6734 23340 7024 23352
rect 6734 23324 6911 23340
rect 6883 22024 7024 22052
rect 6883 22020 6911 22024
rect 6734 21992 6911 22020
rect 6883 21898 7024 21926
rect 6883 21894 6911 21898
rect 6734 21866 6911 21894
rect 6883 21672 7024 21700
rect 6883 21668 6911 21672
rect 6734 21640 6911 21668
rect 6883 20628 7024 20640
rect 6734 20612 7024 20628
rect 6734 20600 6911 20612
rect 6883 20402 7024 20414
rect 6734 20386 7024 20402
rect 6734 20374 6911 20386
rect 6883 20276 7024 20288
rect 6734 20260 7024 20276
rect 6734 20248 6911 20260
rect 6883 18944 7024 18972
rect 6734 18916 6911 18944
rect 6883 18818 7024 18846
rect 6734 18790 6911 18818
rect 6883 18592 7024 18620
rect 6734 18564 6911 18592
rect 6883 17552 7024 17560
rect 6734 17532 7024 17552
rect 6734 17524 6911 17532
rect 6883 17326 7024 17334
rect 6734 17306 7024 17326
rect 6734 17298 6911 17306
rect 6883 17200 7024 17208
rect 6734 17180 7024 17200
rect 6734 17172 6911 17180
rect 6883 15868 7024 15892
rect 6734 15864 7024 15868
rect 6734 15840 6911 15864
rect 6883 15742 7024 15766
rect 6734 15738 7024 15742
rect 6734 15714 6911 15738
rect 6883 15516 7024 15540
rect 6734 15512 7024 15516
rect 6734 15488 6911 15512
rect 6883 14476 7024 14480
rect 6734 14452 7024 14476
rect 6734 14448 6911 14452
rect 6883 14250 7024 14254
rect 6734 14226 7024 14250
rect 6734 14222 6911 14226
rect 6883 14124 7024 14128
rect 6734 14100 7024 14124
rect 6734 14096 6911 14100
rect 6883 12792 7024 12812
rect 6734 12784 7024 12792
rect 6734 12764 6911 12784
rect 6883 12666 7024 12686
rect 6734 12658 7024 12666
rect 6734 12638 6911 12658
rect 6883 12440 7024 12460
rect 6734 12432 7024 12440
rect 6734 12412 6911 12432
rect 6734 11372 7024 11400
rect 6734 11146 7024 11174
rect 6734 11020 7024 11048
rect 6883 9716 7024 9732
rect 6734 9704 7024 9716
rect 6734 9688 6911 9704
rect 6883 9590 7024 9606
rect 6734 9578 7024 9590
rect 6734 9562 6911 9578
rect 6883 9364 7024 9380
rect 6734 9352 7024 9364
rect 6734 9336 6911 9352
rect 6734 8320 6911 8324
rect 6734 8296 7024 8320
rect 6883 8292 7024 8296
rect 6734 8094 6911 8098
rect 6734 8070 7024 8094
rect 6883 8066 7024 8070
rect 6734 7968 6911 7972
rect 6734 7944 7024 7968
rect 6883 7940 7024 7944
rect 6883 6640 7024 6652
rect 6734 6624 7024 6640
rect 6734 6612 6911 6624
rect 6883 6514 7024 6526
rect 6734 6498 7024 6514
rect 6734 6486 6911 6498
rect 6883 6288 7024 6300
rect 6734 6272 7024 6288
rect 6734 6260 6911 6272
rect 6734 5240 6911 5248
rect 6734 5220 7024 5240
rect 6883 5212 7024 5220
rect 6734 5014 6911 5022
rect 6734 4994 7024 5014
rect 6883 4986 7024 4994
rect 6734 4888 6911 4896
rect 6734 4868 7024 4888
rect 6883 4860 7024 4868
rect 6634 3568 6640 3620
rect 6692 3608 6698 3620
rect 6692 3580 8570 3608
rect 6692 3568 6698 3580
rect 10428 1447 10434 1459
rect 8969 1419 10434 1447
rect 10428 1407 10434 1419
rect 10486 1407 10492 1459
<< via1 >>
rect 6640 3568 6692 3620
rect 10434 1407 10486 1459
<< metal2 >>
rect 18 4216 46 28848
rect 102 4216 130 28848
rect 186 4216 214 28848
rect 270 4216 298 28848
rect 354 4216 382 28848
rect 438 4216 466 28848
rect 5530 28810 5558 28838
rect 6652 3626 6680 3796
rect 7220 3664 7274 3692
rect 8018 3664 8072 3692
rect 8816 3664 8870 3692
rect 9614 3664 9668 3692
rect 6640 3620 6692 3626
rect 6640 3562 6692 3568
rect 6652 0 6680 3562
rect 7226 2520 7254 2760
rect 7498 2520 7526 2760
rect 8004 2520 8032 2760
rect 8276 2520 8304 2760
rect 10446 1465 10474 28960
rect 10434 1459 10486 1465
rect 10434 1401 10486 1407
rect 10446 0 10474 1401
<< metal3 >>
rect 792 28811 924 28885
rect 1664 28811 1796 28885
rect 5128 28787 5260 28861
rect 6668 28787 6800 28861
rect 792 27271 924 27345
rect 1664 27271 1796 27345
rect 5128 27249 5260 27323
rect 6668 27249 6800 27323
rect 792 25731 924 25805
rect 1664 25731 1796 25805
rect 5128 25711 5260 25785
rect 6668 25711 6800 25785
rect 792 24191 924 24265
rect 1664 24191 1796 24265
rect 5128 24173 5260 24247
rect 6668 24173 6800 24247
rect 792 22651 924 22725
rect 1664 22651 1796 22725
rect 5128 22635 5260 22709
rect 6668 22635 6800 22709
rect 5128 21097 5260 21171
rect 6668 21097 6800 21171
rect 792 19575 924 19649
rect 1664 19575 1796 19649
rect 5128 19559 5260 19633
rect 6668 19559 6800 19633
rect 792 18035 924 18109
rect 1664 18035 1796 18109
rect 5128 18021 5260 18095
rect 6668 18021 6800 18095
rect 792 16495 924 16569
rect 1664 16495 1796 16569
rect 5128 16483 5260 16557
rect 6668 16483 6800 16557
rect 792 14955 924 15029
rect 1664 14955 1796 15029
rect 5128 14945 5260 15019
rect 6668 14945 6800 15019
rect 792 13415 924 13489
rect 1664 13415 1796 13489
rect 5128 13407 5260 13481
rect 6668 13407 6800 13481
rect 5128 11869 5260 11943
rect 6668 11869 6800 11943
rect 792 10339 924 10413
rect 1664 10339 1796 10413
rect 5128 10331 5260 10405
rect 6668 10331 6800 10405
rect 792 8799 924 8873
rect 1664 8799 1796 8873
rect 5128 8793 5260 8867
rect 6668 8793 6800 8867
rect 792 7259 924 7333
rect 1664 7259 1796 7333
rect 5128 7255 5260 7329
rect 6668 7255 6800 7329
rect 792 5719 924 5793
rect 1664 5719 1796 5793
rect 5128 5717 5260 5791
rect 6668 5717 6800 5791
rect 792 4179 924 4253
rect 1664 4179 1796 4253
rect 5128 4179 5260 4253
rect 6668 4179 6800 4253
rect 7340 3856 7406 3988
rect 8138 3856 8204 3988
rect 8936 3856 9002 3988
rect 9734 3856 9800 3988
rect 7340 3024 7406 3156
rect 8138 3024 8204 3156
rect 8936 3024 9002 3156
rect 9734 3024 9800 3156
rect 7094 2689 7226 2763
rect 7366 2689 7498 2763
rect 7872 2689 8004 2763
rect 8144 2689 8276 2763
rect 8650 2689 8782 2763
rect 8922 2689 9054 2763
rect 9428 2689 9560 2763
rect 9700 2689 9832 2763
rect 7094 1743 7226 1817
rect 7366 1743 7498 1817
rect 7872 1743 8004 1817
rect 8144 1743 8276 1817
rect 8650 1743 8782 1817
rect 8922 1743 9054 1817
rect 9428 1743 9560 1817
rect 9700 1743 9832 1817
rect 7184 464 7250 596
rect 7962 464 8028 596
rect 8740 464 8806 596
rect 9518 464 9584 596
rect 10296 464 10362 596
use contact_17  contact_17_0
timestamp 1644949024
transform 1 0 10428 0 1 1401
box 0 0 1 1
use contact_17  contact_17_1
timestamp 1644949024
transform 1 0 6634 0 1 3562
box 0 0 1 1
use port_address  port_address_0
timestamp 1644949024
transform 1 0 0 0 1 4216
box 0 -42 6800 24669
use port_data  port_data_0
timestamp 1644949024
transform 1 0 7024 0 1 0
box 0 406 3890 3988
use replica_bitcell_array  replica_bitcell_array_0
timestamp 1644949024
transform 1 0 7024 0 1 4216
box 0 -42 3112 24682
<< labels >>
rlabel metal2 s 6652 0 6680 3796 4 w_en
rlabel metal2 s 5530 28810 5558 28838 4 wl_en
rlabel metal2 s 10446 0 10474 28960 4 p_en_bar
rlabel metal2 s 7220 3664 7274 3692 4 din0_0
rlabel metal2 s 8018 3664 8072 3692 4 din0_1
rlabel metal2 s 8816 3664 8870 3692 4 din0_2
rlabel metal2 s 9614 3664 9668 3692 4 din0_3
rlabel metal2 s 7226 2520 7254 2760 4 dout0_0
rlabel metal2 s 7240 2640 7240 2640 4 dout1_0
rlabel metal2 s 7498 2520 7526 2760 4 dout0_1
rlabel metal2 s 7512 2640 7512 2640 4 dout1_1
rlabel metal2 s 8004 2520 8032 2760 4 dout0_2
rlabel metal2 s 8018 2640 8018 2640 4 dout1_2
rlabel metal2 s 8276 2520 8304 2760 4 dout0_3
rlabel metal2 s 8290 2640 8290 2640 4 dout1_3
rlabel metal2 s 18 4216 46 28848 4 addr0
rlabel metal2 s 102 4216 130 28848 4 addr1
rlabel metal2 s 186 4216 214 28848 4 addr2
rlabel metal2 s 270 4216 298 28848 4 addr3
rlabel metal2 s 354 4216 382 28848 4 addr4
rlabel metal2 s 438 4216 466 28848 4 addr5
rlabel metal3 s 6668 21096 6800 21170 4 vdd
rlabel metal3 s 5128 18020 5260 18094 4 vdd
rlabel metal3 s 792 24190 924 24264 4 vdd
rlabel metal3 s 8144 1742 8276 1816 4 vdd
rlabel metal3 s 8922 1742 9054 1816 4 vdd
rlabel metal3 s 8650 1742 8782 1816 4 vdd
rlabel metal3 s 1664 18034 1796 18108 4 vdd
rlabel metal3 s 1664 8798 1796 8872 4 vdd
rlabel metal3 s 5128 24172 5260 24246 4 vdd
rlabel metal3 s 1664 5718 1796 5792 4 vdd
rlabel metal3 s 1664 24190 1796 24264 4 vdd
rlabel metal3 s 1664 27270 1796 27344 4 vdd
rlabel metal3 s 5128 5716 5260 5790 4 vdd
rlabel metal3 s 10296 464 10362 596 4 vdd
rlabel metal3 s 8740 464 8806 596 4 vdd
rlabel metal3 s 5128 27248 5260 27322 4 vdd
rlabel metal3 s 5128 11868 5260 11942 4 vdd
rlabel metal3 s 6668 8792 6800 8866 4 vdd
rlabel metal3 s 6668 14944 6800 15018 4 vdd
rlabel metal3 s 8936 3024 9002 3156 4 vdd
rlabel metal3 s 792 18034 924 18108 4 vdd
rlabel metal3 s 792 5718 924 5792 4 vdd
rlabel metal3 s 6668 24172 6800 24246 4 vdd
rlabel metal3 s 6668 18020 6800 18094 4 vdd
rlabel metal3 s 9518 464 9584 596 4 vdd
rlabel metal3 s 7962 464 8028 596 4 vdd
rlabel metal3 s 6668 11868 6800 11942 4 vdd
rlabel metal3 s 792 27270 924 27344 4 vdd
rlabel metal3 s 7872 1742 8004 1816 4 vdd
rlabel metal3 s 6668 27248 6800 27322 4 vdd
rlabel metal3 s 9734 3024 9800 3156 4 vdd
rlabel metal3 s 8138 3024 8204 3156 4 vdd
rlabel metal3 s 9428 1742 9560 1816 4 vdd
rlabel metal3 s 1664 14954 1796 15028 4 vdd
rlabel metal3 s 7094 1742 7226 1816 4 vdd
rlabel metal3 s 9700 1742 9832 1816 4 vdd
rlabel metal3 s 5128 21096 5260 21170 4 vdd
rlabel metal3 s 5128 14944 5260 15018 4 vdd
rlabel metal3 s 5128 8792 5260 8866 4 vdd
rlabel metal3 s 6668 5716 6800 5790 4 vdd
rlabel metal3 s 792 14954 924 15028 4 vdd
rlabel metal3 s 7366 1742 7498 1816 4 vdd
rlabel metal3 s 7340 3024 7406 3156 4 vdd
rlabel metal3 s 792 8798 924 8872 4 vdd
rlabel metal3 s 7184 464 7250 596 4 vdd
rlabel metal3 s 8144 2688 8276 2762 4 gnd
rlabel metal3 s 792 4178 924 4252 4 gnd
rlabel metal3 s 1664 4178 1796 4252 4 gnd
rlabel metal3 s 7872 2688 8004 2762 4 gnd
rlabel metal3 s 8138 3856 8204 3988 4 gnd
rlabel metal3 s 9428 2688 9560 2762 4 gnd
rlabel metal3 s 792 28810 924 28884 4 gnd
rlabel metal3 s 1664 7258 1796 7332 4 gnd
rlabel metal3 s 6668 10330 6800 10404 4 gnd
rlabel metal3 s 5128 19558 5260 19632 4 gnd
rlabel metal3 s 8922 2688 9054 2762 4 gnd
rlabel metal3 s 792 13414 924 13488 4 gnd
rlabel metal3 s 8936 3856 9002 3988 4 gnd
rlabel metal3 s 792 10338 924 10412 4 gnd
rlabel metal3 s 1664 28810 1796 28884 4 gnd
rlabel metal3 s 5128 10330 5260 10404 4 gnd
rlabel metal3 s 1664 25730 1796 25804 4 gnd
rlabel metal3 s 5128 16482 5260 16556 4 gnd
rlabel metal3 s 6668 19558 6800 19632 4 gnd
rlabel metal3 s 792 25730 924 25804 4 gnd
rlabel metal3 s 9700 2688 9832 2762 4 gnd
rlabel metal3 s 5128 7254 5260 7328 4 gnd
rlabel metal3 s 7366 2688 7498 2762 4 gnd
rlabel metal3 s 8650 2688 8782 2762 4 gnd
rlabel metal3 s 5128 25710 5260 25784 4 gnd
rlabel metal3 s 9734 3856 9800 3988 4 gnd
rlabel metal3 s 1664 16494 1796 16568 4 gnd
rlabel metal3 s 7340 3856 7406 3988 4 gnd
rlabel metal3 s 6668 22634 6800 22708 4 gnd
rlabel metal3 s 792 16494 924 16568 4 gnd
rlabel metal3 s 1664 22650 1796 22724 4 gnd
rlabel metal3 s 6668 28786 6800 28860 4 gnd
rlabel metal3 s 792 7258 924 7332 4 gnd
rlabel metal3 s 6668 13406 6800 13480 4 gnd
rlabel metal3 s 1664 10338 1796 10412 4 gnd
rlabel metal3 s 5128 28786 5260 28860 4 gnd
rlabel metal3 s 5128 4178 5260 4252 4 gnd
rlabel metal3 s 792 19574 924 19648 4 gnd
rlabel metal3 s 6668 4178 6800 4252 4 gnd
rlabel metal3 s 6668 7254 6800 7328 4 gnd
rlabel metal3 s 6668 16482 6800 16556 4 gnd
rlabel metal3 s 7094 2688 7226 2762 4 gnd
rlabel metal3 s 6668 25710 6800 25784 4 gnd
rlabel metal3 s 1664 13414 1796 13488 4 gnd
rlabel metal3 s 5128 13406 5260 13480 4 gnd
rlabel metal3 s 1664 19574 1796 19648 4 gnd
rlabel metal3 s 792 22650 924 22724 4 gnd
rlabel metal3 s 5128 22634 5260 22708 4 gnd
<< properties >>
string FIXED_BBOX 0 0 10998 28960
string GDS_FILE sram_0rw2r1w_4_16_sky130A.gds
string GDS_END 109736
string GDS_START 73216
<< end >>
