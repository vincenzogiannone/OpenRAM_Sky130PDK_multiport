magic
tech sky130A
magscale 1 2
timestamp 1644951705
<< checkpaint >>
rect -1296 -1277 3824 2155
<< nwell >>
rect -36 402 2564 895
<< locali >>
rect 0 821 2528 855
rect 48 338 114 404
rect 1261 354 1295 388
rect 0 -17 2528 17
use pinv_13  pinv_13_0
timestamp 1644951705
transform 1 0 0 0 1 0
box -36 -17 2564 895
<< labels >>
rlabel locali s 1278 371 1278 371 4 Z
rlabel locali s 81 371 81 371 4 A
rlabel locali s 1264 0 1264 0 4 gnd
rlabel locali s 1264 838 1264 838 4 vdd
<< properties >>
string FIXED_BBOX 0 0 2528 838
string GDS_FILE sram_0rw2r1w_16_128_sky130A.gds
string GDS_END 2042522
string GDS_START 2041676
<< end >>
