VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO sram_0rw2r1w_16_128_sky130A
   CLASS BLOCK ;
   SIZE 379.18 BY 321.94 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  98.58 0.0 99.34 1.82 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  104.94 0.0 105.7 1.82 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  112.36 0.0 113.12 1.82 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  120.84 0.0 121.6 1.82 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  128.26 0.0 129.02 1.82 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  135.68 0.0 136.44 1.82 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  143.1 0.0 143.86 1.82 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  149.46 0.0 150.22 1.82 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  156.88 0.0 157.64 1.82 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  164.3 0.0 165.06 1.82 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  171.72 0.0 172.48 1.82 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  180.2 0.0 180.96 1.82 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  186.56 0.0 187.32 1.82 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  193.98 0.0 194.74 1.82 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  201.4 0.0 202.16 1.82 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  208.82 0.0 209.58 1.82 ;
      END
   END din0[15]
   PIN addr[0]
      DIRECTION INPUT ;
      PORT
      END
   END addr[0]
   PIN addr[1]
      DIRECTION INPUT ;
      PORT
      END
   END addr[1]
   PIN addr[2]
      DIRECTION INPUT ;
      PORT
      END
   END addr[2]
   PIN addr[3]
      DIRECTION INPUT ;
      PORT
      END
   END addr[3]
   PIN addr[4]
      DIRECTION INPUT ;
      PORT
      END
   END addr[4]
   PIN addr[5]
      DIRECTION INPUT ;
      PORT
      END
   END addr[5]
   PIN addr[6]
      DIRECTION INPUT ;
      PORT
      END
   END addr[6]
   PIN addr[7]
      DIRECTION INPUT ;
      PORT
      END
   END addr[7]
   PIN addr[8]
      DIRECTION INPUT ;
      PORT
      END
   END addr[8]
   PIN csb
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  14.605 40.815 15.265 41.185 ;
      END
   END csb
   PIN web
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  14.605 34.895 15.265 35.265 ;
      END
   END web
   PIN clk
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  31.8 0.0 32.56 1.82 ;
      END
   END clk
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  116.6 0.0 117.36 1.82 ;
      END
   END dout0[0]
   PIN dout1[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  116.355 56.155 117.015 56.525 ;
      END
   END dout1[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  117.66 0.0 118.42 1.82 ;
      END
   END dout0[1]
   PIN dout1[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  117.715 56.155 118.375 56.525 ;
      END
   END dout1[1]
   PIN dout0[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  131.44 0.0 132.2 1.82 ;
      END
   END dout0[2]
   PIN dout1[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  131.915 56.155 132.575 56.525 ;
      END
   END dout1[2]
   PIN dout0[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  133.56 0.0 134.32 1.82 ;
      END
   END dout0[3]
   PIN dout1[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  133.275 56.155 133.935 56.525 ;
      END
   END dout1[3]
   PIN dout0[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  147.34 0.0 148.1 1.82 ;
      END
   END dout0[4]
   PIN dout1[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  147.475 56.155 148.135 56.525 ;
      END
   END dout1[4]
   PIN dout0[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  150.52 0.0 151.28 1.82 ;
      END
   END dout0[5]
   PIN dout1[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  148.835 56.155 149.495 56.525 ;
      END
   END dout1[5]
   PIN dout0[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  162.18 0.0 162.94 1.82 ;
      END
   END dout0[6]
   PIN dout1[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  163.035 56.155 163.695 56.525 ;
      END
   END dout1[6]
   PIN dout0[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  165.36 0.0 166.12 1.82 ;
      END
   END dout0[7]
   PIN dout1[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  164.395 56.155 165.055 56.525 ;
      END
   END dout1[7]
   PIN dout0[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  178.08 0.0 178.84 1.82 ;
      END
   END dout0[8]
   PIN dout1[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  178.595 56.155 179.255 56.525 ;
      END
   END dout1[8]
   PIN dout0[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  181.26 0.0 182.02 1.82 ;
      END
   END dout0[9]
   PIN dout1[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  179.955 56.155 180.615 56.525 ;
      END
   END dout1[9]
   PIN dout0[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  195.04 0.0 195.8 1.82 ;
      END
   END dout0[10]
   PIN dout1[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  194.155 56.155 194.815 56.525 ;
      END
   END dout1[10]
   PIN dout0[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  196.1 0.0 196.86 1.82 ;
      END
   END dout0[11]
   PIN dout1[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  195.515 56.155 196.175 56.525 ;
      END
   END dout1[11]
   PIN dout0[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  209.88 0.0 210.64 1.82 ;
      END
   END dout0[12]
   PIN dout1[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  209.715 56.155 210.375 56.525 ;
      END
   END dout1[12]
   PIN dout0[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  210.94 0.0 211.7 1.82 ;
      END
   END dout0[13]
   PIN dout1[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  211.075 56.155 211.735 56.525 ;
      END
   END dout1[13]
   PIN dout0[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  224.72 0.0 225.48 1.82 ;
      END
   END dout0[14]
   PIN dout1[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  225.275 56.155 225.935 56.525 ;
      END
   END dout1[14]
   PIN dout0[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  226.84 0.0 227.6 1.82 ;
      END
   END dout0[15]
   PIN dout1[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  226.635 56.155 227.295 56.525 ;
      END
   END dout1[15]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met4 ;
         RECT  371.0 7.42 373.88 316.64 ;
         LAYER met4 ;
         RECT  7.42 7.42 10.3 316.64 ;
         LAYER met3 ;
         RECT  7.42 7.42 373.88 10.3 ;
         LAYER met3 ;
         RECT  7.42 313.76 373.88 316.64 ;
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met3 ;
         RECT  2.12 319.06 379.18 321.94 ;
         LAYER met4 ;
         RECT  376.3 2.12 379.18 321.94 ;
         LAYER met3 ;
         RECT  2.12 2.12 379.18 5.0 ;
         LAYER met4 ;
         RECT  2.12 2.12 5.0 321.94 ;
      END
   END gnd
   OBS
   LAYER  met1 ;
      RECT  0.62 0.62 378.56 321.32 ;
   LAYER  met2 ;
      RECT  0.62 0.62 378.56 321.32 ;
   LAYER  met3 ;
      RECT  0.62 40.215 14.005 41.785 ;
      RECT  15.865 40.215 378.56 41.785 ;
      RECT  14.005 35.865 15.865 40.215 ;
      RECT  15.865 41.785 115.755 55.555 ;
      RECT  15.865 55.555 115.755 57.125 ;
      RECT  115.755 41.785 117.615 55.555 ;
      RECT  117.615 41.785 378.56 55.555 ;
      RECT  118.975 55.555 131.315 57.125 ;
      RECT  134.535 55.555 146.875 57.125 ;
      RECT  150.095 55.555 162.435 57.125 ;
      RECT  165.655 55.555 177.995 57.125 ;
      RECT  181.215 55.555 193.555 57.125 ;
      RECT  196.775 55.555 209.115 57.125 ;
      RECT  212.335 55.555 224.675 57.125 ;
      RECT  227.895 55.555 378.56 57.125 ;
      RECT  0.62 6.82 6.82 10.9 ;
      RECT  0.62 10.9 6.82 40.215 ;
      RECT  6.82 10.9 14.005 40.215 ;
      RECT  15.865 10.9 374.48 40.215 ;
      RECT  374.48 6.82 378.56 10.9 ;
      RECT  374.48 10.9 378.56 40.215 ;
      RECT  14.005 10.9 15.865 34.295 ;
      RECT  0.62 41.785 6.82 313.16 ;
      RECT  0.62 313.16 6.82 317.24 ;
      RECT  6.82 41.785 14.005 313.16 ;
      RECT  14.005 41.785 15.865 313.16 ;
      RECT  15.865 57.125 115.755 313.16 ;
      RECT  115.755 57.125 117.615 313.16 ;
      RECT  117.615 57.125 374.48 313.16 ;
      RECT  374.48 57.125 378.56 313.16 ;
      RECT  374.48 313.16 378.56 317.24 ;
      RECT  0.62 317.24 1.52 318.46 ;
      RECT  0.62 318.46 1.52 321.32 ;
      RECT  1.52 317.24 6.82 318.46 ;
      RECT  6.82 317.24 14.005 318.46 ;
      RECT  14.005 317.24 15.865 318.46 ;
      RECT  15.865 317.24 115.755 318.46 ;
      RECT  115.755 317.24 117.615 318.46 ;
      RECT  117.615 317.24 374.48 318.46 ;
      RECT  374.48 317.24 378.56 318.46 ;
      RECT  0.62 0.62 1.52 1.52 ;
      RECT  0.62 1.52 1.52 5.6 ;
      RECT  0.62 5.6 1.52 6.82 ;
      RECT  1.52 0.62 6.82 1.52 ;
      RECT  1.52 5.6 6.82 6.82 ;
      RECT  6.82 0.62 14.005 1.52 ;
      RECT  6.82 5.6 14.005 6.82 ;
      RECT  15.865 0.62 374.48 1.52 ;
      RECT  15.865 5.6 374.48 6.82 ;
      RECT  374.48 0.62 378.56 1.52 ;
      RECT  374.48 5.6 378.56 6.82 ;
      RECT  14.005 0.62 15.865 1.52 ;
      RECT  14.005 5.6 15.865 6.82 ;
   LAYER  met4 ;
      RECT  97.98 2.42 99.94 321.32 ;
      RECT  99.94 0.62 104.34 2.42 ;
      RECT  106.3 0.62 111.76 2.42 ;
      RECT  122.2 0.62 127.66 2.42 ;
      RECT  137.04 0.62 142.5 2.42 ;
      RECT  187.92 0.62 193.38 2.42 ;
      RECT  202.76 0.62 208.22 2.42 ;
      RECT  33.16 0.62 97.98 2.42 ;
      RECT  113.72 0.62 116.0 2.42 ;
      RECT  119.02 0.62 120.24 2.42 ;
      RECT  129.62 0.62 130.84 2.42 ;
      RECT  132.8 0.62 132.96 2.42 ;
      RECT  134.92 0.62 135.08 2.42 ;
      RECT  144.46 0.62 146.74 2.42 ;
      RECT  148.7 0.62 148.86 2.42 ;
      RECT  151.88 0.62 156.28 2.42 ;
      RECT  158.24 0.62 161.58 2.42 ;
      RECT  163.54 0.62 163.7 2.42 ;
      RECT  166.72 0.62 171.12 2.42 ;
      RECT  173.08 0.62 177.48 2.42 ;
      RECT  179.44 0.62 179.6 2.42 ;
      RECT  182.62 0.62 185.96 2.42 ;
      RECT  197.46 0.62 200.8 2.42 ;
      RECT  212.3 0.62 224.12 2.42 ;
      RECT  226.08 0.62 226.24 2.42 ;
      RECT  99.94 2.42 370.4 6.82 ;
      RECT  99.94 6.82 370.4 317.24 ;
      RECT  99.94 317.24 370.4 321.32 ;
      RECT  370.4 2.42 374.48 6.82 ;
      RECT  370.4 317.24 374.48 321.32 ;
      RECT  6.82 2.42 10.9 6.82 ;
      RECT  6.82 317.24 10.9 321.32 ;
      RECT  10.9 2.42 97.98 6.82 ;
      RECT  10.9 6.82 97.98 317.24 ;
      RECT  10.9 317.24 97.98 321.32 ;
      RECT  228.2 0.62 375.7 1.52 ;
      RECT  228.2 1.52 375.7 2.42 ;
      RECT  375.7 0.62 378.56 1.52 ;
      RECT  374.48 2.42 375.7 6.82 ;
      RECT  374.48 6.82 375.7 317.24 ;
      RECT  374.48 317.24 375.7 321.32 ;
      RECT  0.62 0.62 1.52 1.52 ;
      RECT  0.62 1.52 1.52 2.42 ;
      RECT  1.52 0.62 5.6 1.52 ;
      RECT  5.6 0.62 31.2 1.52 ;
      RECT  5.6 1.52 31.2 2.42 ;
      RECT  0.62 2.42 1.52 6.82 ;
      RECT  5.6 2.42 6.82 6.82 ;
      RECT  0.62 6.82 1.52 317.24 ;
      RECT  5.6 6.82 6.82 317.24 ;
      RECT  0.62 317.24 1.52 321.32 ;
      RECT  5.6 317.24 6.82 321.32 ;
   END
END    sram_0rw2r1w_16_128_sky130A
END    LIBRARY
