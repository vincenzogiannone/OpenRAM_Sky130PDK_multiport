magic
tech sky130A
magscale 1 2
timestamp 1643671299
<< checkpaint >>
rect -1296 -1277 2079 2155
<< nwell >>
rect -36 402 819 895
<< pwell >>
rect 690 51 740 133
<< psubdiff >>
rect 690 109 740 133
rect 690 75 698 109
rect 732 75 740 109
rect 690 51 740 75
<< nsubdiff >>
rect 690 763 740 787
rect 690 729 698 763
rect 732 729 740 763
rect 690 705 740 729
<< psubdiffcont >>
rect 698 75 732 109
<< nsubdiffcont >>
rect 698 729 732 763
<< poly >>
rect 114 410 144 479
rect 48 394 144 410
rect 48 360 64 394
rect 98 360 144 394
rect 48 344 144 360
rect 114 191 144 344
<< polycont >>
rect 64 360 98 394
<< locali >>
rect 0 821 783 855
rect 62 628 96 821
rect 274 628 308 821
rect 490 628 524 821
rect 698 763 732 821
rect 698 713 732 729
rect 48 394 114 410
rect 48 360 64 394
rect 98 360 114 394
rect 48 344 114 360
rect 380 394 414 594
rect 380 360 431 394
rect 380 160 414 360
rect 698 109 732 125
rect 62 17 96 60
rect 274 17 308 60
rect 490 17 524 60
rect 698 17 732 75
rect 0 -17 783 17
use contact_12  contact_12_0
timestamp 1643671299
transform 1 0 48 0 1 344
box 0 0 1 1
use contact_11  contact_11_0
timestamp 1643671299
transform 1 0 690 0 1 51
box 0 0 1 1
use contact_10  contact_10_0
timestamp 1643671299
transform 1 0 690 0 1 705
box 0 0 1 1
use nmos_m5_w0_420_sli_dli_da_p  nmos_m5_w0_420_sli_dli_da_p_0
timestamp 1643671299
transform 1 0 54 0 1 51
box 0 -26 582 143
use pmos_m5_w1_260_sli_dli_da_p  pmos_m5_w1_260_sli_dli_da_p_0
timestamp 1643671299
transform 1 0 54 0 1 535
box -59 -56 641 306
<< labels >>
rlabel locali s 81 377 81 377 4 A
rlabel locali s 414 377 414 377 4 Z
rlabel locali s 391 0 391 0 4 gnd
rlabel locali s 391 838 391 838 4 vdd
<< properties >>
string FIXED_BBOX 0 0 783 662
string GDS_FILE sram_0rw2r1w_16_32_sky130A.gds
string GDS_END 1150940
string GDS_START 1149192
<< end >>
