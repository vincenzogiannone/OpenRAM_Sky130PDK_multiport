magic
tech sky130A
magscale 1 2
timestamp 1643678851
<< checkpaint >>
rect -1296 -1277 3807 2155
<< nwell >>
rect -36 402 2547 895
<< pwell >>
rect 2418 51 2468 133
<< psubdiff >>
rect 2418 109 2468 133
rect 2418 75 2426 109
rect 2460 75 2468 109
rect 2418 51 2468 75
<< nsubdiff >>
rect 2418 763 2468 787
rect 2418 729 2426 763
rect 2460 729 2468 763
rect 2418 705 2468 729
<< psubdiffcont >>
rect 2426 75 2460 109
<< nsubdiffcont >>
rect 2426 729 2460 763
<< poly >>
rect 114 404 144 443
rect 48 388 144 404
rect 48 354 64 388
rect 98 354 144 388
rect 48 338 144 354
rect 114 203 144 338
<< polycont >>
rect 64 354 98 388
<< locali >>
rect 0 821 2511 855
rect 62 610 96 821
rect 274 610 308 821
rect 490 610 524 821
rect 706 610 740 821
rect 922 610 956 821
rect 1138 610 1172 821
rect 1354 610 1388 821
rect 1570 610 1604 821
rect 1786 610 1820 821
rect 2002 610 2036 821
rect 2218 610 2252 821
rect 2426 763 2460 821
rect 2426 713 2460 729
rect 48 388 114 404
rect 48 354 64 388
rect 98 354 114 388
rect 48 338 114 354
rect 1244 388 1278 576
rect 1244 354 1295 388
rect 1244 166 1278 354
rect 2426 109 2460 125
rect 62 17 96 66
rect 274 17 308 66
rect 490 17 524 66
rect 706 17 740 66
rect 922 17 956 66
rect 1138 17 1172 66
rect 1354 17 1388 66
rect 1570 17 1604 66
rect 1786 17 1820 66
rect 2002 17 2036 66
rect 2218 17 2252 66
rect 2426 17 2460 75
rect 0 -17 2511 17
use contact_12  contact_12_0
timestamp 1643678851
transform 1 0 48 0 1 338
box 0 0 1 1
use contact_11  contact_11_0
timestamp 1643678851
transform 1 0 2418 0 1 51
box 0 0 1 1
use contact_10  contact_10_0
timestamp 1643678851
transform 1 0 2418 0 1 705
box 0 0 1 1
use nmos_m21_w0_480_sli_dli_da_p  nmos_m21_w0_480_sli_dli_da_p_0
timestamp 1643678851
transform 1 0 54 0 1 51
box 0 -26 2310 152
use pmos_m21_w1_440_sli_dli_da_p  pmos_m21_w1_440_sli_dli_da_p_0
timestamp 1643678851
transform 1 0 54 0 1 499
box -59 -56 2369 342
<< labels >>
rlabel locali s 81 371 81 371 4 A
rlabel locali s 1278 371 1278 371 4 Z
rlabel locali s 1255 0 1255 0 4 gnd
rlabel locali s 1255 838 1255 838 4 vdd
<< properties >>
string FIXED_BBOX 0 0 2511 662
string GDS_FILE sram_0rw2r1w_16_128_sky130A.gds
string GDS_END 2110360
string GDS_START 2107588
<< end >>
