magic
tech sky130A
magscale 1 2
timestamp 1644951705
<< checkpaint >>
rect -1296 -1277 3068 2155
<< nwell >>
rect -36 402 1808 895
<< pwell >>
rect 1662 51 1712 133
<< psubdiff >>
rect 1662 109 1712 133
rect 1662 75 1670 109
rect 1704 75 1712 109
rect 1662 51 1712 75
<< nsubdiff >>
rect 1662 763 1712 787
rect 1662 729 1670 763
rect 1704 729 1712 763
rect 1662 705 1712 729
<< psubdiffcont >>
rect 1670 75 1704 109
<< nsubdiffcont >>
rect 1670 729 1704 763
<< poly >>
rect 114 404 144 443
rect 48 388 144 404
rect 48 354 64 388
rect 98 354 144 388
rect 48 338 144 354
rect 114 203 144 338
<< polycont >>
rect 64 354 98 388
<< locali >>
rect 0 821 1772 855
rect 62 610 96 821
rect 274 610 308 821
rect 490 610 524 821
rect 706 610 740 821
rect 922 610 956 821
rect 1138 610 1172 821
rect 1354 610 1388 821
rect 1566 610 1600 821
rect 1670 763 1704 821
rect 1670 713 1704 729
rect 48 388 114 404
rect 48 354 64 388
rect 98 354 114 388
rect 48 338 114 354
rect 814 388 848 576
rect 814 354 865 388
rect 814 166 848 354
rect 1670 109 1704 125
rect 62 17 96 66
rect 274 17 308 66
rect 490 17 524 66
rect 706 17 740 66
rect 922 17 956 66
rect 1138 17 1172 66
rect 1354 17 1388 66
rect 1566 17 1600 66
rect 1670 17 1704 75
rect 0 -17 1772 17
use contact_12  contact_12_0
timestamp 1644951705
transform 1 0 48 0 1 338
box 0 0 1 1
use contact_11  contact_11_0
timestamp 1644951705
transform 1 0 1662 0 1 51
box 0 0 1 1
use contact_10  contact_10_0
timestamp 1644951705
transform 1 0 1662 0 1 705
box 0 0 1 1
use nmos_m14_w0_480_sli_dli_da_p  nmos_m14_w0_480_sli_dli_da_p_0
timestamp 1644951705
transform 1 0 54 0 1 51
box 0 -26 1554 152
use pmos_m14_w1_440_sli_dli_da_p  pmos_m14_w1_440_sli_dli_da_p_0
timestamp 1644951705
transform 1 0 54 0 1 499
box -59 -56 1613 342
<< labels >>
rlabel locali s 81 371 81 371 4 A
rlabel locali s 848 371 848 371 4 Z
rlabel locali s 886 0 886 0 4 gnd
rlabel locali s 886 838 886 838 4 vdd
<< properties >>
string FIXED_BBOX 0 0 1772 838
string GDS_FILE sram_0rw2r1w_16_128_sky130A.gds
string GDS_END 1991500
string GDS_START 1989112
<< end >>
