magic
tech sky130A
magscale 1 2
timestamp 1644951705
<< checkpaint >>
rect -1296 -1277 4064 2155
<< nwell >>
rect -36 402 2804 895
<< locali >>
rect 0 821 2768 855
rect 48 344 114 410
rect 196 360 449 394
rect 564 360 817 394
rect 1027 356 1509 390
rect 2043 356 2077 390
rect 0 -17 2768 17
use pinv_12  pinv_12_0
timestamp 1644951705
transform 1 0 1428 0 1 0
box -36 -17 1376 895
use pinv_11  pinv_11_0
timestamp 1644951705
transform 1 0 736 0 1 0
box -36 -17 728 895
use pinv_0  pinv_0_0
timestamp 1644951705
transform 1 0 368 0 1 0
box -36 -17 404 895
use pinv_0  pinv_0_1
timestamp 1644951705
transform 1 0 0 0 1 0
box -36 -17 404 895
<< labels >>
rlabel locali s 2060 373 2060 373 4 Z
rlabel locali s 81 377 81 377 4 A
rlabel locali s 1384 0 1384 0 4 gnd
rlabel locali s 1384 838 1384 838 4 vdd
<< properties >>
string FIXED_BBOX 0 0 2768 838
string GDS_FILE sram_0rw2r1w_16_128_sky130A.gds
string GDS_END 2031076
string GDS_START 2029800
<< end >>
