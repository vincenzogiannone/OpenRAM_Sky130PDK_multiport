magic
tech sky130A
magscale 1 2
timestamp 1643671299
<< checkpaint >>
rect -1271 -1271 1493 1493
<< via1 >>
rect -11 -11 233 233
<< properties >>
string FIXED_BBOX 0 0 222 222
string GDS_FILE sram_0rw2r1w_16_32_sky130A.gds
string GDS_END 1254052
string GDS_START 1252768
<< end >>
