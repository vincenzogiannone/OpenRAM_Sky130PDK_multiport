magic
tech sky130A
magscale 1 2
timestamp 1643593061
<< checkpaint >>
rect -1292 -1302 8384 7162
<< locali >>
rect 3995 4734 4214 4768
rect 4180 4550 4214 4734
rect 3977 2207 4162 2241
rect 3977 2154 4011 2207
rect 3844 2120 4011 2154
<< viali >>
rect 3712 5472 3746 5506
rect 5257 5472 5291 5506
rect 4663 4550 4697 4584
rect 3760 4463 3794 4497
rect 3760 3883 3794 3917
rect 4639 3800 4673 3834
rect 3860 3643 3894 3677
rect 3860 3027 3894 3061
rect 4747 2870 4781 2904
rect 3760 2787 3794 2821
rect 3712 2120 3746 2154
rect 5115 2124 5149 2158
rect 4228 1967 4262 2001
rect 3712 1198 3746 1232
rect 6121 1192 6155 1226
<< metal1 >>
rect 2958 5463 2964 5515
rect 3016 5503 3022 5515
rect 3700 5506 3758 5512
rect 3700 5503 3712 5506
rect 3016 5475 3712 5503
rect 3016 5463 3022 5475
rect 3700 5472 3712 5475
rect 3746 5472 3758 5506
rect 3700 5466 3758 5472
rect 5242 5463 5248 5515
rect 5300 5463 5306 5515
rect 4648 4541 4654 4593
rect 4706 4541 4712 4593
rect 3042 4454 3048 4506
rect 3100 4494 3106 4506
rect 3748 4497 3806 4503
rect 3748 4494 3760 4497
rect 3100 4466 3760 4494
rect 3100 4454 3106 4466
rect 3748 4463 3760 4466
rect 3794 4463 3806 4497
rect 3748 4457 3806 4463
rect 3126 3874 3132 3926
rect 3184 3914 3190 3926
rect 3748 3917 3806 3923
rect 3748 3914 3760 3917
rect 3184 3886 3760 3914
rect 3184 3874 3190 3886
rect 3748 3883 3760 3886
rect 3794 3883 3806 3917
rect 3748 3877 3806 3883
rect 4624 3791 4630 3843
rect 4682 3791 4688 3843
rect 2958 3634 2964 3686
rect 3016 3674 3022 3686
rect 3848 3677 3906 3683
rect 3848 3674 3860 3677
rect 3016 3646 3860 3674
rect 3016 3634 3022 3646
rect 3848 3643 3860 3646
rect 3894 3643 3906 3677
rect 3848 3637 3906 3643
rect -18 3246 -12 3298
rect 40 3286 46 3298
rect 3294 3286 3300 3298
rect 40 3258 3300 3286
rect 40 3246 46 3258
rect 3294 3246 3300 3258
rect 3352 3246 3358 3298
rect 3378 3018 3384 3070
rect 3436 3058 3442 3070
rect 3848 3061 3906 3067
rect 3848 3058 3860 3061
rect 3436 3030 3860 3058
rect 3436 3018 3442 3030
rect 3848 3027 3860 3030
rect 3894 3027 3906 3061
rect 3848 3021 3906 3027
rect 4732 2861 4738 2913
rect 4790 2861 4796 2913
rect 3294 2778 3300 2830
rect 3352 2818 3358 2830
rect 3748 2821 3806 2827
rect 3748 2818 3760 2821
rect 3352 2790 3760 2818
rect 3352 2778 3358 2790
rect 3748 2787 3760 2790
rect 3794 2787 3806 2821
rect 3748 2781 3806 2787
rect 3294 2111 3300 2163
rect 3352 2151 3358 2163
rect 3700 2154 3758 2160
rect 3700 2151 3712 2154
rect 3352 2123 3712 2151
rect 3352 2111 3358 2123
rect 3700 2120 3712 2123
rect 3746 2120 3758 2154
rect 3700 2114 3758 2120
rect 5100 2115 5106 2167
rect 5158 2115 5164 2167
rect 4213 1958 4219 2010
rect 4271 1958 4277 2010
rect 3697 1189 3703 1241
rect 3755 1189 3761 1241
rect 6106 1183 6112 1235
rect 6164 1183 6170 1235
<< via1 >>
rect 2964 5463 3016 5515
rect 5248 5506 5300 5515
rect 5248 5472 5257 5506
rect 5257 5472 5291 5506
rect 5291 5472 5300 5506
rect 5248 5463 5300 5472
rect 4654 4584 4706 4593
rect 4654 4550 4663 4584
rect 4663 4550 4697 4584
rect 4697 4550 4706 4584
rect 4654 4541 4706 4550
rect 3048 4454 3100 4506
rect 3132 3874 3184 3926
rect 4630 3834 4682 3843
rect 4630 3800 4639 3834
rect 4639 3800 4673 3834
rect 4673 3800 4682 3834
rect 4630 3791 4682 3800
rect 2964 3634 3016 3686
rect -12 3246 40 3298
rect 3300 3246 3352 3298
rect 3384 3018 3436 3070
rect 4738 2904 4790 2913
rect 4738 2870 4747 2904
rect 4747 2870 4781 2904
rect 4781 2870 4790 2904
rect 4738 2861 4790 2870
rect 3300 2778 3352 2830
rect 3300 2111 3352 2163
rect 5106 2158 5158 2167
rect 5106 2124 5115 2158
rect 5115 2124 5149 2158
rect 5149 2124 5158 2158
rect 5106 2115 5158 2124
rect 4219 2001 4271 2010
rect 4219 1967 4228 2001
rect 4228 1967 4262 2001
rect 4262 1967 4271 2001
rect 4219 1958 4271 1967
rect 3703 1232 3755 1241
rect 3703 1198 3712 1232
rect 3712 1198 3746 1232
rect 3746 1198 3755 1232
rect 3703 1189 3755 1198
rect 6112 1226 6164 1235
rect 6112 1192 6121 1226
rect 6121 1192 6155 1226
rect 6155 1192 6164 1226
rect 6112 1183 6164 1192
<< metal2 >>
rect 2976 5515 3004 5902
rect 2976 3686 3004 5463
rect 3060 4506 3088 5902
rect 0 1676 28 3246
rect 2976 1834 3004 3634
rect 3060 2915 3088 4454
rect 3144 3926 3172 5902
rect 180 1416 234 1444
rect 180 232 234 260
rect 2976 0 3004 1778
rect 3060 0 3088 2859
rect 3144 573 3172 3874
rect 3144 0 3172 517
rect 3228 237 3256 5902
rect 3312 3298 3340 5902
rect 3312 2830 3340 3246
rect 3396 3070 3424 5902
rect 3312 2163 3340 2778
rect 3312 902 3340 2111
rect 3396 2012 3424 3018
rect 3396 1159 3424 1956
rect 3480 1495 3508 5902
rect 5300 5475 7124 5503
rect 4706 4553 7124 4581
rect 4682 3803 7124 3831
rect 5118 1834 5146 2115
rect 3228 0 3256 181
rect 3312 0 3340 846
rect 3396 0 3424 1103
rect 3480 0 3508 1439
rect 6164 1195 7124 1223
rect 6124 902 6152 1183
<< via2 >>
rect 3046 2859 3102 2915
rect 2962 1778 3018 1834
rect 2648 1439 2704 1495
rect 2158 1103 2214 1159
rect 2158 517 2214 573
rect 2648 181 2704 237
rect 3130 517 3186 573
rect 3382 1956 3438 2012
rect 4736 2913 4792 2915
rect 4736 2861 4738 2913
rect 4738 2861 4790 2913
rect 4790 2861 4792 2913
rect 4736 2859 4792 2861
rect 4217 2010 4273 2012
rect 4217 1958 4219 2010
rect 4219 1958 4271 2010
rect 4271 1958 4273 2010
rect 4217 1956 4273 1958
rect 5104 1778 5160 1834
rect 3466 1439 3522 1495
rect 3382 1103 3438 1159
rect 3298 846 3354 902
rect 3214 181 3270 237
rect 6110 846 6166 902
<< metal3 >>
rect 3044 2915 4794 2917
rect 3044 2859 3046 2915
rect 3102 2859 4736 2915
rect 4792 2859 4794 2915
rect 3044 2857 4794 2859
rect 3380 2012 4275 2014
rect 3380 1956 3382 2012
rect 3438 1956 4217 2012
rect 4273 1956 4275 2012
rect 3380 1954 4275 1956
rect 2960 1834 5162 1836
rect 2960 1778 2962 1834
rect 3018 1778 5104 1834
rect 5160 1778 5162 1834
rect 2960 1776 5162 1778
rect -30 1646 30 1706
rect 2646 1495 3524 1497
rect 2646 1439 2648 1495
rect 2704 1439 3466 1495
rect 3522 1439 3524 1495
rect 2646 1437 3524 1439
rect 2156 1159 3440 1161
rect 2156 1103 2158 1159
rect 2214 1103 3382 1159
rect 3438 1103 3440 1159
rect 2156 1101 3440 1103
rect 3296 902 6168 904
rect -30 808 30 868
rect 3296 846 3298 902
rect 3354 846 6110 902
rect 6166 846 6168 902
rect 3296 844 6168 846
rect 2156 573 3188 575
rect 2156 517 2158 573
rect 2214 517 3130 573
rect 3186 517 3188 573
rect 2156 515 3188 517
rect 2646 237 3272 239
rect 2646 181 2648 237
rect 2704 181 3214 237
rect 3270 181 3272 237
rect 2646 179 3272 181
rect -30 -30 30 30
use contact_17  contact_17_0
timestamp 1643593061
transform 1 0 4732 0 1 2861
box 0 0 1 1
use contact_13  contact_13_0
timestamp 1643593061
transform 1 0 4735 0 1 2864
box 0 0 1 1
use contact_18  contact_18_0
timestamp 1643593061
transform 1 0 4734 0 1 2857
box 0 0 1 1
use contact_17  contact_17_1
timestamp 1643593061
transform 1 0 4732 0 1 2861
box 0 0 1 1
use contact_13  contact_13_1
timestamp 1643593061
transform 1 0 4735 0 1 2864
box 0 0 1 1
use contact_26  contact_26_0
timestamp 1643593061
transform 1 0 3044 0 1 2857
box 0 0 1 1
use contact_13  contact_13_2
timestamp 1643593061
transform 1 0 3848 0 1 3021
box 0 0 1 1
use contact_17  contact_17_2
timestamp 1643593061
transform 1 0 3378 0 1 3018
box 0 0 1 1
use contact_13  contact_13_3
timestamp 1643593061
transform 1 0 3748 0 1 2781
box 0 0 1 1
use contact_17  contact_17_3
timestamp 1643593061
transform 1 0 3294 0 1 2778
box 0 0 1 1
use contact_17  contact_17_4
timestamp 1643593061
transform 1 0 5100 0 1 2115
box 0 0 1 1
use contact_13  contact_13_4
timestamp 1643593061
transform 1 0 5103 0 1 2118
box 0 0 1 1
use contact_26  contact_26_1
timestamp 1643593061
transform 1 0 2960 0 1 1776
box 0 0 1 1
use contact_26  contact_26_2
timestamp 1643593061
transform 1 0 5102 0 1 1776
box 0 0 1 1
use contact_18  contact_18_1
timestamp 1643593061
transform 1 0 4215 0 1 1954
box 0 0 1 1
use contact_17  contact_17_5
timestamp 1643593061
transform 1 0 4213 0 1 1958
box 0 0 1 1
use contact_13  contact_13_5
timestamp 1643593061
transform 1 0 4216 0 1 1961
box 0 0 1 1
use contact_18  contact_18_2
timestamp 1643593061
transform 1 0 4215 0 1 1954
box 0 0 1 1
use contact_17  contact_17_6
timestamp 1643593061
transform 1 0 4213 0 1 1958
box 0 0 1 1
use contact_13  contact_13_6
timestamp 1643593061
transform 1 0 4216 0 1 1961
box 0 0 1 1
use contact_26  contact_26_3
timestamp 1643593061
transform 1 0 3380 0 1 1954
box 0 0 1 1
use contact_13  contact_13_7
timestamp 1643593061
transform 1 0 3700 0 1 2114
box 0 0 1 1
use contact_17  contact_17_7
timestamp 1643593061
transform 1 0 3294 0 1 2111
box 0 0 1 1
use contact_17  contact_17_8
timestamp 1643593061
transform 1 0 6106 0 1 1183
box 0 0 1 1
use contact_13  contact_13_8
timestamp 1643593061
transform 1 0 6109 0 1 1186
box 0 0 1 1
use contact_17  contact_17_9
timestamp 1643593061
transform 1 0 6106 0 1 1183
box 0 0 1 1
use contact_13  contact_13_9
timestamp 1643593061
transform 1 0 6109 0 1 1186
box 0 0 1 1
use contact_26  contact_26_4
timestamp 1643593061
transform 1 0 3296 0 1 844
box 0 0 1 1
use contact_26  contact_26_5
timestamp 1643593061
transform 1 0 6108 0 1 844
box 0 0 1 1
use contact_17  contact_17_10
timestamp 1643593061
transform 1 0 3697 0 1 1189
box 0 0 1 1
use contact_13  contact_13_10
timestamp 1643593061
transform 1 0 3700 0 1 1192
box 0 0 1 1
use contact_17  contact_17_11
timestamp 1643593061
transform 1 0 4648 0 1 4541
box 0 0 1 1
use contact_13  contact_13_11
timestamp 1643593061
transform 1 0 4651 0 1 4544
box 0 0 1 1
use contact_13  contact_13_12
timestamp 1643593061
transform 1 0 3748 0 1 4457
box 0 0 1 1
use contact_17  contact_17_12
timestamp 1643593061
transform 1 0 3042 0 1 4454
box 0 0 1 1
use contact_17  contact_17_13
timestamp 1643593061
transform 1 0 4624 0 1 3791
box 0 0 1 1
use contact_13  contact_13_13
timestamp 1643593061
transform 1 0 4627 0 1 3794
box 0 0 1 1
use contact_13  contact_13_14
timestamp 1643593061
transform 1 0 3848 0 1 3637
box 0 0 1 1
use contact_17  contact_17_14
timestamp 1643593061
transform 1 0 2958 0 1 3634
box 0 0 1 1
use contact_13  contact_13_15
timestamp 1643593061
transform 1 0 3748 0 1 3877
box 0 0 1 1
use contact_17  contact_17_15
timestamp 1643593061
transform 1 0 3126 0 1 3874
box 0 0 1 1
use contact_17  contact_17_16
timestamp 1643593061
transform 1 0 5242 0 1 5463
box 0 0 1 1
use contact_13  contact_13_16
timestamp 1643593061
transform 1 0 5245 0 1 5466
box 0 0 1 1
use contact_13  contact_13_17
timestamp 1643593061
transform 1 0 3700 0 1 5466
box 0 0 1 1
use contact_17  contact_17_17
timestamp 1643593061
transform 1 0 2958 0 1 5463
box 0 0 1 1
use contact_17  contact_17_18
timestamp 1643593061
transform 1 0 3294 0 1 3246
box 0 0 1 1
use contact_17  contact_17_19
timestamp 1643593061
transform 1 0 -18 0 1 3246
box 0 0 1 1
use contact_18  contact_18_3
timestamp 1643593061
transform 1 0 2646 0 1 1437
box 0 0 1 1
use contact_26  contact_26_6
timestamp 1643593061
transform 1 0 3464 0 1 1437
box 0 0 1 1
use contact_18  contact_18_4
timestamp 1643593061
transform 1 0 2156 0 1 1101
box 0 0 1 1
use contact_26  contact_26_7
timestamp 1643593061
transform 1 0 3380 0 1 1101
box 0 0 1 1
use contact_18  contact_18_5
timestamp 1643593061
transform 1 0 2646 0 1 179
box 0 0 1 1
use contact_26  contact_26_8
timestamp 1643593061
transform 1 0 3212 0 1 179
box 0 0 1 1
use contact_18  contact_18_6
timestamp 1643593061
transform 1 0 2156 0 1 515
box 0 0 1 1
use contact_26  contact_26_9
timestamp 1643593061
transform 1 0 3128 0 1 515
box 0 0 1 1
use pdriver_3  pdriver_3_0
timestamp 1643593061
transform 1 0 4116 0 1 4190
box -36 -17 772 895
use pnand2_1  pnand2_1_0
timestamp 1643593061
transform 1 0 3648 0 1 4190
box -36 -17 504 895
use pand2_0  pand2_0_0
timestamp 1643593061
transform 1 0 3648 0 -1 4190
box -36 -17 1646 895
use pdriver_1  pdriver_1_0
timestamp 1643593061
transform 1 0 3648 0 -1 5866
box -36 -17 2048 895
use pand2  pand2_0
timestamp 1643593061
transform 1 0 3648 0 1 2514
box -36 -17 1862 895
use pand2  pand2_1
timestamp 1643593061
transform 1 0 4016 0 -1 2514
box -36 -17 1862 895
use pinv_3  pinv_3_0
timestamp 1643593061
transform 1 0 3648 0 -1 2514
box -36 -17 404 895
use pdriver_0  pdriver_0_0
timestamp 1643593061
transform 1 0 3648 0 1 838
box -36 -17 3344 895
use dff_buf_array  dff_buf_array_0
timestamp 1643593061
transform 1 0 0 0 1 0
box -32 -42 3012 1718
<< labels >>
rlabel metal2 s 180 1416 234 1444 4 csb
rlabel metal2 s 180 232 234 260 4 web
rlabel metal2 s 5274 5475 7124 5503 4 wl_en
rlabel metal2 s 4656 3803 7124 3831 4 w_en
rlabel metal2 s 4680 4553 7124 4581 4 p_en_bar
rlabel metal2 s 3715 1201 3743 1229 4 clk
rlabel metal2 s 6138 1195 7124 1223 4 clk_buf
rlabel metal3 s -30 -30 30 30 4 gnd
rlabel metal3 s -30 1646 30 1706 4 gnd
rlabel metal3 s -30 808 30 868 4 vdd
<< properties >>
string FIXED_BBOX 0 0 7124 160
string GDS_FILE sram_0rw2r1w_2_16_sky130A.gds
string GDS_END 488916
string GDS_START 480206
<< end >>
