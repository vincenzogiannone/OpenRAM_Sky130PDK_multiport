magic
tech sky130A
magscale 1 2
timestamp 1644951705
<< checkpaint >>
rect -1260 -1302 8912 50518
<< metal1 >>
rect 6018 48634 6312 48636
rect 6018 48608 6932 48634
rect 6284 48606 6932 48608
rect 7558 48536 7586 48564
rect 6018 48486 6630 48514
rect 7558 48410 7586 48438
rect 6018 48340 6452 48368
rect 7558 48184 7586 48212
rect 7558 47144 7586 47172
rect 6018 46988 6452 47016
rect 7558 46918 7586 46946
rect 6018 46842 6630 46870
rect 7558 46792 7586 46820
rect 6284 46748 6932 46750
rect 6018 46722 6932 46748
rect 6018 46720 6312 46722
rect 6018 45558 6312 45560
rect 6018 45532 6932 45558
rect 6284 45530 6932 45532
rect 7558 45460 7586 45488
rect 6018 45410 6630 45438
rect 7558 45334 7586 45362
rect 6018 45264 6452 45292
rect 7558 45108 7586 45136
rect 7558 44068 7586 44096
rect 6018 43912 6452 43940
rect 7558 43842 7586 43870
rect 6018 43766 6630 43794
rect 7558 43716 7586 43744
rect 6284 43672 6932 43674
rect 6018 43646 6932 43672
rect 6018 43644 6312 43646
rect 6018 42482 6312 42484
rect 6018 42456 6932 42482
rect 6284 42454 6932 42456
rect 7558 42384 7586 42412
rect 6018 42334 6630 42362
rect 7558 42258 7586 42286
rect 6018 42188 6452 42216
rect 7558 42032 7586 42060
rect 7558 40992 7586 41020
rect 6018 40836 6452 40864
rect 7558 40766 7586 40794
rect 6018 40690 6630 40718
rect 7558 40640 7586 40668
rect 6284 40596 6932 40598
rect 6018 40570 6932 40596
rect 6018 40568 6312 40570
rect 6018 39406 6312 39408
rect 6018 39380 6932 39406
rect 6284 39378 6932 39380
rect 7558 39308 7586 39336
rect 6018 39258 6630 39286
rect 7558 39182 7586 39210
rect 6018 39112 6452 39140
rect 7558 38956 7586 38984
rect 7558 37916 7586 37944
rect 6018 37760 6452 37788
rect 7558 37690 7586 37718
rect 6018 37614 6630 37642
rect 7558 37564 7586 37592
rect 6284 37520 6932 37522
rect 6018 37494 6932 37520
rect 6018 37492 6312 37494
rect 6018 36330 6312 36332
rect 6018 36304 6932 36330
rect 6284 36302 6932 36304
rect 7558 36232 7586 36260
rect 6018 36182 6630 36210
rect 7558 36106 7586 36134
rect 6018 36036 6452 36064
rect 7558 35880 7586 35908
rect 7558 34840 7586 34868
rect 6018 34684 6452 34712
rect 7558 34614 7586 34642
rect 6018 34538 6630 34566
rect 7558 34488 7586 34516
rect 6284 34444 6932 34446
rect 6018 34418 6932 34444
rect 6018 34416 6312 34418
rect 6018 33254 6312 33256
rect 6018 33228 6932 33254
rect 6284 33226 6932 33228
rect 7558 33156 7586 33184
rect 6018 33106 6630 33134
rect 7558 33030 7586 33058
rect 6018 32960 6452 32988
rect 7558 32804 7586 32832
rect 7558 31764 7586 31792
rect 6018 31608 6452 31636
rect 7558 31538 7586 31566
rect 6018 31462 6630 31490
rect 7558 31412 7586 31440
rect 6284 31368 6932 31370
rect 6018 31342 6932 31368
rect 6018 31340 6312 31342
rect 6018 30178 6312 30180
rect 6018 30152 6932 30178
rect 6284 30150 6932 30152
rect 7558 30080 7586 30108
rect 6018 30030 6630 30058
rect 7558 29954 7586 29982
rect 6018 29884 6452 29912
rect 7558 29728 7586 29756
rect 7558 28688 7586 28716
rect 6018 28532 6452 28560
rect 7558 28462 7586 28490
rect 6018 28386 6630 28414
rect 7558 28336 7586 28364
rect 6284 28292 6932 28294
rect 6018 28266 6932 28292
rect 6018 28264 6312 28266
rect 6018 27102 6312 27104
rect 6018 27076 6932 27102
rect 6284 27074 6932 27076
rect 7558 27004 7586 27032
rect 6018 26954 6630 26982
rect 7558 26878 7586 26906
rect 6018 26808 6452 26836
rect 7558 26652 7586 26680
rect 7558 25612 7586 25640
rect 6018 25456 6452 25484
rect 7558 25386 7586 25414
rect 6018 25310 6630 25338
rect 7558 25260 7586 25288
rect 6284 25216 6932 25218
rect 6018 25190 6932 25216
rect 6018 25188 6312 25190
rect 6018 24026 6312 24028
rect 6018 24000 6932 24026
rect 6284 23998 6932 24000
rect 7558 23928 7586 23956
rect 6018 23878 6630 23906
rect 7558 23802 7586 23830
rect 6018 23732 6452 23760
rect 7558 23576 7586 23604
rect 7558 22536 7586 22564
rect 6018 22380 6452 22408
rect 7558 22310 7586 22338
rect 6018 22234 6630 22262
rect 7558 22184 7586 22212
rect 6284 22140 6932 22142
rect 6018 22114 6932 22140
rect 6018 22112 6312 22114
rect 6018 20950 6312 20952
rect 6018 20924 6932 20950
rect 6284 20922 6932 20924
rect 7558 20852 7586 20880
rect 6018 20802 6630 20830
rect 7558 20726 7586 20754
rect 6018 20656 6452 20684
rect 7558 20500 7586 20528
rect 7558 19460 7586 19488
rect 6018 19304 6452 19332
rect 7558 19234 7586 19262
rect 6018 19158 6630 19186
rect 7558 19108 7586 19136
rect 6284 19064 6932 19066
rect 6018 19038 6932 19064
rect 6018 19036 6312 19038
rect 6018 17874 6312 17876
rect 6018 17848 6932 17874
rect 6284 17846 6932 17848
rect 7558 17776 7586 17804
rect 6018 17726 6630 17754
rect 7558 17650 7586 17678
rect 6018 17580 6452 17608
rect 7558 17424 7586 17452
rect 7558 16384 7586 16412
rect 6018 16228 6452 16256
rect 7558 16158 7586 16186
rect 6018 16082 6630 16110
rect 7558 16032 7586 16060
rect 6284 15988 6932 15990
rect 6018 15962 6932 15988
rect 6018 15960 6312 15962
rect 6018 14798 6312 14800
rect 6018 14772 6932 14798
rect 6284 14770 6932 14772
rect 7558 14700 7586 14728
rect 6018 14650 6630 14678
rect 7558 14574 7586 14602
rect 6018 14504 6452 14532
rect 7558 14348 7586 14376
rect 7558 13308 7586 13336
rect 6018 13152 6452 13180
rect 7558 13082 7586 13110
rect 6018 13006 6630 13034
rect 7558 12956 7586 12984
rect 6284 12912 6932 12914
rect 6018 12886 6932 12912
rect 6018 12884 6312 12886
rect 6018 11722 6312 11724
rect 6018 11696 6932 11722
rect 6284 11694 6932 11696
rect 7558 11624 7586 11652
rect 6018 11574 6630 11602
rect 7558 11498 7586 11526
rect 6018 11428 6452 11456
rect 7558 11272 7586 11300
rect 7558 10232 7586 10260
rect 6018 10076 6452 10104
rect 7558 10006 7586 10034
rect 6018 9930 6630 9958
rect 7558 9880 7586 9908
rect 6284 9836 6932 9838
rect 6018 9810 6932 9836
rect 6018 9808 6312 9810
rect 6018 8646 6312 8648
rect 6018 8620 6932 8646
rect 6284 8618 6932 8620
rect 7558 8548 7586 8576
rect 6018 8498 6630 8526
rect 7558 8422 7586 8450
rect 6018 8352 6452 8380
rect 7558 8196 7586 8224
rect 7558 7156 7586 7184
rect 6018 7000 6452 7028
rect 7558 6930 7586 6958
rect 6018 6854 6630 6882
rect 7558 6804 7586 6832
rect 6284 6760 6932 6762
rect 6018 6734 6932 6760
rect 6018 6732 6312 6734
rect 6018 5570 6312 5572
rect 6018 5544 6932 5570
rect 6284 5542 6932 5544
rect 7558 5472 7586 5500
rect 6018 5422 6630 5450
rect 7558 5346 7586 5374
rect 6018 5276 6452 5304
rect 7558 5120 7586 5148
rect 7558 4080 7586 4108
rect 6018 3924 6452 3952
rect 7558 3854 7586 3882
rect 6018 3778 6630 3806
rect 7558 3728 7586 3756
rect 6284 3684 6932 3686
rect 6018 3658 6932 3684
rect 6018 3656 6312 3658
rect 6018 2494 6312 2496
rect 6018 2468 6932 2494
rect 6284 2466 6932 2468
rect 7558 2396 7586 2424
rect 6018 2346 6630 2374
rect 7558 2270 7586 2298
rect 6018 2200 6452 2228
rect 7558 2044 7586 2072
rect 7558 1004 7586 1032
rect 6018 848 6452 876
rect 7558 778 7586 806
rect 6018 702 6630 730
rect 7558 652 7586 680
rect 6284 608 6932 610
rect 6018 582 6932 608
rect 6018 580 6312 582
<< metal2 >>
rect 6196 49202 6410 49230
rect 18 0 46 30792
rect 102 0 130 30792
rect 186 0 214 30792
rect 270 0 298 30792
rect 354 0 382 30792
rect 438 0 466 30792
rect 522 0 550 30792
<< metal3 >>
rect 5980 49179 6112 49253
rect 7520 49179 7652 49253
rect 5980 47641 6112 47715
rect 7520 47641 7652 47715
rect 5980 46103 6112 46177
rect 7520 46103 7652 46177
rect 5980 44565 6112 44639
rect 7520 44565 7652 44639
rect 5980 43027 6112 43101
rect 7520 43027 7652 43101
rect 5980 41489 6112 41563
rect 7520 41489 7652 41563
rect 5980 39951 6112 40025
rect 7520 39951 7652 40025
rect 5980 38413 6112 38487
rect 7520 38413 7652 38487
rect 5980 36875 6112 36949
rect 7520 36875 7652 36949
rect 5980 35337 6112 35411
rect 7520 35337 7652 35411
rect 5980 33799 6112 33873
rect 7520 33799 7652 33873
rect 5980 32261 6112 32335
rect 7520 32261 7652 32335
rect 960 30755 1092 30829
rect 2000 30755 2132 30829
rect 5980 30723 6112 30797
rect 7520 30723 7652 30797
rect 960 29215 1092 29289
rect 2000 29215 2132 29289
rect 5980 29185 6112 29259
rect 7520 29185 7652 29259
rect 960 27675 1092 27749
rect 2000 27675 2132 27749
rect 5980 27647 6112 27721
rect 7520 27647 7652 27721
rect 960 26135 1092 26209
rect 2000 26135 2132 26209
rect 5980 26109 6112 26183
rect 7520 26109 7652 26183
rect 960 24595 1092 24669
rect 2000 24595 2132 24669
rect 5980 24571 6112 24645
rect 7520 24571 7652 24645
rect 960 23055 1092 23129
rect 2000 23055 2132 23129
rect 5980 23033 6112 23107
rect 7520 23033 7652 23107
rect 960 21515 1092 21589
rect 2000 21515 2132 21589
rect 5980 21495 6112 21569
rect 7520 21495 7652 21569
rect 960 19975 1092 20049
rect 2000 19975 2132 20049
rect 5980 19957 6112 20031
rect 7520 19957 7652 20031
rect 960 18435 1092 18509
rect 2000 18435 2132 18509
rect 5980 18419 6112 18493
rect 7520 18419 7652 18493
rect 5980 16881 6112 16955
rect 7520 16881 7652 16955
rect 1308 15359 1440 15433
rect 2180 15359 2312 15433
rect 5980 15343 6112 15417
rect 7520 15343 7652 15417
rect 1308 13819 1440 13893
rect 2180 13819 2312 13893
rect 5980 13805 6112 13879
rect 7520 13805 7652 13879
rect 1308 12279 1440 12353
rect 2180 12279 2312 12353
rect 5980 12267 6112 12341
rect 7520 12267 7652 12341
rect 1308 10739 1440 10813
rect 2180 10739 2312 10813
rect 5980 10729 6112 10803
rect 7520 10729 7652 10803
rect 1308 9199 1440 9273
rect 2180 9199 2312 9273
rect 5980 9191 6112 9265
rect 7520 9191 7652 9265
rect 5980 7653 6112 7727
rect 7520 7653 7652 7727
rect 1308 6123 1440 6197
rect 2180 6123 2312 6197
rect 5980 6115 6112 6189
rect 7520 6115 7652 6189
rect 1308 4583 1440 4657
rect 2180 4583 2312 4657
rect 5980 4577 6112 4651
rect 7520 4577 7652 4651
rect 1308 3043 1440 3117
rect 2180 3043 2312 3117
rect 5980 3039 6112 3113
rect 7520 3039 7652 3113
rect 1308 1503 1440 1577
rect 2180 1503 2312 1577
rect 5980 1501 6112 1575
rect 7520 1501 7652 1575
rect 1308 -37 1440 37
rect 2180 -37 2312 37
rect 5980 -37 6112 37
rect 7520 -37 7652 37
use wordline_driver_array  wordline_driver_array_0
timestamp 1644951705
transform 1 0 6382 0 1 0
box 0 -42 1270 49258
use hierarchical_decoder  hierarchical_decoder_0
timestamp 1644951705
transform 1 0 0 0 1 0
box 0 -42 6112 49258
<< labels >>
rlabel metal2 s 18 0 46 30792 4 addr0
rlabel metal2 s 102 0 130 30792 4 addr1
rlabel metal2 s 186 0 214 30792 4 addr2
rlabel metal2 s 270 0 298 30792 4 addr3
rlabel metal2 s 354 0 382 30792 4 addr4
rlabel metal2 s 438 0 466 30792 4 addr5
rlabel metal2 s 522 0 550 30792 4 addr6
rlabel metal1 s 7558 778 7586 806 4 rwl0_0
rlabel metal1 s 7558 1004 7586 1032 4 rwl1_0
rlabel metal1 s 7558 652 7586 680 4 wwl0_0
rlabel metal1 s 7558 2270 7586 2298 4 rwl0_1
rlabel metal1 s 7558 2044 7586 2072 4 rwl1_1
rlabel metal1 s 7558 2396 7586 2424 4 wwl0_1
rlabel metal1 s 7558 3854 7586 3882 4 rwl0_2
rlabel metal1 s 7558 4080 7586 4108 4 rwl1_2
rlabel metal1 s 7558 3728 7586 3756 4 wwl0_2
rlabel metal1 s 7558 5346 7586 5374 4 rwl0_3
rlabel metal1 s 7558 5120 7586 5148 4 rwl1_3
rlabel metal1 s 7558 5472 7586 5500 4 wwl0_3
rlabel metal1 s 7558 6930 7586 6958 4 rwl0_4
rlabel metal1 s 7558 7156 7586 7184 4 rwl1_4
rlabel metal1 s 7558 6804 7586 6832 4 wwl0_4
rlabel metal1 s 7558 8422 7586 8450 4 rwl0_5
rlabel metal1 s 7558 8196 7586 8224 4 rwl1_5
rlabel metal1 s 7558 8548 7586 8576 4 wwl0_5
rlabel metal1 s 7558 10006 7586 10034 4 rwl0_6
rlabel metal1 s 7558 10232 7586 10260 4 rwl1_6
rlabel metal1 s 7558 9880 7586 9908 4 wwl0_6
rlabel metal1 s 7558 11498 7586 11526 4 rwl0_7
rlabel metal1 s 7558 11272 7586 11300 4 rwl1_7
rlabel metal1 s 7558 11624 7586 11652 4 wwl0_7
rlabel metal1 s 7558 13082 7586 13110 4 rwl0_8
rlabel metal1 s 7558 13308 7586 13336 4 rwl1_8
rlabel metal1 s 7558 12956 7586 12984 4 wwl0_8
rlabel metal1 s 7558 14574 7586 14602 4 rwl0_9
rlabel metal1 s 7558 14348 7586 14376 4 rwl1_9
rlabel metal1 s 7558 14700 7586 14728 4 wwl0_9
rlabel metal1 s 7558 16158 7586 16186 4 rwl0_10
rlabel metal1 s 7558 16384 7586 16412 4 rwl1_10
rlabel metal1 s 7558 16032 7586 16060 4 wwl0_10
rlabel metal1 s 7558 17650 7586 17678 4 rwl0_11
rlabel metal1 s 7558 17424 7586 17452 4 rwl1_11
rlabel metal1 s 7558 17776 7586 17804 4 wwl0_11
rlabel metal1 s 7558 19234 7586 19262 4 rwl0_12
rlabel metal1 s 7558 19460 7586 19488 4 rwl1_12
rlabel metal1 s 7558 19108 7586 19136 4 wwl0_12
rlabel metal1 s 7558 20726 7586 20754 4 rwl0_13
rlabel metal1 s 7558 20500 7586 20528 4 rwl1_13
rlabel metal1 s 7558 20852 7586 20880 4 wwl0_13
rlabel metal1 s 7558 22310 7586 22338 4 rwl0_14
rlabel metal1 s 7558 22536 7586 22564 4 rwl1_14
rlabel metal1 s 7558 22184 7586 22212 4 wwl0_14
rlabel metal1 s 7558 23802 7586 23830 4 rwl0_15
rlabel metal1 s 7558 23576 7586 23604 4 rwl1_15
rlabel metal1 s 7558 23928 7586 23956 4 wwl0_15
rlabel metal1 s 7558 25386 7586 25414 4 rwl0_16
rlabel metal1 s 7558 25612 7586 25640 4 rwl1_16
rlabel metal1 s 7558 25260 7586 25288 4 wwl0_16
rlabel metal1 s 7558 26878 7586 26906 4 rwl0_17
rlabel metal1 s 7558 26652 7586 26680 4 rwl1_17
rlabel metal1 s 7558 27004 7586 27032 4 wwl0_17
rlabel metal1 s 7558 28462 7586 28490 4 rwl0_18
rlabel metal1 s 7558 28688 7586 28716 4 rwl1_18
rlabel metal1 s 7558 28336 7586 28364 4 wwl0_18
rlabel metal1 s 7558 29954 7586 29982 4 rwl0_19
rlabel metal1 s 7558 29728 7586 29756 4 rwl1_19
rlabel metal1 s 7558 30080 7586 30108 4 wwl0_19
rlabel metal1 s 7558 31538 7586 31566 4 rwl0_20
rlabel metal1 s 7558 31764 7586 31792 4 rwl1_20
rlabel metal1 s 7558 31412 7586 31440 4 wwl0_20
rlabel metal1 s 7558 33030 7586 33058 4 rwl0_21
rlabel metal1 s 7558 32804 7586 32832 4 rwl1_21
rlabel metal1 s 7558 33156 7586 33184 4 wwl0_21
rlabel metal1 s 7558 34614 7586 34642 4 rwl0_22
rlabel metal1 s 7558 34840 7586 34868 4 rwl1_22
rlabel metal1 s 7558 34488 7586 34516 4 wwl0_22
rlabel metal1 s 7558 36106 7586 36134 4 rwl0_23
rlabel metal1 s 7558 35880 7586 35908 4 rwl1_23
rlabel metal1 s 7558 36232 7586 36260 4 wwl0_23
rlabel metal1 s 7558 37690 7586 37718 4 rwl0_24
rlabel metal1 s 7558 37916 7586 37944 4 rwl1_24
rlabel metal1 s 7558 37564 7586 37592 4 wwl0_24
rlabel metal1 s 7558 39182 7586 39210 4 rwl0_25
rlabel metal1 s 7558 38956 7586 38984 4 rwl1_25
rlabel metal1 s 7558 39308 7586 39336 4 wwl0_25
rlabel metal1 s 7558 40766 7586 40794 4 rwl0_26
rlabel metal1 s 7558 40992 7586 41020 4 rwl1_26
rlabel metal1 s 7558 40640 7586 40668 4 wwl0_26
rlabel metal1 s 7558 42258 7586 42286 4 rwl0_27
rlabel metal1 s 7558 42032 7586 42060 4 rwl1_27
rlabel metal1 s 7558 42384 7586 42412 4 wwl0_27
rlabel metal1 s 7558 43842 7586 43870 4 rwl0_28
rlabel metal1 s 7558 44068 7586 44096 4 rwl1_28
rlabel metal1 s 7558 43716 7586 43744 4 wwl0_28
rlabel metal1 s 7558 45334 7586 45362 4 rwl0_29
rlabel metal1 s 7558 45108 7586 45136 4 rwl1_29
rlabel metal1 s 7558 45460 7586 45488 4 wwl0_29
rlabel metal1 s 7558 46918 7586 46946 4 rwl0_30
rlabel metal1 s 7558 47144 7586 47172 4 rwl1_30
rlabel metal1 s 7558 46792 7586 46820 4 wwl0_30
rlabel metal1 s 7558 48410 7586 48438 4 rwl0_31
rlabel metal1 s 7558 48184 7586 48212 4 rwl1_31
rlabel metal1 s 7558 48536 7586 48564 4 wwl0_31
rlabel metal2 s 6382 49202 6410 49230 4 wl_en
rlabel metal3 s 7520 32261 7652 32335 4 vdd
rlabel metal3 s 7520 29185 7652 29259 4 vdd
rlabel metal3 s 7520 1501 7652 1575 4 vdd
rlabel metal3 s 7520 26109 7652 26183 4 vdd
rlabel metal3 s 960 29215 1092 29289 4 vdd
rlabel metal3 s 5980 35337 6112 35411 4 vdd
rlabel metal3 s 5980 23033 6112 23107 4 vdd
rlabel metal3 s 5980 41489 6112 41563 4 vdd
rlabel metal3 s 7520 23033 7652 23107 4 vdd
rlabel metal3 s 7520 35337 7652 35411 4 vdd
rlabel metal3 s 7520 44565 7652 44639 4 vdd
rlabel metal3 s 5980 47641 6112 47715 4 vdd
rlabel metal3 s 7520 13805 7652 13879 4 vdd
rlabel metal3 s 5980 29185 6112 29259 4 vdd
rlabel metal3 s 5980 19957 6112 20031 4 vdd
rlabel metal3 s 5980 26109 6112 26183 4 vdd
rlabel metal3 s 1308 1503 1440 1577 4 vdd
rlabel metal3 s 7520 19957 7652 20031 4 vdd
rlabel metal3 s 5980 7653 6112 7727 4 vdd
rlabel metal3 s 2000 29215 2132 29289 4 vdd
rlabel metal3 s 5980 44565 6112 44639 4 vdd
rlabel metal3 s 7520 41489 7652 41563 4 vdd
rlabel metal3 s 5980 16881 6112 16955 4 vdd
rlabel metal3 s 2180 13819 2312 13893 4 vdd
rlabel metal3 s 7520 4577 7652 4651 4 vdd
rlabel metal3 s 5980 32261 6112 32335 4 vdd
rlabel metal3 s 7520 38413 7652 38487 4 vdd
rlabel metal3 s 2000 26135 2132 26209 4 vdd
rlabel metal3 s 5980 1501 6112 1575 4 vdd
rlabel metal3 s 960 19975 1092 20049 4 vdd
rlabel metal3 s 2180 10739 2312 10813 4 vdd
rlabel metal3 s 1308 4583 1440 4657 4 vdd
rlabel metal3 s 5980 10729 6112 10803 4 vdd
rlabel metal3 s 2000 23055 2132 23129 4 vdd
rlabel metal3 s 2000 19975 2132 20049 4 vdd
rlabel metal3 s 5980 13805 6112 13879 4 vdd
rlabel metal3 s 1308 13819 1440 13893 4 vdd
rlabel metal3 s 5980 38413 6112 38487 4 vdd
rlabel metal3 s 7520 47641 7652 47715 4 vdd
rlabel metal3 s 7520 10729 7652 10803 4 vdd
rlabel metal3 s 960 26135 1092 26209 4 vdd
rlabel metal3 s 2180 4583 2312 4657 4 vdd
rlabel metal3 s 5980 4577 6112 4651 4 vdd
rlabel metal3 s 960 23055 1092 23129 4 vdd
rlabel metal3 s 7520 7653 7652 7727 4 vdd
rlabel metal3 s 2180 1503 2312 1577 4 vdd
rlabel metal3 s 1308 10739 1440 10813 4 vdd
rlabel metal3 s 7520 16881 7652 16955 4 vdd
rlabel metal3 s 5980 49179 6112 49253 4 gnd
rlabel metal3 s 7520 43027 7652 43101 4 gnd
rlabel metal3 s 2000 18435 2132 18509 4 gnd
rlabel metal3 s 960 30755 1092 30829 4 gnd
rlabel metal3 s 5980 33799 6112 33873 4 gnd
rlabel metal3 s 5980 39951 6112 40025 4 gnd
rlabel metal3 s 1308 3043 1440 3117 4 gnd
rlabel metal3 s 5980 15343 6112 15417 4 gnd
rlabel metal3 s 2000 30755 2132 30829 4 gnd
rlabel metal3 s 2180 3043 2312 3117 4 gnd
rlabel metal3 s 5980 24571 6112 24645 4 gnd
rlabel metal3 s 7520 15343 7652 15417 4 gnd
rlabel metal3 s 2180 6123 2312 6197 4 gnd
rlabel metal3 s 5980 27647 6112 27721 4 gnd
rlabel metal3 s 5980 -37 6112 37 4 gnd
rlabel metal3 s 7520 18419 7652 18493 4 gnd
rlabel metal3 s 7520 27647 7652 27721 4 gnd
rlabel metal3 s 7520 30723 7652 30797 4 gnd
rlabel metal3 s 2000 27675 2132 27749 4 gnd
rlabel metal3 s 5980 43027 6112 43101 4 gnd
rlabel metal3 s 5980 3039 6112 3113 4 gnd
rlabel metal3 s 7520 3039 7652 3113 4 gnd
rlabel metal3 s 7520 9191 7652 9265 4 gnd
rlabel metal3 s 7520 46103 7652 46177 4 gnd
rlabel metal3 s 7520 49179 7652 49253 4 gnd
rlabel metal3 s 7520 24571 7652 24645 4 gnd
rlabel metal3 s 5980 36875 6112 36949 4 gnd
rlabel metal3 s 5980 12267 6112 12341 4 gnd
rlabel metal3 s 7520 21495 7652 21569 4 gnd
rlabel metal3 s 5980 9191 6112 9265 4 gnd
rlabel metal3 s 7520 39951 7652 40025 4 gnd
rlabel metal3 s 7520 6115 7652 6189 4 gnd
rlabel metal3 s 960 18435 1092 18509 4 gnd
rlabel metal3 s 7520 33799 7652 33873 4 gnd
rlabel metal3 s 1308 12279 1440 12353 4 gnd
rlabel metal3 s 960 24595 1092 24669 4 gnd
rlabel metal3 s 960 27675 1092 27749 4 gnd
rlabel metal3 s 2180 -37 2312 37 4 gnd
rlabel metal3 s 7520 -37 7652 37 4 gnd
rlabel metal3 s 5980 18419 6112 18493 4 gnd
rlabel metal3 s 5980 46103 6112 46177 4 gnd
rlabel metal3 s 1308 -37 1440 37 4 gnd
rlabel metal3 s 2000 24595 2132 24669 4 gnd
rlabel metal3 s 2180 12279 2312 12353 4 gnd
rlabel metal3 s 5980 30723 6112 30797 4 gnd
rlabel metal3 s 960 21515 1092 21589 4 gnd
rlabel metal3 s 2180 9199 2312 9273 4 gnd
rlabel metal3 s 2180 15359 2312 15433 4 gnd
rlabel metal3 s 1308 9199 1440 9273 4 gnd
rlabel metal3 s 5980 21495 6112 21569 4 gnd
rlabel metal3 s 7520 12267 7652 12341 4 gnd
rlabel metal3 s 1308 15359 1440 15433 4 gnd
rlabel metal3 s 1308 6123 1440 6197 4 gnd
rlabel metal3 s 2000 21515 2132 21589 4 gnd
rlabel metal3 s 5980 6115 6112 6189 4 gnd
rlabel metal3 s 7520 36875 7652 36949 4 gnd
<< properties >>
string FIXED_BBOX 0 0 7622 49244
string GDS_FILE sram_0rw2r1w_16_128_sky130A.gds
string GDS_END 1667940
string GDS_START 1597894
<< end >>
