magic
tech sky130A
magscale 1 2
timestamp 1643671299
<< checkpaint >>
rect -1260 -1260 25298 2212
<< metal1 >>
rect 0 356 24038 384
<< via1 >>
rect 323 848 375 900
rect 1879 848 1931 900
rect 3435 848 3487 900
rect 4991 848 5043 900
rect 6547 848 6599 900
rect 8103 848 8155 900
rect 9659 848 9711 900
rect 11215 848 11267 900
rect 12771 848 12823 900
rect 14327 848 14379 900
rect 15883 848 15935 900
rect 17439 848 17491 900
rect 18995 848 19047 900
rect 20551 848 20603 900
rect 22107 848 22159 900
rect 23663 848 23715 900
rect 323 16 375 68
rect 1879 16 1931 68
rect 3435 16 3487 68
rect 4991 16 5043 68
rect 6547 16 6599 68
rect 8103 16 8155 68
rect 9659 16 9711 68
rect 11215 16 11267 68
rect 12771 16 12823 68
rect 14327 16 14379 68
rect 15883 16 15935 68
rect 17439 16 17491 68
rect 18995 16 19047 68
rect 20551 16 20603 68
rect 22107 16 22159 68
rect 23663 16 23715 68
<< metal2 >>
rect 329 902 369 908
rect 329 840 369 846
rect 630 322 658 952
rect 1885 902 1925 908
rect 1885 840 1925 846
rect 2186 322 2214 952
rect 3441 902 3481 908
rect 3441 840 3481 846
rect 3742 322 3770 952
rect 4997 902 5037 908
rect 4997 840 5037 846
rect 5298 322 5326 952
rect 6553 902 6593 908
rect 6553 840 6593 846
rect 6854 322 6882 952
rect 8109 902 8149 908
rect 8109 840 8149 846
rect 8410 322 8438 952
rect 9665 902 9705 908
rect 9665 840 9705 846
rect 9966 322 9994 952
rect 11221 902 11261 908
rect 11221 840 11261 846
rect 11522 322 11550 952
rect 12777 902 12817 908
rect 12777 840 12817 846
rect 13078 322 13106 952
rect 14333 902 14373 908
rect 14333 840 14373 846
rect 14634 322 14662 952
rect 15889 902 15929 908
rect 15889 840 15929 846
rect 16190 322 16218 952
rect 17445 902 17485 908
rect 17445 840 17485 846
rect 17746 322 17774 952
rect 19001 902 19041 908
rect 19001 840 19041 846
rect 19302 322 19330 952
rect 20557 902 20597 908
rect 20557 840 20597 846
rect 20858 322 20886 952
rect 22113 902 22153 908
rect 22113 840 22153 846
rect 22414 322 22442 952
rect 23669 902 23709 908
rect 23669 840 23709 846
rect 23970 322 23998 952
rect 196 272 250 300
rect 1752 272 1806 300
rect 3308 272 3362 300
rect 4864 272 4918 300
rect 6420 272 6474 300
rect 7976 272 8030 300
rect 9532 272 9586 300
rect 11088 272 11142 300
rect 12644 272 12698 300
rect 14200 272 14254 300
rect 15756 272 15810 300
rect 17312 272 17366 300
rect 18868 272 18922 300
rect 20424 272 20478 300
rect 21980 272 22034 300
rect 23536 272 23590 300
rect 329 70 369 76
rect 1885 70 1925 76
rect 3441 70 3481 76
rect 4997 70 5037 76
rect 6553 70 6593 76
rect 8109 70 8149 76
rect 9665 70 9705 76
rect 11221 70 11261 76
rect 12777 70 12817 76
rect 14333 70 14373 76
rect 15889 70 15929 76
rect 17445 70 17485 76
rect 19001 70 19041 76
rect 20557 70 20597 76
rect 22113 70 22153 76
rect 23669 70 23709 76
rect 329 8 369 14
rect 1885 8 1925 14
rect 3441 8 3481 14
rect 4997 8 5037 14
rect 6553 8 6593 14
rect 8109 8 8149 14
rect 9665 8 9705 14
rect 11221 8 11261 14
rect 12777 8 12817 14
rect 14333 8 14373 14
rect 15889 8 15929 14
rect 17445 8 17485 14
rect 19001 8 19041 14
rect 20557 8 20597 14
rect 22113 8 22153 14
rect 23669 8 23709 14
<< via2 >>
rect 321 900 377 902
rect 321 848 323 900
rect 323 848 375 900
rect 375 848 377 900
rect 321 846 377 848
rect 1877 900 1933 902
rect 1877 848 1879 900
rect 1879 848 1931 900
rect 1931 848 1933 900
rect 1877 846 1933 848
rect 3433 900 3489 902
rect 3433 848 3435 900
rect 3435 848 3487 900
rect 3487 848 3489 900
rect 3433 846 3489 848
rect 4989 900 5045 902
rect 4989 848 4991 900
rect 4991 848 5043 900
rect 5043 848 5045 900
rect 4989 846 5045 848
rect 6545 900 6601 902
rect 6545 848 6547 900
rect 6547 848 6599 900
rect 6599 848 6601 900
rect 6545 846 6601 848
rect 8101 900 8157 902
rect 8101 848 8103 900
rect 8103 848 8155 900
rect 8155 848 8157 900
rect 8101 846 8157 848
rect 9657 900 9713 902
rect 9657 848 9659 900
rect 9659 848 9711 900
rect 9711 848 9713 900
rect 9657 846 9713 848
rect 11213 900 11269 902
rect 11213 848 11215 900
rect 11215 848 11267 900
rect 11267 848 11269 900
rect 11213 846 11269 848
rect 12769 900 12825 902
rect 12769 848 12771 900
rect 12771 848 12823 900
rect 12823 848 12825 900
rect 12769 846 12825 848
rect 14325 900 14381 902
rect 14325 848 14327 900
rect 14327 848 14379 900
rect 14379 848 14381 900
rect 14325 846 14381 848
rect 15881 900 15937 902
rect 15881 848 15883 900
rect 15883 848 15935 900
rect 15935 848 15937 900
rect 15881 846 15937 848
rect 17437 900 17493 902
rect 17437 848 17439 900
rect 17439 848 17491 900
rect 17491 848 17493 900
rect 17437 846 17493 848
rect 18993 900 19049 902
rect 18993 848 18995 900
rect 18995 848 19047 900
rect 19047 848 19049 900
rect 18993 846 19049 848
rect 20549 900 20605 902
rect 20549 848 20551 900
rect 20551 848 20603 900
rect 20603 848 20605 900
rect 20549 846 20605 848
rect 22105 900 22161 902
rect 22105 848 22107 900
rect 22107 848 22159 900
rect 22159 848 22161 900
rect 22105 846 22161 848
rect 23661 900 23717 902
rect 23661 848 23663 900
rect 23663 848 23715 900
rect 23715 848 23717 900
rect 23661 846 23717 848
rect 321 68 377 70
rect 321 16 323 68
rect 323 16 375 68
rect 375 16 377 68
rect 321 14 377 16
rect 1877 68 1933 70
rect 1877 16 1879 68
rect 1879 16 1931 68
rect 1931 16 1933 68
rect 1877 14 1933 16
rect 3433 68 3489 70
rect 3433 16 3435 68
rect 3435 16 3487 68
rect 3487 16 3489 68
rect 3433 14 3489 16
rect 4989 68 5045 70
rect 4989 16 4991 68
rect 4991 16 5043 68
rect 5043 16 5045 68
rect 4989 14 5045 16
rect 6545 68 6601 70
rect 6545 16 6547 68
rect 6547 16 6599 68
rect 6599 16 6601 68
rect 6545 14 6601 16
rect 8101 68 8157 70
rect 8101 16 8103 68
rect 8103 16 8155 68
rect 8155 16 8157 68
rect 8101 14 8157 16
rect 9657 68 9713 70
rect 9657 16 9659 68
rect 9659 16 9711 68
rect 9711 16 9713 68
rect 9657 14 9713 16
rect 11213 68 11269 70
rect 11213 16 11215 68
rect 11215 16 11267 68
rect 11267 16 11269 68
rect 11213 14 11269 16
rect 12769 68 12825 70
rect 12769 16 12771 68
rect 12771 16 12823 68
rect 12823 16 12825 68
rect 12769 14 12825 16
rect 14325 68 14381 70
rect 14325 16 14327 68
rect 14327 16 14379 68
rect 14379 16 14381 68
rect 14325 14 14381 16
rect 15881 68 15937 70
rect 15881 16 15883 68
rect 15883 16 15935 68
rect 15935 16 15937 68
rect 15881 14 15937 16
rect 17437 68 17493 70
rect 17437 16 17439 68
rect 17439 16 17491 68
rect 17491 16 17493 68
rect 17437 14 17493 16
rect 18993 68 19049 70
rect 18993 16 18995 68
rect 18995 16 19047 68
rect 19047 16 19049 68
rect 18993 14 19049 16
rect 20549 68 20605 70
rect 20549 16 20551 68
rect 20551 16 20603 68
rect 20603 16 20605 68
rect 20549 14 20605 16
rect 22105 68 22161 70
rect 22105 16 22107 68
rect 22107 16 22159 68
rect 22159 16 22161 68
rect 22105 14 22161 16
rect 23661 68 23717 70
rect 23661 16 23663 68
rect 23663 16 23715 68
rect 23715 16 23717 68
rect 23661 14 23717 16
<< metal3 >>
rect 319 902 379 904
rect 319 846 321 902
rect 377 846 379 902
rect 319 844 379 846
rect 1875 902 1935 904
rect 1875 846 1877 902
rect 1933 846 1935 902
rect 1875 844 1935 846
rect 3431 902 3491 904
rect 3431 846 3433 902
rect 3489 846 3491 902
rect 3431 844 3491 846
rect 4987 902 5047 904
rect 4987 846 4989 902
rect 5045 846 5047 902
rect 4987 844 5047 846
rect 6543 902 6603 904
rect 6543 846 6545 902
rect 6601 846 6603 902
rect 6543 844 6603 846
rect 8099 902 8159 904
rect 8099 846 8101 902
rect 8157 846 8159 902
rect 8099 844 8159 846
rect 9655 902 9715 904
rect 9655 846 9657 902
rect 9713 846 9715 902
rect 9655 844 9715 846
rect 11211 902 11271 904
rect 11211 846 11213 902
rect 11269 846 11271 902
rect 11211 844 11271 846
rect 12767 902 12827 904
rect 12767 846 12769 902
rect 12825 846 12827 902
rect 12767 844 12827 846
rect 14323 902 14383 904
rect 14323 846 14325 902
rect 14381 846 14383 902
rect 14323 844 14383 846
rect 15879 902 15939 904
rect 15879 846 15881 902
rect 15937 846 15939 902
rect 15879 844 15939 846
rect 17435 902 17495 904
rect 17435 846 17437 902
rect 17493 846 17495 902
rect 17435 844 17495 846
rect 18991 902 19051 904
rect 18991 846 18993 902
rect 19049 846 19051 902
rect 18991 844 19051 846
rect 20547 902 20607 904
rect 20547 846 20549 902
rect 20605 846 20607 902
rect 20547 844 20607 846
rect 22103 902 22163 904
rect 22103 846 22105 902
rect 22161 846 22163 902
rect 22103 844 22163 846
rect 23659 902 23719 904
rect 23659 846 23661 902
rect 23717 846 23719 902
rect 23659 844 23719 846
rect 319 70 379 72
rect 319 14 321 70
rect 377 14 379 70
rect 319 12 379 14
rect 1875 70 1935 72
rect 1875 14 1877 70
rect 1933 14 1935 70
rect 1875 12 1935 14
rect 3431 70 3491 72
rect 3431 14 3433 70
rect 3489 14 3491 70
rect 3431 12 3491 14
rect 4987 70 5047 72
rect 4987 14 4989 70
rect 5045 14 5047 70
rect 4987 12 5047 14
rect 6543 70 6603 72
rect 6543 14 6545 70
rect 6601 14 6603 70
rect 6543 12 6603 14
rect 8099 70 8159 72
rect 8099 14 8101 70
rect 8157 14 8159 70
rect 8099 12 8159 14
rect 9655 70 9715 72
rect 9655 14 9657 70
rect 9713 14 9715 70
rect 9655 12 9715 14
rect 11211 70 11271 72
rect 11211 14 11213 70
rect 11269 14 11271 70
rect 11211 12 11271 14
rect 12767 70 12827 72
rect 12767 14 12769 70
rect 12825 14 12827 70
rect 12767 12 12827 14
rect 14323 70 14383 72
rect 14323 14 14325 70
rect 14381 14 14383 70
rect 14323 12 14383 14
rect 15879 70 15939 72
rect 15879 14 15881 70
rect 15937 14 15939 70
rect 15879 12 15939 14
rect 17435 70 17495 72
rect 17435 14 17437 70
rect 17493 14 17495 70
rect 17435 12 17495 14
rect 18991 70 19051 72
rect 18991 14 18993 70
rect 19049 14 19051 70
rect 18991 12 19051 14
rect 20547 70 20607 72
rect 20547 14 20549 70
rect 20605 14 20607 70
rect 20547 12 20607 14
rect 22103 70 22163 72
rect 22103 14 22105 70
rect 22161 14 22163 70
rect 22103 12 22163 14
rect 23659 70 23719 72
rect 23659 14 23661 70
rect 23717 14 23719 70
rect 23659 12 23719 14
use contact_23  contact_23_0
timestamp 1643671299
transform 1 0 23659 0 1 12
box 0 0 1 1
use contact_22  contact_22_0
timestamp 1643671299
transform 1 0 23674 0 1 27
box 0 0 1 1
use contact_23  contact_23_1
timestamp 1643671299
transform 1 0 23659 0 1 844
box 0 0 1 1
use contact_22  contact_22_1
timestamp 1643671299
transform 1 0 23674 0 1 859
box 0 0 1 1
use contact_23  contact_23_2
timestamp 1643671299
transform 1 0 22103 0 1 12
box 0 0 1 1
use contact_22  contact_22_2
timestamp 1643671299
transform 1 0 22118 0 1 27
box 0 0 1 1
use contact_23  contact_23_3
timestamp 1643671299
transform 1 0 22103 0 1 844
box 0 0 1 1
use contact_22  contact_22_3
timestamp 1643671299
transform 1 0 22118 0 1 859
box 0 0 1 1
use contact_23  contact_23_4
timestamp 1643671299
transform 1 0 20547 0 1 12
box 0 0 1 1
use contact_22  contact_22_4
timestamp 1643671299
transform 1 0 20562 0 1 27
box 0 0 1 1
use contact_23  contact_23_5
timestamp 1643671299
transform 1 0 20547 0 1 844
box 0 0 1 1
use contact_22  contact_22_5
timestamp 1643671299
transform 1 0 20562 0 1 859
box 0 0 1 1
use contact_23  contact_23_6
timestamp 1643671299
transform 1 0 18991 0 1 12
box 0 0 1 1
use contact_22  contact_22_6
timestamp 1643671299
transform 1 0 19006 0 1 27
box 0 0 1 1
use contact_23  contact_23_7
timestamp 1643671299
transform 1 0 18991 0 1 844
box 0 0 1 1
use contact_22  contact_22_7
timestamp 1643671299
transform 1 0 19006 0 1 859
box 0 0 1 1
use contact_23  contact_23_8
timestamp 1643671299
transform 1 0 17435 0 1 12
box 0 0 1 1
use contact_22  contact_22_8
timestamp 1643671299
transform 1 0 17450 0 1 27
box 0 0 1 1
use contact_23  contact_23_9
timestamp 1643671299
transform 1 0 17435 0 1 844
box 0 0 1 1
use contact_22  contact_22_9
timestamp 1643671299
transform 1 0 17450 0 1 859
box 0 0 1 1
use contact_23  contact_23_10
timestamp 1643671299
transform 1 0 15879 0 1 12
box 0 0 1 1
use contact_22  contact_22_10
timestamp 1643671299
transform 1 0 15894 0 1 27
box 0 0 1 1
use contact_23  contact_23_11
timestamp 1643671299
transform 1 0 15879 0 1 844
box 0 0 1 1
use contact_22  contact_22_11
timestamp 1643671299
transform 1 0 15894 0 1 859
box 0 0 1 1
use contact_23  contact_23_12
timestamp 1643671299
transform 1 0 14323 0 1 12
box 0 0 1 1
use contact_22  contact_22_12
timestamp 1643671299
transform 1 0 14338 0 1 27
box 0 0 1 1
use contact_23  contact_23_13
timestamp 1643671299
transform 1 0 14323 0 1 844
box 0 0 1 1
use contact_22  contact_22_13
timestamp 1643671299
transform 1 0 14338 0 1 859
box 0 0 1 1
use contact_23  contact_23_14
timestamp 1643671299
transform 1 0 12767 0 1 12
box 0 0 1 1
use contact_22  contact_22_14
timestamp 1643671299
transform 1 0 12782 0 1 27
box 0 0 1 1
use contact_23  contact_23_15
timestamp 1643671299
transform 1 0 12767 0 1 844
box 0 0 1 1
use contact_22  contact_22_15
timestamp 1643671299
transform 1 0 12782 0 1 859
box 0 0 1 1
use contact_23  contact_23_16
timestamp 1643671299
transform 1 0 11211 0 1 12
box 0 0 1 1
use contact_22  contact_22_16
timestamp 1643671299
transform 1 0 11226 0 1 27
box 0 0 1 1
use contact_23  contact_23_17
timestamp 1643671299
transform 1 0 11211 0 1 844
box 0 0 1 1
use contact_22  contact_22_17
timestamp 1643671299
transform 1 0 11226 0 1 859
box 0 0 1 1
use contact_23  contact_23_18
timestamp 1643671299
transform 1 0 9655 0 1 12
box 0 0 1 1
use contact_22  contact_22_18
timestamp 1643671299
transform 1 0 9670 0 1 27
box 0 0 1 1
use contact_23  contact_23_19
timestamp 1643671299
transform 1 0 9655 0 1 844
box 0 0 1 1
use contact_22  contact_22_19
timestamp 1643671299
transform 1 0 9670 0 1 859
box 0 0 1 1
use contact_23  contact_23_20
timestamp 1643671299
transform 1 0 8099 0 1 12
box 0 0 1 1
use contact_22  contact_22_20
timestamp 1643671299
transform 1 0 8114 0 1 27
box 0 0 1 1
use contact_23  contact_23_21
timestamp 1643671299
transform 1 0 8099 0 1 844
box 0 0 1 1
use contact_22  contact_22_21
timestamp 1643671299
transform 1 0 8114 0 1 859
box 0 0 1 1
use contact_23  contact_23_22
timestamp 1643671299
transform 1 0 6543 0 1 12
box 0 0 1 1
use contact_22  contact_22_22
timestamp 1643671299
transform 1 0 6558 0 1 27
box 0 0 1 1
use contact_23  contact_23_23
timestamp 1643671299
transform 1 0 6543 0 1 844
box 0 0 1 1
use contact_22  contact_22_23
timestamp 1643671299
transform 1 0 6558 0 1 859
box 0 0 1 1
use contact_23  contact_23_24
timestamp 1643671299
transform 1 0 4987 0 1 12
box 0 0 1 1
use contact_22  contact_22_24
timestamp 1643671299
transform 1 0 5002 0 1 27
box 0 0 1 1
use contact_23  contact_23_25
timestamp 1643671299
transform 1 0 4987 0 1 844
box 0 0 1 1
use contact_22  contact_22_25
timestamp 1643671299
transform 1 0 5002 0 1 859
box 0 0 1 1
use contact_23  contact_23_26
timestamp 1643671299
transform 1 0 3431 0 1 12
box 0 0 1 1
use contact_22  contact_22_26
timestamp 1643671299
transform 1 0 3446 0 1 27
box 0 0 1 1
use contact_23  contact_23_27
timestamp 1643671299
transform 1 0 3431 0 1 844
box 0 0 1 1
use contact_22  contact_22_27
timestamp 1643671299
transform 1 0 3446 0 1 859
box 0 0 1 1
use contact_23  contact_23_28
timestamp 1643671299
transform 1 0 1875 0 1 12
box 0 0 1 1
use contact_22  contact_22_28
timestamp 1643671299
transform 1 0 1890 0 1 27
box 0 0 1 1
use contact_23  contact_23_29
timestamp 1643671299
transform 1 0 1875 0 1 844
box 0 0 1 1
use contact_22  contact_22_29
timestamp 1643671299
transform 1 0 1890 0 1 859
box 0 0 1 1
use contact_23  contact_23_30
timestamp 1643671299
transform 1 0 319 0 1 12
box 0 0 1 1
use contact_22  contact_22_30
timestamp 1643671299
transform 1 0 334 0 1 27
box 0 0 1 1
use contact_23  contact_23_31
timestamp 1643671299
transform 1 0 319 0 1 844
box 0 0 1 1
use contact_22  contact_22_31
timestamp 1643671299
transform 1 0 334 0 1 859
box 0 0 1 1
use write_driver_multiport  write_driver_multiport_0
timestamp 1643671299
transform 1 0 23340 0 1 0
box 0 0 698 952
use write_driver_multiport  write_driver_multiport_1
timestamp 1643671299
transform 1 0 21784 0 1 0
box 0 0 698 952
use write_driver_multiport  write_driver_multiport_2
timestamp 1643671299
transform 1 0 20228 0 1 0
box 0 0 698 952
use write_driver_multiport  write_driver_multiport_3
timestamp 1643671299
transform 1 0 18672 0 1 0
box 0 0 698 952
use write_driver_multiport  write_driver_multiport_4
timestamp 1643671299
transform 1 0 17116 0 1 0
box 0 0 698 952
use write_driver_multiport  write_driver_multiport_5
timestamp 1643671299
transform 1 0 15560 0 1 0
box 0 0 698 952
use write_driver_multiport  write_driver_multiport_6
timestamp 1643671299
transform 1 0 14004 0 1 0
box 0 0 698 952
use write_driver_multiport  write_driver_multiport_7
timestamp 1643671299
transform 1 0 12448 0 1 0
box 0 0 698 952
use write_driver_multiport  write_driver_multiport_8
timestamp 1643671299
transform 1 0 10892 0 1 0
box 0 0 698 952
use write_driver_multiport  write_driver_multiport_9
timestamp 1643671299
transform 1 0 9336 0 1 0
box 0 0 698 952
use write_driver_multiport  write_driver_multiport_10
timestamp 1643671299
transform 1 0 7780 0 1 0
box 0 0 698 952
use write_driver_multiport  write_driver_multiport_11
timestamp 1643671299
transform 1 0 6224 0 1 0
box 0 0 698 952
use write_driver_multiport  write_driver_multiport_12
timestamp 1643671299
transform 1 0 4668 0 1 0
box 0 0 698 952
use write_driver_multiport  write_driver_multiport_13
timestamp 1643671299
transform 1 0 3112 0 1 0
box 0 0 698 952
use write_driver_multiport  write_driver_multiport_14
timestamp 1643671299
transform 1 0 1556 0 1 0
box 0 0 698 952
use write_driver_multiport  write_driver_multiport_15
timestamp 1643671299
transform 1 0 0 0 1 0
box 0 0 698 952
<< labels >>
rlabel metal2 s 196 272 250 300 4 din_0
rlabel metal2 s 630 322 658 952 4 wbl0_0
rlabel metal3 s 12767 844 12827 904 4 vdd
rlabel metal3 s 11211 844 11271 904 4 vdd
rlabel metal3 s 14323 844 14383 904 4 vdd
rlabel metal3 s 20547 844 20607 904 4 vdd
rlabel metal3 s 9655 844 9715 904 4 vdd
rlabel metal3 s 319 844 379 904 4 vdd
rlabel metal3 s 4987 844 5047 904 4 vdd
rlabel metal3 s 1875 844 1935 904 4 vdd
rlabel metal3 s 8099 844 8159 904 4 vdd
rlabel metal3 s 23659 844 23719 904 4 vdd
rlabel metal3 s 3431 844 3491 904 4 vdd
rlabel metal3 s 17435 844 17495 904 4 vdd
rlabel metal3 s 18991 844 19051 904 4 vdd
rlabel metal3 s 15879 844 15939 904 4 vdd
rlabel metal3 s 6543 844 6603 904 4 vdd
rlabel metal3 s 22103 844 22163 904 4 vdd
rlabel metal3 s 319 12 379 72 4 gnd
rlabel metal3 s 3431 12 3491 72 4 gnd
rlabel metal3 s 8099 12 8159 72 4 gnd
rlabel metal3 s 14323 12 14383 72 4 gnd
rlabel metal3 s 18991 12 19051 72 4 gnd
rlabel metal3 s 1875 12 1935 72 4 gnd
rlabel metal3 s 6543 12 6603 72 4 gnd
rlabel metal3 s 22103 12 22163 72 4 gnd
rlabel metal3 s 9655 12 9715 72 4 gnd
rlabel metal3 s 11211 12 11271 72 4 gnd
rlabel metal3 s 12767 12 12827 72 4 gnd
rlabel metal3 s 20547 12 20607 72 4 gnd
rlabel metal3 s 23659 12 23719 72 4 gnd
rlabel metal3 s 15879 12 15939 72 4 gnd
rlabel metal3 s 17435 12 17495 72 4 gnd
rlabel metal3 s 4987 12 5047 72 4 gnd
rlabel metal2 s 1752 272 1806 300 4 din_1
rlabel metal2 s 2186 322 2214 952 4 wbl0_1
rlabel metal2 s 3308 272 3362 300 4 din_2
rlabel metal2 s 3742 322 3770 952 4 wbl0_2
rlabel metal2 s 4864 272 4918 300 4 din_3
rlabel metal2 s 5298 322 5326 952 4 wbl0_3
rlabel metal2 s 6420 272 6474 300 4 din_4
rlabel metal2 s 6854 322 6882 952 4 wbl0_4
rlabel metal2 s 7976 272 8030 300 4 din_5
rlabel metal2 s 8410 322 8438 952 4 wbl0_5
rlabel metal2 s 9532 272 9586 300 4 din_6
rlabel metal2 s 9966 322 9994 952 4 wbl0_6
rlabel metal2 s 11088 272 11142 300 4 din_7
rlabel metal2 s 11522 322 11550 952 4 wbl0_7
rlabel metal2 s 12644 272 12698 300 4 din_8
rlabel metal2 s 13078 322 13106 952 4 wbl0_8
rlabel metal2 s 14200 272 14254 300 4 din_9
rlabel metal2 s 14634 322 14662 952 4 wbl0_9
rlabel metal2 s 15756 272 15810 300 4 din_10
rlabel metal2 s 16190 322 16218 952 4 wbl0_10
rlabel metal2 s 17312 272 17366 300 4 din_11
rlabel metal2 s 17746 322 17774 952 4 wbl0_11
rlabel metal2 s 18868 272 18922 300 4 din_12
rlabel metal2 s 19302 322 19330 952 4 wbl0_12
rlabel metal2 s 20424 272 20478 300 4 din_13
rlabel metal2 s 20858 322 20886 952 4 wbl0_13
rlabel metal2 s 21980 272 22034 300 4 din_14
rlabel metal2 s 22414 322 22442 952 4 wbl0_14
rlabel metal2 s 23536 272 23590 300 4 din_15
rlabel metal2 s 23970 322 23998 952 4 wbl0_15
rlabel metal1 s 0 356 24038 384 4 en
<< properties >>
string FIXED_BBOX 0 0 24038 952
string GDS_FILE sram_0rw2r1w_16_32_sky130A.gds
string GDS_END 837744
string GDS_START 820008
<< end >>
