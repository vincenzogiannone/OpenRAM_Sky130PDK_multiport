magic
tech sky130A
magscale 1 2
timestamp 1643593061
<< checkpaint >>
rect -1260 -1260 2736 2212
<< metal1 >>
rect 323 900 375 906
rect 323 842 375 848
rect 1101 900 1153 906
rect 1101 842 1153 848
rect 0 356 1476 384
rect 323 68 375 74
rect 323 10 375 16
rect 1101 68 1153 74
rect 1101 10 1153 16
<< via1 >>
rect 323 848 375 900
rect 1101 848 1153 900
rect 323 16 375 68
rect 1101 16 1153 68
<< metal2 >>
rect 630 322 658 952
rect 1408 322 1436 952
rect 196 272 250 300
rect 974 272 1028 300
<< via2 >>
rect 321 900 377 902
rect 321 848 323 900
rect 323 848 375 900
rect 375 848 377 900
rect 321 846 377 848
rect 1099 900 1155 902
rect 1099 848 1101 900
rect 1101 848 1153 900
rect 1153 848 1155 900
rect 1099 846 1155 848
rect 321 68 377 70
rect 321 16 323 68
rect 323 16 375 68
rect 375 16 377 68
rect 321 14 377 16
rect 1099 68 1155 70
rect 1099 16 1101 68
rect 1101 16 1153 68
rect 1153 16 1155 68
rect 1099 14 1155 16
<< metal3 >>
rect 319 902 379 904
rect 319 846 321 902
rect 377 846 379 902
rect 319 844 379 846
rect 1097 902 1157 904
rect 1097 846 1099 902
rect 1155 846 1157 902
rect 1097 844 1157 846
rect 319 70 379 72
rect 319 14 321 70
rect 377 14 379 70
rect 319 12 379 14
rect 1097 70 1157 72
rect 1097 14 1099 70
rect 1155 14 1157 70
rect 1097 12 1157 14
use contact_23  contact_23_0
timestamp 1643593061
transform 1 0 1097 0 1 12
box 0 0 1 1
use contact_22  contact_22_0
timestamp 1643593061
transform 1 0 1101 0 1 10
box 0 0 1 1
use contact_23  contact_23_1
timestamp 1643593061
transform 1 0 1097 0 1 844
box 0 0 1 1
use contact_22  contact_22_1
timestamp 1643593061
transform 1 0 1101 0 1 842
box 0 0 1 1
use contact_23  contact_23_2
timestamp 1643593061
transform 1 0 319 0 1 12
box 0 0 1 1
use contact_22  contact_22_2
timestamp 1643593061
transform 1 0 323 0 1 10
box 0 0 1 1
use contact_23  contact_23_3
timestamp 1643593061
transform 1 0 319 0 1 844
box 0 0 1 1
use contact_22  contact_22_3
timestamp 1643593061
transform 1 0 323 0 1 842
box 0 0 1 1
use write_driver_multiport  write_driver_multiport_0
timestamp 1643593061
transform 1 0 778 0 1 0
box 0 0 698 952
use write_driver_multiport  write_driver_multiport_1
timestamp 1643593061
transform 1 0 0 0 1 0
box 0 0 698 952
<< labels >>
rlabel metal2 s 196 272 250 300 4 din_0
rlabel metal2 s 630 322 658 952 4 wbl0_0
rlabel metal3 s 1097 844 1157 904 4 vdd
rlabel metal3 s 319 844 379 904 4 vdd
rlabel metal3 s 1097 12 1157 72 4 gnd
rlabel metal3 s 319 12 379 72 4 gnd
rlabel metal2 s 974 272 1028 300 4 din_1
rlabel metal2 s 1408 322 1436 952 4 wbl0_1
rlabel metal1 s 0 356 1476 384 4 en
<< properties >>
string FIXED_BBOX 0 0 1476 952
string GDS_FILE sram_0rw2r1w_2_16_sky130A.gds
string GDS_END 263762
string GDS_START 261270
<< end >>
