magic
tech sky130A
magscale 1 2
timestamp 1643678851
<< checkpaint >>
rect -1296 -1277 2098 2857
<< locali >>
rect 0 1523 802 1557
rect 330 745 364 1263
rect 330 711 532 745
rect 630 711 664 745
rect 196 505 262 571
rect 96 257 162 323
rect 0 -17 802 17
use pinv  pinv_0
timestamp 1643678851
transform 1 0 451 0 1 0
box -36 -17 387 1597
use pnand2  pnand2_0
timestamp 1643678851
transform 1 0 0 0 1 0
box -36 -17 487 1597
<< labels >>
rlabel locali s 647 728 647 728 4 Z
rlabel locali s 129 290 129 290 4 A
rlabel locali s 229 538 229 538 4 B
rlabel locali s 401 0 401 0 4 gnd
rlabel locali s 401 1540 401 1540 4 vdd
<< properties >>
string FIXED_BBOX 0 0 802 1540
string GDS_FILE sram_0rw2r1w_16_128_sky130A.gds
string GDS_END 1852922
string GDS_START 1851924
<< end >>
