magic
tech sky130A
magscale 1 2
timestamp 1644951705
<< checkpaint >>
rect -1260 -1260 77096 65648
<< metal2 >>
rect 13657 18230 13713 18239
rect 13657 18165 13713 18174
rect 14737 18226 14793 18235
rect 14737 18161 14793 18170
rect 13657 17738 13713 17747
rect 13657 17673 13713 17682
rect 14737 17742 14793 17751
rect 14737 17677 14793 17686
rect 13657 16554 13713 16563
rect 13657 16489 13713 16498
rect 14737 16550 14793 16559
rect 14737 16485 14793 16494
rect 13657 16062 13713 16071
rect 13657 15997 13713 16006
rect 14737 16066 14793 16075
rect 14737 16001 14793 16010
rect 13657 14878 13713 14887
rect 13657 14813 13713 14822
rect 14737 14874 14793 14883
rect 14737 14809 14793 14818
rect 13657 14386 13713 14395
rect 13657 14321 13713 14330
rect 14737 14390 14793 14399
rect 14737 14325 14793 14334
rect 13366 13264 13422 13273
rect 13366 13199 13422 13208
rect 13657 13202 13713 13211
rect 15146 13207 15174 28156
rect 15230 14399 15258 28156
rect 15314 14883 15342 28156
rect 15398 16075 15426 28156
rect 15482 16559 15510 28156
rect 15566 17751 15594 28156
rect 15650 18235 15678 28156
rect 15636 18226 15692 18235
rect 15636 18161 15692 18170
rect 15552 17742 15608 17751
rect 15552 17677 15608 17686
rect 15468 16550 15524 16559
rect 15468 16485 15524 16494
rect 15384 16066 15440 16075
rect 15384 16001 15440 16010
rect 15300 14874 15356 14883
rect 15300 14809 15356 14818
rect 15216 14390 15272 14399
rect 15216 14325 15272 14334
rect 2959 8228 3015 8237
rect 2959 8163 3015 8172
rect 6481 8013 6537 8022
rect 13380 7991 13408 13199
rect 13657 13137 13713 13146
rect 14737 13198 14793 13207
rect 14737 13133 14793 13142
rect 15132 13198 15188 13207
rect 15132 13133 15188 13142
rect 21510 12300 21538 61976
rect 14932 12291 14988 12300
rect 14932 12226 14988 12235
rect 21496 12291 21552 12300
rect 21496 12226 21552 12235
rect 14932 11358 14988 11367
rect 14932 11293 14988 11302
rect 22632 10626 22660 12354
rect 73092 11358 73148 11367
rect 23309 11296 23365 11305
rect 23309 11231 23365 11240
rect 23581 11296 23637 11305
rect 23581 11231 23637 11240
rect 26421 11296 26477 11305
rect 26421 11231 26477 11240
rect 26693 11296 26749 11305
rect 26693 11231 26749 11240
rect 29533 11296 29589 11305
rect 29533 11231 29589 11240
rect 29805 11296 29861 11305
rect 29805 11231 29861 11240
rect 32645 11296 32701 11305
rect 32645 11231 32701 11240
rect 32917 11296 32973 11305
rect 32917 11231 32973 11240
rect 35757 11296 35813 11305
rect 35757 11231 35813 11240
rect 36029 11296 36085 11305
rect 36029 11231 36085 11240
rect 38869 11296 38925 11305
rect 38869 11231 38925 11240
rect 39141 11296 39197 11305
rect 39141 11231 39197 11240
rect 41981 11296 42037 11305
rect 41981 11231 42037 11240
rect 42253 11296 42309 11305
rect 42253 11231 42309 11240
rect 45093 11296 45149 11305
rect 45093 11231 45149 11240
rect 45365 11296 45421 11305
rect 73092 11293 73148 11302
rect 45365 11231 45421 11240
rect 14932 10617 14988 10626
rect 14932 10552 14988 10561
rect 22618 10617 22674 10626
rect 22618 10552 22674 10561
rect 12464 7977 13408 7991
rect 12464 7963 13460 7977
rect 6481 7948 6537 7957
rect 2959 7044 3015 7053
rect 2959 6979 3015 6988
rect 13328 3038 13460 7963
rect 73106 6210 73134 11293
rect 13328 3010 13366 3038
rect 13422 3010 13460 3038
rect 13366 2973 13422 2982
rect 16621 2976 16677 2985
rect 16621 2911 16677 2920
rect 18103 2976 18159 2985
rect 18103 2911 18159 2920
rect 19585 2976 19641 2985
rect 19585 2911 19641 2920
rect 21067 2976 21123 2985
rect 21067 2911 21123 2920
rect 22549 2976 22605 2985
rect 22549 2911 22605 2920
rect 24031 2976 24087 2985
rect 24031 2911 24087 2920
rect 25513 2976 25569 2985
rect 25513 2911 25569 2920
rect 26995 2976 27051 2985
rect 26995 2911 27051 2920
rect 28477 2976 28533 2985
rect 28477 2911 28533 2920
rect 29959 2976 30015 2985
rect 29959 2911 30015 2920
rect 31441 2976 31497 2985
rect 31441 2911 31497 2920
rect 32923 2976 32979 2985
rect 32923 2911 32979 2920
rect 34405 2976 34461 2985
rect 34405 2911 34461 2920
rect 35887 2976 35943 2985
rect 35887 2911 35943 2920
rect 37369 2976 37425 2985
rect 37369 2911 37425 2920
rect 38851 2976 38907 2985
rect 38851 2911 38907 2920
rect 40333 2976 40389 2985
rect 40333 2911 40389 2920
rect 41815 2976 41871 2985
rect 41815 2911 41871 2920
<< via2 >>
rect 13657 18174 13713 18230
rect 14737 18170 14793 18226
rect 13657 17682 13713 17738
rect 14737 17686 14793 17742
rect 13657 16498 13713 16554
rect 14737 16494 14793 16550
rect 13657 16006 13713 16062
rect 14737 16010 14793 16066
rect 13657 14822 13713 14878
rect 14737 14818 14793 14874
rect 13657 14330 13713 14386
rect 14737 14334 14793 14390
rect 13366 13208 13422 13264
rect 15636 18170 15692 18226
rect 15552 17686 15608 17742
rect 15468 16494 15524 16550
rect 15384 16010 15440 16066
rect 15300 14818 15356 14874
rect 15216 14334 15272 14390
rect 2959 8172 3015 8228
rect 6481 7957 6537 8013
rect 13657 13146 13713 13202
rect 14737 13142 14793 13198
rect 15132 13142 15188 13198
rect 14932 12235 14988 12291
rect 21496 12235 21552 12291
rect 14932 11302 14988 11358
rect 23309 11240 23365 11296
rect 23581 11240 23637 11296
rect 26421 11240 26477 11296
rect 26693 11240 26749 11296
rect 29533 11240 29589 11296
rect 29805 11240 29861 11296
rect 32645 11240 32701 11296
rect 32917 11240 32973 11296
rect 35757 11240 35813 11296
rect 36029 11240 36085 11296
rect 38869 11240 38925 11296
rect 39141 11240 39197 11296
rect 41981 11240 42037 11296
rect 42253 11240 42309 11296
rect 45093 11240 45149 11296
rect 45365 11240 45421 11296
rect 73092 11302 73148 11358
rect 14932 10561 14988 10617
rect 22618 10561 22674 10617
rect 2959 6988 3015 7044
rect 13366 2982 13422 3038
rect 16621 2920 16677 2976
rect 18103 2920 18159 2976
rect 19585 2920 19641 2976
rect 21067 2920 21123 2976
rect 22549 2920 22605 2976
rect 24031 2920 24087 2976
rect 25513 2920 25569 2976
rect 26995 2920 27051 2976
rect 28477 2920 28533 2976
rect 29959 2920 30015 2976
rect 31441 2920 31497 2976
rect 32923 2920 32979 2976
rect 34405 2920 34461 2976
rect 35887 2920 35943 2976
rect 37369 2920 37425 2976
rect 38851 2920 38907 2976
rect 40333 2920 40389 2976
rect 41815 2920 41871 2976
<< metal3 >>
rect 424 64344 75836 64388
rect 424 64280 468 64344
rect 532 64280 680 64344
rect 744 64280 892 64344
rect 956 64280 75304 64344
rect 75368 64280 75516 64344
rect 75580 64280 75728 64344
rect 75792 64280 75836 64344
rect 424 64132 75836 64280
rect 424 64068 468 64132
rect 532 64068 680 64132
rect 744 64068 892 64132
rect 956 64068 75304 64132
rect 75368 64068 75516 64132
rect 75580 64068 75728 64132
rect 75792 64068 75836 64132
rect 424 63920 75836 64068
rect 424 63856 468 63920
rect 532 63856 680 63920
rect 744 63856 892 63920
rect 956 63856 21032 63920
rect 21096 63856 75304 63920
rect 75368 63856 75516 63920
rect 75580 63856 75728 63920
rect 75792 63856 75836 63920
rect 424 63812 75836 63856
rect 1484 63284 74776 63328
rect 1484 63220 1528 63284
rect 1592 63220 1740 63284
rect 1804 63220 1952 63284
rect 2016 63220 74244 63284
rect 74308 63220 74456 63284
rect 74520 63220 74668 63284
rect 74732 63220 74776 63284
rect 1484 63072 74776 63220
rect 1484 63008 1528 63072
rect 1592 63008 1740 63072
rect 1804 63008 1952 63072
rect 2016 63008 74244 63072
rect 74308 63008 74456 63072
rect 74520 63008 74668 63072
rect 74732 63008 74776 63072
rect 1484 62860 74776 63008
rect 1484 62796 1528 62860
rect 1592 62796 1740 62860
rect 1804 62796 1952 62860
rect 2016 62796 22728 62860
rect 22792 62796 74244 62860
rect 74308 62796 74456 62860
rect 74520 62796 74668 62860
rect 74732 62796 74776 62860
rect 1484 62752 74776 62796
rect 20988 62012 22972 62056
rect 20988 61948 21032 62012
rect 21096 61948 22940 62012
rect 23004 61948 23048 62012
rect 20988 61904 22972 61948
rect 20988 60360 21352 60572
rect 22472 60528 22836 60572
rect 22472 60464 22728 60528
rect 22792 60464 22836 60528
rect 22472 60360 22836 60464
rect 20988 60316 22836 60360
rect 20988 60252 22516 60316
rect 22580 60252 22836 60316
rect 20988 60208 22836 60252
rect 20988 59044 23048 59088
rect 20988 58980 22940 59044
rect 23004 58980 23048 59044
rect 20988 58936 23048 58980
rect 20988 58832 21352 58936
rect 20988 58768 21032 58832
rect 21096 58768 21352 58832
rect 20988 58724 21352 58768
rect 22472 58724 22836 58936
rect 20988 57392 21352 57604
rect 22472 57560 22836 57604
rect 22472 57496 22516 57560
rect 22580 57496 22836 57560
rect 22472 57392 22836 57496
rect 20988 57348 22836 57392
rect 20988 57284 21244 57348
rect 21308 57284 22836 57348
rect 20988 57240 22836 57284
rect 20988 55864 22836 55908
rect 20988 55800 21032 55864
rect 21096 55800 22836 55864
rect 20988 55756 22836 55800
rect 20988 55652 21140 55756
rect 20988 55588 21032 55652
rect 21096 55588 21140 55652
rect 20988 55544 21140 55588
rect 20988 54380 22836 54424
rect 20988 54316 21244 54380
rect 21308 54316 22836 54380
rect 20988 54272 22836 54316
rect 20988 54060 21352 54272
rect 22472 54168 22836 54272
rect 22472 54104 22516 54168
rect 22580 54104 22836 54168
rect 22472 54060 22836 54104
rect 20988 52896 21352 52940
rect 20988 52832 21032 52896
rect 21096 52832 21352 52896
rect 20988 52728 21352 52832
rect 22472 52728 22836 52940
rect 20988 52684 22836 52728
rect 20988 52620 21244 52684
rect 21308 52620 22836 52684
rect 20988 52576 22836 52620
rect 20988 51244 21352 51456
rect 22472 51412 22836 51456
rect 22472 51348 22516 51412
rect 22580 51348 22836 51412
rect 22472 51244 22836 51348
rect 20988 51200 22836 51244
rect 20988 51136 21032 51200
rect 21096 51136 22836 51200
rect 20988 51092 22836 51136
rect 21200 49928 21352 49972
rect 21200 49864 21244 49928
rect 21308 49864 21352 49928
rect 21200 49760 21352 49864
rect 20988 49716 22836 49760
rect 20988 49652 21244 49716
rect 21308 49652 22836 49716
rect 20988 49608 22836 49652
rect 20988 48232 22836 48276
rect 20988 48168 21032 48232
rect 21096 48168 22836 48232
rect 20988 48124 22836 48168
rect 20988 47912 21352 48124
rect 22472 48020 22836 48124
rect 22472 47956 22516 48020
rect 22580 47956 22836 48020
rect 22472 47912 22836 47956
rect 20988 46748 21352 46792
rect 20988 46684 21244 46748
rect 21308 46684 21352 46748
rect 20988 46580 21352 46684
rect 22472 46580 22836 46792
rect 20988 46536 22836 46580
rect 20988 46472 21244 46536
rect 21308 46472 22836 46536
rect 20988 46428 22836 46472
rect 20988 45052 22836 45096
rect 20988 44988 21032 45052
rect 21096 44988 22516 45052
rect 22580 44988 22836 45052
rect 20988 44944 22836 44988
rect 15900 43568 17324 43612
rect 15900 43504 16156 43568
rect 16220 43504 17324 43568
rect 15900 43460 17324 43504
rect 20988 43568 22836 43612
rect 20988 43504 21244 43568
rect 21308 43504 22728 43568
rect 22792 43504 22836 43568
rect 20988 43460 22836 43504
rect 15900 41916 16264 42128
rect 16960 41916 17324 42128
rect 15900 41872 17324 41916
rect 15900 41808 17216 41872
rect 17280 41808 17324 41872
rect 15900 41764 17324 41808
rect 20988 42084 22836 42128
rect 20988 42020 21032 42084
rect 21096 42020 22836 42084
rect 20988 41976 22836 42020
rect 20988 41764 21352 41976
rect 22472 41872 22836 41976
rect 22472 41808 22516 41872
rect 22580 41808 22836 41872
rect 22472 41764 22836 41808
rect 15900 40600 17324 40644
rect 15900 40536 16156 40600
rect 16220 40536 17324 40600
rect 15900 40492 17324 40536
rect 15900 40388 16264 40492
rect 15900 40324 15944 40388
rect 16008 40324 16264 40388
rect 15900 40280 16264 40324
rect 16960 40280 17324 40492
rect 20988 40432 21352 40644
rect 22472 40600 22836 40644
rect 22472 40536 22728 40600
rect 22792 40536 22836 40600
rect 22472 40432 22836 40536
rect 20988 40388 22972 40432
rect 20988 40324 22940 40388
rect 23004 40324 23048 40388
rect 20988 40280 22972 40324
rect 15900 39116 17324 39160
rect 15900 39052 17216 39116
rect 17280 39052 17324 39116
rect 15900 39008 17324 39052
rect 15900 38796 16264 39008
rect 16960 38904 17324 39008
rect 16960 38840 17216 38904
rect 17280 38840 17324 38904
rect 16960 38796 17324 38840
rect 20988 38904 22836 38948
rect 20988 38840 22516 38904
rect 22580 38840 22728 38904
rect 22792 38840 22836 38904
rect 20988 38796 22836 38840
rect 16112 37524 17112 37676
rect 16112 37464 16264 37524
rect 16960 37464 17112 37524
rect 15900 37420 16688 37464
rect 15900 37356 15944 37420
rect 16008 37356 16580 37420
rect 16644 37356 16688 37420
rect 15900 37312 16688 37356
rect 16960 37312 17324 37464
rect 20988 37420 23048 37464
rect 20988 37356 21032 37420
rect 21096 37356 22940 37420
rect 23004 37356 23048 37420
rect 20988 37312 23048 37356
rect 15900 35936 17324 35980
rect 15900 35872 17216 35936
rect 17280 35872 17324 35936
rect 15900 35828 17324 35872
rect 15900 35616 16264 35828
rect 16960 35768 17324 35828
rect 20988 35768 21352 35980
rect 22472 35936 22836 35980
rect 22472 35872 22728 35936
rect 22792 35872 22836 35936
rect 22472 35768 22836 35872
rect 16824 35724 17960 35768
rect 16748 35660 16792 35724
rect 16856 35660 17960 35724
rect 16824 35616 17960 35660
rect 17808 35556 17960 35616
rect 20988 35724 22836 35768
rect 20988 35660 22516 35724
rect 22580 35660 22836 35724
rect 20988 35616 22836 35660
rect 20988 35556 21140 35616
rect 17808 35404 21140 35556
rect 15900 34284 16264 34496
rect 16612 34452 17324 34496
rect 16536 34388 16580 34452
rect 16644 34388 17324 34452
rect 16612 34344 17324 34388
rect 16960 34284 17324 34344
rect 15900 34240 17324 34284
rect 15900 34176 16156 34240
rect 16220 34176 17324 34240
rect 15900 34132 17324 34176
rect 20988 34452 22836 34496
rect 20988 34388 21032 34452
rect 21096 34388 22836 34452
rect 20988 34344 22836 34388
rect 20988 34132 21352 34344
rect 22472 34284 22836 34344
rect 22336 34240 22836 34284
rect 22260 34176 22304 34240
rect 22368 34176 22836 34240
rect 22336 34132 22836 34176
rect 15900 32860 17324 33012
rect 15900 32800 16264 32860
rect 15900 32756 16900 32800
rect 15900 32692 16792 32756
rect 16856 32692 16900 32756
rect 15900 32648 16900 32692
rect 16960 32648 17324 32860
rect 20988 32756 22836 32800
rect 20988 32692 22516 32756
rect 22580 32692 22728 32756
rect 22792 32692 22836 32756
rect 20988 32648 22836 32692
rect 15900 31272 17324 31316
rect 15900 31208 16156 31272
rect 16220 31208 17216 31272
rect 17280 31208 17324 31272
rect 15900 31164 17324 31208
rect 20988 31272 22972 31316
rect 20988 31208 22516 31272
rect 22580 31208 22940 31272
rect 23004 31208 23048 31272
rect 20988 31164 22972 31208
rect 20988 29788 22836 29832
rect 20988 29724 22728 29788
rect 22792 29724 22836 29788
rect 20988 29680 22836 29724
rect 20988 29468 21352 29680
rect 22472 29576 22836 29680
rect 22472 29512 22516 29576
rect 22580 29512 22836 29576
rect 22472 29468 22836 29512
rect 16324 28136 16688 28348
rect 17172 28304 17536 28348
rect 17172 28240 17216 28304
rect 17280 28240 17536 28304
rect 17172 28136 17536 28240
rect 16324 28092 17536 28136
rect 16324 28028 17428 28092
rect 17492 28028 17536 28092
rect 16324 27984 17536 28028
rect 20988 28136 21352 28348
rect 22472 28304 23048 28348
rect 22472 28240 22940 28304
rect 23004 28240 23048 28304
rect 22472 28196 23048 28240
rect 22472 28136 22836 28196
rect 20988 28092 23048 28136
rect 20988 28028 22940 28092
rect 23004 28028 23048 28092
rect 20988 27984 23048 28028
rect 16324 26712 17536 26864
rect 16324 26652 16688 26712
rect 16324 26608 17112 26652
rect 16324 26544 17004 26608
rect 17068 26544 17112 26608
rect 16324 26500 17112 26544
rect 17172 26500 17536 26712
rect 20988 26608 22836 26652
rect 20988 26544 22516 26608
rect 22580 26544 22728 26608
rect 22792 26544 22836 26608
rect 20988 26500 22836 26544
rect 16324 25124 17536 25168
rect 16324 25060 17216 25124
rect 17280 25060 17428 25124
rect 17492 25060 17536 25124
rect 16324 25016 17536 25060
rect 20988 25124 22972 25168
rect 20988 25060 21032 25124
rect 21096 25060 22940 25124
rect 23004 25060 23048 25124
rect 20988 25016 22972 25060
rect 16324 23472 16688 23684
rect 17036 23640 17536 23684
rect 16960 23576 17004 23640
rect 17068 23576 17536 23640
rect 17036 23532 17536 23576
rect 17172 23472 17536 23532
rect 20988 23472 21352 23684
rect 22472 23640 22836 23684
rect 22472 23576 22728 23640
rect 22792 23576 22836 23640
rect 22472 23472 22836 23576
rect 16324 23428 17960 23472
rect 16324 23364 16368 23428
rect 16432 23364 17960 23428
rect 16324 23320 17960 23364
rect 17808 23260 17960 23320
rect 20988 23428 22836 23472
rect 20988 23364 21244 23428
rect 21308 23364 22836 23428
rect 20988 23320 22836 23364
rect 20988 23260 21140 23320
rect 17808 23108 21140 23260
rect 16324 22156 17536 22200
rect 16324 22092 17216 22156
rect 17280 22092 17536 22156
rect 16324 22048 17536 22092
rect 16324 21836 16688 22048
rect 17172 21944 17536 22048
rect 17172 21880 17216 21944
rect 17280 21880 17536 21944
rect 17172 21836 17536 21880
rect 20988 22156 22836 22200
rect 20988 22092 21032 22156
rect 21096 22092 22836 22156
rect 20988 22048 22836 22092
rect 20988 21944 21352 22048
rect 20988 21880 21032 21944
rect 21096 21880 21352 21944
rect 20988 21836 21352 21880
rect 22472 21836 22836 22048
rect 13992 20672 16476 20716
rect 13992 20608 16368 20672
rect 16432 20608 16476 20672
rect 13992 20564 16476 20608
rect 13992 20460 14356 20564
rect 13992 20396 14036 20460
rect 14100 20396 14356 20460
rect 13992 20352 14356 20396
rect 20988 20460 22836 20504
rect 20988 20396 21244 20460
rect 21308 20396 22516 20460
rect 22580 20396 22836 20460
rect 20988 20352 22836 20396
rect 13992 19612 14356 19868
rect 13992 19548 14248 19612
rect 14312 19548 14356 19612
rect 13992 19504 14356 19548
rect 16536 19188 17324 19232
rect 16536 19124 17216 19188
rect 17280 19124 17324 19188
rect 16536 19080 17324 19124
rect 16536 19020 16688 19080
rect 13992 18976 14356 19020
rect 13992 18912 14036 18976
rect 14100 18912 14356 18976
rect 13992 18764 14356 18912
rect 16324 18976 17536 19020
rect 16324 18912 16368 18976
rect 16432 18912 17536 18976
rect 16324 18868 17536 18912
rect 20988 18976 22836 19020
rect 20988 18912 21032 18976
rect 21096 18912 21244 18976
rect 21308 18912 22836 18976
rect 20988 18868 22836 18912
rect 13992 18700 14036 18764
rect 14100 18700 14356 18764
rect 13992 18656 14356 18700
rect 13568 18230 13932 18384
rect 13568 18174 13657 18230
rect 13713 18174 13932 18230
rect 13568 18172 13932 18174
rect 14699 18228 14831 18231
rect 15598 18228 15730 18231
rect 14699 18226 15730 18228
rect 0 18020 13932 18172
rect 14204 18128 14356 18172
rect 14699 18170 14737 18226
rect 14793 18170 15636 18226
rect 15692 18170 15730 18226
rect 14699 18168 15730 18170
rect 14699 18165 14831 18168
rect 15598 18165 15730 18168
rect 14204 18064 14248 18128
rect 14312 18064 14356 18128
rect 14204 17993 14356 18064
rect 14153 17960 14356 17993
rect 14153 17919 16476 17960
rect 14204 17916 16476 17919
rect 14204 17852 14248 17916
rect 14312 17852 16368 17916
rect 16432 17852 16476 17916
rect 14204 17808 16476 17852
rect 0 17738 13932 17748
rect 0 17682 13657 17738
rect 13713 17682 13932 17738
rect 0 17596 13932 17682
rect 14699 17744 14831 17747
rect 15514 17744 15646 17747
rect 14699 17742 15646 17744
rect 14699 17686 14737 17742
rect 14793 17686 15552 17742
rect 15608 17686 15646 17742
rect 14699 17684 15646 17686
rect 14699 17681 14831 17684
rect 15514 17681 15646 17684
rect 16324 17384 17536 17536
rect 16324 17324 16688 17384
rect 13992 17280 16688 17324
rect 13992 17216 14036 17280
rect 14100 17216 16688 17280
rect 13992 17172 16688 17216
rect 17172 17172 17536 17384
rect 20988 17324 21352 17536
rect 22472 17492 22836 17536
rect 22472 17428 22516 17492
rect 22580 17428 22836 17492
rect 22472 17324 22836 17428
rect 20988 17280 22836 17324
rect 20988 17216 21032 17280
rect 21096 17216 22836 17280
rect 20988 17172 22836 17216
rect 13992 17068 14356 17172
rect 13992 17004 14036 17068
rect 14100 17004 14356 17068
rect 13992 16960 14356 17004
rect 13568 16554 13932 16688
rect 13568 16498 13657 16554
rect 13713 16498 13932 16554
rect 13568 16476 13932 16498
rect 14699 16552 14831 16555
rect 15430 16552 15562 16555
rect 14699 16550 15562 16552
rect 14699 16494 14737 16550
rect 14793 16494 15468 16550
rect 15524 16494 15562 16550
rect 14699 16492 15562 16494
rect 14699 16489 14831 16492
rect 15430 16489 15562 16492
rect 0 16324 13932 16476
rect 14204 16432 14356 16476
rect 14204 16368 14248 16432
rect 14312 16368 14356 16432
rect 14204 16317 14356 16368
rect 14153 16264 14356 16317
rect 13568 16062 13932 16264
rect 14153 16243 14568 16264
rect 14204 16220 14568 16243
rect 14204 16156 14248 16220
rect 14312 16156 14460 16220
rect 14524 16156 14568 16220
rect 14204 16112 14568 16156
rect 13568 16052 13657 16062
rect 0 16006 13657 16052
rect 13713 16006 13932 16062
rect 0 15900 13932 16006
rect 14699 16068 14831 16071
rect 15346 16068 15478 16071
rect 14699 16066 15478 16068
rect 14699 16010 14737 16066
rect 14793 16010 15384 16066
rect 15440 16010 15478 16066
rect 14699 16008 15478 16010
rect 14699 16005 14831 16008
rect 15346 16005 15478 16008
rect 16324 15840 16688 16052
rect 17172 15840 17536 16052
rect 14492 15796 17536 15840
rect 14416 15732 14460 15796
rect 14524 15732 17536 15796
rect 14492 15688 17536 15732
rect 20988 16008 22836 16052
rect 20988 15944 21244 16008
rect 21308 15944 22836 16008
rect 20988 15900 22836 15944
rect 20988 15688 21352 15900
rect 22472 15796 22836 15900
rect 22472 15732 22516 15796
rect 22580 15732 22836 15796
rect 22472 15688 22836 15732
rect 13992 15584 14356 15628
rect 13992 15520 14036 15584
rect 14100 15520 14356 15584
rect 13992 15372 14356 15520
rect 13992 15308 14036 15372
rect 14100 15308 14356 15372
rect 13992 15264 14356 15308
rect 13568 14878 13932 14992
rect 13568 14822 13657 14878
rect 13713 14822 13932 14878
rect 13568 14780 13932 14822
rect 14699 14876 14831 14879
rect 15262 14876 15394 14879
rect 14699 14874 15394 14876
rect 14699 14818 14737 14874
rect 14793 14818 15300 14874
rect 15356 14818 15394 14874
rect 14699 14816 15394 14818
rect 14699 14813 14831 14816
rect 15262 14813 15394 14816
rect 0 14628 13932 14780
rect 14204 14736 14356 14780
rect 14204 14672 14248 14736
rect 14312 14672 14356 14736
rect 14204 14641 14356 14672
rect 13568 14386 13932 14568
rect 14153 14567 14356 14641
rect 14204 14524 14356 14567
rect 14204 14460 14248 14524
rect 14312 14460 14356 14524
rect 14204 14416 14356 14460
rect 13568 14356 13657 14386
rect 0 14330 13657 14356
rect 13713 14330 13932 14386
rect 0 14204 13932 14330
rect 14699 14392 14831 14395
rect 15178 14392 15310 14395
rect 14699 14390 15310 14392
rect 14699 14334 14737 14390
rect 14793 14334 15216 14390
rect 15272 14334 15310 14390
rect 14699 14332 15310 14334
rect 14699 14329 14831 14332
rect 15178 14329 15310 14332
rect 16324 14312 17536 14356
rect 16324 14248 16368 14312
rect 16432 14248 17536 14312
rect 16324 14204 17536 14248
rect 20988 14312 23684 14356
rect 20988 14248 21032 14312
rect 21096 14248 23576 14312
rect 23640 14248 23684 14312
rect 20988 14204 23684 14248
rect 13992 13888 16476 13932
rect 13992 13824 14036 13888
rect 14100 13824 16368 13888
rect 16432 13824 16476 13888
rect 13992 13780 16476 13824
rect 13992 13568 14356 13780
rect 13394 13269 13478 13273
rect 13328 13264 13478 13269
rect 13328 13208 13366 13264
rect 13422 13208 13478 13264
rect 13328 13203 13478 13208
rect 13394 13199 13478 13203
rect 13619 13202 13751 13211
rect 13619 13146 13657 13202
rect 13713 13146 13751 13202
rect 13619 13084 13751 13146
rect 14699 13200 14831 13203
rect 15094 13200 15226 13203
rect 14699 13198 15226 13200
rect 14699 13142 14737 13198
rect 14793 13142 15132 13198
rect 15188 13142 15226 13198
rect 14699 13140 15226 13142
rect 14699 13137 14831 13140
rect 15094 13137 15226 13140
rect 13568 13040 13932 13084
rect 13568 12976 13612 13040
rect 13676 12976 13932 13040
rect 13568 12932 13932 12976
rect 14204 13040 14356 13084
rect 14204 12976 14248 13040
rect 14312 12976 14356 13040
rect 14204 12965 14356 12976
rect 14153 12891 14356 12965
rect 14204 12872 14356 12891
rect 14204 12828 17960 12872
rect 14204 12764 17852 12828
rect 17916 12764 17960 12828
rect 14204 12720 17960 12764
rect 20988 12828 23684 12872
rect 20988 12764 21032 12828
rect 21096 12764 22516 12828
rect 22580 12764 23684 12828
rect 20988 12720 23684 12764
rect 23532 12660 23684 12720
rect 23532 12448 23896 12660
rect 26712 12448 27076 12660
rect 29892 12508 33224 12660
rect 29892 12448 30044 12508
rect 23532 12296 30044 12448
rect 32860 12296 33224 12508
rect 36040 12448 36404 12660
rect 39220 12508 45732 12660
rect 39220 12448 39372 12508
rect 36040 12296 39372 12448
rect 42188 12296 42552 12508
rect 45368 12448 45732 12508
rect 48548 12508 58028 12660
rect 48548 12448 48700 12508
rect 45368 12296 48700 12448
rect 51516 12296 51880 12508
rect 54696 12296 55060 12508
rect 57876 12404 58028 12508
rect 60844 12508 70536 12660
rect 60844 12448 61208 12508
rect 60496 12404 61208 12448
rect 57876 12340 57920 12404
rect 57984 12340 58028 12404
rect 60420 12340 60464 12404
rect 60528 12340 61208 12404
rect 57876 12296 58028 12340
rect 60496 12296 61208 12340
rect 64024 12296 64388 12508
rect 67204 12296 67356 12508
rect 70384 12296 70536 12508
rect 14894 12293 15026 12296
rect 21458 12293 21590 12296
rect 14894 12291 21590 12293
rect 14894 12235 14932 12291
rect 14988 12235 21496 12291
rect 21552 12235 21590 12291
rect 14894 12233 21590 12235
rect 14894 12230 15026 12233
rect 21458 12230 21590 12233
rect 17884 11768 21140 11812
rect 17808 11704 17852 11768
rect 17916 11704 19124 11768
rect 19188 11704 21032 11768
rect 21096 11704 21140 11768
rect 17884 11660 21140 11704
rect 23532 11768 26016 11812
rect 23532 11704 23576 11768
rect 23640 11704 25908 11768
rect 25972 11704 26016 11768
rect 23532 11660 26016 11704
rect 23532 11600 23896 11660
rect 23108 11524 23472 11600
rect 23532 11556 24032 11600
rect 26712 11556 27076 11812
rect 29892 11768 32800 11812
rect 29892 11704 32692 11768
rect 32756 11704 32800 11768
rect 29892 11660 32800 11704
rect 32860 11768 35344 11812
rect 32860 11704 35236 11768
rect 35300 11704 35344 11768
rect 32860 11660 35344 11704
rect 23532 11524 23788 11556
rect 23108 11492 23788 11524
rect 23852 11492 24000 11556
rect 24064 11524 24108 11556
rect 24064 11492 25708 11524
rect 23108 11448 25708 11492
rect 26712 11492 26968 11556
rect 27032 11492 27076 11556
rect 26712 11448 27076 11492
rect 29256 11524 29832 11600
rect 29892 11556 30044 11660
rect 32860 11600 33224 11660
rect 36040 11600 36404 11812
rect 39220 11768 41704 11812
rect 39220 11704 41596 11768
rect 41660 11704 41704 11768
rect 39220 11660 41704 11704
rect 39220 11600 39372 11660
rect 42188 11600 42552 11812
rect 44596 11768 48064 11812
rect 44520 11704 44564 11768
rect 44628 11704 47956 11768
rect 48020 11704 48064 11768
rect 44596 11660 48064 11704
rect 45368 11600 45732 11660
rect 29892 11524 29936 11556
rect 29256 11492 29936 11524
rect 30000 11524 30044 11556
rect 32436 11524 32800 11600
rect 32860 11556 33360 11600
rect 32860 11524 33328 11556
rect 30000 11492 33328 11524
rect 33392 11524 33436 11556
rect 35616 11524 35980 11600
rect 36040 11556 36540 11600
rect 36040 11524 36508 11556
rect 33392 11492 36508 11524
rect 36572 11524 36616 11556
rect 38584 11524 39160 11600
rect 36572 11492 39160 11524
rect 29256 11448 39160 11492
rect 39220 11556 39508 11600
rect 42188 11556 42688 11600
rect 45368 11556 45868 11600
rect 39220 11492 39476 11556
rect 39540 11492 39584 11556
rect 42188 11492 42444 11556
rect 42508 11492 42656 11556
rect 42720 11492 42764 11556
rect 45368 11492 45836 11556
rect 45900 11492 45944 11556
rect 39220 11448 39508 11492
rect 42188 11448 42688 11492
rect 45368 11448 45868 11492
rect 23191 11391 25708 11448
rect 29256 11391 38736 11448
rect 47912 11391 48488 11600
rect 48548 11556 48700 11812
rect 48548 11492 48592 11556
rect 48656 11492 48700 11556
rect 48548 11448 48700 11492
rect 51092 11391 51456 11600
rect 51516 11556 51880 11812
rect 51516 11492 51560 11556
rect 51624 11492 51880 11556
rect 51516 11448 51880 11492
rect 54272 11391 54636 11600
rect 54696 11556 55060 11812
rect 57528 11768 58028 11812
rect 57452 11704 57496 11768
rect 57560 11704 58028 11768
rect 57528 11660 58028 11704
rect 54696 11492 54740 11556
rect 54804 11492 55060 11556
rect 54696 11448 55060 11492
rect 57240 11391 57816 11600
rect 57876 11448 58028 11660
rect 60844 11768 63964 11812
rect 60844 11704 63856 11768
rect 63920 11704 63964 11768
rect 60844 11660 63964 11704
rect 64024 11768 66720 11812
rect 66856 11768 67356 11812
rect 64024 11704 66612 11768
rect 66676 11704 66720 11768
rect 66780 11704 66824 11768
rect 66888 11704 67356 11768
rect 64024 11660 66720 11704
rect 66856 11660 67356 11704
rect 59572 11556 60784 11600
rect 59572 11492 59616 11556
rect 59680 11492 60464 11556
rect 60528 11492 60784 11556
rect 59572 11448 60784 11492
rect 60844 11556 61208 11660
rect 60844 11492 60888 11556
rect 60952 11492 61100 11556
rect 61164 11492 61208 11556
rect 60844 11448 61208 11492
rect 60420 11391 60784 11448
rect 63600 11391 63964 11600
rect 64024 11556 64388 11660
rect 64024 11492 64068 11556
rect 64132 11492 64388 11556
rect 64024 11448 64388 11492
rect 66568 11391 67144 11600
rect 67204 11448 67356 11660
rect 69748 11391 70324 11600
rect 70384 11556 70536 11812
rect 70384 11492 70428 11556
rect 70492 11492 70536 11556
rect 70384 11448 70536 11492
rect 14894 11360 15026 11363
rect 23191 11360 70324 11391
rect 73054 11360 73186 11363
rect 14894 11358 73186 11360
rect 14894 11302 14932 11358
rect 14988 11344 73092 11358
rect 14988 11302 57920 11344
rect 14894 11300 57920 11302
rect 14894 11297 15026 11300
rect 23271 11296 23403 11300
rect 23271 11240 23309 11296
rect 23365 11240 23403 11296
rect 23271 11176 23403 11240
rect 23543 11296 23675 11300
rect 23543 11240 23581 11296
rect 23637 11240 23675 11296
rect 23543 11176 23675 11240
rect 26383 11296 26515 11300
rect 26383 11240 26421 11296
rect 26477 11240 26515 11296
rect 26383 11176 26515 11240
rect 26655 11296 26787 11300
rect 26655 11240 26693 11296
rect 26749 11240 26787 11296
rect 26655 11176 26787 11240
rect 29256 11236 29408 11300
rect 29495 11296 29627 11300
rect 29495 11240 29533 11296
rect 29589 11240 29627 11296
rect 29495 11176 29627 11240
rect 23108 11132 23472 11176
rect 23108 11068 23364 11132
rect 23428 11068 23472 11132
rect 23108 11024 23472 11068
rect 23532 11132 23684 11176
rect 23532 11068 23576 11132
rect 23640 11068 23684 11132
rect 23532 11024 23684 11068
rect 26288 11132 26652 11176
rect 26288 11068 26332 11132
rect 26396 11100 26652 11132
rect 26655 11132 26864 11176
rect 26655 11100 26756 11132
rect 26396 11068 26440 11100
rect 26288 11024 26440 11068
rect 26500 11024 26652 11100
rect 26712 11068 26756 11100
rect 26820 11068 26864 11132
rect 26712 11024 26864 11068
rect 29468 11132 29627 11176
rect 29468 11068 29512 11132
rect 29576 11100 29627 11132
rect 29767 11296 29899 11300
rect 29767 11240 29805 11296
rect 29861 11240 29899 11296
rect 29767 11176 29899 11240
rect 32607 11296 32739 11300
rect 32607 11240 32645 11296
rect 32701 11240 32739 11296
rect 32607 11176 32739 11240
rect 32879 11296 33011 11300
rect 32879 11240 32917 11296
rect 32973 11240 33011 11296
rect 32879 11176 33011 11240
rect 35719 11296 35851 11300
rect 35719 11240 35757 11296
rect 35813 11240 35851 11296
rect 35719 11176 35851 11240
rect 35991 11296 36123 11300
rect 35991 11240 36029 11296
rect 36085 11240 36123 11296
rect 35991 11176 36123 11240
rect 38584 11236 38736 11300
rect 38831 11296 38963 11300
rect 38831 11240 38869 11296
rect 38925 11240 38963 11296
rect 38831 11176 38963 11240
rect 39103 11296 39235 11300
rect 39103 11240 39141 11296
rect 39197 11240 39235 11296
rect 39103 11176 39235 11240
rect 41943 11296 42075 11300
rect 41943 11240 41981 11296
rect 42037 11240 42075 11296
rect 41943 11176 42075 11240
rect 42215 11296 42347 11300
rect 42215 11240 42253 11296
rect 42309 11240 42347 11296
rect 42215 11176 42347 11240
rect 45055 11296 45187 11300
rect 45055 11240 45093 11296
rect 45149 11240 45187 11296
rect 45055 11176 45187 11240
rect 45327 11296 45459 11300
rect 45327 11240 45365 11296
rect 45421 11240 45459 11296
rect 45327 11176 45459 11240
rect 47912 11236 48700 11300
rect 51092 11236 51668 11300
rect 54272 11236 54848 11300
rect 57240 11280 57920 11300
rect 57984 11302 73092 11344
rect 73148 11302 73186 11358
rect 57984 11300 73186 11302
rect 57984 11280 58028 11300
rect 57240 11236 58028 11280
rect 60420 11236 60996 11300
rect 63600 11236 64176 11300
rect 66568 11236 67356 11300
rect 69748 11236 70324 11300
rect 73054 11297 73186 11300
rect 29767 11132 30256 11176
rect 29767 11100 30148 11132
rect 29576 11068 29620 11100
rect 29468 11024 29620 11068
rect 29892 11068 30148 11100
rect 30212 11068 30256 11132
rect 29892 11024 30256 11068
rect 32436 11132 32800 11176
rect 32436 11068 32480 11132
rect 32544 11068 32800 11132
rect 32436 11024 32800 11068
rect 32860 11132 33224 11176
rect 32860 11068 33116 11132
rect 33180 11068 33224 11132
rect 32860 11024 33224 11068
rect 35616 11132 35980 11176
rect 35616 11068 35660 11132
rect 35724 11100 35980 11132
rect 35991 11132 36404 11176
rect 35991 11100 36296 11132
rect 35724 11068 35768 11100
rect 35616 11024 35768 11068
rect 35828 11024 35980 11100
rect 36040 11068 36296 11100
rect 36360 11068 36404 11132
rect 36040 11024 36404 11068
rect 38796 11132 39372 11176
rect 38796 11068 39052 11132
rect 39116 11100 39264 11132
rect 39116 11068 39160 11100
rect 38796 11024 39160 11068
rect 39220 11068 39264 11100
rect 39328 11068 39372 11132
rect 39220 11024 39372 11068
rect 41764 11132 42128 11176
rect 41764 11068 42020 11132
rect 42084 11068 42128 11132
rect 41764 11024 42128 11068
rect 42188 11132 42552 11176
rect 42188 11068 42232 11132
rect 42296 11068 42552 11132
rect 42188 11024 42552 11068
rect 44944 11132 45308 11176
rect 44944 11068 44988 11132
rect 45052 11100 45308 11132
rect 45327 11132 45520 11176
rect 45327 11100 45412 11132
rect 45052 11068 45096 11100
rect 44944 11024 45096 11068
rect 45156 11024 45308 11100
rect 45368 11068 45412 11100
rect 45476 11068 45520 11132
rect 45368 11024 45520 11068
rect 19080 10920 22836 10964
rect 19080 10856 19336 10920
rect 19400 10856 22728 10920
rect 22792 10856 22836 10920
rect 19080 10812 22836 10856
rect 23320 10708 23896 10752
rect 23320 10644 23788 10708
rect 23852 10644 23896 10708
rect 14894 10619 15026 10622
rect 22580 10619 22712 10622
rect 14894 10617 22712 10619
rect 14894 10561 14932 10617
rect 14988 10561 22618 10617
rect 22674 10561 22712 10617
rect 14894 10559 22712 10561
rect 14894 10556 15026 10559
rect 22580 10556 22712 10559
rect 23320 10600 23896 10644
rect 26288 10708 27076 10752
rect 26288 10644 26968 10708
rect 27032 10644 27076 10708
rect 26288 10600 27076 10644
rect 29468 10708 29832 10752
rect 35268 10708 35980 10752
rect 41628 10708 42128 10752
rect 29468 10644 29724 10708
rect 29788 10644 29832 10708
rect 35192 10644 35236 10708
rect 35300 10644 35980 10708
rect 41552 10644 41596 10708
rect 41660 10644 42128 10708
rect 29468 10600 29832 10644
rect 35268 10600 35980 10644
rect 41628 10600 42128 10644
rect 23320 10540 23472 10600
rect 26288 10540 26440 10600
rect 29468 10540 29620 10600
rect 35828 10540 35980 10600
rect 41976 10540 42128 10600
rect 23108 10496 24108 10540
rect 25940 10496 26864 10540
rect 23108 10432 24000 10496
rect 24064 10432 24108 10496
rect 25864 10432 25908 10496
rect 25972 10432 26864 10496
rect 23108 10388 24108 10432
rect 25940 10388 26864 10432
rect 23108 10328 23684 10388
rect 22760 10284 23684 10328
rect 22684 10220 22728 10284
rect 22792 10220 23684 10284
rect 22760 10176 23684 10220
rect 26288 10176 26440 10388
rect 26500 10328 26864 10388
rect 29256 10388 29832 10540
rect 29256 10328 29620 10388
rect 26500 10176 29620 10328
rect 29680 10176 29832 10388
rect 32436 10496 33436 10540
rect 32436 10432 32692 10496
rect 32756 10432 33328 10496
rect 33392 10432 33436 10496
rect 32436 10388 33436 10432
rect 35616 10496 36616 10540
rect 35616 10432 36508 10496
rect 36572 10432 36616 10496
rect 35616 10388 36616 10432
rect 32436 10176 33012 10388
rect 35616 10328 36192 10388
rect 38584 10328 38948 10540
rect 39008 10496 39584 10540
rect 39008 10432 39476 10496
rect 39540 10432 39584 10496
rect 39008 10388 39584 10432
rect 41764 10496 42764 10540
rect 41764 10432 42656 10496
rect 42720 10432 42764 10496
rect 41764 10388 42764 10432
rect 44520 10496 45944 10540
rect 44520 10432 44564 10496
rect 44628 10432 45836 10496
rect 45900 10432 45944 10496
rect 44520 10388 45944 10432
rect 47912 10496 48276 10540
rect 47912 10432 47956 10496
rect 48020 10432 48276 10496
rect 39008 10328 39160 10388
rect 35616 10176 39160 10328
rect 41764 10328 42340 10388
rect 44944 10328 45520 10388
rect 41764 10176 45520 10328
rect 47912 10328 48276 10432
rect 48336 10496 48700 10540
rect 48336 10432 48592 10496
rect 48656 10432 48700 10496
rect 48336 10328 48700 10432
rect 51092 10496 54848 10540
rect 51092 10432 51560 10496
rect 51624 10432 54528 10496
rect 54592 10432 54848 10496
rect 51092 10388 54848 10432
rect 51092 10328 51668 10388
rect 47912 10176 51668 10328
rect 54272 10328 54848 10388
rect 57240 10496 57604 10540
rect 57240 10432 57496 10496
rect 57560 10432 57604 10496
rect 57240 10328 57604 10432
rect 57664 10328 58028 10540
rect 60420 10496 61208 10540
rect 60420 10432 60676 10496
rect 60740 10432 61100 10496
rect 61164 10432 61208 10496
rect 60420 10388 61208 10432
rect 63600 10496 64176 10540
rect 63600 10432 63856 10496
rect 63920 10432 64068 10496
rect 64132 10432 64176 10496
rect 60420 10328 60996 10388
rect 54272 10176 60996 10328
rect 63600 10176 64176 10432
rect 66568 10496 67356 10540
rect 66568 10432 66612 10496
rect 66676 10432 66824 10496
rect 66888 10432 67356 10496
rect 66568 10388 67356 10432
rect 66568 10176 66932 10388
rect 66992 10328 67356 10388
rect 69748 10496 70536 10540
rect 69748 10432 70428 10496
rect 70492 10432 70536 10496
rect 69748 10388 70536 10432
rect 69748 10328 70324 10388
rect 66992 10176 70324 10328
rect 41976 10116 42128 10176
rect 19080 10072 20716 10116
rect 19080 10008 19124 10072
rect 19188 10008 20608 10072
rect 20672 10008 20716 10072
rect 19080 9964 20716 10008
rect 41976 10072 42552 10116
rect 41976 10008 42444 10072
rect 42508 10008 42552 10072
rect 41976 9964 42552 10008
rect 19080 9224 20716 9268
rect 19080 9160 19336 9224
rect 19400 9160 20716 9224
rect 19080 9116 20716 9160
rect 23532 8800 75412 8844
rect 23532 8736 59616 8800
rect 59680 8736 75304 8800
rect 75368 8736 75412 8800
rect 23532 8692 75412 8736
rect 2544 8480 2908 8632
rect 2544 8420 2846 8480
rect 848 8409 2846 8420
rect 848 8376 2696 8409
rect 848 8312 892 8376
rect 956 8312 2588 8376
rect 2652 8312 2696 8376
rect 848 8268 2696 8312
rect 19080 8376 20716 8420
rect 19080 8312 20608 8376
rect 20672 8312 20716 8376
rect 19080 8268 20716 8312
rect 2921 8228 3053 8237
rect 2921 8172 2959 8228
rect 3015 8172 3053 8228
rect 2921 8163 3053 8172
rect 6572 8022 6724 8208
rect 6443 8013 6724 8022
rect 6443 7996 6481 8013
rect 6360 7957 6481 7996
rect 6537 7957 6724 8013
rect 6360 7952 6724 7957
rect 6360 7888 6404 7952
rect 6468 7888 6724 7952
rect 6360 7844 6724 7888
rect 1908 7740 2908 7784
rect 1908 7676 1952 7740
rect 2016 7676 2908 7740
rect 1908 7632 2908 7676
rect 2544 7420 2908 7632
rect 2921 7044 3053 7053
rect 2921 6988 2959 7044
rect 3015 6988 3053 7044
rect 2921 6979 3053 6988
rect 2544 6892 2696 6936
rect 2544 6828 2588 6892
rect 2652 6828 2696 6892
rect 2544 6807 2696 6828
rect 2544 6724 2846 6807
rect 23108 6724 23260 6936
rect 23744 6724 24108 6936
rect 24592 6724 24956 6936
rect 25440 6724 25592 6936
rect 26076 6724 26440 6936
rect 26924 6784 28772 6936
rect 26924 6724 27288 6784
rect 2544 6572 2908 6724
rect 23108 6572 27288 6724
rect 27772 6572 27924 6784
rect 28408 6724 28772 6784
rect 29256 6784 30256 6936
rect 29256 6724 29620 6784
rect 28408 6572 29620 6724
rect 30104 6724 30256 6784
rect 30740 6784 34284 6936
rect 30740 6724 31104 6784
rect 30104 6572 31104 6724
rect 31588 6572 31952 6784
rect 32436 6572 32588 6784
rect 33072 6572 33436 6784
rect 33920 6724 34284 6784
rect 34768 6724 34920 6936
rect 35404 6784 36616 6936
rect 35404 6724 35768 6784
rect 33920 6572 35768 6724
rect 36252 6724 36616 6784
rect 37100 6784 38100 6936
rect 37100 6724 37252 6784
rect 36252 6572 37252 6724
rect 37736 6724 38100 6784
rect 38584 6724 38948 6936
rect 39432 6724 39584 6936
rect 40068 6784 41280 6936
rect 40068 6772 40346 6784
rect 40068 6724 40220 6772
rect 37736 6572 40220 6724
rect 40916 6724 41280 6784
rect 41764 6784 42764 6936
rect 41764 6724 41916 6784
rect 40916 6572 41916 6724
rect 42612 6724 42764 6784
rect 43248 6724 43612 6936
rect 44096 6724 44248 6936
rect 44944 6724 45096 6936
rect 45580 6784 46580 6936
rect 45580 6724 45944 6784
rect 42612 6572 45944 6724
rect 46428 6724 46580 6784
rect 47276 6724 47428 6936
rect 47912 6784 48912 6936
rect 47912 6724 48276 6784
rect 46428 6572 48276 6724
rect 48760 6724 48912 6784
rect 49608 6784 52092 6936
rect 49608 6724 49760 6784
rect 48760 6572 49760 6724
rect 50244 6572 50608 6784
rect 51092 6572 51244 6784
rect 51940 6724 52092 6784
rect 52576 6724 52940 6936
rect 53424 6724 53576 6936
rect 54272 6784 55272 6936
rect 54272 6724 54424 6784
rect 51940 6572 54424 6724
rect 54908 6724 55272 6784
rect 55756 6784 56756 6936
rect 55756 6724 55908 6784
rect 54908 6572 55908 6724
rect 56604 6724 56756 6784
rect 57240 6784 59088 6936
rect 57240 6724 57604 6784
rect 58174 6772 58452 6784
rect 56604 6572 57604 6724
rect 58300 6572 58452 6772
rect 58936 6724 59088 6784
rect 59572 6724 59936 6936
rect 60420 6724 60784 6936
rect 61268 6724 61420 6936
rect 61904 6724 62268 6936
rect 62752 6724 63116 6936
rect 63600 6784 64600 6936
rect 63600 6724 63752 6784
rect 58936 6572 63752 6724
rect 64236 6724 64600 6784
rect 65084 6784 66084 6936
rect 65084 6724 65448 6784
rect 64236 6572 65448 6724
rect 65932 6724 66084 6784
rect 66568 6784 67780 6936
rect 66568 6724 66932 6784
rect 65932 6572 66932 6724
rect 67416 6724 67780 6784
rect 68264 6784 69264 6936
rect 68264 6724 68416 6784
rect 67416 6572 68416 6724
rect 68900 6724 69264 6784
rect 69748 6724 70112 6936
rect 70596 6724 70748 6936
rect 71232 6724 71596 6936
rect 72080 6892 74352 6936
rect 72080 6828 74244 6892
rect 74308 6828 74352 6892
rect 72080 6784 74352 6828
rect 72080 6724 72444 6784
rect 68900 6572 72444 6724
rect 72928 6572 73080 6784
rect 16960 3544 17324 3756
rect 18444 3544 18808 3756
rect 16960 3500 18808 3544
rect 16960 3436 18488 3500
rect 18552 3436 18808 3500
rect 16960 3392 18808 3436
rect 19928 3604 21776 3756
rect 19928 3500 20292 3604
rect 19928 3436 19972 3500
rect 20036 3436 20292 3500
rect 19928 3392 20292 3436
rect 21412 3544 21776 3604
rect 22896 3604 24744 3756
rect 22896 3544 23260 3604
rect 21412 3392 23260 3544
rect 24380 3544 24744 3604
rect 25864 3544 26228 3756
rect 27348 3544 27712 3756
rect 28832 3604 30680 3756
rect 28832 3544 29196 3604
rect 24380 3392 29196 3544
rect 30316 3544 30680 3604
rect 31800 3544 32164 3756
rect 30316 3392 32164 3544
rect 33284 3544 33648 3756
rect 34768 3544 35132 3756
rect 36252 3604 38100 3756
rect 36252 3544 36616 3604
rect 33284 3500 36616 3544
rect 33284 3436 36508 3500
rect 36572 3436 36616 3500
rect 33284 3392 36616 3436
rect 37736 3392 38100 3604
rect 39220 3544 39584 3756
rect 40704 3544 41068 3756
rect 39220 3500 41068 3544
rect 39220 3436 40748 3500
rect 40812 3436 41068 3500
rect 39220 3392 41068 3436
rect 42188 3500 42552 3756
rect 42188 3436 42444 3500
rect 42508 3436 42552 3500
rect 42188 3392 42552 3436
rect 13328 3040 13460 3043
rect 13328 3038 31262 3040
rect 13328 2982 13366 3038
rect 13422 2982 31262 3038
rect 13328 2980 31262 2982
rect 13328 2977 13460 2980
rect 16583 2976 16715 2980
rect 16583 2920 16621 2976
rect 16677 2920 16715 2976
rect 16583 2908 16715 2920
rect 18065 2976 18197 2980
rect 18065 2920 18103 2976
rect 18159 2920 18197 2976
rect 18065 2908 18197 2920
rect 19547 2976 19679 2980
rect 19547 2920 19585 2976
rect 19641 2920 19679 2976
rect 19547 2908 19679 2920
rect 21029 2976 21161 2980
rect 21029 2920 21067 2976
rect 21123 2920 21161 2976
rect 21029 2908 21161 2920
rect 22511 2976 22643 2980
rect 22511 2920 22549 2976
rect 22605 2920 22643 2976
rect 22511 2908 22643 2920
rect 23993 2976 24125 2980
rect 23993 2920 24031 2976
rect 24087 2920 24125 2976
rect 23993 2908 24125 2920
rect 25475 2976 25607 2980
rect 25475 2920 25513 2976
rect 25569 2920 25607 2976
rect 25475 2908 25607 2920
rect 26957 2976 27089 2980
rect 26957 2920 26995 2976
rect 27051 2920 27089 2976
rect 26957 2908 27089 2920
rect 28439 2976 28571 2980
rect 28439 2920 28477 2976
rect 28533 2920 28571 2976
rect 28439 2908 28571 2920
rect 29921 2976 30053 2980
rect 29921 2920 29959 2976
rect 30015 2920 30053 2976
rect 29921 2908 30053 2920
rect 31403 2976 31535 2985
rect 31403 2920 31441 2976
rect 31497 2920 31535 2976
rect 31403 2908 31535 2920
rect 32885 2976 33017 2985
rect 32885 2920 32923 2976
rect 32979 2920 33017 2976
rect 32885 2908 33017 2920
rect 34367 2976 34499 2985
rect 34367 2920 34405 2976
rect 34461 2920 34499 2976
rect 34367 2908 34499 2920
rect 35849 2976 35981 2985
rect 35849 2920 35887 2976
rect 35943 2920 35981 2976
rect 35849 2908 35981 2920
rect 37331 2976 37463 2985
rect 37331 2920 37369 2976
rect 37425 2920 37463 2976
rect 37331 2908 37463 2920
rect 38813 2976 38945 2985
rect 38813 2920 38851 2976
rect 38907 2920 38945 2976
rect 38813 2908 38945 2920
rect 40295 2976 40427 2985
rect 40295 2920 40333 2976
rect 40389 2920 40427 2976
rect 40295 2908 40427 2920
rect 41777 2976 41909 2985
rect 41777 2920 41815 2976
rect 41871 2920 41909 2976
rect 41777 2908 41909 2920
rect 16536 2864 16900 2908
rect 16536 2800 16580 2864
rect 16644 2800 16900 2864
rect 16536 2756 16900 2800
rect 16960 2696 17324 2908
rect 18020 2864 18384 2908
rect 18020 2800 18064 2864
rect 18128 2800 18384 2864
rect 18020 2756 18384 2800
rect 18444 2696 18808 2908
rect 19504 2864 19868 2908
rect 19504 2800 19760 2864
rect 19824 2800 19868 2864
rect 19504 2756 19868 2800
rect 19928 2696 20292 2908
rect 20988 2864 21352 2908
rect 20988 2800 21032 2864
rect 21096 2800 21352 2864
rect 20988 2756 21352 2800
rect 21412 2696 21776 2908
rect 22472 2864 22836 2908
rect 22472 2800 22516 2864
rect 22580 2800 22836 2864
rect 22472 2756 22836 2800
rect 22896 2696 23260 2908
rect 23956 2864 24320 2908
rect 23956 2800 24212 2864
rect 24276 2800 24320 2864
rect 23956 2756 24320 2800
rect 24380 2696 24744 2908
rect 25440 2864 25804 2908
rect 25440 2800 25696 2864
rect 25760 2800 25804 2864
rect 25440 2756 25804 2800
rect 25864 2696 26228 2908
rect 26924 2864 27288 2908
rect 26924 2800 27180 2864
rect 27244 2800 27288 2864
rect 26924 2756 27288 2800
rect 27560 2739 27712 2908
rect 28408 2864 28772 2908
rect 28408 2800 28664 2864
rect 28728 2800 28772 2864
rect 28408 2756 28772 2800
rect 27491 2696 27712 2739
rect 28832 2696 29196 2908
rect 29892 2864 30256 2908
rect 29892 2800 29936 2864
rect 30000 2800 30256 2864
rect 29892 2756 30256 2800
rect 30528 2739 30680 2908
rect 31376 2864 31740 2908
rect 31376 2800 31420 2864
rect 31484 2800 31740 2864
rect 31376 2756 31740 2800
rect 30455 2696 30680 2739
rect 31800 2696 32164 2908
rect 32860 2864 33224 2908
rect 32860 2800 32904 2864
rect 32968 2800 33224 2864
rect 32860 2756 33224 2800
rect 33284 2696 33648 2908
rect 34344 2864 34708 2908
rect 34344 2800 34388 2864
rect 34452 2800 34708 2864
rect 34344 2756 34708 2800
rect 34768 2696 35132 2908
rect 35828 2864 36192 2908
rect 35828 2800 36084 2864
rect 36148 2800 36192 2864
rect 35828 2756 36192 2800
rect 36252 2696 36616 2908
rect 37312 2864 37464 2908
rect 37312 2800 37356 2864
rect 37420 2800 37464 2864
rect 37312 2756 37464 2800
rect 37736 2696 38100 2908
rect 38796 2864 38948 2908
rect 38796 2800 38840 2864
rect 38904 2800 38948 2864
rect 38796 2756 38948 2800
rect 39220 2696 39584 2908
rect 40280 2864 40432 2908
rect 40280 2800 40324 2864
rect 40388 2800 40432 2864
rect 40280 2756 40432 2800
rect 40704 2696 41068 2908
rect 41764 2864 41916 2908
rect 41764 2800 41808 2864
rect 41872 2800 41916 2864
rect 41764 2756 41916 2800
rect 42188 2696 42552 2908
rect 16960 2652 42552 2696
rect 16960 2588 29088 2652
rect 29152 2588 42552 2652
rect 16960 2544 42552 2588
rect 1484 2016 74776 2060
rect 1484 1952 1528 2016
rect 1592 1952 1740 2016
rect 1804 1952 1952 2016
rect 2016 1952 18488 2016
rect 18552 1952 19972 2016
rect 20036 1952 36508 2016
rect 36572 1952 40748 2016
rect 40812 1952 42444 2016
rect 42508 1952 74244 2016
rect 74308 1952 74456 2016
rect 74520 1952 74668 2016
rect 74732 1952 74776 2016
rect 1484 1804 74776 1952
rect 1484 1740 1528 1804
rect 1592 1740 1740 1804
rect 1804 1740 1952 1804
rect 2016 1740 74244 1804
rect 74308 1740 74456 1804
rect 74520 1740 74668 1804
rect 74732 1740 74776 1804
rect 1484 1592 74776 1740
rect 1484 1528 1528 1592
rect 1592 1528 1740 1592
rect 1804 1528 1952 1592
rect 2016 1528 74244 1592
rect 74308 1528 74456 1592
rect 74520 1528 74668 1592
rect 74732 1528 74776 1592
rect 1484 1484 74776 1528
rect 424 956 75836 1000
rect 424 892 468 956
rect 532 892 680 956
rect 744 892 892 956
rect 956 892 29088 956
rect 29152 892 75304 956
rect 75368 892 75516 956
rect 75580 892 75728 956
rect 75792 892 75836 956
rect 424 744 75836 892
rect 424 680 468 744
rect 532 680 680 744
rect 744 680 892 744
rect 956 680 75304 744
rect 75368 680 75516 744
rect 75580 680 75728 744
rect 75792 680 75836 744
rect 424 532 75836 680
rect 424 468 468 532
rect 532 468 680 532
rect 744 468 892 532
rect 956 468 75304 532
rect 75368 468 75516 532
rect 75580 468 75728 532
rect 75792 468 75836 532
rect 424 424 75836 468
<< via3 >>
rect 468 64280 532 64344
rect 680 64280 744 64344
rect 892 64280 956 64344
rect 75304 64280 75368 64344
rect 75516 64280 75580 64344
rect 75728 64280 75792 64344
rect 468 64068 532 64132
rect 680 64068 744 64132
rect 892 64068 956 64132
rect 75304 64068 75368 64132
rect 75516 64068 75580 64132
rect 75728 64068 75792 64132
rect 468 63856 532 63920
rect 680 63856 744 63920
rect 892 63856 956 63920
rect 21032 63856 21096 63920
rect 75304 63856 75368 63920
rect 75516 63856 75580 63920
rect 75728 63856 75792 63920
rect 1528 63220 1592 63284
rect 1740 63220 1804 63284
rect 1952 63220 2016 63284
rect 74244 63220 74308 63284
rect 74456 63220 74520 63284
rect 74668 63220 74732 63284
rect 1528 63008 1592 63072
rect 1740 63008 1804 63072
rect 1952 63008 2016 63072
rect 74244 63008 74308 63072
rect 74456 63008 74520 63072
rect 74668 63008 74732 63072
rect 1528 62796 1592 62860
rect 1740 62796 1804 62860
rect 1952 62796 2016 62860
rect 22728 62796 22792 62860
rect 74244 62796 74308 62860
rect 74456 62796 74520 62860
rect 74668 62796 74732 62860
rect 21032 61948 21096 62012
rect 22940 61948 23004 62012
rect 22728 60464 22792 60528
rect 22516 60252 22580 60316
rect 22940 58980 23004 59044
rect 21032 58768 21096 58832
rect 22516 57496 22580 57560
rect 21244 57284 21308 57348
rect 21032 55800 21096 55864
rect 21032 55588 21096 55652
rect 21244 54316 21308 54380
rect 22516 54104 22580 54168
rect 21032 52832 21096 52896
rect 21244 52620 21308 52684
rect 22516 51348 22580 51412
rect 21032 51136 21096 51200
rect 21244 49864 21308 49928
rect 21244 49652 21308 49716
rect 21032 48168 21096 48232
rect 22516 47956 22580 48020
rect 21244 46684 21308 46748
rect 21244 46472 21308 46536
rect 21032 44988 21096 45052
rect 22516 44988 22580 45052
rect 16156 43504 16220 43568
rect 21244 43504 21308 43568
rect 22728 43504 22792 43568
rect 17216 41808 17280 41872
rect 21032 42020 21096 42084
rect 22516 41808 22580 41872
rect 16156 40536 16220 40600
rect 15944 40324 16008 40388
rect 22728 40536 22792 40600
rect 22940 40324 23004 40388
rect 17216 39052 17280 39116
rect 17216 38840 17280 38904
rect 22516 38840 22580 38904
rect 22728 38840 22792 38904
rect 15944 37356 16008 37420
rect 16580 37356 16644 37420
rect 21032 37356 21096 37420
rect 22940 37356 23004 37420
rect 17216 35872 17280 35936
rect 22728 35872 22792 35936
rect 16792 35660 16856 35724
rect 22516 35660 22580 35724
rect 16580 34388 16644 34452
rect 16156 34176 16220 34240
rect 21032 34388 21096 34452
rect 22304 34176 22368 34240
rect 16792 32692 16856 32756
rect 22516 32692 22580 32756
rect 22728 32692 22792 32756
rect 16156 31208 16220 31272
rect 17216 31208 17280 31272
rect 22516 31208 22580 31272
rect 22940 31208 23004 31272
rect 22728 29724 22792 29788
rect 22516 29512 22580 29576
rect 17216 28240 17280 28304
rect 17428 28028 17492 28092
rect 22940 28240 23004 28304
rect 22940 28028 23004 28092
rect 17004 26544 17068 26608
rect 22516 26544 22580 26608
rect 22728 26544 22792 26608
rect 17216 25060 17280 25124
rect 17428 25060 17492 25124
rect 21032 25060 21096 25124
rect 22940 25060 23004 25124
rect 17004 23576 17068 23640
rect 22728 23576 22792 23640
rect 16368 23364 16432 23428
rect 21244 23364 21308 23428
rect 17216 22092 17280 22156
rect 17216 21880 17280 21944
rect 21032 22092 21096 22156
rect 21032 21880 21096 21944
rect 16368 20608 16432 20672
rect 14036 20396 14100 20460
rect 21244 20396 21308 20460
rect 22516 20396 22580 20460
rect 14248 19548 14312 19612
rect 17216 19124 17280 19188
rect 14036 18912 14100 18976
rect 16368 18912 16432 18976
rect 21032 18912 21096 18976
rect 21244 18912 21308 18976
rect 14036 18700 14100 18764
rect 14248 18064 14312 18128
rect 14248 17852 14312 17916
rect 16368 17852 16432 17916
rect 14036 17216 14100 17280
rect 22516 17428 22580 17492
rect 21032 17216 21096 17280
rect 14036 17004 14100 17068
rect 14248 16368 14312 16432
rect 14248 16156 14312 16220
rect 14460 16156 14524 16220
rect 14460 15732 14524 15796
rect 21244 15944 21308 16008
rect 22516 15732 22580 15796
rect 14036 15520 14100 15584
rect 14036 15308 14100 15372
rect 14248 14672 14312 14736
rect 14248 14460 14312 14524
rect 16368 14248 16432 14312
rect 21032 14248 21096 14312
rect 23576 14248 23640 14312
rect 14036 13824 14100 13888
rect 16368 13824 16432 13888
rect 13612 12976 13676 13040
rect 14248 12976 14312 13040
rect 17852 12764 17916 12828
rect 21032 12764 21096 12828
rect 22516 12764 22580 12828
rect 57920 12340 57984 12404
rect 60464 12340 60528 12404
rect 17852 11704 17916 11768
rect 19124 11704 19188 11768
rect 21032 11704 21096 11768
rect 23576 11704 23640 11768
rect 25908 11704 25972 11768
rect 32692 11704 32756 11768
rect 35236 11704 35300 11768
rect 23788 11492 23852 11556
rect 24000 11492 24064 11556
rect 26968 11492 27032 11556
rect 41596 11704 41660 11768
rect 44564 11704 44628 11768
rect 47956 11704 48020 11768
rect 29936 11492 30000 11556
rect 33328 11492 33392 11556
rect 36508 11492 36572 11556
rect 39476 11492 39540 11556
rect 42444 11492 42508 11556
rect 42656 11492 42720 11556
rect 45836 11492 45900 11556
rect 48592 11492 48656 11556
rect 51560 11492 51624 11556
rect 57496 11704 57560 11768
rect 54740 11492 54804 11556
rect 63856 11704 63920 11768
rect 66612 11704 66676 11768
rect 66824 11704 66888 11768
rect 59616 11492 59680 11556
rect 60464 11492 60528 11556
rect 60888 11492 60952 11556
rect 61100 11492 61164 11556
rect 64068 11492 64132 11556
rect 70428 11492 70492 11556
rect 23364 11068 23428 11132
rect 23576 11068 23640 11132
rect 26332 11068 26396 11132
rect 26756 11068 26820 11132
rect 29512 11068 29576 11132
rect 57920 11280 57984 11344
rect 30148 11068 30212 11132
rect 32480 11068 32544 11132
rect 33116 11068 33180 11132
rect 35660 11068 35724 11132
rect 36296 11068 36360 11132
rect 39052 11068 39116 11132
rect 39264 11068 39328 11132
rect 42020 11068 42084 11132
rect 42232 11068 42296 11132
rect 44988 11068 45052 11132
rect 45412 11068 45476 11132
rect 19336 10856 19400 10920
rect 22728 10856 22792 10920
rect 23788 10644 23852 10708
rect 26968 10644 27032 10708
rect 29724 10644 29788 10708
rect 35236 10644 35300 10708
rect 41596 10644 41660 10708
rect 24000 10432 24064 10496
rect 25908 10432 25972 10496
rect 22728 10220 22792 10284
rect 32692 10432 32756 10496
rect 33328 10432 33392 10496
rect 36508 10432 36572 10496
rect 39476 10432 39540 10496
rect 42656 10432 42720 10496
rect 44564 10432 44628 10496
rect 45836 10432 45900 10496
rect 47956 10432 48020 10496
rect 48592 10432 48656 10496
rect 51560 10432 51624 10496
rect 54528 10432 54592 10496
rect 57496 10432 57560 10496
rect 60676 10432 60740 10496
rect 61100 10432 61164 10496
rect 63856 10432 63920 10496
rect 64068 10432 64132 10496
rect 66612 10432 66676 10496
rect 66824 10432 66888 10496
rect 70428 10432 70492 10496
rect 19124 10008 19188 10072
rect 20608 10008 20672 10072
rect 42444 10008 42508 10072
rect 19336 9160 19400 9224
rect 59616 8736 59680 8800
rect 75304 8736 75368 8800
rect 892 8312 956 8376
rect 2588 8312 2652 8376
rect 20608 8312 20672 8376
rect 6404 7888 6468 7952
rect 1952 7676 2016 7740
rect 2588 6828 2652 6892
rect 74244 6828 74308 6892
rect 18488 3436 18552 3500
rect 19972 3436 20036 3500
rect 36508 3436 36572 3500
rect 40748 3436 40812 3500
rect 42444 3436 42508 3500
rect 16580 2800 16644 2864
rect 18064 2800 18128 2864
rect 19760 2800 19824 2864
rect 21032 2800 21096 2864
rect 22516 2800 22580 2864
rect 24212 2800 24276 2864
rect 25696 2800 25760 2864
rect 27180 2800 27244 2864
rect 28664 2800 28728 2864
rect 29936 2800 30000 2864
rect 31420 2800 31484 2864
rect 32904 2800 32968 2864
rect 34388 2800 34452 2864
rect 36084 2800 36148 2864
rect 37356 2800 37420 2864
rect 38840 2800 38904 2864
rect 40324 2800 40388 2864
rect 41808 2800 41872 2864
rect 29088 2588 29152 2652
rect 1528 1952 1592 2016
rect 1740 1952 1804 2016
rect 1952 1952 2016 2016
rect 18488 1952 18552 2016
rect 19972 1952 20036 2016
rect 36508 1952 36572 2016
rect 40748 1952 40812 2016
rect 42444 1952 42508 2016
rect 74244 1952 74308 2016
rect 74456 1952 74520 2016
rect 74668 1952 74732 2016
rect 1528 1740 1592 1804
rect 1740 1740 1804 1804
rect 1952 1740 2016 1804
rect 74244 1740 74308 1804
rect 74456 1740 74520 1804
rect 74668 1740 74732 1804
rect 1528 1528 1592 1592
rect 1740 1528 1804 1592
rect 1952 1528 2016 1592
rect 74244 1528 74308 1592
rect 74456 1528 74520 1592
rect 74668 1528 74732 1592
rect 468 892 532 956
rect 680 892 744 956
rect 892 892 956 956
rect 29088 892 29152 956
rect 75304 892 75368 956
rect 75516 892 75580 956
rect 75728 892 75792 956
rect 468 680 532 744
rect 680 680 744 744
rect 892 680 956 744
rect 75304 680 75368 744
rect 75516 680 75580 744
rect 75728 680 75792 744
rect 468 468 532 532
rect 680 468 744 532
rect 892 468 956 532
rect 75304 468 75368 532
rect 75516 468 75580 532
rect 75728 468 75792 532
<< metal4 >>
rect 424 64344 1000 64388
rect 424 64280 468 64344
rect 532 64280 680 64344
rect 744 64280 892 64344
rect 956 64280 1000 64344
rect 424 64132 1000 64280
rect 424 64068 468 64132
rect 532 64068 680 64132
rect 744 64068 892 64132
rect 956 64068 1000 64132
rect 424 63920 1000 64068
rect 75260 64344 75836 64388
rect 75260 64280 75304 64344
rect 75368 64280 75516 64344
rect 75580 64280 75728 64344
rect 75792 64280 75836 64344
rect 75260 64132 75836 64280
rect 75260 64068 75304 64132
rect 75368 64068 75516 64132
rect 75580 64068 75728 64132
rect 75792 64068 75836 64132
rect 424 63856 468 63920
rect 532 63856 680 63920
rect 744 63856 892 63920
rect 956 63856 1000 63920
rect 424 8376 1000 63856
rect 20988 63920 21140 63964
rect 20988 63856 21032 63920
rect 21096 63856 21140 63920
rect 424 8312 892 8376
rect 956 8312 1000 8376
rect 424 956 1000 8312
rect 1484 63284 2060 63328
rect 1484 63220 1528 63284
rect 1592 63220 1740 63284
rect 1804 63220 1952 63284
rect 2016 63220 2060 63284
rect 1484 63072 2060 63220
rect 1484 63008 1528 63072
rect 1592 63008 1740 63072
rect 1804 63008 1952 63072
rect 2016 63008 2060 63072
rect 1484 62860 2060 63008
rect 1484 62796 1528 62860
rect 1592 62796 1740 62860
rect 1804 62796 1952 62860
rect 2016 62796 2060 62860
rect 1484 7740 2060 62796
rect 20988 62012 21140 63856
rect 75260 63920 75836 64068
rect 75260 63856 75304 63920
rect 75368 63856 75516 63920
rect 75580 63856 75728 63920
rect 75792 63856 75836 63920
rect 74200 63284 74776 63328
rect 74200 63220 74244 63284
rect 74308 63220 74456 63284
rect 74520 63220 74668 63284
rect 74732 63220 74776 63284
rect 74200 63072 74776 63220
rect 74200 63008 74244 63072
rect 74308 63008 74456 63072
rect 74520 63008 74668 63072
rect 74732 63008 74776 63072
rect 20988 61980 21032 62012
rect 21018 61948 21032 61980
rect 21096 61980 21140 62012
rect 22684 62860 22836 62904
rect 22684 62796 22728 62860
rect 22792 62796 22836 62860
rect 21096 61948 21110 61980
rect 21018 61934 21110 61948
rect 22684 60528 22836 62796
rect 74200 62860 74776 63008
rect 74200 62796 74244 62860
rect 74308 62796 74456 62860
rect 74520 62796 74668 62860
rect 74732 62796 74776 62860
rect 22684 60496 22728 60528
rect 22714 60464 22728 60496
rect 22792 60496 22836 60528
rect 22896 62012 23048 62056
rect 22896 61948 22940 62012
rect 23004 61948 23048 62012
rect 22792 60464 22806 60496
rect 22714 60450 22806 60464
rect 22502 60316 22594 60330
rect 22502 60284 22516 60316
rect 22472 60252 22516 60284
rect 22580 60284 22594 60316
rect 22580 60252 22624 60284
rect 20988 58832 21140 58876
rect 20988 58768 21032 58832
rect 21096 58768 21140 58832
rect 20988 55864 21140 58768
rect 22472 57560 22624 60252
rect 22896 59044 23048 61948
rect 22896 59012 22940 59044
rect 22926 58980 22940 59012
rect 23004 59012 23048 59044
rect 23004 58980 23018 59012
rect 22926 58966 23018 58980
rect 22472 57496 22516 57560
rect 22580 57496 22624 57560
rect 22472 57452 22624 57496
rect 20988 55832 21032 55864
rect 21018 55800 21032 55832
rect 21096 55832 21140 55864
rect 21200 57348 21352 57392
rect 21200 57284 21244 57348
rect 21308 57284 21352 57348
rect 21096 55800 21110 55832
rect 21018 55786 21110 55800
rect 21018 55652 21110 55666
rect 21018 55620 21032 55652
rect 20988 55588 21032 55620
rect 21096 55620 21110 55652
rect 21096 55588 21140 55620
rect 20988 52896 21140 55588
rect 21200 54380 21352 57284
rect 21200 54348 21244 54380
rect 21230 54316 21244 54348
rect 21308 54348 21352 54380
rect 21308 54316 21322 54348
rect 21230 54302 21322 54316
rect 22502 54168 22594 54182
rect 22502 54136 22516 54168
rect 20988 52832 21032 52896
rect 21096 52832 21140 52896
rect 20988 52788 21140 52832
rect 22472 54104 22516 54136
rect 22580 54136 22594 54168
rect 22580 54104 22624 54136
rect 21200 52684 21352 52728
rect 21200 52620 21244 52684
rect 21308 52620 21352 52684
rect 21018 51200 21110 51214
rect 21018 51168 21032 51200
rect 20988 51136 21032 51168
rect 21096 51168 21110 51200
rect 21096 51136 21140 51168
rect 20988 48232 21140 51136
rect 21200 49928 21352 52620
rect 22472 51412 22624 54104
rect 22472 51348 22516 51412
rect 22580 51348 22624 51412
rect 22472 51304 22624 51348
rect 21200 49896 21244 49928
rect 21230 49864 21244 49896
rect 21308 49896 21352 49928
rect 21308 49864 21322 49896
rect 21230 49850 21322 49864
rect 21230 49716 21322 49730
rect 21230 49684 21244 49716
rect 20988 48168 21032 48232
rect 21096 48168 21140 48232
rect 20988 48124 21140 48168
rect 21200 49652 21244 49684
rect 21308 49684 21322 49716
rect 21308 49652 21352 49684
rect 21200 46748 21352 49652
rect 22502 48020 22594 48034
rect 22502 47988 22516 48020
rect 21200 46684 21244 46748
rect 21308 46684 21352 46748
rect 21200 46640 21352 46684
rect 22472 47956 22516 47988
rect 22580 47988 22594 48020
rect 22580 47956 22624 47988
rect 21230 46536 21322 46550
rect 21230 46504 21244 46536
rect 21200 46472 21244 46504
rect 21308 46504 21322 46536
rect 21308 46472 21352 46504
rect 21018 45052 21110 45066
rect 21018 45020 21032 45052
rect 20988 44988 21032 45020
rect 21096 45020 21110 45052
rect 21096 44988 21140 45020
rect 16142 43568 16234 43582
rect 16142 43536 16156 43568
rect 16112 43504 16156 43536
rect 16220 43536 16234 43568
rect 16220 43504 16264 43536
rect 16112 40600 16264 43504
rect 20988 42084 21140 44988
rect 21200 43568 21352 46472
rect 22472 45052 22624 47956
rect 22472 44988 22516 45052
rect 22580 44988 22624 45052
rect 22472 44944 22624 44988
rect 21200 43504 21244 43568
rect 21308 43504 21352 43568
rect 21200 43460 21352 43504
rect 22684 43568 22836 43612
rect 22684 43504 22728 43568
rect 22792 43504 22836 43568
rect 20988 42020 21032 42084
rect 21096 42020 21140 42084
rect 20988 41976 21140 42020
rect 17202 41872 17294 41886
rect 17202 41840 17216 41872
rect 16112 40536 16156 40600
rect 16220 40536 16264 40600
rect 16112 40492 16264 40536
rect 17172 41808 17216 41840
rect 17280 41840 17294 41872
rect 22472 41872 22624 41916
rect 17280 41808 17324 41840
rect 15900 40388 16052 40432
rect 15900 40324 15944 40388
rect 16008 40324 16052 40388
rect 15900 37420 16052 40324
rect 17172 39116 17324 41808
rect 17172 39052 17216 39116
rect 17280 39052 17324 39116
rect 17172 39008 17324 39052
rect 22472 41808 22516 41872
rect 22580 41808 22624 41872
rect 17202 38904 17294 38918
rect 17202 38872 17216 38904
rect 17172 38840 17216 38872
rect 17280 38872 17294 38904
rect 22472 38904 22624 41808
rect 22684 40600 22836 43504
rect 22684 40568 22728 40600
rect 22714 40536 22728 40568
rect 22792 40568 22836 40600
rect 22792 40536 22806 40568
rect 22714 40522 22806 40536
rect 22896 40388 23048 40432
rect 22896 40324 22940 40388
rect 23004 40324 23048 40388
rect 22472 38872 22516 38904
rect 17280 38840 17324 38872
rect 15900 37388 15944 37420
rect 15930 37356 15944 37388
rect 16008 37388 16052 37420
rect 16566 37420 16658 37434
rect 16566 37388 16580 37420
rect 16008 37356 16022 37388
rect 15930 37342 16022 37356
rect 16536 37356 16580 37388
rect 16644 37388 16658 37420
rect 16644 37356 16688 37388
rect 16536 34452 16688 37356
rect 17172 35936 17324 38840
rect 22502 38840 22516 38872
rect 22580 38872 22624 38904
rect 22714 38904 22806 38918
rect 22714 38872 22728 38904
rect 22580 38840 22594 38872
rect 22502 38826 22594 38840
rect 22684 38840 22728 38872
rect 22792 38872 22806 38904
rect 22792 38840 22836 38872
rect 17172 35872 17216 35936
rect 17280 35872 17324 35936
rect 17172 35828 17324 35872
rect 20988 37420 21140 37464
rect 20988 37356 21032 37420
rect 21096 37356 21140 37420
rect 16536 34388 16580 34452
rect 16644 34388 16688 34452
rect 16536 34344 16688 34388
rect 16748 35724 16900 35768
rect 16748 35660 16792 35724
rect 16856 35660 16900 35724
rect 16142 34240 16234 34254
rect 16142 34208 16156 34240
rect 16112 34176 16156 34208
rect 16220 34208 16234 34240
rect 16220 34176 16264 34208
rect 16112 31272 16264 34176
rect 16748 32756 16900 35660
rect 20988 34452 21140 37356
rect 22684 35936 22836 38840
rect 22896 37420 23048 40324
rect 22896 37388 22940 37420
rect 22926 37356 22940 37388
rect 23004 37388 23048 37420
rect 23004 37356 23018 37388
rect 22926 37342 23018 37356
rect 22684 35872 22728 35936
rect 22792 35872 22836 35936
rect 22684 35828 22836 35872
rect 20988 34420 21032 34452
rect 21018 34388 21032 34420
rect 21096 34420 21140 34452
rect 22472 35724 22624 35768
rect 22472 35660 22516 35724
rect 22580 35660 22624 35724
rect 21096 34388 21110 34420
rect 21018 34374 21110 34388
rect 16748 32724 16792 32756
rect 16778 32692 16792 32724
rect 16856 32724 16900 32756
rect 22260 34240 22412 34284
rect 22260 34176 22304 34240
rect 22368 34176 22412 34240
rect 16856 32692 16870 32724
rect 16778 32678 16870 32692
rect 22260 32588 22412 34176
rect 22472 32756 22624 35660
rect 22472 32724 22516 32756
rect 22502 32692 22516 32724
rect 22580 32724 22624 32756
rect 22714 32756 22806 32770
rect 22714 32724 22728 32756
rect 22580 32692 22594 32724
rect 22502 32678 22594 32692
rect 22684 32692 22728 32724
rect 22792 32724 22806 32756
rect 22792 32692 22836 32724
rect 22260 32436 22624 32588
rect 16112 31208 16156 31272
rect 16220 31208 16264 31272
rect 17202 31272 17294 31286
rect 17202 31240 17216 31272
rect 16112 31164 16264 31208
rect 17172 31208 17216 31240
rect 17280 31240 17294 31272
rect 22472 31272 22624 32436
rect 22472 31240 22516 31272
rect 17280 31208 17324 31240
rect 17172 28304 17324 31208
rect 22502 31208 22516 31240
rect 22580 31240 22624 31272
rect 22580 31208 22594 31240
rect 22502 31194 22594 31208
rect 22684 29788 22836 32692
rect 22684 29724 22728 29788
rect 22792 29724 22836 29788
rect 22684 29680 22836 29724
rect 22896 31272 23048 31316
rect 22896 31208 22940 31272
rect 23004 31208 23048 31272
rect 17172 28240 17216 28304
rect 17280 28240 17324 28304
rect 17172 28196 17324 28240
rect 22472 29576 22624 29620
rect 22472 29512 22516 29576
rect 22580 29512 22624 29576
rect 17414 28092 17506 28106
rect 17414 28060 17428 28092
rect 17384 28028 17428 28060
rect 17492 28060 17506 28092
rect 17492 28028 17536 28060
rect 16990 26608 17082 26622
rect 16990 26576 17004 26608
rect 16960 26544 17004 26576
rect 17068 26576 17082 26608
rect 17068 26544 17112 26576
rect 16960 23640 17112 26544
rect 16960 23576 17004 23640
rect 17068 23576 17112 23640
rect 16960 23532 17112 23576
rect 17172 25124 17324 25168
rect 17172 25060 17216 25124
rect 17280 25060 17324 25124
rect 16324 23428 16476 23472
rect 16324 23364 16368 23428
rect 16432 23364 16476 23428
rect 16324 20672 16476 23364
rect 17172 22156 17324 25060
rect 17384 25124 17536 28028
rect 22472 26608 22624 29512
rect 22896 28304 23048 31208
rect 22896 28272 22940 28304
rect 22926 28240 22940 28272
rect 23004 28272 23048 28304
rect 23004 28240 23018 28272
rect 22926 28226 23018 28240
rect 22926 28092 23018 28106
rect 22926 28060 22940 28092
rect 22896 28028 22940 28060
rect 23004 28060 23018 28092
rect 23004 28028 23048 28060
rect 22472 26576 22516 26608
rect 22502 26544 22516 26576
rect 22580 26576 22624 26608
rect 22714 26608 22806 26622
rect 22714 26576 22728 26608
rect 22580 26544 22594 26576
rect 22502 26530 22594 26544
rect 22684 26544 22728 26576
rect 22792 26576 22806 26608
rect 22792 26544 22836 26576
rect 17384 25060 17428 25124
rect 17492 25060 17536 25124
rect 21018 25124 21110 25138
rect 21018 25092 21032 25124
rect 17384 25016 17536 25060
rect 20988 25060 21032 25092
rect 21096 25092 21110 25124
rect 21096 25060 21140 25092
rect 17172 22124 17216 22156
rect 17202 22092 17216 22124
rect 17280 22124 17324 22156
rect 20988 22156 21140 25060
rect 22684 23640 22836 26544
rect 22896 25124 23048 28028
rect 22896 25060 22940 25124
rect 23004 25060 23048 25124
rect 22896 25016 23048 25060
rect 22684 23576 22728 23640
rect 22792 23576 22836 23640
rect 22684 23532 22836 23576
rect 21230 23428 21322 23442
rect 21230 23396 21244 23428
rect 17280 22092 17294 22124
rect 17202 22078 17294 22092
rect 20988 22092 21032 22156
rect 21096 22092 21140 22156
rect 20988 22048 21140 22092
rect 21200 23364 21244 23396
rect 21308 23396 21322 23428
rect 21308 23364 21352 23396
rect 16324 20640 16368 20672
rect 16354 20608 16368 20640
rect 16432 20640 16476 20672
rect 17172 21944 17324 21988
rect 17172 21880 17216 21944
rect 17280 21880 17324 21944
rect 16432 20608 16446 20640
rect 16354 20594 16446 20608
rect 13992 20460 14144 20504
rect 13992 20396 14036 20460
rect 14100 20396 14144 20460
rect 13992 18976 14144 20396
rect 14234 19612 14326 19626
rect 14234 19580 14248 19612
rect 13992 18944 14036 18976
rect 14022 18912 14036 18944
rect 14100 18944 14144 18976
rect 14204 19548 14248 19580
rect 14312 19580 14326 19612
rect 14312 19548 14356 19580
rect 14100 18912 14114 18944
rect 14022 18898 14114 18912
rect 14022 18764 14114 18778
rect 14022 18732 14036 18764
rect 13992 18700 14036 18732
rect 14100 18732 14114 18764
rect 14100 18700 14144 18732
rect 13992 17280 14144 18700
rect 14204 18128 14356 19548
rect 17172 19188 17324 21880
rect 17172 19156 17216 19188
rect 17202 19124 17216 19156
rect 17280 19156 17324 19188
rect 20988 21944 21140 21988
rect 20988 21880 21032 21944
rect 21096 21880 21140 21944
rect 17280 19124 17294 19156
rect 17202 19110 17294 19124
rect 14204 18064 14248 18128
rect 14312 18064 14356 18128
rect 14204 18020 14356 18064
rect 16324 18976 16476 19020
rect 16324 18912 16368 18976
rect 16432 18912 16476 18976
rect 20988 18976 21140 21880
rect 21200 20460 21352 23364
rect 21200 20396 21244 20460
rect 21308 20396 21352 20460
rect 22502 20460 22594 20474
rect 22502 20428 22516 20460
rect 21200 20352 21352 20396
rect 22472 20396 22516 20428
rect 22580 20428 22594 20460
rect 22580 20396 22624 20428
rect 20988 18944 21032 18976
rect 13992 17216 14036 17280
rect 14100 17216 14144 17280
rect 13992 17172 14144 17216
rect 14204 17916 14356 17960
rect 14204 17852 14248 17916
rect 14312 17852 14356 17916
rect 16324 17916 16476 18912
rect 21018 18912 21032 18944
rect 21096 18944 21140 18976
rect 21200 18976 21352 19020
rect 21096 18912 21110 18944
rect 21018 18898 21110 18912
rect 21200 18912 21244 18976
rect 21308 18912 21352 18976
rect 16324 17884 16368 17916
rect 13992 17068 14144 17112
rect 13992 17004 14036 17068
rect 14100 17004 14144 17068
rect 13992 15584 14144 17004
rect 14204 16432 14356 17852
rect 16354 17852 16368 17884
rect 16432 17884 16476 17916
rect 16432 17852 16446 17884
rect 16354 17838 16446 17852
rect 21018 17280 21110 17294
rect 21018 17248 21032 17280
rect 14204 16400 14248 16432
rect 14234 16368 14248 16400
rect 14312 16400 14356 16432
rect 20988 17216 21032 17248
rect 21096 17248 21110 17280
rect 21096 17216 21140 17248
rect 14312 16368 14326 16400
rect 14234 16354 14326 16368
rect 14234 16220 14326 16234
rect 14234 16188 14248 16220
rect 13992 15552 14036 15584
rect 14022 15520 14036 15552
rect 14100 15552 14144 15584
rect 14204 16156 14248 16188
rect 14312 16188 14326 16220
rect 14446 16220 14538 16234
rect 14446 16188 14460 16220
rect 14312 16156 14356 16188
rect 14100 15520 14114 15552
rect 14022 15506 14114 15520
rect 14022 15372 14114 15386
rect 14022 15340 14036 15372
rect 13992 15308 14036 15340
rect 14100 15340 14114 15372
rect 14100 15308 14144 15340
rect 13992 13888 14144 15308
rect 14204 14736 14356 16156
rect 14416 16156 14460 16188
rect 14524 16188 14538 16220
rect 14524 16156 14568 16188
rect 14416 15796 14568 16156
rect 14416 15732 14460 15796
rect 14524 15732 14568 15796
rect 14416 15688 14568 15732
rect 14204 14672 14248 14736
rect 14312 14672 14356 14736
rect 14204 14628 14356 14672
rect 14234 14524 14326 14538
rect 14234 14492 14248 14524
rect 13992 13824 14036 13888
rect 14100 13824 14144 13888
rect 13992 13780 14144 13824
rect 14204 14460 14248 14492
rect 14312 14492 14326 14524
rect 14312 14460 14356 14492
rect 13598 13040 13690 13054
rect 13598 13008 13612 13040
rect 13568 12976 13612 13008
rect 13676 13008 13690 13040
rect 14204 13040 14356 14460
rect 16324 14312 16476 14356
rect 16324 14248 16368 14312
rect 16432 14248 16476 14312
rect 16324 13888 16476 14248
rect 20988 14312 21140 17216
rect 21200 16008 21352 18912
rect 22472 17492 22624 20396
rect 22472 17428 22516 17492
rect 22580 17428 22624 17492
rect 22472 17384 22624 17428
rect 21200 15976 21244 16008
rect 21230 15944 21244 15976
rect 21308 15976 21352 16008
rect 21308 15944 21322 15976
rect 21230 15930 21322 15944
rect 22502 15796 22594 15810
rect 22502 15764 22516 15796
rect 20988 14248 21032 14312
rect 21096 14248 21140 14312
rect 20988 14204 21140 14248
rect 22472 15732 22516 15764
rect 22580 15764 22594 15796
rect 22580 15732 22624 15764
rect 16324 13856 16368 13888
rect 16354 13824 16368 13856
rect 16432 13856 16476 13888
rect 16432 13824 16446 13856
rect 16354 13810 16446 13824
rect 13676 12976 13720 13008
rect 1484 7676 1952 7740
rect 2016 7676 2060 7740
rect 1484 2016 2060 7676
rect 2544 8376 2696 8420
rect 2544 8312 2588 8376
rect 2652 8312 2696 8376
rect 2544 6892 2696 8312
rect 6390 7952 6482 7966
rect 6390 7920 6404 7952
rect 2544 6860 2588 6892
rect 2574 6828 2588 6860
rect 2652 6860 2696 6892
rect 6360 7888 6404 7920
rect 6468 7920 6482 7952
rect 6468 7888 6512 7920
rect 2652 6828 2666 6860
rect 2574 6814 2666 6828
rect 1484 1952 1528 2016
rect 1592 1952 1740 2016
rect 1804 1952 1952 2016
rect 2016 1952 2060 2016
rect 1484 1804 2060 1952
rect 1484 1740 1528 1804
rect 1592 1740 1740 1804
rect 1804 1740 1952 1804
rect 2016 1740 2060 1804
rect 1484 1592 2060 1740
rect 1484 1528 1528 1592
rect 1592 1528 1740 1592
rect 1804 1528 1952 1592
rect 2016 1528 2060 1592
rect 1484 1484 2060 1528
rect 424 892 468 956
rect 532 892 680 956
rect 744 892 892 956
rect 956 892 1000 956
rect 424 744 1000 892
rect 424 680 468 744
rect 532 680 680 744
rect 744 680 892 744
rect 956 680 1000 744
rect 424 532 1000 680
rect 424 468 468 532
rect 532 468 680 532
rect 744 468 892 532
rect 956 468 1000 532
rect 424 424 1000 468
rect 6360 0 6512 7888
rect 13568 0 13720 12976
rect 14204 12976 14248 13040
rect 14312 12976 14356 13040
rect 14204 12932 14356 12976
rect 17838 12828 17930 12842
rect 17838 12796 17852 12828
rect 17808 12764 17852 12796
rect 17916 12796 17930 12828
rect 20988 12828 21140 12872
rect 17916 12764 17960 12796
rect 17808 11768 17960 12764
rect 20988 12764 21032 12828
rect 21096 12764 21140 12828
rect 17808 11704 17852 11768
rect 17916 11704 17960 11768
rect 17808 11660 17960 11704
rect 19080 11768 19232 11812
rect 19080 11704 19124 11768
rect 19188 11704 19232 11768
rect 20988 11768 21140 12764
rect 22472 12828 22624 15732
rect 23562 14312 23654 14326
rect 23562 14280 23576 14312
rect 22472 12764 22516 12828
rect 22580 12764 22624 12828
rect 22472 12720 22624 12764
rect 23532 14248 23576 14280
rect 23640 14280 23654 14312
rect 23640 14248 23684 14280
rect 20988 11736 21032 11768
rect 19080 10072 19232 11704
rect 21018 11704 21032 11736
rect 21096 11736 21140 11768
rect 23532 11768 23684 14248
rect 57876 12404 58028 12448
rect 57876 12340 57920 12404
rect 57984 12340 58028 12404
rect 21096 11704 21110 11736
rect 21018 11690 21110 11704
rect 23532 11704 23576 11768
rect 23640 11704 23684 11768
rect 25894 11768 25986 11782
rect 25894 11736 25908 11768
rect 23532 11660 23684 11704
rect 25864 11704 25908 11736
rect 25972 11736 25986 11768
rect 32678 11768 32770 11782
rect 32678 11736 32692 11768
rect 25972 11704 26016 11736
rect 23744 11556 23896 11600
rect 23744 11492 23788 11556
rect 23852 11492 23896 11556
rect 23350 11132 23442 11146
rect 23350 11100 23364 11132
rect 23320 11068 23364 11100
rect 23428 11100 23442 11132
rect 23562 11132 23654 11146
rect 23562 11100 23576 11132
rect 23428 11068 23472 11100
rect 19322 10920 19414 10934
rect 19322 10888 19336 10920
rect 19080 10040 19124 10072
rect 19110 10008 19124 10040
rect 19188 10040 19232 10072
rect 19292 10856 19336 10888
rect 19400 10888 19414 10920
rect 22714 10920 22806 10934
rect 22714 10888 22728 10920
rect 19400 10856 19444 10888
rect 19188 10008 19202 10040
rect 19110 9994 19202 10008
rect 19292 9224 19444 10856
rect 22684 10856 22728 10888
rect 22792 10888 22806 10920
rect 22792 10856 22836 10888
rect 22684 10284 22836 10856
rect 22684 10220 22728 10284
rect 22792 10220 22836 10284
rect 22684 10176 22836 10220
rect 20594 10072 20686 10086
rect 20594 10040 20608 10072
rect 19292 9160 19336 9224
rect 19400 9160 19444 9224
rect 19292 9116 19444 9160
rect 20564 10008 20608 10040
rect 20672 10040 20686 10072
rect 20672 10008 20716 10040
rect 20564 8376 20716 10008
rect 20564 8312 20608 8376
rect 20672 8312 20716 8376
rect 20564 8268 20716 8312
rect 18474 3500 18566 3514
rect 18474 3468 18488 3500
rect 18444 3436 18488 3468
rect 18552 3468 18566 3500
rect 19958 3500 20050 3514
rect 19958 3468 19972 3500
rect 18552 3436 18596 3468
rect 16566 2864 16658 2878
rect 16566 2832 16580 2864
rect 16536 2800 16580 2832
rect 16644 2832 16658 2864
rect 18050 2864 18142 2878
rect 18050 2832 18064 2864
rect 16644 2800 16688 2832
rect 16536 0 16688 2800
rect 18020 2800 18064 2832
rect 18128 2832 18142 2864
rect 18128 2800 18172 2832
rect 18020 0 18172 2800
rect 18444 2016 18596 3436
rect 19928 3436 19972 3468
rect 20036 3468 20050 3500
rect 20036 3436 20080 3468
rect 19746 2864 19838 2878
rect 19746 2832 19760 2864
rect 18444 1952 18488 2016
rect 18552 1952 18596 2016
rect 18444 1908 18596 1952
rect 19716 2800 19760 2832
rect 19824 2832 19838 2864
rect 19824 2800 19868 2832
rect 19716 0 19868 2800
rect 19928 2016 20080 3436
rect 21018 2864 21110 2878
rect 21018 2832 21032 2864
rect 19928 1952 19972 2016
rect 20036 1952 20080 2016
rect 19928 1908 20080 1952
rect 20988 2800 21032 2832
rect 21096 2832 21110 2864
rect 22502 2864 22594 2878
rect 22502 2832 22516 2864
rect 21096 2800 21140 2832
rect 20988 0 21140 2800
rect 22472 2800 22516 2832
rect 22580 2832 22594 2864
rect 22580 2800 22624 2832
rect 22472 0 22624 2800
rect 23320 0 23472 11068
rect 23532 11068 23576 11100
rect 23640 11100 23654 11132
rect 23640 11068 23684 11100
rect 23532 0 23684 11068
rect 23744 10708 23896 11492
rect 23744 10676 23788 10708
rect 23774 10644 23788 10676
rect 23852 10676 23896 10708
rect 23956 11556 24108 11600
rect 23956 11492 24000 11556
rect 24064 11492 24108 11556
rect 23852 10644 23866 10676
rect 23774 10630 23866 10644
rect 23956 10496 24108 11492
rect 23956 10464 24000 10496
rect 23986 10432 24000 10464
rect 24064 10464 24108 10496
rect 25864 10496 26016 11704
rect 32648 11704 32692 11736
rect 32756 11736 32770 11768
rect 35222 11768 35314 11782
rect 35222 11736 35236 11768
rect 32756 11704 32800 11736
rect 26924 11556 27076 11600
rect 26924 11492 26968 11556
rect 27032 11492 27076 11556
rect 26318 11132 26410 11146
rect 26318 11100 26332 11132
rect 24064 10432 24078 10464
rect 23986 10418 24078 10432
rect 25864 10432 25908 10496
rect 25972 10432 26016 10496
rect 25864 10388 26016 10432
rect 26288 11068 26332 11100
rect 26396 11100 26410 11132
rect 26742 11132 26834 11146
rect 26742 11100 26756 11132
rect 26396 11068 26440 11100
rect 24198 2864 24290 2878
rect 24198 2832 24212 2864
rect 24168 2800 24212 2832
rect 24276 2832 24290 2864
rect 25682 2864 25774 2878
rect 25682 2832 25696 2864
rect 24276 2800 24320 2832
rect 24168 0 24320 2800
rect 25652 2800 25696 2832
rect 25760 2832 25774 2864
rect 25760 2800 25804 2832
rect 25652 0 25804 2800
rect 26288 0 26440 11068
rect 26712 11068 26756 11100
rect 26820 11100 26834 11132
rect 26820 11068 26864 11100
rect 26712 0 26864 11068
rect 26924 10708 27076 11492
rect 29680 11556 30044 11600
rect 29680 11492 29936 11556
rect 30000 11492 30044 11556
rect 29680 11448 30044 11492
rect 29498 11132 29590 11146
rect 29498 11100 29512 11132
rect 26924 10676 26968 10708
rect 26954 10644 26968 10676
rect 27032 10676 27076 10708
rect 29468 11068 29512 11100
rect 29576 11100 29590 11132
rect 29576 11068 29620 11100
rect 27032 10644 27046 10676
rect 26954 10630 27046 10644
rect 27166 2864 27258 2878
rect 27166 2832 27180 2864
rect 27136 2800 27180 2832
rect 27244 2832 27258 2864
rect 28650 2864 28742 2878
rect 28650 2832 28664 2864
rect 27244 2800 27288 2832
rect 27136 0 27288 2800
rect 28620 2800 28664 2832
rect 28728 2832 28742 2864
rect 28728 2800 28772 2832
rect 28620 0 28772 2800
rect 29074 2652 29166 2666
rect 29074 2620 29088 2652
rect 29044 2588 29088 2620
rect 29152 2620 29166 2652
rect 29152 2588 29196 2620
rect 29044 956 29196 2588
rect 29044 892 29088 956
rect 29152 892 29196 956
rect 29044 848 29196 892
rect 29468 0 29620 11068
rect 29680 10708 29832 11448
rect 30134 11132 30226 11146
rect 30134 11100 30148 11132
rect 29680 10676 29724 10708
rect 29710 10644 29724 10676
rect 29788 10676 29832 10708
rect 30104 11068 30148 11100
rect 30212 11100 30226 11132
rect 32466 11132 32558 11146
rect 32466 11100 32480 11132
rect 30212 11068 30256 11100
rect 29788 10644 29802 10676
rect 29710 10630 29802 10644
rect 29922 2864 30014 2878
rect 29922 2832 29936 2864
rect 29892 2800 29936 2832
rect 30000 2832 30014 2864
rect 30000 2800 30044 2832
rect 29892 0 30044 2800
rect 30104 0 30256 11068
rect 32436 11068 32480 11100
rect 32544 11100 32558 11132
rect 32544 11068 32588 11100
rect 31406 2864 31498 2878
rect 31406 2832 31420 2864
rect 31376 2800 31420 2832
rect 31484 2832 31498 2864
rect 31484 2800 31528 2832
rect 31376 0 31528 2800
rect 32436 0 32588 11068
rect 32648 10496 32800 11704
rect 35192 11704 35236 11736
rect 35300 11736 35314 11768
rect 41582 11768 41674 11782
rect 41582 11736 41596 11768
rect 35300 11704 35344 11736
rect 33284 11556 33436 11600
rect 33284 11492 33328 11556
rect 33392 11492 33436 11556
rect 33102 11132 33194 11146
rect 33102 11100 33116 11132
rect 32648 10432 32692 10496
rect 32756 10432 32800 10496
rect 32648 10388 32800 10432
rect 33072 11068 33116 11100
rect 33180 11100 33194 11132
rect 33180 11068 33224 11100
rect 32890 2864 32982 2878
rect 32890 2832 32904 2864
rect 32860 2800 32904 2832
rect 32968 2832 32982 2864
rect 32968 2800 33012 2832
rect 32860 0 33012 2800
rect 33072 0 33224 11068
rect 33284 10496 33436 11492
rect 35192 10708 35344 11704
rect 41552 11704 41596 11736
rect 41660 11736 41674 11768
rect 44520 11768 44672 11812
rect 41660 11704 41704 11736
rect 36464 11556 36616 11600
rect 36464 11492 36508 11556
rect 36572 11492 36616 11556
rect 35646 11132 35738 11146
rect 35646 11100 35660 11132
rect 35192 10644 35236 10708
rect 35300 10644 35344 10708
rect 35192 10600 35344 10644
rect 35616 11068 35660 11100
rect 35724 11100 35738 11132
rect 36282 11132 36374 11146
rect 36282 11100 36296 11132
rect 35724 11068 35768 11100
rect 33284 10464 33328 10496
rect 33314 10432 33328 10464
rect 33392 10464 33436 10496
rect 33392 10432 33406 10464
rect 33314 10418 33406 10432
rect 34374 2864 34466 2878
rect 34374 2832 34388 2864
rect 34344 2800 34388 2832
rect 34452 2832 34466 2864
rect 34452 2800 34496 2832
rect 34344 0 34496 2800
rect 35616 0 35768 11068
rect 36252 11068 36296 11100
rect 36360 11100 36374 11132
rect 36360 11068 36404 11100
rect 36070 2864 36162 2878
rect 36070 2832 36084 2864
rect 36040 2800 36084 2832
rect 36148 2832 36162 2864
rect 36148 2800 36192 2832
rect 36040 0 36192 2800
rect 36252 0 36404 11068
rect 36464 10496 36616 11492
rect 39432 11556 39584 11600
rect 39432 11492 39476 11556
rect 39540 11492 39584 11556
rect 39038 11132 39130 11146
rect 39038 11100 39052 11132
rect 36464 10464 36508 10496
rect 36494 10432 36508 10464
rect 36572 10464 36616 10496
rect 39008 11068 39052 11100
rect 39116 11100 39130 11132
rect 39250 11132 39342 11146
rect 39250 11100 39264 11132
rect 39116 11068 39160 11100
rect 36572 10432 36586 10464
rect 36494 10418 36586 10432
rect 36494 3500 36586 3514
rect 36494 3468 36508 3500
rect 36464 3436 36508 3468
rect 36572 3468 36586 3500
rect 36572 3436 36616 3468
rect 36464 2016 36616 3436
rect 37342 2864 37434 2878
rect 37342 2832 37356 2864
rect 36464 1952 36508 2016
rect 36572 1952 36616 2016
rect 36464 1908 36616 1952
rect 37312 2800 37356 2832
rect 37420 2832 37434 2864
rect 38826 2864 38918 2878
rect 38826 2832 38840 2864
rect 37420 2800 37464 2832
rect 37312 0 37464 2800
rect 38796 2800 38840 2832
rect 38904 2832 38918 2864
rect 38904 2800 38948 2832
rect 38796 0 38948 2800
rect 39008 0 39160 11068
rect 39220 11068 39264 11100
rect 39328 11100 39342 11132
rect 39328 11068 39372 11100
rect 39220 0 39372 11068
rect 39432 10496 39584 11492
rect 41552 10708 41704 11704
rect 44520 11704 44564 11768
rect 44628 11704 44672 11768
rect 47942 11768 48034 11782
rect 47942 11736 47956 11768
rect 42400 11556 42552 11600
rect 42400 11492 42444 11556
rect 42508 11492 42552 11556
rect 42006 11132 42098 11146
rect 42006 11100 42020 11132
rect 41552 10644 41596 10708
rect 41660 10644 41704 10708
rect 41552 10600 41704 10644
rect 41976 11068 42020 11100
rect 42084 11100 42098 11132
rect 42218 11132 42310 11146
rect 42218 11100 42232 11132
rect 42084 11068 42128 11100
rect 39432 10464 39476 10496
rect 39462 10432 39476 10464
rect 39540 10464 39584 10496
rect 39540 10432 39554 10464
rect 39462 10418 39554 10432
rect 40734 3500 40826 3514
rect 40734 3468 40748 3500
rect 40704 3436 40748 3468
rect 40812 3468 40826 3500
rect 40812 3436 40856 3468
rect 40310 2864 40402 2878
rect 40310 2832 40324 2864
rect 40280 2800 40324 2832
rect 40388 2832 40402 2864
rect 40388 2800 40432 2832
rect 40280 0 40432 2800
rect 40704 2016 40856 3436
rect 41794 2864 41886 2878
rect 41794 2832 41808 2864
rect 40704 1952 40748 2016
rect 40812 1952 40856 2016
rect 40704 1908 40856 1952
rect 41764 2800 41808 2832
rect 41872 2832 41886 2864
rect 41872 2800 41916 2832
rect 41764 0 41916 2800
rect 41976 0 42128 11068
rect 42188 11068 42232 11100
rect 42296 11100 42310 11132
rect 42296 11068 42340 11100
rect 42188 0 42340 11068
rect 42400 10072 42552 11492
rect 42612 11556 42764 11600
rect 42612 11492 42656 11556
rect 42720 11492 42764 11556
rect 42612 10496 42764 11492
rect 42612 10464 42656 10496
rect 42642 10432 42656 10464
rect 42720 10464 42764 10496
rect 44520 10496 44672 11704
rect 47912 11704 47956 11736
rect 48020 11736 48034 11768
rect 57452 11768 57604 11812
rect 48020 11704 48064 11736
rect 45792 11556 45944 11600
rect 45792 11492 45836 11556
rect 45900 11492 45944 11556
rect 44974 11132 45066 11146
rect 44974 11100 44988 11132
rect 44520 10464 44564 10496
rect 42720 10432 42734 10464
rect 42642 10418 42734 10432
rect 44550 10432 44564 10464
rect 44628 10464 44672 10496
rect 44944 11068 44988 11100
rect 45052 11100 45066 11132
rect 45398 11132 45490 11146
rect 45398 11100 45412 11132
rect 45052 11068 45096 11100
rect 44628 10432 44642 10464
rect 44550 10418 44642 10432
rect 42400 10040 42444 10072
rect 42430 10008 42444 10040
rect 42508 10040 42552 10072
rect 42508 10008 42522 10040
rect 42430 9994 42522 10008
rect 42430 3500 42522 3514
rect 42430 3468 42444 3500
rect 42400 3436 42444 3468
rect 42508 3468 42522 3500
rect 42508 3436 42552 3468
rect 42400 2016 42552 3436
rect 42400 1952 42444 2016
rect 42508 1952 42552 2016
rect 42400 1908 42552 1952
rect 44944 0 45096 11068
rect 45368 11068 45412 11100
rect 45476 11100 45490 11132
rect 45476 11068 45520 11100
rect 45368 0 45520 11068
rect 45792 10496 45944 11492
rect 45792 10464 45836 10496
rect 45822 10432 45836 10464
rect 45900 10464 45944 10496
rect 47912 10496 48064 11704
rect 57452 11704 57496 11768
rect 57560 11704 57604 11768
rect 45900 10432 45914 10464
rect 45822 10418 45914 10432
rect 47912 10432 47956 10496
rect 48020 10432 48064 10496
rect 48548 11556 48700 11600
rect 48548 11492 48592 11556
rect 48656 11492 48700 11556
rect 48548 10496 48700 11492
rect 48548 10464 48592 10496
rect 47912 10388 48064 10432
rect 48578 10432 48592 10464
rect 48656 10464 48700 10496
rect 51516 11556 51668 11600
rect 51516 11492 51560 11556
rect 51624 11492 51668 11556
rect 51516 10496 51668 11492
rect 51516 10464 51560 10496
rect 48656 10432 48670 10464
rect 48578 10418 48670 10432
rect 51546 10432 51560 10464
rect 51624 10464 51668 10496
rect 54484 11556 54848 11600
rect 54484 11492 54740 11556
rect 54804 11492 54848 11556
rect 54484 11448 54848 11492
rect 54484 10496 54636 11448
rect 54484 10464 54528 10496
rect 51624 10432 51638 10464
rect 51546 10418 51638 10432
rect 54514 10432 54528 10464
rect 54592 10464 54636 10496
rect 57452 10496 57604 11704
rect 57876 11344 58028 12340
rect 60420 12404 60572 12448
rect 60420 12340 60464 12404
rect 60528 12340 60572 12404
rect 59602 11556 59694 11570
rect 59602 11524 59616 11556
rect 57876 11312 57920 11344
rect 57906 11280 57920 11312
rect 57984 11312 58028 11344
rect 59572 11492 59616 11524
rect 59680 11524 59694 11556
rect 60420 11556 60572 12340
rect 63842 11768 63934 11782
rect 63842 11736 63856 11768
rect 63812 11704 63856 11736
rect 63920 11736 63934 11768
rect 66598 11768 66690 11782
rect 66598 11736 66612 11768
rect 63920 11704 63964 11736
rect 60420 11524 60464 11556
rect 59680 11492 59724 11524
rect 57984 11280 57998 11312
rect 57906 11266 57998 11280
rect 57452 10464 57496 10496
rect 54592 10432 54606 10464
rect 54514 10418 54606 10432
rect 57482 10432 57496 10464
rect 57560 10464 57604 10496
rect 57560 10432 57574 10464
rect 57482 10418 57574 10432
rect 59572 8800 59724 11492
rect 60450 11492 60464 11524
rect 60528 11524 60572 11556
rect 60632 11556 60996 11600
rect 60528 11492 60542 11524
rect 60450 11478 60542 11492
rect 60632 11492 60888 11556
rect 60952 11492 60996 11556
rect 60632 11448 60996 11492
rect 61056 11556 61208 11600
rect 61056 11492 61100 11556
rect 61164 11492 61208 11556
rect 60632 10496 60784 11448
rect 60632 10464 60676 10496
rect 60662 10432 60676 10464
rect 60740 10464 60784 10496
rect 61056 10496 61208 11492
rect 61056 10464 61100 10496
rect 60740 10432 60754 10464
rect 60662 10418 60754 10432
rect 61086 10432 61100 10464
rect 61164 10464 61208 10496
rect 63812 10496 63964 11704
rect 66568 11704 66612 11736
rect 66676 11736 66690 11768
rect 66780 11768 66932 11812
rect 66676 11704 66720 11736
rect 61164 10432 61178 10464
rect 61086 10418 61178 10432
rect 63812 10432 63856 10496
rect 63920 10432 63964 10496
rect 64024 11556 64176 11600
rect 64024 11492 64068 11556
rect 64132 11492 64176 11556
rect 64024 10496 64176 11492
rect 64024 10464 64068 10496
rect 63812 10388 63964 10432
rect 64054 10432 64068 10464
rect 64132 10464 64176 10496
rect 66568 10496 66720 11704
rect 64132 10432 64146 10464
rect 64054 10418 64146 10432
rect 66568 10432 66612 10496
rect 66676 10432 66720 10496
rect 66780 11704 66824 11768
rect 66888 11704 66932 11768
rect 66780 10496 66932 11704
rect 66780 10464 66824 10496
rect 66568 10388 66720 10432
rect 66810 10432 66824 10464
rect 66888 10464 66932 10496
rect 70384 11556 70536 11600
rect 70384 11492 70428 11556
rect 70492 11492 70536 11556
rect 70384 10496 70536 11492
rect 70384 10464 70428 10496
rect 66888 10432 66902 10464
rect 66810 10418 66902 10432
rect 70414 10432 70428 10464
rect 70492 10464 70536 10496
rect 70492 10432 70506 10464
rect 70414 10418 70506 10432
rect 59572 8736 59616 8800
rect 59680 8736 59724 8800
rect 59572 8692 59724 8736
rect 74200 6892 74776 62796
rect 74200 6828 74244 6892
rect 74308 6828 74776 6892
rect 74200 2016 74776 6828
rect 74200 1952 74244 2016
rect 74308 1952 74456 2016
rect 74520 1952 74668 2016
rect 74732 1952 74776 2016
rect 74200 1804 74776 1952
rect 74200 1740 74244 1804
rect 74308 1740 74456 1804
rect 74520 1740 74668 1804
rect 74732 1740 74776 1804
rect 74200 1592 74776 1740
rect 74200 1528 74244 1592
rect 74308 1528 74456 1592
rect 74520 1528 74668 1592
rect 74732 1528 74776 1592
rect 74200 1484 74776 1528
rect 75260 8800 75836 63856
rect 75260 8736 75304 8800
rect 75368 8736 75836 8800
rect 75260 956 75836 8736
rect 75260 892 75304 956
rect 75368 892 75516 956
rect 75580 892 75728 956
rect 75792 892 75836 956
rect 75260 744 75836 892
rect 75260 680 75304 744
rect 75368 680 75516 744
rect 75580 680 75728 744
rect 75792 680 75836 744
rect 75260 532 75836 680
rect 75260 468 75304 532
rect 75368 468 75516 532
rect 75580 468 75728 532
rect 75792 468 75836 532
rect 75260 424 75836 468
use contact_31  contact_31_0
timestamp 1644951705
transform 1 0 75260 0 1 8722
box 0 0 1 1
use contact_31  contact_31_1
timestamp 1644951705
transform 1 0 29044 0 1 878
box 0 0 1 1
use contact_31  contact_31_2
timestamp 1644951705
transform 1 0 29044 0 1 2574
box 0 0 1 1
use contact_31  contact_31_3
timestamp 1644951705
transform 1 0 22260 0 1 34162
box 0 0 1 1
use contact_31  contact_31_4
timestamp 1644951705
transform 1 0 22472 0 1 31194
box 0 0 1 1
use contact_31  contact_31_5
timestamp 1644951705
transform 1 0 22472 0 1 12750
box 0 0 1 1
use contact_31  contact_31_6
timestamp 1644951705
transform 1 0 22472 0 1 15718
box 0 0 1 1
use contact_31  contact_31_7
timestamp 1644951705
transform 1 0 22684 0 1 43490
box 0 0 1 1
use contact_31  contact_31_8
timestamp 1644951705
transform 1 0 22684 0 1 40522
box 0 0 1 1
use contact_31  contact_31_9
timestamp 1644951705
transform 1 0 22896 0 1 61934
box 0 0 1 1
use contact_31  contact_31_10
timestamp 1644951705
transform 1 0 22896 0 1 58966
box 0 0 1 1
use contact_31  contact_31_11
timestamp 1644951705
transform 1 0 22896 0 1 31194
box 0 0 1 1
use contact_31  contact_31_12
timestamp 1644951705
transform 1 0 22896 0 1 28226
box 0 0 1 1
use contact_31  contact_31_13
timestamp 1644951705
transform 1 0 22896 0 1 25046
box 0 0 1 1
use contact_31  contact_31_14
timestamp 1644951705
transform 1 0 22896 0 1 28014
box 0 0 1 1
use contact_31  contact_31_15
timestamp 1644951705
transform 1 0 22896 0 1 40310
box 0 0 1 1
use contact_31  contact_31_16
timestamp 1644951705
transform 1 0 22896 0 1 37342
box 0 0 1 1
use contact_31  contact_31_17
timestamp 1644951705
transform 1 0 20988 0 1 63842
box 0 0 1 1
use contact_31  contact_31_18
timestamp 1644951705
transform 1 0 20988 0 1 61934
box 0 0 1 1
use contact_31  contact_31_19
timestamp 1644951705
transform 1 0 21200 0 1 43490
box 0 0 1 1
use contact_31  contact_31_20
timestamp 1644951705
transform 1 0 21200 0 1 46458
box 0 0 1 1
use contact_31  contact_31_21
timestamp 1644951705
transform 1 0 21200 0 1 52606
box 0 0 1 1
use contact_31  contact_31_22
timestamp 1644951705
transform 1 0 21200 0 1 49850
box 0 0 1 1
use contact_31  contact_31_23
timestamp 1644951705
transform 1 0 21200 0 1 46670
box 0 0 1 1
use contact_31  contact_31_24
timestamp 1644951705
transform 1 0 21200 0 1 49638
box 0 0 1 1
use contact_31  contact_31_25
timestamp 1644951705
transform 1 0 20988 0 1 21866
box 0 0 1 1
use contact_31  contact_31_26
timestamp 1644951705
transform 1 0 20988 0 1 18898
box 0 0 1 1
use contact_31  contact_31_27
timestamp 1644951705
transform 1 0 21200 0 1 18898
box 0 0 1 1
use contact_31  contact_31_28
timestamp 1644951705
transform 1 0 21200 0 1 15930
box 0 0 1 1
use contact_31  contact_31_29
timestamp 1644951705
transform 1 0 20988 0 1 22078
box 0 0 1 1
use contact_31  contact_31_30
timestamp 1644951705
transform 1 0 20988 0 1 25046
box 0 0 1 1
use contact_31  contact_31_31
timestamp 1644951705
transform 1 0 20988 0 1 37342
box 0 0 1 1
use contact_31  contact_31_32
timestamp 1644951705
transform 1 0 20988 0 1 34374
box 0 0 1 1
use contact_31  contact_31_33
timestamp 1644951705
transform 1 0 20988 0 1 52818
box 0 0 1 1
use contact_31  contact_31_34
timestamp 1644951705
transform 1 0 20988 0 1 55574
box 0 0 1 1
use contact_31  contact_31_35
timestamp 1644951705
transform 1 0 20988 0 1 58754
box 0 0 1 1
use contact_31  contact_31_36
timestamp 1644951705
transform 1 0 20988 0 1 55786
box 0 0 1 1
use contact_31  contact_31_37
timestamp 1644951705
transform 1 0 20564 0 1 8298
box 0 0 1 1
use contact_31  contact_31_38
timestamp 1644951705
transform 1 0 20564 0 1 9994
box 0 0 1 1
use contact_31  contact_31_39
timestamp 1644951705
transform 1 0 20988 0 1 12750
box 0 0 1 1
use contact_31  contact_31_40
timestamp 1644951705
transform 1 0 20988 0 1 11690
box 0 0 1 1
use contact_31  contact_31_41
timestamp 1644951705
transform 1 0 19080 0 1 11690
box 0 0 1 1
use contact_31  contact_31_42
timestamp 1644951705
transform 1 0 19080 0 1 9994
box 0 0 1 1
use contact_31  contact_31_43
timestamp 1644951705
transform 1 0 17172 0 1 25046
box 0 0 1 1
use contact_31  contact_31_44
timestamp 1644951705
transform 1 0 17172 0 1 22078
box 0 0 1 1
use contact_31  contact_31_45
timestamp 1644951705
transform 1 0 17384 0 1 25046
box 0 0 1 1
use contact_31  contact_31_46
timestamp 1644951705
transform 1 0 17384 0 1 28014
box 0 0 1 1
use contact_31  contact_31_47
timestamp 1644951705
transform 1 0 17808 0 1 11690
box 0 0 1 1
use contact_31  contact_31_48
timestamp 1644951705
transform 1 0 17808 0 1 12750
box 0 0 1 1
use contact_31  contact_31_49
timestamp 1644951705
transform 1 0 17172 0 1 28226
box 0 0 1 1
use contact_31  contact_31_50
timestamp 1644951705
transform 1 0 17172 0 1 31194
box 0 0 1 1
use contact_31  contact_31_51
timestamp 1644951705
transform 1 0 17172 0 1 21866
box 0 0 1 1
use contact_31  contact_31_52
timestamp 1644951705
transform 1 0 17172 0 1 19110
box 0 0 1 1
use contact_31  contact_31_53
timestamp 1644951705
transform 1 0 16112 0 1 40522
box 0 0 1 1
use contact_31  contact_31_54
timestamp 1644951705
transform 1 0 16112 0 1 43490
box 0 0 1 1
use contact_31  contact_31_55
timestamp 1644951705
transform 1 0 16536 0 1 34374
box 0 0 1 1
use contact_31  contact_31_56
timestamp 1644951705
transform 1 0 16536 0 1 37342
box 0 0 1 1
use contact_31  contact_31_57
timestamp 1644951705
transform 1 0 15900 0 1 40310
box 0 0 1 1
use contact_31  contact_31_58
timestamp 1644951705
transform 1 0 15900 0 1 37342
box 0 0 1 1
use contact_31  contact_31_59
timestamp 1644951705
transform 1 0 16112 0 1 31194
box 0 0 1 1
use contact_31  contact_31_60
timestamp 1644951705
transform 1 0 16112 0 1 34162
box 0 0 1 1
use contact_31  contact_31_61
timestamp 1644951705
transform 1 0 60420 0 1 12326
box 0 0 1 1
use contact_31  contact_31_62
timestamp 1644951705
transform 1 0 60420 0 1 11478
box 0 0 1 1
use contact_31  contact_31_63
timestamp 1644951705
transform 1 0 59572 0 1 8722
box 0 0 1 1
use contact_31  contact_31_64
timestamp 1644951705
transform 1 0 59572 0 1 11478
box 0 0 1 1
use contact_31  contact_31_65
timestamp 1644951705
transform 1 0 57876 0 1 12326
box 0 0 1 1
use contact_31  contact_31_66
timestamp 1644951705
transform 1 0 57876 0 1 11266
box 0 0 1 1
use contact_31  contact_31_67
timestamp 1644951705
transform 1 0 16324 0 1 18898
box 0 0 1 1
use contact_31  contact_31_68
timestamp 1644951705
transform 1 0 16324 0 1 17838
box 0 0 1 1
use contact_31  contact_31_69
timestamp 1644951705
transform 1 0 14204 0 1 12962
box 0 0 1 1
use contact_31  contact_31_70
timestamp 1644951705
transform 1 0 14204 0 1 14446
box 0 0 1 1
use contact_31  contact_31_71
timestamp 1644951705
transform 1 0 14204 0 1 18050
box 0 0 1 1
use contact_31  contact_31_72
timestamp 1644951705
transform 1 0 14204 0 1 19534
box 0 0 1 1
use contact_31  contact_31_73
timestamp 1644951705
transform 1 0 14416 0 1 15718
box 0 0 1 1
use contact_31  contact_31_74
timestamp 1644951705
transform 1 0 14416 0 1 16142
box 0 0 1 1
use contact_31  contact_31_75
timestamp 1644951705
transform 1 0 14204 0 1 17838
box 0 0 1 1
use contact_31  contact_31_76
timestamp 1644951705
transform 1 0 14204 0 1 16354
box 0 0 1 1
use contact_31  contact_31_77
timestamp 1644951705
transform 1 0 14204 0 1 14658
box 0 0 1 1
use contact_31  contact_31_78
timestamp 1644951705
transform 1 0 14204 0 1 16142
box 0 0 1 1
use contact_31  contact_31_79
timestamp 1644951705
transform 1 0 848 0 1 8298
box 0 0 1 1
use contact_31  contact_31_80
timestamp 1644951705
transform 1 0 2544 0 1 8298
box 0 0 1 1
use contact_31  contact_31_81
timestamp 1644951705
transform 1 0 2544 0 1 6814
box 0 0 1 1
use contact_31  contact_31_82
timestamp 1644951705
transform 1 0 74200 0 1 6814
box 0 0 1 1
use contact_31  contact_31_83
timestamp 1644951705
transform 1 0 70384 0 1 11478
box 0 0 1 1
use contact_31  contact_31_84
timestamp 1644951705
transform 1 0 70384 0 1 10418
box 0 0 1 1
use contact_31  contact_31_85
timestamp 1644951705
transform 1 0 66780 0 1 11690
box 0 0 1 1
use contact_31  contact_31_86
timestamp 1644951705
transform 1 0 66780 0 1 10418
box 0 0 1 1
use contact_31  contact_31_87
timestamp 1644951705
transform 1 0 66568 0 1 10418
box 0 0 1 1
use contact_31  contact_31_88
timestamp 1644951705
transform 1 0 66568 0 1 11690
box 0 0 1 1
use contact_31  contact_31_89
timestamp 1644951705
transform 1 0 64024 0 1 11478
box 0 0 1 1
use contact_31  contact_31_90
timestamp 1644951705
transform 1 0 64024 0 1 10418
box 0 0 1 1
use contact_31  contact_31_91
timestamp 1644951705
transform 1 0 63812 0 1 10418
box 0 0 1 1
use contact_31  contact_31_92
timestamp 1644951705
transform 1 0 63812 0 1 11690
box 0 0 1 1
use contact_31  contact_31_93
timestamp 1644951705
transform 1 0 61056 0 1 11478
box 0 0 1 1
use contact_31  contact_31_94
timestamp 1644951705
transform 1 0 61056 0 1 10418
box 0 0 1 1
use contact_31  contact_31_95
timestamp 1644951705
transform 1 0 60844 0 1 11478
box 0 0 1 1
use contact_31  contact_31_96
timestamp 1644951705
transform 1 0 60632 0 1 10418
box 0 0 1 1
use contact_31  contact_31_97
timestamp 1644951705
transform 1 0 57452 0 1 11690
box 0 0 1 1
use contact_31  contact_31_98
timestamp 1644951705
transform 1 0 57452 0 1 10418
box 0 0 1 1
use contact_31  contact_31_99
timestamp 1644951705
transform 1 0 54696 0 1 11478
box 0 0 1 1
use contact_31  contact_31_100
timestamp 1644951705
transform 1 0 54484 0 1 10418
box 0 0 1 1
use contact_31  contact_31_101
timestamp 1644951705
transform 1 0 51516 0 1 11478
box 0 0 1 1
use contact_31  contact_31_102
timestamp 1644951705
transform 1 0 51516 0 1 10418
box 0 0 1 1
use contact_31  contact_31_103
timestamp 1644951705
transform 1 0 48548 0 1 11478
box 0 0 1 1
use contact_31  contact_31_104
timestamp 1644951705
transform 1 0 48548 0 1 10418
box 0 0 1 1
use contact_31  contact_31_105
timestamp 1644951705
transform 1 0 47912 0 1 10418
box 0 0 1 1
use contact_31  contact_31_106
timestamp 1644951705
transform 1 0 47912 0 1 11690
box 0 0 1 1
use contact_31  contact_31_107
timestamp 1644951705
transform 1 0 45792 0 1 11478
box 0 0 1 1
use contact_31  contact_31_108
timestamp 1644951705
transform 1 0 45792 0 1 10418
box 0 0 1 1
use contact_31  contact_31_109
timestamp 1644951705
transform 1 0 44520 0 1 11690
box 0 0 1 1
use contact_31  contact_31_110
timestamp 1644951705
transform 1 0 44520 0 1 10418
box 0 0 1 1
use contact_31  contact_31_111
timestamp 1644951705
transform 1 0 42400 0 1 1938
box 0 0 1 1
use contact_31  contact_31_112
timestamp 1644951705
transform 1 0 42400 0 1 3422
box 0 0 1 1
use contact_31  contact_31_113
timestamp 1644951705
transform 1 0 42612 0 1 11478
box 0 0 1 1
use contact_31  contact_31_114
timestamp 1644951705
transform 1 0 42612 0 1 10418
box 0 0 1 1
use contact_31  contact_31_115
timestamp 1644951705
transform 1 0 42400 0 1 11478
box 0 0 1 1
use contact_31  contact_31_116
timestamp 1644951705
transform 1 0 42400 0 1 9994
box 0 0 1 1
use contact_31  contact_31_117
timestamp 1644951705
transform 1 0 40704 0 1 1938
box 0 0 1 1
use contact_31  contact_31_118
timestamp 1644951705
transform 1 0 40704 0 1 3422
box 0 0 1 1
use contact_31  contact_31_119
timestamp 1644951705
transform 1 0 41552 0 1 10630
box 0 0 1 1
use contact_31  contact_31_120
timestamp 1644951705
transform 1 0 41552 0 1 11690
box 0 0 1 1
use contact_31  contact_31_121
timestamp 1644951705
transform 1 0 39432 0 1 11478
box 0 0 1 1
use contact_31  contact_31_122
timestamp 1644951705
transform 1 0 39432 0 1 10418
box 0 0 1 1
use contact_31  contact_31_123
timestamp 1644951705
transform 1 0 36464 0 1 1938
box 0 0 1 1
use contact_31  contact_31_124
timestamp 1644951705
transform 1 0 36464 0 1 3422
box 0 0 1 1
use contact_31  contact_31_125
timestamp 1644951705
transform 1 0 36464 0 1 11478
box 0 0 1 1
use contact_31  contact_31_126
timestamp 1644951705
transform 1 0 36464 0 1 10418
box 0 0 1 1
use contact_31  contact_31_127
timestamp 1644951705
transform 1 0 35192 0 1 10630
box 0 0 1 1
use contact_31  contact_31_128
timestamp 1644951705
transform 1 0 35192 0 1 11690
box 0 0 1 1
use contact_31  contact_31_129
timestamp 1644951705
transform 1 0 33284 0 1 11478
box 0 0 1 1
use contact_31  contact_31_130
timestamp 1644951705
transform 1 0 33284 0 1 10418
box 0 0 1 1
use contact_31  contact_31_131
timestamp 1644951705
transform 1 0 32648 0 1 10418
box 0 0 1 1
use contact_31  contact_31_132
timestamp 1644951705
transform 1 0 32648 0 1 11690
box 0 0 1 1
use contact_31  contact_31_133
timestamp 1644951705
transform 1 0 29892 0 1 11478
box 0 0 1 1
use contact_31  contact_31_134
timestamp 1644951705
transform 1 0 29680 0 1 10630
box 0 0 1 1
use contact_31  contact_31_135
timestamp 1644951705
transform 1 0 26924 0 1 11478
box 0 0 1 1
use contact_31  contact_31_136
timestamp 1644951705
transform 1 0 26924 0 1 10630
box 0 0 1 1
use contact_31  contact_31_137
timestamp 1644951705
transform 1 0 25864 0 1 10418
box 0 0 1 1
use contact_31  contact_31_138
timestamp 1644951705
transform 1 0 25864 0 1 11690
box 0 0 1 1
use contact_31  contact_31_139
timestamp 1644951705
transform 1 0 23956 0 1 11478
box 0 0 1 1
use contact_31  contact_31_140
timestamp 1644951705
transform 1 0 23956 0 1 10418
box 0 0 1 1
use contact_31  contact_31_141
timestamp 1644951705
transform 1 0 23744 0 1 11478
box 0 0 1 1
use contact_31  contact_31_142
timestamp 1644951705
transform 1 0 23744 0 1 10630
box 0 0 1 1
use contact_31  contact_31_143
timestamp 1644951705
transform 1 0 22472 0 1 17414
box 0 0 1 1
use contact_31  contact_31_144
timestamp 1644951705
transform 1 0 22472 0 1 20382
box 0 0 1 1
use contact_31  contact_31_145
timestamp 1644951705
transform 1 0 22684 0 1 29710
box 0 0 1 1
use contact_31  contact_31_146
timestamp 1644951705
transform 1 0 22684 0 1 32678
box 0 0 1 1
use contact_31  contact_31_147
timestamp 1644951705
transform 1 0 22472 0 1 35646
box 0 0 1 1
use contact_31  contact_31_148
timestamp 1644951705
transform 1 0 22472 0 1 32678
box 0 0 1 1
use contact_31  contact_31_149
timestamp 1644951705
transform 1 0 22684 0 1 62782
box 0 0 1 1
use contact_31  contact_31_150
timestamp 1644951705
transform 1 0 22684 0 1 60450
box 0 0 1 1
use contact_31  contact_31_151
timestamp 1644951705
transform 1 0 22472 0 1 57482
box 0 0 1 1
use contact_31  contact_31_152
timestamp 1644951705
transform 1 0 22472 0 1 60238
box 0 0 1 1
use contact_31  contact_31_153
timestamp 1644951705
transform 1 0 22472 0 1 44974
box 0 0 1 1
use contact_31  contact_31_154
timestamp 1644951705
transform 1 0 22472 0 1 47942
box 0 0 1 1
use contact_31  contact_31_155
timestamp 1644951705
transform 1 0 23532 0 1 11690
box 0 0 1 1
use contact_31  contact_31_156
timestamp 1644951705
transform 1 0 23532 0 1 14234
box 0 0 1 1
use contact_31  contact_31_157
timestamp 1644951705
transform 1 0 22472 0 1 29498
box 0 0 1 1
use contact_31  contact_31_158
timestamp 1644951705
transform 1 0 22472 0 1 26530
box 0 0 1 1
use contact_31  contact_31_159
timestamp 1644951705
transform 1 0 22684 0 1 23562
box 0 0 1 1
use contact_31  contact_31_160
timestamp 1644951705
transform 1 0 22684 0 1 26530
box 0 0 1 1
use contact_31  contact_31_161
timestamp 1644951705
transform 1 0 22472 0 1 51334
box 0 0 1 1
use contact_31  contact_31_162
timestamp 1644951705
transform 1 0 22472 0 1 54090
box 0 0 1 1
use contact_31  contact_31_163
timestamp 1644951705
transform 1 0 22684 0 1 35858
box 0 0 1 1
use contact_31  contact_31_164
timestamp 1644951705
transform 1 0 22684 0 1 38826
box 0 0 1 1
use contact_31  contact_31_165
timestamp 1644951705
transform 1 0 22472 0 1 41794
box 0 0 1 1
use contact_31  contact_31_166
timestamp 1644951705
transform 1 0 22472 0 1 38826
box 0 0 1 1
use contact_31  contact_31_167
timestamp 1644951705
transform 1 0 20988 0 1 14234
box 0 0 1 1
use contact_31  contact_31_168
timestamp 1644951705
transform 1 0 20988 0 1 17202
box 0 0 1 1
use contact_31  contact_31_169
timestamp 1644951705
transform 1 0 21200 0 1 20382
box 0 0 1 1
use contact_31  contact_31_170
timestamp 1644951705
transform 1 0 21200 0 1 23350
box 0 0 1 1
use contact_31  contact_31_171
timestamp 1644951705
transform 1 0 20988 0 1 42006
box 0 0 1 1
use contact_31  contact_31_172
timestamp 1644951705
transform 1 0 20988 0 1 44974
box 0 0 1 1
use contact_31  contact_31_173
timestamp 1644951705
transform 1 0 20988 0 1 48154
box 0 0 1 1
use contact_31  contact_31_174
timestamp 1644951705
transform 1 0 20988 0 1 51122
box 0 0 1 1
use contact_31  contact_31_175
timestamp 1644951705
transform 1 0 21200 0 1 57270
box 0 0 1 1
use contact_31  contact_31_176
timestamp 1644951705
transform 1 0 21200 0 1 54302
box 0 0 1 1
use contact_31  contact_31_177
timestamp 1644951705
transform 1 0 22684 0 1 10206
box 0 0 1 1
use contact_31  contact_31_178
timestamp 1644951705
transform 1 0 22684 0 1 10842
box 0 0 1 1
use contact_31  contact_31_179
timestamp 1644951705
transform 1 0 19928 0 1 1938
box 0 0 1 1
use contact_31  contact_31_180
timestamp 1644951705
transform 1 0 19928 0 1 3422
box 0 0 1 1
use contact_31  contact_31_181
timestamp 1644951705
transform 1 0 19292 0 1 9146
box 0 0 1 1
use contact_31  contact_31_182
timestamp 1644951705
transform 1 0 19292 0 1 10842
box 0 0 1 1
use contact_31  contact_31_183
timestamp 1644951705
transform 1 0 18444 0 1 1938
box 0 0 1 1
use contact_31  contact_31_184
timestamp 1644951705
transform 1 0 18444 0 1 3422
box 0 0 1 1
use contact_31  contact_31_185
timestamp 1644951705
transform 1 0 17172 0 1 35858
box 0 0 1 1
use contact_31  contact_31_186
timestamp 1644951705
transform 1 0 17172 0 1 38826
box 0 0 1 1
use contact_31  contact_31_187
timestamp 1644951705
transform 1 0 17172 0 1 39038
box 0 0 1 1
use contact_31  contact_31_188
timestamp 1644951705
transform 1 0 17172 0 1 41794
box 0 0 1 1
use contact_31  contact_31_189
timestamp 1644951705
transform 1 0 16960 0 1 23562
box 0 0 1 1
use contact_31  contact_31_190
timestamp 1644951705
transform 1 0 16960 0 1 26530
box 0 0 1 1
use contact_31  contact_31_191
timestamp 1644951705
transform 1 0 16748 0 1 35646
box 0 0 1 1
use contact_31  contact_31_192
timestamp 1644951705
transform 1 0 16748 0 1 32678
box 0 0 1 1
use contact_31  contact_31_193
timestamp 1644951705
transform 1 0 16324 0 1 14234
box 0 0 1 1
use contact_31  contact_31_194
timestamp 1644951705
transform 1 0 16324 0 1 13810
box 0 0 1 1
use contact_31  contact_31_195
timestamp 1644951705
transform 1 0 16324 0 1 23350
box 0 0 1 1
use contact_31  contact_31_196
timestamp 1644951705
transform 1 0 16324 0 1 20594
box 0 0 1 1
use contact_31  contact_31_197
timestamp 1644951705
transform 1 0 13992 0 1 17202
box 0 0 1 1
use contact_31  contact_31_198
timestamp 1644951705
transform 1 0 13992 0 1 18686
box 0 0 1 1
use contact_31  contact_31_199
timestamp 1644951705
transform 1 0 13992 0 1 20382
box 0 0 1 1
use contact_31  contact_31_200
timestamp 1644951705
transform 1 0 13992 0 1 18898
box 0 0 1 1
use contact_31  contact_31_201
timestamp 1644951705
transform 1 0 13992 0 1 16990
box 0 0 1 1
use contact_31  contact_31_202
timestamp 1644951705
transform 1 0 13992 0 1 15506
box 0 0 1 1
use contact_31  contact_31_203
timestamp 1644951705
transform 1 0 13992 0 1 13810
box 0 0 1 1
use contact_31  contact_31_204
timestamp 1644951705
transform 1 0 13992 0 1 15294
box 0 0 1 1
use contact_31  contact_31_205
timestamp 1644951705
transform 1 0 1908 0 1 7662
box 0 0 1 1
use contact_33  contact_33_0
timestamp 1644951705
transform 1 0 75684 0 1 64266
box 0 0 1 1
use contact_33  contact_33_1
timestamp 1644951705
transform 1 0 636 0 1 454
box 0 0 1 1
use contact_33  contact_33_2
timestamp 1644951705
transform 1 0 75472 0 1 64266
box 0 0 1 1
use contact_33  contact_33_3
timestamp 1644951705
transform 1 0 75472 0 1 63842
box 0 0 1 1
use contact_33  contact_33_4
timestamp 1644951705
transform 1 0 424 0 1 666
box 0 0 1 1
use contact_33  contact_33_5
timestamp 1644951705
transform 1 0 75472 0 1 878
box 0 0 1 1
use contact_33  contact_33_6
timestamp 1644951705
transform 1 0 75260 0 1 63842
box 0 0 1 1
use contact_33  contact_33_7
timestamp 1644951705
transform 1 0 75684 0 1 63842
box 0 0 1 1
use contact_33  contact_33_8
timestamp 1644951705
transform 1 0 75684 0 1 878
box 0 0 1 1
use contact_33  contact_33_9
timestamp 1644951705
transform 1 0 848 0 1 64054
box 0 0 1 1
use contact_33  contact_33_10
timestamp 1644951705
transform 1 0 848 0 1 666
box 0 0 1 1
use contact_33  contact_33_11
timestamp 1644951705
transform 1 0 75260 0 1 64266
box 0 0 1 1
use contact_33  contact_33_12
timestamp 1644951705
transform 1 0 75472 0 1 454
box 0 0 1 1
use contact_33  contact_33_13
timestamp 1644951705
transform 1 0 636 0 1 64054
box 0 0 1 1
use contact_33  contact_33_14
timestamp 1644951705
transform 1 0 636 0 1 666
box 0 0 1 1
use contact_33  contact_33_15
timestamp 1644951705
transform 1 0 75260 0 1 878
box 0 0 1 1
use contact_33  contact_33_16
timestamp 1644951705
transform 1 0 75684 0 1 454
box 0 0 1 1
use contact_33  contact_33_17
timestamp 1644951705
transform 1 0 424 0 1 64266
box 0 0 1 1
use contact_33  contact_33_18
timestamp 1644951705
transform 1 0 75260 0 1 454
box 0 0 1 1
use contact_33  contact_33_19
timestamp 1644951705
transform 1 0 424 0 1 63842
box 0 0 1 1
use contact_33  contact_33_20
timestamp 1644951705
transform 1 0 424 0 1 878
box 0 0 1 1
use contact_33  contact_33_21
timestamp 1644951705
transform 1 0 424 0 1 454
box 0 0 1 1
use contact_33  contact_33_22
timestamp 1644951705
transform 1 0 75684 0 1 64054
box 0 0 1 1
use contact_33  contact_33_23
timestamp 1644951705
transform 1 0 848 0 1 64266
box 0 0 1 1
use contact_33  contact_33_24
timestamp 1644951705
transform 1 0 75472 0 1 64054
box 0 0 1 1
use contact_33  contact_33_25
timestamp 1644951705
transform 1 0 75684 0 1 666
box 0 0 1 1
use contact_33  contact_33_26
timestamp 1644951705
transform 1 0 75472 0 1 666
box 0 0 1 1
use contact_33  contact_33_27
timestamp 1644951705
transform 1 0 636 0 1 64266
box 0 0 1 1
use contact_33  contact_33_28
timestamp 1644951705
transform 1 0 75260 0 1 64054
box 0 0 1 1
use contact_33  contact_33_29
timestamp 1644951705
transform 1 0 636 0 1 878
box 0 0 1 1
use contact_33  contact_33_30
timestamp 1644951705
transform 1 0 636 0 1 63842
box 0 0 1 1
use contact_33  contact_33_31
timestamp 1644951705
transform 1 0 75260 0 1 666
box 0 0 1 1
use contact_33  contact_33_32
timestamp 1644951705
transform 1 0 848 0 1 63842
box 0 0 1 1
use contact_33  contact_33_33
timestamp 1644951705
transform 1 0 848 0 1 878
box 0 0 1 1
use contact_33  contact_33_34
timestamp 1644951705
transform 1 0 424 0 1 64054
box 0 0 1 1
use contact_33  contact_33_35
timestamp 1644951705
transform 1 0 848 0 1 454
box 0 0 1 1
use contact_33  contact_33_36
timestamp 1644951705
transform 1 0 74200 0 1 62994
box 0 0 1 1
use contact_33  contact_33_37
timestamp 1644951705
transform 1 0 74624 0 1 1938
box 0 0 1 1
use contact_33  contact_33_38
timestamp 1644951705
transform 1 0 1908 0 1 63206
box 0 0 1 1
use contact_33  contact_33_39
timestamp 1644951705
transform 1 0 1908 0 1 62782
box 0 0 1 1
use contact_33  contact_33_40
timestamp 1644951705
transform 1 0 1696 0 1 62782
box 0 0 1 1
use contact_33  contact_33_41
timestamp 1644951705
transform 1 0 1908 0 1 1726
box 0 0 1 1
use contact_33  contact_33_42
timestamp 1644951705
transform 1 0 1696 0 1 63206
box 0 0 1 1
use contact_33  contact_33_43
timestamp 1644951705
transform 1 0 74200 0 1 1938
box 0 0 1 1
use contact_33  contact_33_44
timestamp 1644951705
transform 1 0 1696 0 1 1726
box 0 0 1 1
use contact_33  contact_33_45
timestamp 1644951705
transform 1 0 74412 0 1 62994
box 0 0 1 1
use contact_33  contact_33_46
timestamp 1644951705
transform 1 0 74200 0 1 1514
box 0 0 1 1
use contact_33  contact_33_47
timestamp 1644951705
transform 1 0 1484 0 1 62994
box 0 0 1 1
use contact_33  contact_33_48
timestamp 1644951705
transform 1 0 74624 0 1 63206
box 0 0 1 1
use contact_33  contact_33_49
timestamp 1644951705
transform 1 0 74624 0 1 62782
box 0 0 1 1
use contact_33  contact_33_50
timestamp 1644951705
transform 1 0 74412 0 1 1938
box 0 0 1 1
use contact_33  contact_33_51
timestamp 1644951705
transform 1 0 1484 0 1 1938
box 0 0 1 1
use contact_33  contact_33_52
timestamp 1644951705
transform 1 0 74412 0 1 1514
box 0 0 1 1
use contact_33  contact_33_53
timestamp 1644951705
transform 1 0 74200 0 1 63206
box 0 0 1 1
use contact_33  contact_33_54
timestamp 1644951705
transform 1 0 1696 0 1 62994
box 0 0 1 1
use contact_33  contact_33_55
timestamp 1644951705
transform 1 0 1484 0 1 1514
box 0 0 1 1
use contact_33  contact_33_56
timestamp 1644951705
transform 1 0 74200 0 1 62782
box 0 0 1 1
use contact_33  contact_33_57
timestamp 1644951705
transform 1 0 74624 0 1 1726
box 0 0 1 1
use contact_33  contact_33_58
timestamp 1644951705
transform 1 0 1908 0 1 62994
box 0 0 1 1
use contact_33  contact_33_59
timestamp 1644951705
transform 1 0 1696 0 1 1938
box 0 0 1 1
use contact_33  contact_33_60
timestamp 1644951705
transform 1 0 74200 0 1 1726
box 0 0 1 1
use contact_33  contact_33_61
timestamp 1644951705
transform 1 0 1484 0 1 63206
box 0 0 1 1
use contact_33  contact_33_62
timestamp 1644951705
transform 1 0 74412 0 1 62782
box 0 0 1 1
use contact_33  contact_33_63
timestamp 1644951705
transform 1 0 1908 0 1 1938
box 0 0 1 1
use contact_33  contact_33_64
timestamp 1644951705
transform 1 0 1484 0 1 62782
box 0 0 1 1
use contact_33  contact_33_65
timestamp 1644951705
transform 1 0 1908 0 1 1514
box 0 0 1 1
use contact_33  contact_33_66
timestamp 1644951705
transform 1 0 1484 0 1 1726
box 0 0 1 1
use contact_33  contact_33_67
timestamp 1644951705
transform 1 0 74412 0 1 63206
box 0 0 1 1
use contact_33  contact_33_68
timestamp 1644951705
transform 1 0 74624 0 1 62994
box 0 0 1 1
use contact_33  contact_33_69
timestamp 1644951705
transform 1 0 1696 0 1 1514
box 0 0 1 1
use contact_33  contact_33_70
timestamp 1644951705
transform 1 0 74412 0 1 1726
box 0 0 1 1
use contact_33  contact_33_71
timestamp 1644951705
transform 1 0 74624 0 1 1514
box 0 0 1 1
use contact_31  contact_31_206
timestamp 1644951705
transform 1 0 13568 0 1 12962
box 0 0 1 1
use contact_31  contact_31_207
timestamp 1644951705
transform 1 0 45368 0 1 11054
box 0 0 1 1
use contact_31  contact_31_208
timestamp 1644951705
transform 1 0 44944 0 1 11054
box 0 0 1 1
use contact_31  contact_31_209
timestamp 1644951705
transform 1 0 42188 0 1 11054
box 0 0 1 1
use contact_31  contact_31_210
timestamp 1644951705
transform 1 0 41976 0 1 11054
box 0 0 1 1
use contact_31  contact_31_211
timestamp 1644951705
transform 1 0 39220 0 1 11054
box 0 0 1 1
use contact_31  contact_31_212
timestamp 1644951705
transform 1 0 39008 0 1 11054
box 0 0 1 1
use contact_31  contact_31_213
timestamp 1644951705
transform 1 0 36252 0 1 11054
box 0 0 1 1
use contact_31  contact_31_214
timestamp 1644951705
transform 1 0 35616 0 1 11054
box 0 0 1 1
use contact_31  contact_31_215
timestamp 1644951705
transform 1 0 33072 0 1 11054
box 0 0 1 1
use contact_31  contact_31_216
timestamp 1644951705
transform 1 0 32436 0 1 11054
box 0 0 1 1
use contact_31  contact_31_217
timestamp 1644951705
transform 1 0 30104 0 1 11054
box 0 0 1 1
use contact_31  contact_31_218
timestamp 1644951705
transform 1 0 29468 0 1 11054
box 0 0 1 1
use contact_31  contact_31_219
timestamp 1644951705
transform 1 0 26712 0 1 11054
box 0 0 1 1
use contact_31  contact_31_220
timestamp 1644951705
transform 1 0 26288 0 1 11054
box 0 0 1 1
use contact_31  contact_31_221
timestamp 1644951705
transform 1 0 23532 0 1 11054
box 0 0 1 1
use contact_31  contact_31_222
timestamp 1644951705
transform 1 0 23320 0 1 11054
box 0 0 1 1
use contact_31  contact_31_223
timestamp 1644951705
transform 1 0 6360 0 1 7874
box 0 0 1 1
use contact_31  contact_31_224
timestamp 1644951705
transform 1 0 18020 0 1 2786
box 0 0 1 1
use contact_31  contact_31_225
timestamp 1644951705
transform 1 0 16536 0 1 2786
box 0 0 1 1
use contact_31  contact_31_226
timestamp 1644951705
transform 1 0 41764 0 1 2786
box 0 0 1 1
use contact_31  contact_31_227
timestamp 1644951705
transform 1 0 40280 0 1 2786
box 0 0 1 1
use contact_31  contact_31_228
timestamp 1644951705
transform 1 0 38796 0 1 2786
box 0 0 1 1
use contact_31  contact_31_229
timestamp 1644951705
transform 1 0 37312 0 1 2786
box 0 0 1 1
use contact_31  contact_31_230
timestamp 1644951705
transform 1 0 36040 0 1 2786
box 0 0 1 1
use contact_31  contact_31_231
timestamp 1644951705
transform 1 0 34344 0 1 2786
box 0 0 1 1
use contact_31  contact_31_232
timestamp 1644951705
transform 1 0 32860 0 1 2786
box 0 0 1 1
use contact_31  contact_31_233
timestamp 1644951705
transform 1 0 31376 0 1 2786
box 0 0 1 1
use contact_31  contact_31_234
timestamp 1644951705
transform 1 0 29892 0 1 2786
box 0 0 1 1
use contact_31  contact_31_235
timestamp 1644951705
transform 1 0 28620 0 1 2786
box 0 0 1 1
use contact_31  contact_31_236
timestamp 1644951705
transform 1 0 27136 0 1 2786
box 0 0 1 1
use contact_31  contact_31_237
timestamp 1644951705
transform 1 0 25652 0 1 2786
box 0 0 1 1
use contact_31  contact_31_238
timestamp 1644951705
transform 1 0 24168 0 1 2786
box 0 0 1 1
use contact_31  contact_31_239
timestamp 1644951705
transform 1 0 22472 0 1 2786
box 0 0 1 1
use contact_31  contact_31_240
timestamp 1644951705
transform 1 0 20988 0 1 2786
box 0 0 1 1
use contact_31  contact_31_241
timestamp 1644951705
transform 1 0 19716 0 1 2786
box 0 0 1 1
use contact_18  contact_18_0
timestamp 1644951705
transform 1 0 13619 0 1 18165
box 0 0 1 1
use contact_18  contact_18_1
timestamp 1644951705
transform 1 0 13619 0 1 17673
box 0 0 1 1
use contact_18  contact_18_2
timestamp 1644951705
transform 1 0 13619 0 1 16489
box 0 0 1 1
use contact_18  contact_18_3
timestamp 1644951705
transform 1 0 13619 0 1 15997
box 0 0 1 1
use contact_18  contact_18_4
timestamp 1644951705
transform 1 0 13619 0 1 14813
box 0 0 1 1
use contact_18  contact_18_5
timestamp 1644951705
transform 1 0 13619 0 1 14321
box 0 0 1 1
use contact_18  contact_18_6
timestamp 1644951705
transform 1 0 13619 0 1 13137
box 0 0 1 1
use contact_18  contact_18_7
timestamp 1644951705
transform 1 0 18065 0 1 2911
box 0 0 1 1
use contact_18  contact_18_8
timestamp 1644951705
transform 1 0 16583 0 1 2911
box 0 0 1 1
use contact_18  contact_18_9
timestamp 1644951705
transform 1 0 45327 0 1 11231
box 0 0 1 1
use contact_18  contact_18_10
timestamp 1644951705
transform 1 0 45327 0 1 11231
box 0 0 1 1
use contact_18  contact_18_11
timestamp 1644951705
transform 1 0 45055 0 1 11231
box 0 0 1 1
use contact_18  contact_18_12
timestamp 1644951705
transform 1 0 45055 0 1 11231
box 0 0 1 1
use contact_18  contact_18_13
timestamp 1644951705
transform 1 0 42215 0 1 11231
box 0 0 1 1
use contact_18  contact_18_14
timestamp 1644951705
transform 1 0 42215 0 1 11231
box 0 0 1 1
use contact_18  contact_18_15
timestamp 1644951705
transform 1 0 41943 0 1 11231
box 0 0 1 1
use contact_18  contact_18_16
timestamp 1644951705
transform 1 0 41943 0 1 11231
box 0 0 1 1
use contact_18  contact_18_17
timestamp 1644951705
transform 1 0 39103 0 1 11231
box 0 0 1 1
use contact_18  contact_18_18
timestamp 1644951705
transform 1 0 39103 0 1 11231
box 0 0 1 1
use contact_18  contact_18_19
timestamp 1644951705
transform 1 0 38831 0 1 11231
box 0 0 1 1
use contact_18  contact_18_20
timestamp 1644951705
transform 1 0 38831 0 1 11231
box 0 0 1 1
use contact_18  contact_18_21
timestamp 1644951705
transform 1 0 35991 0 1 11231
box 0 0 1 1
use contact_18  contact_18_22
timestamp 1644951705
transform 1 0 35991 0 1 11231
box 0 0 1 1
use contact_18  contact_18_23
timestamp 1644951705
transform 1 0 35719 0 1 11231
box 0 0 1 1
use contact_18  contact_18_24
timestamp 1644951705
transform 1 0 35719 0 1 11231
box 0 0 1 1
use contact_18  contact_18_25
timestamp 1644951705
transform 1 0 32879 0 1 11231
box 0 0 1 1
use contact_18  contact_18_26
timestamp 1644951705
transform 1 0 32879 0 1 11231
box 0 0 1 1
use contact_18  contact_18_27
timestamp 1644951705
transform 1 0 32607 0 1 11231
box 0 0 1 1
use contact_18  contact_18_28
timestamp 1644951705
transform 1 0 32607 0 1 11231
box 0 0 1 1
use contact_18  contact_18_29
timestamp 1644951705
transform 1 0 29767 0 1 11231
box 0 0 1 1
use contact_18  contact_18_30
timestamp 1644951705
transform 1 0 29767 0 1 11231
box 0 0 1 1
use contact_18  contact_18_31
timestamp 1644951705
transform 1 0 29495 0 1 11231
box 0 0 1 1
use contact_18  contact_18_32
timestamp 1644951705
transform 1 0 29495 0 1 11231
box 0 0 1 1
use contact_18  contact_18_33
timestamp 1644951705
transform 1 0 26655 0 1 11231
box 0 0 1 1
use contact_18  contact_18_34
timestamp 1644951705
transform 1 0 26655 0 1 11231
box 0 0 1 1
use contact_18  contact_18_35
timestamp 1644951705
transform 1 0 26383 0 1 11231
box 0 0 1 1
use contact_18  contact_18_36
timestamp 1644951705
transform 1 0 26383 0 1 11231
box 0 0 1 1
use contact_18  contact_18_37
timestamp 1644951705
transform 1 0 23543 0 1 11231
box 0 0 1 1
use contact_18  contact_18_38
timestamp 1644951705
transform 1 0 23543 0 1 11231
box 0 0 1 1
use contact_18  contact_18_39
timestamp 1644951705
transform 1 0 23271 0 1 11231
box 0 0 1 1
use contact_18  contact_18_40
timestamp 1644951705
transform 1 0 23271 0 1 11231
box 0 0 1 1
use contact_18  contact_18_41
timestamp 1644951705
transform 1 0 41777 0 1 2911
box 0 0 1 1
use contact_18  contact_18_42
timestamp 1644951705
transform 1 0 40295 0 1 2911
box 0 0 1 1
use contact_18  contact_18_43
timestamp 1644951705
transform 1 0 38813 0 1 2911
box 0 0 1 1
use contact_18  contact_18_44
timestamp 1644951705
transform 1 0 37331 0 1 2911
box 0 0 1 1
use contact_18  contact_18_45
timestamp 1644951705
transform 1 0 35849 0 1 2911
box 0 0 1 1
use contact_18  contact_18_46
timestamp 1644951705
transform 1 0 34367 0 1 2911
box 0 0 1 1
use contact_18  contact_18_47
timestamp 1644951705
transform 1 0 32885 0 1 2911
box 0 0 1 1
use contact_18  contact_18_48
timestamp 1644951705
transform 1 0 31403 0 1 2911
box 0 0 1 1
use contact_18  contact_18_49
timestamp 1644951705
transform 1 0 29921 0 1 2911
box 0 0 1 1
use contact_18  contact_18_50
timestamp 1644951705
transform 1 0 28439 0 1 2911
box 0 0 1 1
use contact_18  contact_18_51
timestamp 1644951705
transform 1 0 26957 0 1 2911
box 0 0 1 1
use contact_18  contact_18_52
timestamp 1644951705
transform 1 0 25475 0 1 2911
box 0 0 1 1
use contact_18  contact_18_53
timestamp 1644951705
transform 1 0 23993 0 1 2911
box 0 0 1 1
use contact_18  contact_18_54
timestamp 1644951705
transform 1 0 22511 0 1 2911
box 0 0 1 1
use contact_18  contact_18_55
timestamp 1644951705
transform 1 0 21029 0 1 2911
box 0 0 1 1
use contact_18  contact_18_56
timestamp 1644951705
transform 1 0 19547 0 1 2911
box 0 0 1 1
use contact_18  contact_18_57
timestamp 1644951705
transform 1 0 6443 0 1 7948
box 0 0 1 1
use contact_18  contact_18_58
timestamp 1644951705
transform 1 0 2921 0 1 8163
box 0 0 1 1
use contact_18  contact_18_59
timestamp 1644951705
transform 1 0 2921 0 1 6979
box 0 0 1 1
use contact_18  contact_18_60
timestamp 1644951705
transform 1 0 15598 0 1 18161
box 0 0 1 1
use contact_18  contact_18_61
timestamp 1644951705
transform 1 0 14699 0 1 18161
box 0 0 1 1
use contact_18  contact_18_62
timestamp 1644951705
transform 1 0 15514 0 1 17677
box 0 0 1 1
use contact_18  contact_18_63
timestamp 1644951705
transform 1 0 14699 0 1 17677
box 0 0 1 1
use contact_18  contact_18_64
timestamp 1644951705
transform 1 0 15430 0 1 16485
box 0 0 1 1
use contact_18  contact_18_65
timestamp 1644951705
transform 1 0 14699 0 1 16485
box 0 0 1 1
use contact_18  contact_18_66
timestamp 1644951705
transform 1 0 15346 0 1 16001
box 0 0 1 1
use contact_18  contact_18_67
timestamp 1644951705
transform 1 0 14699 0 1 16001
box 0 0 1 1
use contact_18  contact_18_68
timestamp 1644951705
transform 1 0 15262 0 1 14809
box 0 0 1 1
use contact_18  contact_18_69
timestamp 1644951705
transform 1 0 14699 0 1 14809
box 0 0 1 1
use contact_18  contact_18_70
timestamp 1644951705
transform 1 0 15178 0 1 14325
box 0 0 1 1
use contact_18  contact_18_71
timestamp 1644951705
transform 1 0 14699 0 1 14325
box 0 0 1 1
use contact_18  contact_18_72
timestamp 1644951705
transform 1 0 15094 0 1 13133
box 0 0 1 1
use contact_18  contact_18_73
timestamp 1644951705
transform 1 0 14699 0 1 13133
box 0 0 1 1
use contact_18  contact_18_74
timestamp 1644951705
transform 1 0 21458 0 1 12226
box 0 0 1 1
use contact_18  contact_18_75
timestamp 1644951705
transform 1 0 14894 0 1 12226
box 0 0 1 1
use contact_18  contact_18_76
timestamp 1644951705
transform 1 0 73054 0 1 11293
box 0 0 1 1
use contact_18  contact_18_77
timestamp 1644951705
transform 1 0 14894 0 1 11293
box 0 0 1 1
use contact_18  contact_18_78
timestamp 1644951705
transform 1 0 22580 0 1 10552
box 0 0 1 1
use contact_18  contact_18_79
timestamp 1644951705
transform 1 0 14894 0 1 10552
box 0 0 1 1
use contact_29  contact_29_0
timestamp 1644951705
transform 1 0 13328 0 1 2973
box 0 0 1 1
use contact_29  contact_29_1
timestamp 1644951705
transform 1 0 13328 0 1 2973
box 0 0 1 1
use contact_29  contact_29_2
timestamp 1644951705
transform 1 0 13328 0 1 13199
box 0 0 1 1
use data_dff  data_dff_0
timestamp 1644951705
transform 1 0 19406 0 1 2702
box -39 -42 23712 916
use col_addr_dff  col_addr_dff_0
timestamp 1644951705
transform 1 0 16442 0 1 2702
box -39 -42 2964 916
use row_addr_dff  row_addr_dff_0
timestamp 1644951705
transform 1 0 13478 0 1 12928
box -39 -42 1482 7620
use control_logic_multiport  control_logic_multiport_0
timestamp 1644951705
transform 1 0 2780 0 1 6770
box -66 -42 12180 5906
use bank  bank_0
timestamp 1644951705
transform 1 0 15128 0 1 6224
box 0 0 58446 55900
<< labels >>
rlabel metal3 s 2920 6978 3052 7052 4 web
rlabel metal3 s 2920 8162 3052 8236 4 csb
rlabel metal4 s 6360 0 6512 364 4 clk
rlabel metal4 s 19716 0 19868 364 4 din0[0]
rlabel metal4 s 20988 0 21140 364 4 din0[1]
rlabel metal4 s 22472 0 22624 364 4 din0[2]
rlabel metal4 s 24168 0 24320 364 4 din0[3]
rlabel metal4 s 25652 0 25804 364 4 din0[4]
rlabel metal4 s 27136 0 27288 364 4 din0[5]
rlabel metal4 s 28620 0 28772 364 4 din0[6]
rlabel metal4 s 29892 0 30044 364 4 din0[7]
rlabel metal4 s 31376 0 31528 364 4 din0[8]
rlabel metal4 s 32860 0 33012 364 4 din0[9]
rlabel metal4 s 34344 0 34496 364 4 din0[10]
rlabel metal4 s 36040 0 36192 364 4 din0[11]
rlabel metal4 s 37312 0 37464 364 4 din0[12]
rlabel metal4 s 38796 0 38948 364 4 din0[13]
rlabel metal4 s 40280 0 40432 364 4 din0[14]
rlabel metal4 s 41764 0 41916 364 4 din0[15]
rlabel metal4 s 23320 0 23472 364 4 dout0[0]
rlabel metal3 s 23270 11230 23402 11304 4 dout1[0]
rlabel metal4 s 23532 0 23684 364 4 dout0[1]
rlabel metal3 s 23542 11230 23674 11304 4 dout1[1]
rlabel metal4 s 26288 0 26440 364 4 dout0[2]
rlabel metal3 s 26382 11230 26514 11304 4 dout1[2]
rlabel metal4 s 26712 0 26864 364 4 dout0[3]
rlabel metal3 s 26654 11230 26786 11304 4 dout1[3]
rlabel metal4 s 29468 0 29620 364 4 dout0[4]
rlabel metal3 s 29494 11230 29626 11304 4 dout1[4]
rlabel metal4 s 30104 0 30256 364 4 dout0[5]
rlabel metal3 s 29766 11230 29898 11304 4 dout1[5]
rlabel metal4 s 32436 0 32588 364 4 dout0[6]
rlabel metal3 s 32606 11230 32738 11304 4 dout1[6]
rlabel metal4 s 33072 0 33224 364 4 dout0[7]
rlabel metal3 s 32878 11230 33010 11304 4 dout1[7]
rlabel metal4 s 35616 0 35768 364 4 dout0[8]
rlabel metal3 s 35718 11230 35850 11304 4 dout1[8]
rlabel metal4 s 36252 0 36404 364 4 dout0[9]
rlabel metal3 s 35990 11230 36122 11304 4 dout1[9]
rlabel metal4 s 39008 0 39160 364 4 dout0[10]
rlabel metal3 s 38830 11230 38962 11304 4 dout1[10]
rlabel metal4 s 39220 0 39372 364 4 dout0[11]
rlabel metal3 s 39102 11230 39234 11304 4 dout1[11]
rlabel metal4 s 41976 0 42128 364 4 dout0[12]
rlabel metal3 s 41942 11230 42074 11304 4 dout1[12]
rlabel metal4 s 42188 0 42340 364 4 dout0[13]
rlabel metal3 s 42214 11230 42346 11304 4 dout1[13]
rlabel metal4 s 44944 0 45096 364 4 dout0[14]
rlabel metal3 s 45054 11230 45186 11304 4 dout1[14]
rlabel metal4 s 45368 0 45520 364 4 dout0[15]
rlabel metal3 s 45326 11230 45458 11304 4 dout1[15]
rlabel metal4 s 16536 0 16688 364 4 addr0
rlabel metal4 s 18020 0 18172 364 4 addr1
rlabel metal4 s 13568 0 13720 364 4 addr1[2]
rlabel metal3 s 0 14204 364 14356 4 addr1[3]
rlabel metal3 s 0 14628 364 14780 4 addr1[4]
rlabel metal3 s 0 15900 364 16052 4 addr1[5]
rlabel metal3 s 0 16324 364 16476 4 addr1[6]
rlabel metal3 s 0 17596 364 17748 4 addr1[7]
rlabel metal3 s 0 18020 364 18172 4 addr1[8]
rlabel metal4 s 74200 1484 74776 63328 4 vdd
rlabel metal4 s 1484 1484 2060 63328 4 vdd
rlabel metal3 s 1484 1484 74776 2060 4 vdd
rlabel metal3 s 1484 62752 74776 63328 4 vdd
rlabel metal3 s 424 63812 75836 64388 4 gnd
rlabel metal4 s 75260 424 75836 64388 4 gnd
rlabel metal3 s 424 424 75836 1000 4 gnd
rlabel metal4 s 424 424 1000 64388 4 gnd
<< properties >>
string FIXED_BBOX 0 0 75836 64388
string GDS_FILE sram_0rw2r1w_16_128_sky130A.gds
string GDS_END 201790
string GDS_START 128
<< end >>
