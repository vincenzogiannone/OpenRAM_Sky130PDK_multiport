magic
tech sky130A
magscale 1 2
timestamp 1644969367
<< checkpaint >>
rect -1296 -1277 2744 2155
<< nwell >>
rect -36 402 1484 895
<< pwell >>
rect 1338 51 1388 133
<< psubdiff >>
rect 1338 109 1388 133
rect 1338 75 1346 109
rect 1380 75 1388 109
rect 1338 51 1388 75
<< nsubdiff >>
rect 1338 763 1388 787
rect 1338 729 1346 763
rect 1380 729 1388 763
rect 1338 705 1388 729
<< psubdiffcont >>
rect 1346 75 1380 109
<< nsubdiffcont >>
rect 1346 729 1380 763
<< poly >>
rect 114 406 144 456
rect 48 390 144 406
rect 48 356 64 390
rect 98 356 144 390
rect 48 340 144 356
rect 114 199 144 340
<< polycont >>
rect 64 356 98 390
<< locali >>
rect 0 821 1448 855
rect 62 616 96 821
rect 274 616 308 821
rect 490 616 524 821
rect 706 616 740 821
rect 922 616 956 821
rect 1138 616 1172 821
rect 1346 763 1380 821
rect 1346 713 1380 729
rect 48 390 114 406
rect 48 356 64 390
rect 98 356 114 390
rect 48 340 114 356
rect 704 390 738 582
rect 704 356 755 390
rect 704 164 738 356
rect 1346 109 1380 125
rect 62 17 96 64
rect 274 17 308 64
rect 490 17 524 64
rect 706 17 740 64
rect 922 17 956 64
rect 1138 17 1172 64
rect 1346 17 1380 75
rect 0 -17 1448 17
use contact_12  contact_12_0
timestamp 1644969367
transform 1 0 48 0 1 340
box 0 0 1 1
use contact_11  contact_11_0
timestamp 1644969367
transform 1 0 1338 0 1 51
box 0 0 1 1
use contact_10  contact_10_0
timestamp 1644969367
transform 1 0 1338 0 1 705
box 0 0 1 1
use nmos_m11_w0_460_sli_dli_da_p  nmos_m11_w0_460_sli_dli_da_p_0
timestamp 1644969367
transform 1 0 54 0 1 51
box 0 -26 1230 148
use pmos_m11_w1_375_sli_dli_da_p  pmos_m11_w1_375_sli_dli_da_p_0
timestamp 1644969367
transform 1 0 54 0 1 512
box -59 -56 1289 329
<< labels >>
rlabel locali s 81 373 81 373 4 A
rlabel locali s 738 373 738 373 4 Z
rlabel locali s 724 0 724 0 4 gnd
rlabel locali s 724 838 724 838 4 vdd
<< properties >>
string FIXED_BBOX 0 0 1448 838
string GDS_FILE sram_0rw2r1w_32_128_sky130A.gds
string GDS_END 3366828
string GDS_START 3364696
<< end >>
