magic
tech sky130A
magscale 1 2
timestamp 1644949024
<< checkpaint >>
rect -1260 -1286 1842 1403
<< scnmos >>
rect 60 0 90 84
rect 168 0 198 84
rect 276 0 306 84
rect 384 0 414 84
rect 492 0 522 84
<< ndiff >>
rect 0 59 60 84
rect 0 25 8 59
rect 42 25 60 59
rect 0 0 60 25
rect 90 59 168 84
rect 90 25 112 59
rect 146 25 168 59
rect 90 0 168 25
rect 198 59 276 84
rect 198 25 220 59
rect 254 25 276 59
rect 198 0 276 25
rect 306 59 384 84
rect 306 25 328 59
rect 362 25 384 59
rect 306 0 384 25
rect 414 59 492 84
rect 414 25 436 59
rect 470 25 492 59
rect 414 0 492 25
rect 522 59 582 84
rect 522 25 540 59
rect 574 25 582 59
rect 522 0 582 25
<< ndiffc >>
rect 8 25 42 59
rect 112 25 146 59
rect 220 25 254 59
rect 328 25 362 59
rect 436 25 470 59
rect 540 25 574 59
<< poly >>
rect 60 110 522 140
rect 60 84 90 110
rect 168 84 198 110
rect 276 84 306 110
rect 384 84 414 110
rect 492 84 522 110
rect 60 -26 90 0
rect 168 -26 198 0
rect 276 -26 306 0
rect 384 -26 414 0
rect 492 -26 522 0
<< locali >>
rect 112 109 574 143
rect 8 59 42 75
rect 8 9 42 25
rect 112 59 146 109
rect 112 9 146 25
rect 220 59 254 75
rect 220 9 254 25
rect 328 59 362 109
rect 328 9 362 25
rect 436 59 470 75
rect 436 9 470 25
rect 540 59 574 109
rect 540 9 574 25
use contact_8  contact_8_0
timestamp 1644949024
transform 1 0 532 0 1 1
box 0 0 1 1
use contact_8  contact_8_1
timestamp 1644949024
transform 1 0 428 0 1 1
box 0 0 1 1
use contact_8  contact_8_2
timestamp 1644949024
transform 1 0 320 0 1 1
box 0 0 1 1
use contact_8  contact_8_3
timestamp 1644949024
transform 1 0 212 0 1 1
box 0 0 1 1
use contact_8  contact_8_4
timestamp 1644949024
transform 1 0 104 0 1 1
box 0 0 1 1
use contact_8  contact_8_5
timestamp 1644949024
transform 1 0 0 0 1 1
box 0 0 1 1
<< labels >>
rlabel mvvaractor s 291 125 291 125 4 G
rlabel locali s 237 42 237 42 4 S
rlabel locali s 453 42 453 42 4 S
rlabel locali s 25 42 25 42 4 S
rlabel locali s 343 126 343 126 4 D
<< properties >>
string FIXED_BBOX -25 -26 607 143
string GDS_FILE sram_0rw2r1w_4_16_sky130A.gds
string GDS_END 504532
string GDS_START 502920
<< end >>
