magic
tech sky130A
magscale 1 2
timestamp 1644969367
<< checkpaint >>
rect -1260 -1212 51118 3168
<< poly >>
rect 374 287 404 428
rect 1152 367 1182 428
rect 1134 351 1200 367
rect 1134 317 1150 351
rect 1184 317 1200 351
rect 1134 301 1200 317
rect 1930 287 1960 428
rect 2708 367 2738 428
rect 2690 351 2756 367
rect 2690 317 2706 351
rect 2740 317 2756 351
rect 2690 301 2756 317
rect 3486 287 3516 428
rect 4264 367 4294 428
rect 4246 351 4312 367
rect 4246 317 4262 351
rect 4296 317 4312 351
rect 4246 301 4312 317
rect 5042 287 5072 428
rect 5820 367 5850 428
rect 5802 351 5868 367
rect 5802 317 5818 351
rect 5852 317 5868 351
rect 5802 301 5868 317
rect 6598 287 6628 428
rect 7376 367 7406 428
rect 7358 351 7424 367
rect 7358 317 7374 351
rect 7408 317 7424 351
rect 7358 301 7424 317
rect 8154 287 8184 428
rect 8932 367 8962 428
rect 8914 351 8980 367
rect 8914 317 8930 351
rect 8964 317 8980 351
rect 8914 301 8980 317
rect 9710 287 9740 428
rect 10488 367 10518 428
rect 10470 351 10536 367
rect 10470 317 10486 351
rect 10520 317 10536 351
rect 10470 301 10536 317
rect 11266 287 11296 428
rect 12044 367 12074 428
rect 12026 351 12092 367
rect 12026 317 12042 351
rect 12076 317 12092 351
rect 12026 301 12092 317
rect 12822 287 12852 428
rect 13600 367 13630 428
rect 13582 351 13648 367
rect 13582 317 13598 351
rect 13632 317 13648 351
rect 13582 301 13648 317
rect 14378 287 14408 428
rect 15156 367 15186 428
rect 15138 351 15204 367
rect 15138 317 15154 351
rect 15188 317 15204 351
rect 15138 301 15204 317
rect 15934 287 15964 428
rect 16712 367 16742 428
rect 16694 351 16760 367
rect 16694 317 16710 351
rect 16744 317 16760 351
rect 16694 301 16760 317
rect 17490 287 17520 428
rect 18268 367 18298 428
rect 18250 351 18316 367
rect 18250 317 18266 351
rect 18300 317 18316 351
rect 18250 301 18316 317
rect 19046 287 19076 428
rect 19824 367 19854 428
rect 19806 351 19872 367
rect 19806 317 19822 351
rect 19856 317 19872 351
rect 19806 301 19872 317
rect 20602 287 20632 428
rect 21380 367 21410 428
rect 21362 351 21428 367
rect 21362 317 21378 351
rect 21412 317 21428 351
rect 21362 301 21428 317
rect 22158 287 22188 428
rect 22936 367 22966 428
rect 22918 351 22984 367
rect 22918 317 22934 351
rect 22968 317 22984 351
rect 22918 301 22984 317
rect 23714 287 23744 428
rect 24492 367 24522 428
rect 24474 351 24540 367
rect 24474 317 24490 351
rect 24524 317 24540 351
rect 24474 301 24540 317
rect 25270 287 25300 428
rect 26048 367 26078 428
rect 26030 351 26096 367
rect 26030 317 26046 351
rect 26080 317 26096 351
rect 26030 301 26096 317
rect 26826 287 26856 428
rect 27604 367 27634 428
rect 27586 351 27652 367
rect 27586 317 27602 351
rect 27636 317 27652 351
rect 27586 301 27652 317
rect 28382 287 28412 428
rect 29160 367 29190 428
rect 29142 351 29208 367
rect 29142 317 29158 351
rect 29192 317 29208 351
rect 29142 301 29208 317
rect 29938 287 29968 428
rect 30716 367 30746 428
rect 30698 351 30764 367
rect 30698 317 30714 351
rect 30748 317 30764 351
rect 30698 301 30764 317
rect 31494 287 31524 428
rect 32272 367 32302 428
rect 32254 351 32320 367
rect 32254 317 32270 351
rect 32304 317 32320 351
rect 32254 301 32320 317
rect 33050 287 33080 428
rect 33828 367 33858 428
rect 33810 351 33876 367
rect 33810 317 33826 351
rect 33860 317 33876 351
rect 33810 301 33876 317
rect 34606 287 34636 428
rect 35384 367 35414 428
rect 35366 351 35432 367
rect 35366 317 35382 351
rect 35416 317 35432 351
rect 35366 301 35432 317
rect 36162 287 36192 428
rect 36940 367 36970 428
rect 36922 351 36988 367
rect 36922 317 36938 351
rect 36972 317 36988 351
rect 36922 301 36988 317
rect 37718 287 37748 428
rect 38496 367 38526 428
rect 38478 351 38544 367
rect 38478 317 38494 351
rect 38528 317 38544 351
rect 38478 301 38544 317
rect 39274 287 39304 428
rect 40052 367 40082 428
rect 40034 351 40100 367
rect 40034 317 40050 351
rect 40084 317 40100 351
rect 40034 301 40100 317
rect 40830 287 40860 428
rect 41608 367 41638 428
rect 41590 351 41656 367
rect 41590 317 41606 351
rect 41640 317 41656 351
rect 41590 301 41656 317
rect 42386 287 42416 428
rect 43164 367 43194 428
rect 43146 351 43212 367
rect 43146 317 43162 351
rect 43196 317 43212 351
rect 43146 301 43212 317
rect 43942 287 43972 428
rect 44720 367 44750 428
rect 44702 351 44768 367
rect 44702 317 44718 351
rect 44752 317 44768 351
rect 44702 301 44768 317
rect 45498 287 45528 428
rect 46276 367 46306 428
rect 46258 351 46324 367
rect 46258 317 46274 351
rect 46308 317 46324 351
rect 46258 301 46324 317
rect 47054 287 47084 428
rect 47832 367 47862 428
rect 47814 351 47880 367
rect 47814 317 47830 351
rect 47864 317 47880 351
rect 47814 301 47880 317
rect 48610 287 48640 428
rect 49388 367 49418 428
rect 49370 351 49436 367
rect 49370 317 49386 351
rect 49420 317 49436 351
rect 49370 301 49436 317
rect 356 271 422 287
rect 356 237 372 271
rect 406 237 422 271
rect 356 221 422 237
rect 1912 271 1978 287
rect 1912 237 1928 271
rect 1962 237 1978 271
rect 1912 221 1978 237
rect 3468 271 3534 287
rect 3468 237 3484 271
rect 3518 237 3534 271
rect 3468 221 3534 237
rect 5024 271 5090 287
rect 5024 237 5040 271
rect 5074 237 5090 271
rect 5024 221 5090 237
rect 6580 271 6646 287
rect 6580 237 6596 271
rect 6630 237 6646 271
rect 6580 221 6646 237
rect 8136 271 8202 287
rect 8136 237 8152 271
rect 8186 237 8202 271
rect 8136 221 8202 237
rect 9692 271 9758 287
rect 9692 237 9708 271
rect 9742 237 9758 271
rect 9692 221 9758 237
rect 11248 271 11314 287
rect 11248 237 11264 271
rect 11298 237 11314 271
rect 11248 221 11314 237
rect 12804 271 12870 287
rect 12804 237 12820 271
rect 12854 237 12870 271
rect 12804 221 12870 237
rect 14360 271 14426 287
rect 14360 237 14376 271
rect 14410 237 14426 271
rect 14360 221 14426 237
rect 15916 271 15982 287
rect 15916 237 15932 271
rect 15966 237 15982 271
rect 15916 221 15982 237
rect 17472 271 17538 287
rect 17472 237 17488 271
rect 17522 237 17538 271
rect 17472 221 17538 237
rect 19028 271 19094 287
rect 19028 237 19044 271
rect 19078 237 19094 271
rect 19028 221 19094 237
rect 20584 271 20650 287
rect 20584 237 20600 271
rect 20634 237 20650 271
rect 20584 221 20650 237
rect 22140 271 22206 287
rect 22140 237 22156 271
rect 22190 237 22206 271
rect 22140 221 22206 237
rect 23696 271 23762 287
rect 23696 237 23712 271
rect 23746 237 23762 271
rect 23696 221 23762 237
rect 25252 271 25318 287
rect 25252 237 25268 271
rect 25302 237 25318 271
rect 25252 221 25318 237
rect 26808 271 26874 287
rect 26808 237 26824 271
rect 26858 237 26874 271
rect 26808 221 26874 237
rect 28364 271 28430 287
rect 28364 237 28380 271
rect 28414 237 28430 271
rect 28364 221 28430 237
rect 29920 271 29986 287
rect 29920 237 29936 271
rect 29970 237 29986 271
rect 29920 221 29986 237
rect 31476 271 31542 287
rect 31476 237 31492 271
rect 31526 237 31542 271
rect 31476 221 31542 237
rect 33032 271 33098 287
rect 33032 237 33048 271
rect 33082 237 33098 271
rect 33032 221 33098 237
rect 34588 271 34654 287
rect 34588 237 34604 271
rect 34638 237 34654 271
rect 34588 221 34654 237
rect 36144 271 36210 287
rect 36144 237 36160 271
rect 36194 237 36210 271
rect 36144 221 36210 237
rect 37700 271 37766 287
rect 37700 237 37716 271
rect 37750 237 37766 271
rect 37700 221 37766 237
rect 39256 271 39322 287
rect 39256 237 39272 271
rect 39306 237 39322 271
rect 39256 221 39322 237
rect 40812 271 40878 287
rect 40812 237 40828 271
rect 40862 237 40878 271
rect 40812 221 40878 237
rect 42368 271 42434 287
rect 42368 237 42384 271
rect 42418 237 42434 271
rect 42368 221 42434 237
rect 43924 271 43990 287
rect 43924 237 43940 271
rect 43974 237 43990 271
rect 43924 221 43990 237
rect 45480 271 45546 287
rect 45480 237 45496 271
rect 45530 237 45546 271
rect 45480 221 45546 237
rect 47036 271 47102 287
rect 47036 237 47052 271
rect 47086 237 47102 271
rect 47036 221 47102 237
rect 48592 271 48658 287
rect 48592 237 48608 271
rect 48642 237 48658 271
rect 48592 221 48658 237
<< polycont >>
rect 1150 317 1184 351
rect 2706 317 2740 351
rect 4262 317 4296 351
rect 5818 317 5852 351
rect 7374 317 7408 351
rect 8930 317 8964 351
rect 10486 317 10520 351
rect 12042 317 12076 351
rect 13598 317 13632 351
rect 15154 317 15188 351
rect 16710 317 16744 351
rect 18266 317 18300 351
rect 19822 317 19856 351
rect 21378 317 21412 351
rect 22934 317 22968 351
rect 24490 317 24524 351
rect 26046 317 26080 351
rect 27602 317 27636 351
rect 29158 317 29192 351
rect 30714 317 30748 351
rect 32270 317 32304 351
rect 33826 317 33860 351
rect 35382 317 35416 351
rect 36938 317 36972 351
rect 38494 317 38528 351
rect 40050 317 40084 351
rect 41606 317 41640 351
rect 43162 317 43196 351
rect 44718 317 44752 351
rect 46274 317 46308 351
rect 47830 317 47864 351
rect 49386 317 49420 351
rect 372 237 406 271
rect 1928 237 1962 271
rect 3484 237 3518 271
rect 5040 237 5074 271
rect 6596 237 6630 271
rect 8152 237 8186 271
rect 9708 237 9742 271
rect 11264 237 11298 271
rect 12820 237 12854 271
rect 14376 237 14410 271
rect 15932 237 15966 271
rect 17488 237 17522 271
rect 19044 237 19078 271
rect 20600 237 20634 271
rect 22156 237 22190 271
rect 23712 237 23746 271
rect 25268 237 25302 271
rect 26824 237 26858 271
rect 28380 237 28414 271
rect 29936 237 29970 271
rect 31492 237 31526 271
rect 33048 237 33082 271
rect 34604 237 34638 271
rect 36160 237 36194 271
rect 37716 237 37750 271
rect 39272 237 39306 271
rect 40828 237 40862 271
rect 42384 237 42418 271
rect 43940 237 43974 271
rect 45496 237 45530 271
rect 47052 237 47086 271
rect 48608 237 48642 271
<< locali >>
rect 1134 351 1200 367
rect 1134 317 1150 351
rect 1184 317 1200 351
rect 1134 301 1200 317
rect 2690 351 2756 367
rect 2690 317 2706 351
rect 2740 317 2756 351
rect 2690 301 2756 317
rect 4246 351 4312 367
rect 4246 317 4262 351
rect 4296 317 4312 351
rect 4246 301 4312 317
rect 5802 351 5868 367
rect 5802 317 5818 351
rect 5852 317 5868 351
rect 5802 301 5868 317
rect 7358 351 7424 367
rect 7358 317 7374 351
rect 7408 317 7424 351
rect 7358 301 7424 317
rect 8914 351 8980 367
rect 8914 317 8930 351
rect 8964 317 8980 351
rect 8914 301 8980 317
rect 10470 351 10536 367
rect 10470 317 10486 351
rect 10520 317 10536 351
rect 10470 301 10536 317
rect 12026 351 12092 367
rect 12026 317 12042 351
rect 12076 317 12092 351
rect 12026 301 12092 317
rect 13582 351 13648 367
rect 13582 317 13598 351
rect 13632 317 13648 351
rect 13582 301 13648 317
rect 15138 351 15204 367
rect 15138 317 15154 351
rect 15188 317 15204 351
rect 15138 301 15204 317
rect 16694 351 16760 367
rect 16694 317 16710 351
rect 16744 317 16760 351
rect 16694 301 16760 317
rect 18250 351 18316 367
rect 18250 317 18266 351
rect 18300 317 18316 351
rect 18250 301 18316 317
rect 19806 351 19872 367
rect 19806 317 19822 351
rect 19856 317 19872 351
rect 19806 301 19872 317
rect 21362 351 21428 367
rect 21362 317 21378 351
rect 21412 317 21428 351
rect 21362 301 21428 317
rect 22918 351 22984 367
rect 22918 317 22934 351
rect 22968 317 22984 351
rect 22918 301 22984 317
rect 24474 351 24540 367
rect 24474 317 24490 351
rect 24524 317 24540 351
rect 24474 301 24540 317
rect 26030 351 26096 367
rect 26030 317 26046 351
rect 26080 317 26096 351
rect 26030 301 26096 317
rect 27586 351 27652 367
rect 27586 317 27602 351
rect 27636 317 27652 351
rect 27586 301 27652 317
rect 29142 351 29208 367
rect 29142 317 29158 351
rect 29192 317 29208 351
rect 29142 301 29208 317
rect 30698 351 30764 367
rect 30698 317 30714 351
rect 30748 317 30764 351
rect 30698 301 30764 317
rect 32254 351 32320 367
rect 32254 317 32270 351
rect 32304 317 32320 351
rect 32254 301 32320 317
rect 33810 351 33876 367
rect 33810 317 33826 351
rect 33860 317 33876 351
rect 33810 301 33876 317
rect 35366 351 35432 367
rect 35366 317 35382 351
rect 35416 317 35432 351
rect 35366 301 35432 317
rect 36922 351 36988 367
rect 36922 317 36938 351
rect 36972 317 36988 351
rect 36922 301 36988 317
rect 38478 351 38544 367
rect 38478 317 38494 351
rect 38528 317 38544 351
rect 38478 301 38544 317
rect 40034 351 40100 367
rect 40034 317 40050 351
rect 40084 317 40100 351
rect 40034 301 40100 317
rect 41590 351 41656 367
rect 41590 317 41606 351
rect 41640 317 41656 351
rect 41590 301 41656 317
rect 43146 351 43212 367
rect 43146 317 43162 351
rect 43196 317 43212 351
rect 43146 301 43212 317
rect 44702 351 44768 367
rect 44702 317 44718 351
rect 44752 317 44768 351
rect 44702 301 44768 317
rect 46258 351 46324 367
rect 46258 317 46274 351
rect 46308 317 46324 351
rect 46258 301 46324 317
rect 47814 351 47880 367
rect 47814 317 47830 351
rect 47864 317 47880 351
rect 47814 301 47880 317
rect 49370 351 49436 367
rect 49370 317 49386 351
rect 49420 317 49436 351
rect 49370 301 49436 317
rect 356 271 422 287
rect 356 237 372 271
rect 406 237 422 271
rect 356 221 422 237
rect 1912 271 1978 287
rect 1912 237 1928 271
rect 1962 237 1978 271
rect 1912 221 1978 237
rect 3468 271 3534 287
rect 3468 237 3484 271
rect 3518 237 3534 271
rect 3468 221 3534 237
rect 5024 271 5090 287
rect 5024 237 5040 271
rect 5074 237 5090 271
rect 5024 221 5090 237
rect 6580 271 6646 287
rect 6580 237 6596 271
rect 6630 237 6646 271
rect 6580 221 6646 237
rect 8136 271 8202 287
rect 8136 237 8152 271
rect 8186 237 8202 271
rect 8136 221 8202 237
rect 9692 271 9758 287
rect 9692 237 9708 271
rect 9742 237 9758 271
rect 9692 221 9758 237
rect 11248 271 11314 287
rect 11248 237 11264 271
rect 11298 237 11314 271
rect 11248 221 11314 237
rect 12804 271 12870 287
rect 12804 237 12820 271
rect 12854 237 12870 271
rect 12804 221 12870 237
rect 14360 271 14426 287
rect 14360 237 14376 271
rect 14410 237 14426 271
rect 14360 221 14426 237
rect 15916 271 15982 287
rect 15916 237 15932 271
rect 15966 237 15982 271
rect 15916 221 15982 237
rect 17472 271 17538 287
rect 17472 237 17488 271
rect 17522 237 17538 271
rect 17472 221 17538 237
rect 19028 271 19094 287
rect 19028 237 19044 271
rect 19078 237 19094 271
rect 19028 221 19094 237
rect 20584 271 20650 287
rect 20584 237 20600 271
rect 20634 237 20650 271
rect 20584 221 20650 237
rect 22140 271 22206 287
rect 22140 237 22156 271
rect 22190 237 22206 271
rect 22140 221 22206 237
rect 23696 271 23762 287
rect 23696 237 23712 271
rect 23746 237 23762 271
rect 23696 221 23762 237
rect 25252 271 25318 287
rect 25252 237 25268 271
rect 25302 237 25318 271
rect 25252 221 25318 237
rect 26808 271 26874 287
rect 26808 237 26824 271
rect 26858 237 26874 271
rect 26808 221 26874 237
rect 28364 271 28430 287
rect 28364 237 28380 271
rect 28414 237 28430 271
rect 28364 221 28430 237
rect 29920 271 29986 287
rect 29920 237 29936 271
rect 29970 237 29986 271
rect 29920 221 29986 237
rect 31476 271 31542 287
rect 31476 237 31492 271
rect 31526 237 31542 271
rect 31476 221 31542 237
rect 33032 271 33098 287
rect 33032 237 33048 271
rect 33082 237 33098 271
rect 33032 221 33098 237
rect 34588 271 34654 287
rect 34588 237 34604 271
rect 34638 237 34654 271
rect 34588 221 34654 237
rect 36144 271 36210 287
rect 36144 237 36160 271
rect 36194 237 36210 271
rect 36144 221 36210 237
rect 37700 271 37766 287
rect 37700 237 37716 271
rect 37750 237 37766 271
rect 37700 221 37766 237
rect 39256 271 39322 287
rect 39256 237 39272 271
rect 39306 237 39322 271
rect 39256 221 39322 237
rect 40812 271 40878 287
rect 40812 237 40828 271
rect 40862 237 40878 271
rect 40812 221 40878 237
rect 42368 271 42434 287
rect 42368 237 42384 271
rect 42418 237 42434 271
rect 42368 221 42434 237
rect 43924 271 43990 287
rect 43924 237 43940 271
rect 43974 237 43990 271
rect 43924 221 43990 237
rect 45480 271 45546 287
rect 45480 237 45496 271
rect 45530 237 45546 271
rect 45480 221 45546 237
rect 47036 271 47102 287
rect 47036 237 47052 271
rect 47086 237 47102 271
rect 47036 221 47102 237
rect 48592 271 48658 287
rect 48592 237 48608 271
rect 48642 237 48658 271
rect 48592 221 48658 237
<< viali >>
rect 1150 317 1184 351
rect 2706 317 2740 351
rect 4262 317 4296 351
rect 5818 317 5852 351
rect 7374 317 7408 351
rect 8930 317 8964 351
rect 10486 317 10520 351
rect 12042 317 12076 351
rect 13598 317 13632 351
rect 15154 317 15188 351
rect 16710 317 16744 351
rect 18266 317 18300 351
rect 19822 317 19856 351
rect 21378 317 21412 351
rect 22934 317 22968 351
rect 24490 317 24524 351
rect 26046 317 26080 351
rect 27602 317 27636 351
rect 29158 317 29192 351
rect 30714 317 30748 351
rect 32270 317 32304 351
rect 33826 317 33860 351
rect 35382 317 35416 351
rect 36938 317 36972 351
rect 38494 317 38528 351
rect 40050 317 40084 351
rect 41606 317 41640 351
rect 43162 317 43196 351
rect 44718 317 44752 351
rect 46274 317 46308 351
rect 47830 317 47864 351
rect 49386 317 49420 351
rect 372 237 406 271
rect 1928 237 1962 271
rect 3484 237 3518 271
rect 5040 237 5074 271
rect 6596 237 6630 271
rect 8152 237 8186 271
rect 9708 237 9742 271
rect 11264 237 11298 271
rect 12820 237 12854 271
rect 14376 237 14410 271
rect 15932 237 15966 271
rect 17488 237 17522 271
rect 19044 237 19078 271
rect 20600 237 20634 271
rect 22156 237 22190 271
rect 23712 237 23746 271
rect 25268 237 25302 271
rect 26824 237 26858 271
rect 28380 237 28414 271
rect 29936 237 29970 271
rect 31492 237 31526 271
rect 33048 237 33082 271
rect 34604 237 34638 271
rect 36160 237 36194 271
rect 37716 237 37750 271
rect 39272 237 39306 271
rect 40828 237 40862 271
rect 42384 237 42418 271
rect 43940 237 43974 271
rect 45496 237 45530 271
rect 47052 237 47086 271
rect 48608 237 48642 271
<< metal1 >>
rect 1138 351 1196 357
rect 1138 348 1150 351
rect 0 320 1150 348
rect 1138 317 1150 320
rect 1184 348 1196 351
rect 2694 351 2752 357
rect 2694 348 2706 351
rect 1184 320 2706 348
rect 1184 317 1196 320
rect 1138 311 1196 317
rect 2694 317 2706 320
rect 2740 348 2752 351
rect 4250 351 4308 357
rect 4250 348 4262 351
rect 2740 320 4262 348
rect 2740 317 2752 320
rect 2694 311 2752 317
rect 4250 317 4262 320
rect 4296 348 4308 351
rect 5806 351 5864 357
rect 5806 348 5818 351
rect 4296 320 5818 348
rect 4296 317 4308 320
rect 4250 311 4308 317
rect 5806 317 5818 320
rect 5852 348 5864 351
rect 7362 351 7420 357
rect 7362 348 7374 351
rect 5852 320 7374 348
rect 5852 317 5864 320
rect 5806 311 5864 317
rect 7362 317 7374 320
rect 7408 348 7420 351
rect 8918 351 8976 357
rect 8918 348 8930 351
rect 7408 320 8930 348
rect 7408 317 7420 320
rect 7362 311 7420 317
rect 8918 317 8930 320
rect 8964 348 8976 351
rect 10474 351 10532 357
rect 10474 348 10486 351
rect 8964 320 10486 348
rect 8964 317 8976 320
rect 8918 311 8976 317
rect 10474 317 10486 320
rect 10520 348 10532 351
rect 12030 351 12088 357
rect 12030 348 12042 351
rect 10520 320 12042 348
rect 10520 317 10532 320
rect 10474 311 10532 317
rect 12030 317 12042 320
rect 12076 348 12088 351
rect 13586 351 13644 357
rect 13586 348 13598 351
rect 12076 320 13598 348
rect 12076 317 12088 320
rect 12030 311 12088 317
rect 13586 317 13598 320
rect 13632 348 13644 351
rect 15142 351 15200 357
rect 15142 348 15154 351
rect 13632 320 15154 348
rect 13632 317 13644 320
rect 13586 311 13644 317
rect 15142 317 15154 320
rect 15188 348 15200 351
rect 16698 351 16756 357
rect 16698 348 16710 351
rect 15188 320 16710 348
rect 15188 317 15200 320
rect 15142 311 15200 317
rect 16698 317 16710 320
rect 16744 348 16756 351
rect 18254 351 18312 357
rect 18254 348 18266 351
rect 16744 320 18266 348
rect 16744 317 16756 320
rect 16698 311 16756 317
rect 18254 317 18266 320
rect 18300 348 18312 351
rect 19810 351 19868 357
rect 19810 348 19822 351
rect 18300 320 19822 348
rect 18300 317 18312 320
rect 18254 311 18312 317
rect 19810 317 19822 320
rect 19856 348 19868 351
rect 21366 351 21424 357
rect 21366 348 21378 351
rect 19856 320 21378 348
rect 19856 317 19868 320
rect 19810 311 19868 317
rect 21366 317 21378 320
rect 21412 348 21424 351
rect 22922 351 22980 357
rect 22922 348 22934 351
rect 21412 320 22934 348
rect 21412 317 21424 320
rect 21366 311 21424 317
rect 22922 317 22934 320
rect 22968 348 22980 351
rect 24478 351 24536 357
rect 24478 348 24490 351
rect 22968 320 24490 348
rect 22968 317 22980 320
rect 22922 311 22980 317
rect 24478 317 24490 320
rect 24524 348 24536 351
rect 26034 351 26092 357
rect 26034 348 26046 351
rect 24524 320 26046 348
rect 24524 317 24536 320
rect 24478 311 24536 317
rect 26034 317 26046 320
rect 26080 348 26092 351
rect 27590 351 27648 357
rect 27590 348 27602 351
rect 26080 320 27602 348
rect 26080 317 26092 320
rect 26034 311 26092 317
rect 27590 317 27602 320
rect 27636 348 27648 351
rect 29146 351 29204 357
rect 29146 348 29158 351
rect 27636 320 29158 348
rect 27636 317 27648 320
rect 27590 311 27648 317
rect 29146 317 29158 320
rect 29192 348 29204 351
rect 30702 351 30760 357
rect 30702 348 30714 351
rect 29192 320 30714 348
rect 29192 317 29204 320
rect 29146 311 29204 317
rect 30702 317 30714 320
rect 30748 348 30760 351
rect 32258 351 32316 357
rect 32258 348 32270 351
rect 30748 320 32270 348
rect 30748 317 30760 320
rect 30702 311 30760 317
rect 32258 317 32270 320
rect 32304 348 32316 351
rect 33814 351 33872 357
rect 33814 348 33826 351
rect 32304 320 33826 348
rect 32304 317 32316 320
rect 32258 311 32316 317
rect 33814 317 33826 320
rect 33860 348 33872 351
rect 35370 351 35428 357
rect 35370 348 35382 351
rect 33860 320 35382 348
rect 33860 317 33872 320
rect 33814 311 33872 317
rect 35370 317 35382 320
rect 35416 348 35428 351
rect 36926 351 36984 357
rect 36926 348 36938 351
rect 35416 320 36938 348
rect 35416 317 35428 320
rect 35370 311 35428 317
rect 36926 317 36938 320
rect 36972 348 36984 351
rect 38482 351 38540 357
rect 38482 348 38494 351
rect 36972 320 38494 348
rect 36972 317 36984 320
rect 36926 311 36984 317
rect 38482 317 38494 320
rect 38528 348 38540 351
rect 40038 351 40096 357
rect 40038 348 40050 351
rect 38528 320 40050 348
rect 38528 317 38540 320
rect 38482 311 38540 317
rect 40038 317 40050 320
rect 40084 348 40096 351
rect 41594 351 41652 357
rect 41594 348 41606 351
rect 40084 320 41606 348
rect 40084 317 40096 320
rect 40038 311 40096 317
rect 41594 317 41606 320
rect 41640 348 41652 351
rect 43150 351 43208 357
rect 43150 348 43162 351
rect 41640 320 43162 348
rect 41640 317 41652 320
rect 41594 311 41652 317
rect 43150 317 43162 320
rect 43196 348 43208 351
rect 44706 351 44764 357
rect 44706 348 44718 351
rect 43196 320 44718 348
rect 43196 317 43208 320
rect 43150 311 43208 317
rect 44706 317 44718 320
rect 44752 348 44764 351
rect 46262 351 46320 357
rect 46262 348 46274 351
rect 44752 320 46274 348
rect 44752 317 44764 320
rect 44706 311 44764 317
rect 46262 317 46274 320
rect 46308 348 46320 351
rect 47818 351 47876 357
rect 47818 348 47830 351
rect 46308 320 47830 348
rect 46308 317 46320 320
rect 46262 311 46320 317
rect 47818 317 47830 320
rect 47864 348 47876 351
rect 49374 351 49432 357
rect 49374 348 49386 351
rect 47864 320 49386 348
rect 47864 317 47876 320
rect 47818 311 47876 317
rect 49374 317 49386 320
rect 49420 348 49432 351
rect 49420 320 49792 348
rect 49420 317 49432 320
rect 49374 311 49432 317
rect 360 271 418 277
rect 360 268 372 271
rect 0 240 372 268
rect 360 237 372 240
rect 406 268 418 271
rect 1916 271 1974 277
rect 1916 268 1928 271
rect 406 240 1928 268
rect 406 237 418 240
rect 360 231 418 237
rect 1916 237 1928 240
rect 1962 268 1974 271
rect 3472 271 3530 277
rect 3472 268 3484 271
rect 1962 240 3484 268
rect 1962 237 1974 240
rect 1916 231 1974 237
rect 3472 237 3484 240
rect 3518 268 3530 271
rect 5028 271 5086 277
rect 5028 268 5040 271
rect 3518 240 5040 268
rect 3518 237 3530 240
rect 3472 231 3530 237
rect 5028 237 5040 240
rect 5074 268 5086 271
rect 6584 271 6642 277
rect 6584 268 6596 271
rect 5074 240 6596 268
rect 5074 237 5086 240
rect 5028 231 5086 237
rect 6584 237 6596 240
rect 6630 268 6642 271
rect 8140 271 8198 277
rect 8140 268 8152 271
rect 6630 240 8152 268
rect 6630 237 6642 240
rect 6584 231 6642 237
rect 8140 237 8152 240
rect 8186 268 8198 271
rect 9696 271 9754 277
rect 9696 268 9708 271
rect 8186 240 9708 268
rect 8186 237 8198 240
rect 8140 231 8198 237
rect 9696 237 9708 240
rect 9742 268 9754 271
rect 11252 271 11310 277
rect 11252 268 11264 271
rect 9742 240 11264 268
rect 9742 237 9754 240
rect 9696 231 9754 237
rect 11252 237 11264 240
rect 11298 268 11310 271
rect 12808 271 12866 277
rect 12808 268 12820 271
rect 11298 240 12820 268
rect 11298 237 11310 240
rect 11252 231 11310 237
rect 12808 237 12820 240
rect 12854 268 12866 271
rect 14364 271 14422 277
rect 14364 268 14376 271
rect 12854 240 14376 268
rect 12854 237 12866 240
rect 12808 231 12866 237
rect 14364 237 14376 240
rect 14410 268 14422 271
rect 15920 271 15978 277
rect 15920 268 15932 271
rect 14410 240 15932 268
rect 14410 237 14422 240
rect 14364 231 14422 237
rect 15920 237 15932 240
rect 15966 268 15978 271
rect 17476 271 17534 277
rect 17476 268 17488 271
rect 15966 240 17488 268
rect 15966 237 15978 240
rect 15920 231 15978 237
rect 17476 237 17488 240
rect 17522 268 17534 271
rect 19032 271 19090 277
rect 19032 268 19044 271
rect 17522 240 19044 268
rect 17522 237 17534 240
rect 17476 231 17534 237
rect 19032 237 19044 240
rect 19078 268 19090 271
rect 20588 271 20646 277
rect 20588 268 20600 271
rect 19078 240 20600 268
rect 19078 237 19090 240
rect 19032 231 19090 237
rect 20588 237 20600 240
rect 20634 268 20646 271
rect 22144 271 22202 277
rect 22144 268 22156 271
rect 20634 240 22156 268
rect 20634 237 20646 240
rect 20588 231 20646 237
rect 22144 237 22156 240
rect 22190 268 22202 271
rect 23700 271 23758 277
rect 23700 268 23712 271
rect 22190 240 23712 268
rect 22190 237 22202 240
rect 22144 231 22202 237
rect 23700 237 23712 240
rect 23746 268 23758 271
rect 25256 271 25314 277
rect 25256 268 25268 271
rect 23746 240 25268 268
rect 23746 237 23758 240
rect 23700 231 23758 237
rect 25256 237 25268 240
rect 25302 268 25314 271
rect 26812 271 26870 277
rect 26812 268 26824 271
rect 25302 240 26824 268
rect 25302 237 25314 240
rect 25256 231 25314 237
rect 26812 237 26824 240
rect 26858 268 26870 271
rect 28368 271 28426 277
rect 28368 268 28380 271
rect 26858 240 28380 268
rect 26858 237 26870 240
rect 26812 231 26870 237
rect 28368 237 28380 240
rect 28414 268 28426 271
rect 29924 271 29982 277
rect 29924 268 29936 271
rect 28414 240 29936 268
rect 28414 237 28426 240
rect 28368 231 28426 237
rect 29924 237 29936 240
rect 29970 268 29982 271
rect 31480 271 31538 277
rect 31480 268 31492 271
rect 29970 240 31492 268
rect 29970 237 29982 240
rect 29924 231 29982 237
rect 31480 237 31492 240
rect 31526 268 31538 271
rect 33036 271 33094 277
rect 33036 268 33048 271
rect 31526 240 33048 268
rect 31526 237 31538 240
rect 31480 231 31538 237
rect 33036 237 33048 240
rect 33082 268 33094 271
rect 34592 271 34650 277
rect 34592 268 34604 271
rect 33082 240 34604 268
rect 33082 237 33094 240
rect 33036 231 33094 237
rect 34592 237 34604 240
rect 34638 268 34650 271
rect 36148 271 36206 277
rect 36148 268 36160 271
rect 34638 240 36160 268
rect 34638 237 34650 240
rect 34592 231 34650 237
rect 36148 237 36160 240
rect 36194 268 36206 271
rect 37704 271 37762 277
rect 37704 268 37716 271
rect 36194 240 37716 268
rect 36194 237 36206 240
rect 36148 231 36206 237
rect 37704 237 37716 240
rect 37750 268 37762 271
rect 39260 271 39318 277
rect 39260 268 39272 271
rect 37750 240 39272 268
rect 37750 237 37762 240
rect 37704 231 37762 237
rect 39260 237 39272 240
rect 39306 268 39318 271
rect 40816 271 40874 277
rect 40816 268 40828 271
rect 39306 240 40828 268
rect 39306 237 39318 240
rect 39260 231 39318 237
rect 40816 237 40828 240
rect 40862 268 40874 271
rect 42372 271 42430 277
rect 42372 268 42384 271
rect 40862 240 42384 268
rect 40862 237 40874 240
rect 40816 231 40874 237
rect 42372 237 42384 240
rect 42418 268 42430 271
rect 43928 271 43986 277
rect 43928 268 43940 271
rect 42418 240 43940 268
rect 42418 237 42430 240
rect 42372 231 42430 237
rect 43928 237 43940 240
rect 43974 268 43986 271
rect 45484 271 45542 277
rect 45484 268 45496 271
rect 43974 240 45496 268
rect 43974 237 43986 240
rect 43928 231 43986 237
rect 45484 237 45496 240
rect 45530 268 45542 271
rect 47040 271 47098 277
rect 47040 268 47052 271
rect 45530 240 47052 268
rect 45530 237 45542 240
rect 45484 231 45542 237
rect 47040 237 47052 240
rect 47086 268 47098 271
rect 48596 271 48654 277
rect 48596 268 48608 271
rect 47086 240 48608 268
rect 47086 237 47098 240
rect 47040 231 47098 237
rect 48596 237 48608 240
rect 48642 268 48654 271
rect 48642 240 49792 268
rect 48642 237 48654 240
rect 48596 231 48654 237
rect 66 134 72 186
rect 124 174 130 186
rect 844 174 850 186
rect 124 146 850 174
rect 124 134 130 146
rect 844 134 850 146
rect 902 134 908 186
rect 1622 134 1628 186
rect 1680 174 1686 186
rect 2400 174 2406 186
rect 1680 146 2406 174
rect 1680 134 1686 146
rect 2400 134 2406 146
rect 2458 134 2464 186
rect 3178 134 3184 186
rect 3236 174 3242 186
rect 3956 174 3962 186
rect 3236 146 3962 174
rect 3236 134 3242 146
rect 3956 134 3962 146
rect 4014 134 4020 186
rect 4734 134 4740 186
rect 4792 174 4798 186
rect 5512 174 5518 186
rect 4792 146 5518 174
rect 4792 134 4798 146
rect 5512 134 5518 146
rect 5570 134 5576 186
rect 6290 134 6296 186
rect 6348 174 6354 186
rect 7068 174 7074 186
rect 6348 146 7074 174
rect 6348 134 6354 146
rect 7068 134 7074 146
rect 7126 134 7132 186
rect 7846 134 7852 186
rect 7904 174 7910 186
rect 8624 174 8630 186
rect 7904 146 8630 174
rect 7904 134 7910 146
rect 8624 134 8630 146
rect 8682 134 8688 186
rect 9402 134 9408 186
rect 9460 174 9466 186
rect 10180 174 10186 186
rect 9460 146 10186 174
rect 9460 134 9466 146
rect 10180 134 10186 146
rect 10238 134 10244 186
rect 10958 134 10964 186
rect 11016 174 11022 186
rect 11736 174 11742 186
rect 11016 146 11742 174
rect 11016 134 11022 146
rect 11736 134 11742 146
rect 11794 134 11800 186
rect 12514 134 12520 186
rect 12572 174 12578 186
rect 13292 174 13298 186
rect 12572 146 13298 174
rect 12572 134 12578 146
rect 13292 134 13298 146
rect 13350 134 13356 186
rect 14070 134 14076 186
rect 14128 174 14134 186
rect 14848 174 14854 186
rect 14128 146 14854 174
rect 14128 134 14134 146
rect 14848 134 14854 146
rect 14906 134 14912 186
rect 15626 134 15632 186
rect 15684 174 15690 186
rect 16404 174 16410 186
rect 15684 146 16410 174
rect 15684 134 15690 146
rect 16404 134 16410 146
rect 16462 134 16468 186
rect 17182 134 17188 186
rect 17240 174 17246 186
rect 17960 174 17966 186
rect 17240 146 17966 174
rect 17240 134 17246 146
rect 17960 134 17966 146
rect 18018 134 18024 186
rect 18738 134 18744 186
rect 18796 174 18802 186
rect 19516 174 19522 186
rect 18796 146 19522 174
rect 18796 134 18802 146
rect 19516 134 19522 146
rect 19574 134 19580 186
rect 20294 134 20300 186
rect 20352 174 20358 186
rect 21072 174 21078 186
rect 20352 146 21078 174
rect 20352 134 20358 146
rect 21072 134 21078 146
rect 21130 134 21136 186
rect 21850 134 21856 186
rect 21908 174 21914 186
rect 22628 174 22634 186
rect 21908 146 22634 174
rect 21908 134 21914 146
rect 22628 134 22634 146
rect 22686 134 22692 186
rect 23406 134 23412 186
rect 23464 174 23470 186
rect 24184 174 24190 186
rect 23464 146 24190 174
rect 23464 134 23470 146
rect 24184 134 24190 146
rect 24242 134 24248 186
rect 24962 134 24968 186
rect 25020 174 25026 186
rect 25740 174 25746 186
rect 25020 146 25746 174
rect 25020 134 25026 146
rect 25740 134 25746 146
rect 25798 134 25804 186
rect 26518 134 26524 186
rect 26576 174 26582 186
rect 27296 174 27302 186
rect 26576 146 27302 174
rect 26576 134 26582 146
rect 27296 134 27302 146
rect 27354 134 27360 186
rect 28074 134 28080 186
rect 28132 174 28138 186
rect 28852 174 28858 186
rect 28132 146 28858 174
rect 28132 134 28138 146
rect 28852 134 28858 146
rect 28910 134 28916 186
rect 29630 134 29636 186
rect 29688 174 29694 186
rect 30408 174 30414 186
rect 29688 146 30414 174
rect 29688 134 29694 146
rect 30408 134 30414 146
rect 30466 134 30472 186
rect 31186 134 31192 186
rect 31244 174 31250 186
rect 31964 174 31970 186
rect 31244 146 31970 174
rect 31244 134 31250 146
rect 31964 134 31970 146
rect 32022 134 32028 186
rect 32742 134 32748 186
rect 32800 174 32806 186
rect 33520 174 33526 186
rect 32800 146 33526 174
rect 32800 134 32806 146
rect 33520 134 33526 146
rect 33578 134 33584 186
rect 34298 134 34304 186
rect 34356 174 34362 186
rect 35076 174 35082 186
rect 34356 146 35082 174
rect 34356 134 34362 146
rect 35076 134 35082 146
rect 35134 134 35140 186
rect 35854 134 35860 186
rect 35912 174 35918 186
rect 36632 174 36638 186
rect 35912 146 36638 174
rect 35912 134 35918 146
rect 36632 134 36638 146
rect 36690 134 36696 186
rect 37410 134 37416 186
rect 37468 174 37474 186
rect 38188 174 38194 186
rect 37468 146 38194 174
rect 37468 134 37474 146
rect 38188 134 38194 146
rect 38246 134 38252 186
rect 38966 134 38972 186
rect 39024 174 39030 186
rect 39744 174 39750 186
rect 39024 146 39750 174
rect 39024 134 39030 146
rect 39744 134 39750 146
rect 39802 134 39808 186
rect 40522 134 40528 186
rect 40580 174 40586 186
rect 41300 174 41306 186
rect 40580 146 41306 174
rect 40580 134 40586 146
rect 41300 134 41306 146
rect 41358 134 41364 186
rect 42078 134 42084 186
rect 42136 174 42142 186
rect 42856 174 42862 186
rect 42136 146 42862 174
rect 42136 134 42142 146
rect 42856 134 42862 146
rect 42914 134 42920 186
rect 43634 134 43640 186
rect 43692 174 43698 186
rect 44412 174 44418 186
rect 43692 146 44418 174
rect 43692 134 43698 146
rect 44412 134 44418 146
rect 44470 134 44476 186
rect 45190 134 45196 186
rect 45248 174 45254 186
rect 45968 174 45974 186
rect 45248 146 45974 174
rect 45248 134 45254 146
rect 45968 134 45974 146
rect 46026 134 46032 186
rect 46746 134 46752 186
rect 46804 174 46810 186
rect 47524 174 47530 186
rect 46804 146 47530 174
rect 46804 134 46810 146
rect 47524 134 47530 146
rect 47582 134 47588 186
rect 48302 134 48308 186
rect 48360 174 48366 186
rect 49080 174 49086 186
rect 48360 146 49086 174
rect 48360 134 48366 146
rect 49080 134 49086 146
rect 49138 134 49144 186
rect 676 54 682 106
rect 734 94 740 106
rect 1454 94 1460 106
rect 734 66 1460 94
rect 734 54 740 66
rect 1454 54 1460 66
rect 1512 54 1518 106
rect 2232 54 2238 106
rect 2290 94 2296 106
rect 3010 94 3016 106
rect 2290 66 3016 94
rect 2290 54 2296 66
rect 3010 54 3016 66
rect 3068 54 3074 106
rect 3788 54 3794 106
rect 3846 94 3852 106
rect 4566 94 4572 106
rect 3846 66 4572 94
rect 3846 54 3852 66
rect 4566 54 4572 66
rect 4624 54 4630 106
rect 5344 54 5350 106
rect 5402 94 5408 106
rect 6122 94 6128 106
rect 5402 66 6128 94
rect 5402 54 5408 66
rect 6122 54 6128 66
rect 6180 54 6186 106
rect 6900 54 6906 106
rect 6958 94 6964 106
rect 7678 94 7684 106
rect 6958 66 7684 94
rect 6958 54 6964 66
rect 7678 54 7684 66
rect 7736 54 7742 106
rect 8456 54 8462 106
rect 8514 94 8520 106
rect 9234 94 9240 106
rect 8514 66 9240 94
rect 8514 54 8520 66
rect 9234 54 9240 66
rect 9292 54 9298 106
rect 10012 54 10018 106
rect 10070 94 10076 106
rect 10790 94 10796 106
rect 10070 66 10796 94
rect 10070 54 10076 66
rect 10790 54 10796 66
rect 10848 54 10854 106
rect 11568 54 11574 106
rect 11626 94 11632 106
rect 12346 94 12352 106
rect 11626 66 12352 94
rect 11626 54 11632 66
rect 12346 54 12352 66
rect 12404 54 12410 106
rect 13124 54 13130 106
rect 13182 94 13188 106
rect 13902 94 13908 106
rect 13182 66 13908 94
rect 13182 54 13188 66
rect 13902 54 13908 66
rect 13960 54 13966 106
rect 14680 54 14686 106
rect 14738 94 14744 106
rect 15458 94 15464 106
rect 14738 66 15464 94
rect 14738 54 14744 66
rect 15458 54 15464 66
rect 15516 54 15522 106
rect 16236 54 16242 106
rect 16294 94 16300 106
rect 17014 94 17020 106
rect 16294 66 17020 94
rect 16294 54 16300 66
rect 17014 54 17020 66
rect 17072 54 17078 106
rect 17792 54 17798 106
rect 17850 94 17856 106
rect 18570 94 18576 106
rect 17850 66 18576 94
rect 17850 54 17856 66
rect 18570 54 18576 66
rect 18628 54 18634 106
rect 19348 54 19354 106
rect 19406 94 19412 106
rect 20126 94 20132 106
rect 19406 66 20132 94
rect 19406 54 19412 66
rect 20126 54 20132 66
rect 20184 54 20190 106
rect 20904 54 20910 106
rect 20962 94 20968 106
rect 21682 94 21688 106
rect 20962 66 21688 94
rect 20962 54 20968 66
rect 21682 54 21688 66
rect 21740 54 21746 106
rect 22460 54 22466 106
rect 22518 94 22524 106
rect 23238 94 23244 106
rect 22518 66 23244 94
rect 22518 54 22524 66
rect 23238 54 23244 66
rect 23296 54 23302 106
rect 24016 54 24022 106
rect 24074 94 24080 106
rect 24794 94 24800 106
rect 24074 66 24800 94
rect 24074 54 24080 66
rect 24794 54 24800 66
rect 24852 54 24858 106
rect 25572 54 25578 106
rect 25630 94 25636 106
rect 26350 94 26356 106
rect 25630 66 26356 94
rect 25630 54 25636 66
rect 26350 54 26356 66
rect 26408 54 26414 106
rect 27128 54 27134 106
rect 27186 94 27192 106
rect 27906 94 27912 106
rect 27186 66 27912 94
rect 27186 54 27192 66
rect 27906 54 27912 66
rect 27964 54 27970 106
rect 28684 54 28690 106
rect 28742 94 28748 106
rect 29462 94 29468 106
rect 28742 66 29468 94
rect 28742 54 28748 66
rect 29462 54 29468 66
rect 29520 54 29526 106
rect 30240 54 30246 106
rect 30298 94 30304 106
rect 31018 94 31024 106
rect 30298 66 31024 94
rect 30298 54 30304 66
rect 31018 54 31024 66
rect 31076 54 31082 106
rect 31796 54 31802 106
rect 31854 94 31860 106
rect 32574 94 32580 106
rect 31854 66 32580 94
rect 31854 54 31860 66
rect 32574 54 32580 66
rect 32632 54 32638 106
rect 33352 54 33358 106
rect 33410 94 33416 106
rect 34130 94 34136 106
rect 33410 66 34136 94
rect 33410 54 33416 66
rect 34130 54 34136 66
rect 34188 54 34194 106
rect 34908 54 34914 106
rect 34966 94 34972 106
rect 35686 94 35692 106
rect 34966 66 35692 94
rect 34966 54 34972 66
rect 35686 54 35692 66
rect 35744 54 35750 106
rect 36464 54 36470 106
rect 36522 94 36528 106
rect 37242 94 37248 106
rect 36522 66 37248 94
rect 36522 54 36528 66
rect 37242 54 37248 66
rect 37300 54 37306 106
rect 38020 54 38026 106
rect 38078 94 38084 106
rect 38798 94 38804 106
rect 38078 66 38804 94
rect 38078 54 38084 66
rect 38798 54 38804 66
rect 38856 54 38862 106
rect 39576 54 39582 106
rect 39634 94 39640 106
rect 40354 94 40360 106
rect 39634 66 40360 94
rect 39634 54 39640 66
rect 40354 54 40360 66
rect 40412 54 40418 106
rect 41132 54 41138 106
rect 41190 94 41196 106
rect 41910 94 41916 106
rect 41190 66 41916 94
rect 41190 54 41196 66
rect 41910 54 41916 66
rect 41968 54 41974 106
rect 42688 54 42694 106
rect 42746 94 42752 106
rect 43466 94 43472 106
rect 42746 66 43472 94
rect 42746 54 42752 66
rect 43466 54 43472 66
rect 43524 54 43530 106
rect 44244 54 44250 106
rect 44302 94 44308 106
rect 45022 94 45028 106
rect 44302 66 45028 94
rect 44302 54 44308 66
rect 45022 54 45028 66
rect 45080 54 45086 106
rect 45800 54 45806 106
rect 45858 94 45864 106
rect 46578 94 46584 106
rect 45858 66 46584 94
rect 45858 54 45864 66
rect 46578 54 46584 66
rect 46636 54 46642 106
rect 47356 54 47362 106
rect 47414 94 47420 106
rect 48134 94 48140 106
rect 47414 66 48140 94
rect 47414 54 47420 66
rect 48134 54 48140 66
rect 48192 54 48198 106
rect 48912 54 48918 106
rect 48970 94 48976 106
rect 49690 94 49696 106
rect 48970 66 49696 94
rect 48970 54 48976 66
rect 49690 54 49696 66
rect 49748 54 49754 106
<< via1 >>
rect 72 134 124 186
rect 850 134 902 186
rect 1628 134 1680 186
rect 2406 134 2458 186
rect 3184 134 3236 186
rect 3962 134 4014 186
rect 4740 134 4792 186
rect 5518 134 5570 186
rect 6296 134 6348 186
rect 7074 134 7126 186
rect 7852 134 7904 186
rect 8630 134 8682 186
rect 9408 134 9460 186
rect 10186 134 10238 186
rect 10964 134 11016 186
rect 11742 134 11794 186
rect 12520 134 12572 186
rect 13298 134 13350 186
rect 14076 134 14128 186
rect 14854 134 14906 186
rect 15632 134 15684 186
rect 16410 134 16462 186
rect 17188 134 17240 186
rect 17966 134 18018 186
rect 18744 134 18796 186
rect 19522 134 19574 186
rect 20300 134 20352 186
rect 21078 134 21130 186
rect 21856 134 21908 186
rect 22634 134 22686 186
rect 23412 134 23464 186
rect 24190 134 24242 186
rect 24968 134 25020 186
rect 25746 134 25798 186
rect 26524 134 26576 186
rect 27302 134 27354 186
rect 28080 134 28132 186
rect 28858 134 28910 186
rect 29636 134 29688 186
rect 30414 134 30466 186
rect 31192 134 31244 186
rect 31970 134 32022 186
rect 32748 134 32800 186
rect 33526 134 33578 186
rect 34304 134 34356 186
rect 35082 134 35134 186
rect 35860 134 35912 186
rect 36638 134 36690 186
rect 37416 134 37468 186
rect 38194 134 38246 186
rect 38972 134 39024 186
rect 39750 134 39802 186
rect 40528 134 40580 186
rect 41306 134 41358 186
rect 42084 134 42136 186
rect 42862 134 42914 186
rect 43640 134 43692 186
rect 44418 134 44470 186
rect 45196 134 45248 186
rect 45974 134 46026 186
rect 46752 134 46804 186
rect 47530 134 47582 186
rect 48308 134 48360 186
rect 49086 134 49138 186
rect 682 54 734 106
rect 1460 54 1512 106
rect 2238 54 2290 106
rect 3016 54 3068 106
rect 3794 54 3846 106
rect 4572 54 4624 106
rect 5350 54 5402 106
rect 6128 54 6180 106
rect 6906 54 6958 106
rect 7684 54 7736 106
rect 8462 54 8514 106
rect 9240 54 9292 106
rect 10018 54 10070 106
rect 10796 54 10848 106
rect 11574 54 11626 106
rect 12352 54 12404 106
rect 13130 54 13182 106
rect 13908 54 13960 106
rect 14686 54 14738 106
rect 15464 54 15516 106
rect 16242 54 16294 106
rect 17020 54 17072 106
rect 17798 54 17850 106
rect 18576 54 18628 106
rect 19354 54 19406 106
rect 20132 54 20184 106
rect 20910 54 20962 106
rect 21688 54 21740 106
rect 22466 54 22518 106
rect 23244 54 23296 106
rect 24022 54 24074 106
rect 24800 54 24852 106
rect 25578 54 25630 106
rect 26356 54 26408 106
rect 27134 54 27186 106
rect 27912 54 27964 106
rect 28690 54 28742 106
rect 29468 54 29520 106
rect 30246 54 30298 106
rect 31024 54 31076 106
rect 31802 54 31854 106
rect 32580 54 32632 106
rect 33358 54 33410 106
rect 34136 54 34188 106
rect 34914 54 34966 106
rect 35692 54 35744 106
rect 36470 54 36522 106
rect 37248 54 37300 106
rect 38026 54 38078 106
rect 38804 54 38856 106
rect 39582 54 39634 106
rect 40360 54 40412 106
rect 41138 54 41190 106
rect 41916 54 41968 106
rect 42694 54 42746 106
rect 43472 54 43524 106
rect 44250 54 44302 106
rect 45028 54 45080 106
rect 45806 54 45858 106
rect 46584 54 46636 106
rect 47362 54 47414 106
rect 48140 54 48192 106
rect 48918 54 48970 106
rect 49696 54 49748 106
<< metal2 >>
rect 84 1852 112 1908
rect 694 1852 722 1908
rect 862 1852 890 1908
rect 1472 1852 1500 1908
rect 1640 1852 1668 1908
rect 2250 1852 2278 1908
rect 2418 1852 2446 1908
rect 3028 1852 3056 1908
rect 3196 1852 3224 1908
rect 3806 1852 3834 1908
rect 3974 1852 4002 1908
rect 4584 1852 4612 1908
rect 4752 1852 4780 1908
rect 5362 1852 5390 1908
rect 5530 1852 5558 1908
rect 6140 1852 6168 1908
rect 6308 1852 6336 1908
rect 6918 1852 6946 1908
rect 7086 1852 7114 1908
rect 7696 1852 7724 1908
rect 7864 1852 7892 1908
rect 8474 1852 8502 1908
rect 8642 1852 8670 1908
rect 9252 1852 9280 1908
rect 9420 1852 9448 1908
rect 10030 1852 10058 1908
rect 10198 1852 10226 1908
rect 10808 1852 10836 1908
rect 10976 1852 11004 1908
rect 11586 1852 11614 1908
rect 11754 1852 11782 1908
rect 12364 1852 12392 1908
rect 12532 1852 12560 1908
rect 13142 1852 13170 1908
rect 13310 1852 13338 1908
rect 13920 1852 13948 1908
rect 14088 1852 14116 1908
rect 14698 1852 14726 1908
rect 14866 1852 14894 1908
rect 15476 1852 15504 1908
rect 15644 1852 15672 1908
rect 16254 1852 16282 1908
rect 16422 1852 16450 1908
rect 17032 1852 17060 1908
rect 17200 1852 17228 1908
rect 17810 1852 17838 1908
rect 17978 1852 18006 1908
rect 18588 1852 18616 1908
rect 18756 1852 18784 1908
rect 19366 1852 19394 1908
rect 19534 1852 19562 1908
rect 20144 1852 20172 1908
rect 20312 1852 20340 1908
rect 20922 1852 20950 1908
rect 21090 1852 21118 1908
rect 21700 1852 21728 1908
rect 21868 1852 21896 1908
rect 22478 1852 22506 1908
rect 22646 1852 22674 1908
rect 23256 1852 23284 1908
rect 23424 1852 23452 1908
rect 24034 1852 24062 1908
rect 24202 1852 24230 1908
rect 24812 1852 24840 1908
rect 24980 1852 25008 1908
rect 25590 1852 25618 1908
rect 25758 1852 25786 1908
rect 26368 1852 26396 1908
rect 26536 1852 26564 1908
rect 27146 1852 27174 1908
rect 27314 1852 27342 1908
rect 27924 1852 27952 1908
rect 28092 1852 28120 1908
rect 28702 1852 28730 1908
rect 28870 1852 28898 1908
rect 29480 1852 29508 1908
rect 29648 1852 29676 1908
rect 30258 1852 30286 1908
rect 30426 1852 30454 1908
rect 31036 1852 31064 1908
rect 31204 1852 31232 1908
rect 31814 1852 31842 1908
rect 31982 1852 32010 1908
rect 32592 1852 32620 1908
rect 32760 1852 32788 1908
rect 33370 1852 33398 1908
rect 33538 1852 33566 1908
rect 34148 1852 34176 1908
rect 34316 1852 34344 1908
rect 34926 1852 34954 1908
rect 35094 1852 35122 1908
rect 35704 1852 35732 1908
rect 35872 1852 35900 1908
rect 36482 1852 36510 1908
rect 36650 1852 36678 1908
rect 37260 1852 37288 1908
rect 37428 1852 37456 1908
rect 38038 1852 38066 1908
rect 38206 1852 38234 1908
rect 38816 1852 38844 1908
rect 38984 1852 39012 1908
rect 39594 1852 39622 1908
rect 39762 1852 39790 1908
rect 40372 1852 40400 1908
rect 40540 1852 40568 1908
rect 41150 1852 41178 1908
rect 41318 1852 41346 1908
rect 41928 1852 41956 1908
rect 42096 1852 42124 1908
rect 42706 1852 42734 1908
rect 42874 1852 42902 1908
rect 43484 1852 43512 1908
rect 43652 1852 43680 1908
rect 44262 1852 44290 1908
rect 44430 1852 44458 1908
rect 45040 1852 45068 1908
rect 45208 1852 45236 1908
rect 45818 1852 45846 1908
rect 45986 1852 46014 1908
rect 46596 1852 46624 1908
rect 46764 1852 46792 1908
rect 47374 1852 47402 1908
rect 47542 1852 47570 1908
rect 48152 1852 48180 1908
rect 48320 1852 48348 1908
rect 48930 1852 48958 1908
rect 49098 1852 49126 1908
rect 49708 1852 49736 1908
rect 84 192 112 400
rect 72 186 124 192
rect 72 128 124 134
rect 694 112 722 400
rect 862 192 890 400
rect 850 186 902 192
rect 850 128 902 134
rect 1472 112 1500 400
rect 1640 192 1668 400
rect 1628 186 1680 192
rect 1628 128 1680 134
rect 2250 112 2278 400
rect 2418 192 2446 400
rect 2406 186 2458 192
rect 2406 128 2458 134
rect 3028 112 3056 400
rect 3196 192 3224 400
rect 3184 186 3236 192
rect 3184 128 3236 134
rect 3806 112 3834 400
rect 3974 192 4002 400
rect 3962 186 4014 192
rect 3962 128 4014 134
rect 4584 112 4612 400
rect 4752 192 4780 400
rect 4740 186 4792 192
rect 4740 128 4792 134
rect 5362 112 5390 400
rect 5530 192 5558 400
rect 5518 186 5570 192
rect 5518 128 5570 134
rect 6140 112 6168 400
rect 6308 192 6336 400
rect 6296 186 6348 192
rect 6296 128 6348 134
rect 6918 112 6946 400
rect 7086 192 7114 400
rect 7074 186 7126 192
rect 7074 128 7126 134
rect 7696 112 7724 400
rect 7864 192 7892 400
rect 7852 186 7904 192
rect 7852 128 7904 134
rect 8474 112 8502 400
rect 8642 192 8670 400
rect 8630 186 8682 192
rect 8630 128 8682 134
rect 9252 112 9280 400
rect 9420 192 9448 400
rect 9408 186 9460 192
rect 9408 128 9460 134
rect 10030 112 10058 400
rect 10198 192 10226 400
rect 10186 186 10238 192
rect 10186 128 10238 134
rect 10808 112 10836 400
rect 10976 192 11004 400
rect 10964 186 11016 192
rect 10964 128 11016 134
rect 11586 112 11614 400
rect 11754 192 11782 400
rect 11742 186 11794 192
rect 11742 128 11794 134
rect 12364 112 12392 400
rect 12532 192 12560 400
rect 12520 186 12572 192
rect 12520 128 12572 134
rect 13142 112 13170 400
rect 13310 192 13338 400
rect 13298 186 13350 192
rect 13298 128 13350 134
rect 13920 112 13948 400
rect 14088 192 14116 400
rect 14076 186 14128 192
rect 14076 128 14128 134
rect 14698 112 14726 400
rect 14866 192 14894 400
rect 14854 186 14906 192
rect 14854 128 14906 134
rect 15476 112 15504 400
rect 15644 192 15672 400
rect 15632 186 15684 192
rect 15632 128 15684 134
rect 16254 112 16282 400
rect 16422 192 16450 400
rect 16410 186 16462 192
rect 16410 128 16462 134
rect 17032 112 17060 400
rect 17200 192 17228 400
rect 17188 186 17240 192
rect 17188 128 17240 134
rect 17810 112 17838 400
rect 17978 192 18006 400
rect 17966 186 18018 192
rect 17966 128 18018 134
rect 18588 112 18616 400
rect 18756 192 18784 400
rect 18744 186 18796 192
rect 18744 128 18796 134
rect 19366 112 19394 400
rect 19534 192 19562 400
rect 19522 186 19574 192
rect 19522 128 19574 134
rect 20144 112 20172 400
rect 20312 192 20340 400
rect 20300 186 20352 192
rect 20300 128 20352 134
rect 20922 112 20950 400
rect 21090 192 21118 400
rect 21078 186 21130 192
rect 21078 128 21130 134
rect 21700 112 21728 400
rect 21868 192 21896 400
rect 21856 186 21908 192
rect 21856 128 21908 134
rect 22478 112 22506 400
rect 22646 192 22674 400
rect 22634 186 22686 192
rect 22634 128 22686 134
rect 23256 112 23284 400
rect 23424 192 23452 400
rect 23412 186 23464 192
rect 23412 128 23464 134
rect 24034 112 24062 400
rect 24202 192 24230 400
rect 24190 186 24242 192
rect 24190 128 24242 134
rect 24812 112 24840 400
rect 24980 192 25008 400
rect 24968 186 25020 192
rect 24968 128 25020 134
rect 25590 112 25618 400
rect 25758 192 25786 400
rect 25746 186 25798 192
rect 25746 128 25798 134
rect 26368 112 26396 400
rect 26536 192 26564 400
rect 26524 186 26576 192
rect 26524 128 26576 134
rect 27146 112 27174 400
rect 27314 192 27342 400
rect 27302 186 27354 192
rect 27302 128 27354 134
rect 27924 112 27952 400
rect 28092 192 28120 400
rect 28080 186 28132 192
rect 28080 128 28132 134
rect 28702 112 28730 400
rect 28870 192 28898 400
rect 28858 186 28910 192
rect 28858 128 28910 134
rect 29480 112 29508 400
rect 29648 192 29676 400
rect 29636 186 29688 192
rect 29636 128 29688 134
rect 30258 112 30286 400
rect 30426 192 30454 400
rect 30414 186 30466 192
rect 30414 128 30466 134
rect 31036 112 31064 400
rect 31204 192 31232 400
rect 31192 186 31244 192
rect 31192 128 31244 134
rect 31814 112 31842 400
rect 31982 192 32010 400
rect 31970 186 32022 192
rect 31970 128 32022 134
rect 32592 112 32620 400
rect 32760 192 32788 400
rect 32748 186 32800 192
rect 32748 128 32800 134
rect 33370 112 33398 400
rect 33538 192 33566 400
rect 33526 186 33578 192
rect 33526 128 33578 134
rect 34148 112 34176 400
rect 34316 192 34344 400
rect 34304 186 34356 192
rect 34304 128 34356 134
rect 34926 112 34954 400
rect 35094 192 35122 400
rect 35082 186 35134 192
rect 35082 128 35134 134
rect 35704 112 35732 400
rect 35872 192 35900 400
rect 35860 186 35912 192
rect 35860 128 35912 134
rect 36482 112 36510 400
rect 36650 192 36678 400
rect 36638 186 36690 192
rect 36638 128 36690 134
rect 37260 112 37288 400
rect 37428 192 37456 400
rect 37416 186 37468 192
rect 37416 128 37468 134
rect 38038 112 38066 400
rect 38206 192 38234 400
rect 38194 186 38246 192
rect 38194 128 38246 134
rect 38816 112 38844 400
rect 38984 192 39012 400
rect 38972 186 39024 192
rect 38972 128 39024 134
rect 39594 112 39622 400
rect 39762 192 39790 400
rect 39750 186 39802 192
rect 39750 128 39802 134
rect 40372 112 40400 400
rect 40540 192 40568 400
rect 40528 186 40580 192
rect 40528 128 40580 134
rect 41150 112 41178 400
rect 41318 192 41346 400
rect 41306 186 41358 192
rect 41306 128 41358 134
rect 41928 112 41956 400
rect 42096 192 42124 400
rect 42084 186 42136 192
rect 42084 128 42136 134
rect 42706 112 42734 400
rect 42874 192 42902 400
rect 42862 186 42914 192
rect 42862 128 42914 134
rect 43484 112 43512 400
rect 43652 192 43680 400
rect 43640 186 43692 192
rect 43640 128 43692 134
rect 44262 112 44290 400
rect 44430 192 44458 400
rect 44418 186 44470 192
rect 44418 128 44470 134
rect 45040 112 45068 400
rect 45208 192 45236 400
rect 45196 186 45248 192
rect 45196 128 45248 134
rect 45818 112 45846 400
rect 45986 192 46014 400
rect 45974 186 46026 192
rect 45974 128 46026 134
rect 46596 112 46624 400
rect 46764 192 46792 400
rect 46752 186 46804 192
rect 46752 128 46804 134
rect 47374 112 47402 400
rect 47542 192 47570 400
rect 47530 186 47582 192
rect 47530 128 47582 134
rect 48152 112 48180 400
rect 48320 192 48348 400
rect 48308 186 48360 192
rect 48308 128 48360 134
rect 48930 112 48958 400
rect 49098 192 49126 400
rect 49086 186 49138 192
rect 49086 128 49138 134
rect 49708 112 49736 400
rect 682 106 734 112
rect 682 48 734 54
rect 1460 106 1512 112
rect 1460 48 1512 54
rect 2238 106 2290 112
rect 2238 48 2290 54
rect 3016 106 3068 112
rect 3016 48 3068 54
rect 3794 106 3846 112
rect 3794 48 3846 54
rect 4572 106 4624 112
rect 4572 48 4624 54
rect 5350 106 5402 112
rect 5350 48 5402 54
rect 6128 106 6180 112
rect 6128 48 6180 54
rect 6906 106 6958 112
rect 6906 48 6958 54
rect 7684 106 7736 112
rect 7684 48 7736 54
rect 8462 106 8514 112
rect 8462 48 8514 54
rect 9240 106 9292 112
rect 9240 48 9292 54
rect 10018 106 10070 112
rect 10018 48 10070 54
rect 10796 106 10848 112
rect 10796 48 10848 54
rect 11574 106 11626 112
rect 11574 48 11626 54
rect 12352 106 12404 112
rect 12352 48 12404 54
rect 13130 106 13182 112
rect 13130 48 13182 54
rect 13908 106 13960 112
rect 13908 48 13960 54
rect 14686 106 14738 112
rect 14686 48 14738 54
rect 15464 106 15516 112
rect 15464 48 15516 54
rect 16242 106 16294 112
rect 16242 48 16294 54
rect 17020 106 17072 112
rect 17020 48 17072 54
rect 17798 106 17850 112
rect 17798 48 17850 54
rect 18576 106 18628 112
rect 18576 48 18628 54
rect 19354 106 19406 112
rect 19354 48 19406 54
rect 20132 106 20184 112
rect 20132 48 20184 54
rect 20910 106 20962 112
rect 20910 48 20962 54
rect 21688 106 21740 112
rect 21688 48 21740 54
rect 22466 106 22518 112
rect 22466 48 22518 54
rect 23244 106 23296 112
rect 23244 48 23296 54
rect 24022 106 24074 112
rect 24022 48 24074 54
rect 24800 106 24852 112
rect 24800 48 24852 54
rect 25578 106 25630 112
rect 25578 48 25630 54
rect 26356 106 26408 112
rect 26356 48 26408 54
rect 27134 106 27186 112
rect 27134 48 27186 54
rect 27912 106 27964 112
rect 27912 48 27964 54
rect 28690 106 28742 112
rect 28690 48 28742 54
rect 29468 106 29520 112
rect 29468 48 29520 54
rect 30246 106 30298 112
rect 30246 48 30298 54
rect 31024 106 31076 112
rect 31024 48 31076 54
rect 31802 106 31854 112
rect 31802 48 31854 54
rect 32580 106 32632 112
rect 32580 48 32632 54
rect 33358 106 33410 112
rect 33358 48 33410 54
rect 34136 106 34188 112
rect 34136 48 34188 54
rect 34914 106 34966 112
rect 34914 48 34966 54
rect 35692 106 35744 112
rect 35692 48 35744 54
rect 36470 106 36522 112
rect 36470 48 36522 54
rect 37248 106 37300 112
rect 37248 48 37300 54
rect 38026 106 38078 112
rect 38026 48 38078 54
rect 38804 106 38856 112
rect 38804 48 38856 54
rect 39582 106 39634 112
rect 39582 48 39634 54
rect 40360 106 40412 112
rect 40360 48 40412 54
rect 41138 106 41190 112
rect 41138 48 41190 54
rect 41916 106 41968 112
rect 41916 48 41968 54
rect 42694 106 42746 112
rect 42694 48 42746 54
rect 43472 106 43524 112
rect 43472 48 43524 54
rect 44250 106 44302 112
rect 44250 48 44302 54
rect 45028 106 45080 112
rect 45028 48 45080 54
rect 45806 106 45858 112
rect 45806 48 45858 54
rect 46584 106 46636 112
rect 46584 48 46636 54
rect 47362 106 47414 112
rect 47362 48 47414 54
rect 48140 106 48192 112
rect 48140 48 48192 54
rect 48918 106 48970 112
rect 48918 48 48970 54
rect 49696 106 49748 112
rect 49696 48 49748 54
<< metal3 >>
rect 712 1122 844 1196
rect 1490 1122 1622 1196
rect 2268 1122 2400 1196
rect 3046 1122 3178 1196
rect 3824 1122 3956 1196
rect 4602 1122 4734 1196
rect 5380 1122 5512 1196
rect 6158 1122 6290 1196
rect 6936 1122 7068 1196
rect 7714 1122 7846 1196
rect 8492 1122 8624 1196
rect 9270 1122 9402 1196
rect 10048 1122 10180 1196
rect 10826 1122 10958 1196
rect 11604 1122 11736 1196
rect 12382 1122 12514 1196
rect 13160 1122 13292 1196
rect 13938 1122 14070 1196
rect 14716 1122 14848 1196
rect 15494 1122 15626 1196
rect 16272 1122 16404 1196
rect 17050 1122 17182 1196
rect 17828 1122 17960 1196
rect 18606 1122 18738 1196
rect 19384 1122 19516 1196
rect 20162 1122 20294 1196
rect 20940 1122 21072 1196
rect 21718 1122 21850 1196
rect 22496 1122 22628 1196
rect 23274 1122 23406 1196
rect 24052 1122 24184 1196
rect 24830 1122 24962 1196
rect 25608 1122 25740 1196
rect 26386 1122 26518 1196
rect 27164 1122 27296 1196
rect 27942 1122 28074 1196
rect 28720 1122 28852 1196
rect 29498 1122 29630 1196
rect 30276 1122 30408 1196
rect 31054 1122 31186 1196
rect 31832 1122 31964 1196
rect 32610 1122 32742 1196
rect 33388 1122 33520 1196
rect 34166 1122 34298 1196
rect 34944 1122 35076 1196
rect 35722 1122 35854 1196
rect 36500 1122 36632 1196
rect 37278 1122 37410 1196
rect 38056 1122 38188 1196
rect 38834 1122 38966 1196
rect 39612 1122 39744 1196
rect 40390 1122 40522 1196
rect 41168 1122 41300 1196
rect 41946 1122 42078 1196
rect 42724 1122 42856 1196
rect 43502 1122 43634 1196
rect 44280 1122 44412 1196
rect 45058 1122 45190 1196
rect 45836 1122 45968 1196
rect 46614 1122 46746 1196
rect 47392 1122 47524 1196
rect 48170 1122 48302 1196
rect 48948 1122 49080 1196
rect 49726 1122 49858 1196
use contact_14  contact_14_0
timestamp 1644969367
transform 1 0 49690 0 1 48
box 0 0 1 1
use contact_14  contact_14_1
timestamp 1644969367
transform 1 0 49080 0 1 128
box 0 0 1 1
use contact_14  contact_14_2
timestamp 1644969367
transform 1 0 48912 0 1 48
box 0 0 1 1
use contact_14  contact_14_3
timestamp 1644969367
transform 1 0 48302 0 1 128
box 0 0 1 1
use contact_14  contact_14_4
timestamp 1644969367
transform 1 0 48134 0 1 48
box 0 0 1 1
use contact_14  contact_14_5
timestamp 1644969367
transform 1 0 47524 0 1 128
box 0 0 1 1
use contact_14  contact_14_6
timestamp 1644969367
transform 1 0 47356 0 1 48
box 0 0 1 1
use contact_14  contact_14_7
timestamp 1644969367
transform 1 0 46746 0 1 128
box 0 0 1 1
use contact_14  contact_14_8
timestamp 1644969367
transform 1 0 46578 0 1 48
box 0 0 1 1
use contact_14  contact_14_9
timestamp 1644969367
transform 1 0 45968 0 1 128
box 0 0 1 1
use contact_14  contact_14_10
timestamp 1644969367
transform 1 0 45800 0 1 48
box 0 0 1 1
use contact_14  contact_14_11
timestamp 1644969367
transform 1 0 45190 0 1 128
box 0 0 1 1
use contact_14  contact_14_12
timestamp 1644969367
transform 1 0 45022 0 1 48
box 0 0 1 1
use contact_14  contact_14_13
timestamp 1644969367
transform 1 0 44412 0 1 128
box 0 0 1 1
use contact_14  contact_14_14
timestamp 1644969367
transform 1 0 44244 0 1 48
box 0 0 1 1
use contact_14  contact_14_15
timestamp 1644969367
transform 1 0 43634 0 1 128
box 0 0 1 1
use contact_14  contact_14_16
timestamp 1644969367
transform 1 0 43466 0 1 48
box 0 0 1 1
use contact_14  contact_14_17
timestamp 1644969367
transform 1 0 42856 0 1 128
box 0 0 1 1
use contact_14  contact_14_18
timestamp 1644969367
transform 1 0 42688 0 1 48
box 0 0 1 1
use contact_14  contact_14_19
timestamp 1644969367
transform 1 0 42078 0 1 128
box 0 0 1 1
use contact_14  contact_14_20
timestamp 1644969367
transform 1 0 41910 0 1 48
box 0 0 1 1
use contact_14  contact_14_21
timestamp 1644969367
transform 1 0 41300 0 1 128
box 0 0 1 1
use contact_14  contact_14_22
timestamp 1644969367
transform 1 0 41132 0 1 48
box 0 0 1 1
use contact_14  contact_14_23
timestamp 1644969367
transform 1 0 40522 0 1 128
box 0 0 1 1
use contact_14  contact_14_24
timestamp 1644969367
transform 1 0 40354 0 1 48
box 0 0 1 1
use contact_14  contact_14_25
timestamp 1644969367
transform 1 0 39744 0 1 128
box 0 0 1 1
use contact_14  contact_14_26
timestamp 1644969367
transform 1 0 39576 0 1 48
box 0 0 1 1
use contact_14  contact_14_27
timestamp 1644969367
transform 1 0 38966 0 1 128
box 0 0 1 1
use contact_14  contact_14_28
timestamp 1644969367
transform 1 0 38798 0 1 48
box 0 0 1 1
use contact_14  contact_14_29
timestamp 1644969367
transform 1 0 38188 0 1 128
box 0 0 1 1
use contact_14  contact_14_30
timestamp 1644969367
transform 1 0 38020 0 1 48
box 0 0 1 1
use contact_14  contact_14_31
timestamp 1644969367
transform 1 0 37410 0 1 128
box 0 0 1 1
use contact_14  contact_14_32
timestamp 1644969367
transform 1 0 37242 0 1 48
box 0 0 1 1
use contact_14  contact_14_33
timestamp 1644969367
transform 1 0 36632 0 1 128
box 0 0 1 1
use contact_14  contact_14_34
timestamp 1644969367
transform 1 0 36464 0 1 48
box 0 0 1 1
use contact_14  contact_14_35
timestamp 1644969367
transform 1 0 35854 0 1 128
box 0 0 1 1
use contact_14  contact_14_36
timestamp 1644969367
transform 1 0 35686 0 1 48
box 0 0 1 1
use contact_14  contact_14_37
timestamp 1644969367
transform 1 0 35076 0 1 128
box 0 0 1 1
use contact_14  contact_14_38
timestamp 1644969367
transform 1 0 34908 0 1 48
box 0 0 1 1
use contact_14  contact_14_39
timestamp 1644969367
transform 1 0 34298 0 1 128
box 0 0 1 1
use contact_14  contact_14_40
timestamp 1644969367
transform 1 0 34130 0 1 48
box 0 0 1 1
use contact_14  contact_14_41
timestamp 1644969367
transform 1 0 33520 0 1 128
box 0 0 1 1
use contact_14  contact_14_42
timestamp 1644969367
transform 1 0 33352 0 1 48
box 0 0 1 1
use contact_14  contact_14_43
timestamp 1644969367
transform 1 0 32742 0 1 128
box 0 0 1 1
use contact_14  contact_14_44
timestamp 1644969367
transform 1 0 32574 0 1 48
box 0 0 1 1
use contact_14  contact_14_45
timestamp 1644969367
transform 1 0 31964 0 1 128
box 0 0 1 1
use contact_14  contact_14_46
timestamp 1644969367
transform 1 0 31796 0 1 48
box 0 0 1 1
use contact_14  contact_14_47
timestamp 1644969367
transform 1 0 31186 0 1 128
box 0 0 1 1
use contact_14  contact_14_48
timestamp 1644969367
transform 1 0 31018 0 1 48
box 0 0 1 1
use contact_14  contact_14_49
timestamp 1644969367
transform 1 0 30408 0 1 128
box 0 0 1 1
use contact_14  contact_14_50
timestamp 1644969367
transform 1 0 30240 0 1 48
box 0 0 1 1
use contact_14  contact_14_51
timestamp 1644969367
transform 1 0 29630 0 1 128
box 0 0 1 1
use contact_14  contact_14_52
timestamp 1644969367
transform 1 0 29462 0 1 48
box 0 0 1 1
use contact_14  contact_14_53
timestamp 1644969367
transform 1 0 28852 0 1 128
box 0 0 1 1
use contact_14  contact_14_54
timestamp 1644969367
transform 1 0 28684 0 1 48
box 0 0 1 1
use contact_14  contact_14_55
timestamp 1644969367
transform 1 0 28074 0 1 128
box 0 0 1 1
use contact_14  contact_14_56
timestamp 1644969367
transform 1 0 27906 0 1 48
box 0 0 1 1
use contact_14  contact_14_57
timestamp 1644969367
transform 1 0 27296 0 1 128
box 0 0 1 1
use contact_14  contact_14_58
timestamp 1644969367
transform 1 0 27128 0 1 48
box 0 0 1 1
use contact_14  contact_14_59
timestamp 1644969367
transform 1 0 26518 0 1 128
box 0 0 1 1
use contact_14  contact_14_60
timestamp 1644969367
transform 1 0 26350 0 1 48
box 0 0 1 1
use contact_14  contact_14_61
timestamp 1644969367
transform 1 0 25740 0 1 128
box 0 0 1 1
use contact_14  contact_14_62
timestamp 1644969367
transform 1 0 25572 0 1 48
box 0 0 1 1
use contact_14  contact_14_63
timestamp 1644969367
transform 1 0 24962 0 1 128
box 0 0 1 1
use contact_14  contact_14_64
timestamp 1644969367
transform 1 0 24794 0 1 48
box 0 0 1 1
use contact_14  contact_14_65
timestamp 1644969367
transform 1 0 24184 0 1 128
box 0 0 1 1
use contact_14  contact_14_66
timestamp 1644969367
transform 1 0 24016 0 1 48
box 0 0 1 1
use contact_14  contact_14_67
timestamp 1644969367
transform 1 0 23406 0 1 128
box 0 0 1 1
use contact_14  contact_14_68
timestamp 1644969367
transform 1 0 23238 0 1 48
box 0 0 1 1
use contact_14  contact_14_69
timestamp 1644969367
transform 1 0 22628 0 1 128
box 0 0 1 1
use contact_14  contact_14_70
timestamp 1644969367
transform 1 0 22460 0 1 48
box 0 0 1 1
use contact_14  contact_14_71
timestamp 1644969367
transform 1 0 21850 0 1 128
box 0 0 1 1
use contact_14  contact_14_72
timestamp 1644969367
transform 1 0 21682 0 1 48
box 0 0 1 1
use contact_14  contact_14_73
timestamp 1644969367
transform 1 0 21072 0 1 128
box 0 0 1 1
use contact_14  contact_14_74
timestamp 1644969367
transform 1 0 20904 0 1 48
box 0 0 1 1
use contact_14  contact_14_75
timestamp 1644969367
transform 1 0 20294 0 1 128
box 0 0 1 1
use contact_14  contact_14_76
timestamp 1644969367
transform 1 0 20126 0 1 48
box 0 0 1 1
use contact_14  contact_14_77
timestamp 1644969367
transform 1 0 19516 0 1 128
box 0 0 1 1
use contact_14  contact_14_78
timestamp 1644969367
transform 1 0 19348 0 1 48
box 0 0 1 1
use contact_14  contact_14_79
timestamp 1644969367
transform 1 0 18738 0 1 128
box 0 0 1 1
use contact_14  contact_14_80
timestamp 1644969367
transform 1 0 18570 0 1 48
box 0 0 1 1
use contact_14  contact_14_81
timestamp 1644969367
transform 1 0 17960 0 1 128
box 0 0 1 1
use contact_14  contact_14_82
timestamp 1644969367
transform 1 0 17792 0 1 48
box 0 0 1 1
use contact_14  contact_14_83
timestamp 1644969367
transform 1 0 17182 0 1 128
box 0 0 1 1
use contact_14  contact_14_84
timestamp 1644969367
transform 1 0 17014 0 1 48
box 0 0 1 1
use contact_14  contact_14_85
timestamp 1644969367
transform 1 0 16404 0 1 128
box 0 0 1 1
use contact_14  contact_14_86
timestamp 1644969367
transform 1 0 16236 0 1 48
box 0 0 1 1
use contact_14  contact_14_87
timestamp 1644969367
transform 1 0 15626 0 1 128
box 0 0 1 1
use contact_14  contact_14_88
timestamp 1644969367
transform 1 0 15458 0 1 48
box 0 0 1 1
use contact_14  contact_14_89
timestamp 1644969367
transform 1 0 14848 0 1 128
box 0 0 1 1
use contact_14  contact_14_90
timestamp 1644969367
transform 1 0 14680 0 1 48
box 0 0 1 1
use contact_14  contact_14_91
timestamp 1644969367
transform 1 0 14070 0 1 128
box 0 0 1 1
use contact_14  contact_14_92
timestamp 1644969367
transform 1 0 13902 0 1 48
box 0 0 1 1
use contact_14  contact_14_93
timestamp 1644969367
transform 1 0 13292 0 1 128
box 0 0 1 1
use contact_14  contact_14_94
timestamp 1644969367
transform 1 0 13124 0 1 48
box 0 0 1 1
use contact_14  contact_14_95
timestamp 1644969367
transform 1 0 12514 0 1 128
box 0 0 1 1
use contact_14  contact_14_96
timestamp 1644969367
transform 1 0 12346 0 1 48
box 0 0 1 1
use contact_14  contact_14_97
timestamp 1644969367
transform 1 0 11736 0 1 128
box 0 0 1 1
use contact_14  contact_14_98
timestamp 1644969367
transform 1 0 11568 0 1 48
box 0 0 1 1
use contact_14  contact_14_99
timestamp 1644969367
transform 1 0 10958 0 1 128
box 0 0 1 1
use contact_14  contact_14_100
timestamp 1644969367
transform 1 0 10790 0 1 48
box 0 0 1 1
use contact_14  contact_14_101
timestamp 1644969367
transform 1 0 10180 0 1 128
box 0 0 1 1
use contact_14  contact_14_102
timestamp 1644969367
transform 1 0 10012 0 1 48
box 0 0 1 1
use contact_14  contact_14_103
timestamp 1644969367
transform 1 0 9402 0 1 128
box 0 0 1 1
use contact_14  contact_14_104
timestamp 1644969367
transform 1 0 9234 0 1 48
box 0 0 1 1
use contact_14  contact_14_105
timestamp 1644969367
transform 1 0 8624 0 1 128
box 0 0 1 1
use contact_14  contact_14_106
timestamp 1644969367
transform 1 0 8456 0 1 48
box 0 0 1 1
use contact_14  contact_14_107
timestamp 1644969367
transform 1 0 7846 0 1 128
box 0 0 1 1
use contact_14  contact_14_108
timestamp 1644969367
transform 1 0 7678 0 1 48
box 0 0 1 1
use contact_14  contact_14_109
timestamp 1644969367
transform 1 0 7068 0 1 128
box 0 0 1 1
use contact_14  contact_14_110
timestamp 1644969367
transform 1 0 6900 0 1 48
box 0 0 1 1
use contact_14  contact_14_111
timestamp 1644969367
transform 1 0 6290 0 1 128
box 0 0 1 1
use contact_14  contact_14_112
timestamp 1644969367
transform 1 0 6122 0 1 48
box 0 0 1 1
use contact_14  contact_14_113
timestamp 1644969367
transform 1 0 5512 0 1 128
box 0 0 1 1
use contact_14  contact_14_114
timestamp 1644969367
transform 1 0 5344 0 1 48
box 0 0 1 1
use contact_14  contact_14_115
timestamp 1644969367
transform 1 0 4734 0 1 128
box 0 0 1 1
use contact_14  contact_14_116
timestamp 1644969367
transform 1 0 4566 0 1 48
box 0 0 1 1
use contact_14  contact_14_117
timestamp 1644969367
transform 1 0 3956 0 1 128
box 0 0 1 1
use contact_14  contact_14_118
timestamp 1644969367
transform 1 0 3788 0 1 48
box 0 0 1 1
use contact_14  contact_14_119
timestamp 1644969367
transform 1 0 3178 0 1 128
box 0 0 1 1
use contact_14  contact_14_120
timestamp 1644969367
transform 1 0 3010 0 1 48
box 0 0 1 1
use contact_14  contact_14_121
timestamp 1644969367
transform 1 0 2400 0 1 128
box 0 0 1 1
use contact_14  contact_14_122
timestamp 1644969367
transform 1 0 2232 0 1 48
box 0 0 1 1
use contact_14  contact_14_123
timestamp 1644969367
transform 1 0 1622 0 1 128
box 0 0 1 1
use contact_14  contact_14_124
timestamp 1644969367
transform 1 0 1454 0 1 48
box 0 0 1 1
use contact_14  contact_14_125
timestamp 1644969367
transform 1 0 844 0 1 128
box 0 0 1 1
use contact_14  contact_14_126
timestamp 1644969367
transform 1 0 676 0 1 48
box 0 0 1 1
use contact_14  contact_14_127
timestamp 1644969367
transform 1 0 66 0 1 128
box 0 0 1 1
use contact_27  contact_27_0
timestamp 1644969367
transform 1 0 49374 0 1 311
box 0 0 1 1
use contact_26  contact_26_0
timestamp 1644969367
transform 1 0 49370 0 1 301
box 0 0 1 1
use contact_27  contact_27_1
timestamp 1644969367
transform 1 0 48596 0 1 231
box 0 0 1 1
use contact_26  contact_26_1
timestamp 1644969367
transform 1 0 48592 0 1 221
box 0 0 1 1
use contact_27  contact_27_2
timestamp 1644969367
transform 1 0 47818 0 1 311
box 0 0 1 1
use contact_26  contact_26_2
timestamp 1644969367
transform 1 0 47814 0 1 301
box 0 0 1 1
use contact_27  contact_27_3
timestamp 1644969367
transform 1 0 47040 0 1 231
box 0 0 1 1
use contact_26  contact_26_3
timestamp 1644969367
transform 1 0 47036 0 1 221
box 0 0 1 1
use contact_27  contact_27_4
timestamp 1644969367
transform 1 0 46262 0 1 311
box 0 0 1 1
use contact_26  contact_26_4
timestamp 1644969367
transform 1 0 46258 0 1 301
box 0 0 1 1
use contact_27  contact_27_5
timestamp 1644969367
transform 1 0 45484 0 1 231
box 0 0 1 1
use contact_26  contact_26_5
timestamp 1644969367
transform 1 0 45480 0 1 221
box 0 0 1 1
use contact_27  contact_27_6
timestamp 1644969367
transform 1 0 44706 0 1 311
box 0 0 1 1
use contact_26  contact_26_6
timestamp 1644969367
transform 1 0 44702 0 1 301
box 0 0 1 1
use contact_27  contact_27_7
timestamp 1644969367
transform 1 0 43928 0 1 231
box 0 0 1 1
use contact_26  contact_26_7
timestamp 1644969367
transform 1 0 43924 0 1 221
box 0 0 1 1
use contact_27  contact_27_8
timestamp 1644969367
transform 1 0 43150 0 1 311
box 0 0 1 1
use contact_26  contact_26_8
timestamp 1644969367
transform 1 0 43146 0 1 301
box 0 0 1 1
use contact_27  contact_27_9
timestamp 1644969367
transform 1 0 42372 0 1 231
box 0 0 1 1
use contact_26  contact_26_9
timestamp 1644969367
transform 1 0 42368 0 1 221
box 0 0 1 1
use contact_27  contact_27_10
timestamp 1644969367
transform 1 0 41594 0 1 311
box 0 0 1 1
use contact_26  contact_26_10
timestamp 1644969367
transform 1 0 41590 0 1 301
box 0 0 1 1
use contact_27  contact_27_11
timestamp 1644969367
transform 1 0 40816 0 1 231
box 0 0 1 1
use contact_26  contact_26_11
timestamp 1644969367
transform 1 0 40812 0 1 221
box 0 0 1 1
use contact_27  contact_27_12
timestamp 1644969367
transform 1 0 40038 0 1 311
box 0 0 1 1
use contact_26  contact_26_12
timestamp 1644969367
transform 1 0 40034 0 1 301
box 0 0 1 1
use contact_27  contact_27_13
timestamp 1644969367
transform 1 0 39260 0 1 231
box 0 0 1 1
use contact_26  contact_26_13
timestamp 1644969367
transform 1 0 39256 0 1 221
box 0 0 1 1
use contact_27  contact_27_14
timestamp 1644969367
transform 1 0 38482 0 1 311
box 0 0 1 1
use contact_26  contact_26_14
timestamp 1644969367
transform 1 0 38478 0 1 301
box 0 0 1 1
use contact_27  contact_27_15
timestamp 1644969367
transform 1 0 37704 0 1 231
box 0 0 1 1
use contact_26  contact_26_15
timestamp 1644969367
transform 1 0 37700 0 1 221
box 0 0 1 1
use contact_27  contact_27_16
timestamp 1644969367
transform 1 0 36926 0 1 311
box 0 0 1 1
use contact_26  contact_26_16
timestamp 1644969367
transform 1 0 36922 0 1 301
box 0 0 1 1
use contact_27  contact_27_17
timestamp 1644969367
transform 1 0 36148 0 1 231
box 0 0 1 1
use contact_26  contact_26_17
timestamp 1644969367
transform 1 0 36144 0 1 221
box 0 0 1 1
use contact_27  contact_27_18
timestamp 1644969367
transform 1 0 35370 0 1 311
box 0 0 1 1
use contact_26  contact_26_18
timestamp 1644969367
transform 1 0 35366 0 1 301
box 0 0 1 1
use contact_27  contact_27_19
timestamp 1644969367
transform 1 0 34592 0 1 231
box 0 0 1 1
use contact_26  contact_26_19
timestamp 1644969367
transform 1 0 34588 0 1 221
box 0 0 1 1
use contact_27  contact_27_20
timestamp 1644969367
transform 1 0 33814 0 1 311
box 0 0 1 1
use contact_26  contact_26_20
timestamp 1644969367
transform 1 0 33810 0 1 301
box 0 0 1 1
use contact_27  contact_27_21
timestamp 1644969367
transform 1 0 33036 0 1 231
box 0 0 1 1
use contact_26  contact_26_21
timestamp 1644969367
transform 1 0 33032 0 1 221
box 0 0 1 1
use contact_27  contact_27_22
timestamp 1644969367
transform 1 0 32258 0 1 311
box 0 0 1 1
use contact_26  contact_26_22
timestamp 1644969367
transform 1 0 32254 0 1 301
box 0 0 1 1
use contact_27  contact_27_23
timestamp 1644969367
transform 1 0 31480 0 1 231
box 0 0 1 1
use contact_26  contact_26_23
timestamp 1644969367
transform 1 0 31476 0 1 221
box 0 0 1 1
use contact_27  contact_27_24
timestamp 1644969367
transform 1 0 30702 0 1 311
box 0 0 1 1
use contact_26  contact_26_24
timestamp 1644969367
transform 1 0 30698 0 1 301
box 0 0 1 1
use contact_27  contact_27_25
timestamp 1644969367
transform 1 0 29924 0 1 231
box 0 0 1 1
use contact_26  contact_26_25
timestamp 1644969367
transform 1 0 29920 0 1 221
box 0 0 1 1
use contact_27  contact_27_26
timestamp 1644969367
transform 1 0 29146 0 1 311
box 0 0 1 1
use contact_26  contact_26_26
timestamp 1644969367
transform 1 0 29142 0 1 301
box 0 0 1 1
use contact_27  contact_27_27
timestamp 1644969367
transform 1 0 28368 0 1 231
box 0 0 1 1
use contact_26  contact_26_27
timestamp 1644969367
transform 1 0 28364 0 1 221
box 0 0 1 1
use contact_27  contact_27_28
timestamp 1644969367
transform 1 0 27590 0 1 311
box 0 0 1 1
use contact_26  contact_26_28
timestamp 1644969367
transform 1 0 27586 0 1 301
box 0 0 1 1
use contact_27  contact_27_29
timestamp 1644969367
transform 1 0 26812 0 1 231
box 0 0 1 1
use contact_26  contact_26_29
timestamp 1644969367
transform 1 0 26808 0 1 221
box 0 0 1 1
use contact_27  contact_27_30
timestamp 1644969367
transform 1 0 26034 0 1 311
box 0 0 1 1
use contact_26  contact_26_30
timestamp 1644969367
transform 1 0 26030 0 1 301
box 0 0 1 1
use contact_27  contact_27_31
timestamp 1644969367
transform 1 0 25256 0 1 231
box 0 0 1 1
use contact_26  contact_26_31
timestamp 1644969367
transform 1 0 25252 0 1 221
box 0 0 1 1
use contact_27  contact_27_32
timestamp 1644969367
transform 1 0 24478 0 1 311
box 0 0 1 1
use contact_26  contact_26_32
timestamp 1644969367
transform 1 0 24474 0 1 301
box 0 0 1 1
use contact_27  contact_27_33
timestamp 1644969367
transform 1 0 23700 0 1 231
box 0 0 1 1
use contact_26  contact_26_33
timestamp 1644969367
transform 1 0 23696 0 1 221
box 0 0 1 1
use contact_27  contact_27_34
timestamp 1644969367
transform 1 0 22922 0 1 311
box 0 0 1 1
use contact_26  contact_26_34
timestamp 1644969367
transform 1 0 22918 0 1 301
box 0 0 1 1
use contact_27  contact_27_35
timestamp 1644969367
transform 1 0 22144 0 1 231
box 0 0 1 1
use contact_26  contact_26_35
timestamp 1644969367
transform 1 0 22140 0 1 221
box 0 0 1 1
use contact_27  contact_27_36
timestamp 1644969367
transform 1 0 21366 0 1 311
box 0 0 1 1
use contact_26  contact_26_36
timestamp 1644969367
transform 1 0 21362 0 1 301
box 0 0 1 1
use contact_27  contact_27_37
timestamp 1644969367
transform 1 0 20588 0 1 231
box 0 0 1 1
use contact_26  contact_26_37
timestamp 1644969367
transform 1 0 20584 0 1 221
box 0 0 1 1
use contact_27  contact_27_38
timestamp 1644969367
transform 1 0 19810 0 1 311
box 0 0 1 1
use contact_26  contact_26_38
timestamp 1644969367
transform 1 0 19806 0 1 301
box 0 0 1 1
use contact_27  contact_27_39
timestamp 1644969367
transform 1 0 19032 0 1 231
box 0 0 1 1
use contact_26  contact_26_39
timestamp 1644969367
transform 1 0 19028 0 1 221
box 0 0 1 1
use contact_27  contact_27_40
timestamp 1644969367
transform 1 0 18254 0 1 311
box 0 0 1 1
use contact_26  contact_26_40
timestamp 1644969367
transform 1 0 18250 0 1 301
box 0 0 1 1
use contact_27  contact_27_41
timestamp 1644969367
transform 1 0 17476 0 1 231
box 0 0 1 1
use contact_26  contact_26_41
timestamp 1644969367
transform 1 0 17472 0 1 221
box 0 0 1 1
use contact_27  contact_27_42
timestamp 1644969367
transform 1 0 16698 0 1 311
box 0 0 1 1
use contact_26  contact_26_42
timestamp 1644969367
transform 1 0 16694 0 1 301
box 0 0 1 1
use contact_27  contact_27_43
timestamp 1644969367
transform 1 0 15920 0 1 231
box 0 0 1 1
use contact_26  contact_26_43
timestamp 1644969367
transform 1 0 15916 0 1 221
box 0 0 1 1
use contact_27  contact_27_44
timestamp 1644969367
transform 1 0 15142 0 1 311
box 0 0 1 1
use contact_26  contact_26_44
timestamp 1644969367
transform 1 0 15138 0 1 301
box 0 0 1 1
use contact_27  contact_27_45
timestamp 1644969367
transform 1 0 14364 0 1 231
box 0 0 1 1
use contact_26  contact_26_45
timestamp 1644969367
transform 1 0 14360 0 1 221
box 0 0 1 1
use contact_27  contact_27_46
timestamp 1644969367
transform 1 0 13586 0 1 311
box 0 0 1 1
use contact_26  contact_26_46
timestamp 1644969367
transform 1 0 13582 0 1 301
box 0 0 1 1
use contact_27  contact_27_47
timestamp 1644969367
transform 1 0 12808 0 1 231
box 0 0 1 1
use contact_26  contact_26_47
timestamp 1644969367
transform 1 0 12804 0 1 221
box 0 0 1 1
use contact_27  contact_27_48
timestamp 1644969367
transform 1 0 12030 0 1 311
box 0 0 1 1
use contact_26  contact_26_48
timestamp 1644969367
transform 1 0 12026 0 1 301
box 0 0 1 1
use contact_27  contact_27_49
timestamp 1644969367
transform 1 0 11252 0 1 231
box 0 0 1 1
use contact_26  contact_26_49
timestamp 1644969367
transform 1 0 11248 0 1 221
box 0 0 1 1
use contact_27  contact_27_50
timestamp 1644969367
transform 1 0 10474 0 1 311
box 0 0 1 1
use contact_26  contact_26_50
timestamp 1644969367
transform 1 0 10470 0 1 301
box 0 0 1 1
use contact_27  contact_27_51
timestamp 1644969367
transform 1 0 9696 0 1 231
box 0 0 1 1
use contact_26  contact_26_51
timestamp 1644969367
transform 1 0 9692 0 1 221
box 0 0 1 1
use contact_27  contact_27_52
timestamp 1644969367
transform 1 0 8918 0 1 311
box 0 0 1 1
use contact_26  contact_26_52
timestamp 1644969367
transform 1 0 8914 0 1 301
box 0 0 1 1
use contact_27  contact_27_53
timestamp 1644969367
transform 1 0 8140 0 1 231
box 0 0 1 1
use contact_26  contact_26_53
timestamp 1644969367
transform 1 0 8136 0 1 221
box 0 0 1 1
use contact_27  contact_27_54
timestamp 1644969367
transform 1 0 7362 0 1 311
box 0 0 1 1
use contact_26  contact_26_54
timestamp 1644969367
transform 1 0 7358 0 1 301
box 0 0 1 1
use contact_27  contact_27_55
timestamp 1644969367
transform 1 0 6584 0 1 231
box 0 0 1 1
use contact_26  contact_26_55
timestamp 1644969367
transform 1 0 6580 0 1 221
box 0 0 1 1
use contact_27  contact_27_56
timestamp 1644969367
transform 1 0 5806 0 1 311
box 0 0 1 1
use contact_26  contact_26_56
timestamp 1644969367
transform 1 0 5802 0 1 301
box 0 0 1 1
use contact_27  contact_27_57
timestamp 1644969367
transform 1 0 5028 0 1 231
box 0 0 1 1
use contact_26  contact_26_57
timestamp 1644969367
transform 1 0 5024 0 1 221
box 0 0 1 1
use contact_27  contact_27_58
timestamp 1644969367
transform 1 0 4250 0 1 311
box 0 0 1 1
use contact_26  contact_26_58
timestamp 1644969367
transform 1 0 4246 0 1 301
box 0 0 1 1
use contact_27  contact_27_59
timestamp 1644969367
transform 1 0 3472 0 1 231
box 0 0 1 1
use contact_26  contact_26_59
timestamp 1644969367
transform 1 0 3468 0 1 221
box 0 0 1 1
use contact_27  contact_27_60
timestamp 1644969367
transform 1 0 2694 0 1 311
box 0 0 1 1
use contact_26  contact_26_60
timestamp 1644969367
transform 1 0 2690 0 1 301
box 0 0 1 1
use contact_27  contact_27_61
timestamp 1644969367
transform 1 0 1916 0 1 231
box 0 0 1 1
use contact_26  contact_26_61
timestamp 1644969367
transform 1 0 1912 0 1 221
box 0 0 1 1
use contact_27  contact_27_62
timestamp 1644969367
transform 1 0 1138 0 1 311
box 0 0 1 1
use contact_26  contact_26_62
timestamp 1644969367
transform 1 0 1134 0 1 301
box 0 0 1 1
use contact_27  contact_27_63
timestamp 1644969367
transform 1 0 360 0 1 231
box 0 0 1 1
use contact_26  contact_26_63
timestamp 1644969367
transform 1 0 356 0 1 221
box 0 0 1 1
use column_mux_multiport  column_mux_multiport_0
timestamp 1644969367
transform 1 0 49014 0 1 400
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_1
timestamp 1644969367
transform 1 0 48236 0 1 400
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_2
timestamp 1644969367
transform 1 0 47458 0 1 400
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_3
timestamp 1644969367
transform 1 0 46680 0 1 400
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_4
timestamp 1644969367
transform 1 0 45902 0 1 400
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_5
timestamp 1644969367
transform 1 0 45124 0 1 400
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_6
timestamp 1644969367
transform 1 0 44346 0 1 400
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_7
timestamp 1644969367
transform 1 0 43568 0 1 400
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_8
timestamp 1644969367
transform 1 0 42790 0 1 400
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_9
timestamp 1644969367
transform 1 0 42012 0 1 400
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_10
timestamp 1644969367
transform 1 0 41234 0 1 400
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_11
timestamp 1644969367
transform 1 0 40456 0 1 400
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_12
timestamp 1644969367
transform 1 0 39678 0 1 400
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_13
timestamp 1644969367
transform 1 0 38900 0 1 400
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_14
timestamp 1644969367
transform 1 0 38122 0 1 400
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_15
timestamp 1644969367
transform 1 0 37344 0 1 400
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_16
timestamp 1644969367
transform 1 0 36566 0 1 400
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_17
timestamp 1644969367
transform 1 0 35788 0 1 400
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_18
timestamp 1644969367
transform 1 0 35010 0 1 400
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_19
timestamp 1644969367
transform 1 0 34232 0 1 400
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_20
timestamp 1644969367
transform 1 0 33454 0 1 400
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_21
timestamp 1644969367
transform 1 0 32676 0 1 400
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_22
timestamp 1644969367
transform 1 0 31898 0 1 400
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_23
timestamp 1644969367
transform 1 0 31120 0 1 400
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_24
timestamp 1644969367
transform 1 0 30342 0 1 400
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_25
timestamp 1644969367
transform 1 0 29564 0 1 400
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_26
timestamp 1644969367
transform 1 0 28786 0 1 400
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_27
timestamp 1644969367
transform 1 0 28008 0 1 400
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_28
timestamp 1644969367
transform 1 0 27230 0 1 400
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_29
timestamp 1644969367
transform 1 0 26452 0 1 400
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_30
timestamp 1644969367
transform 1 0 25674 0 1 400
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_31
timestamp 1644969367
transform 1 0 24896 0 1 400
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_32
timestamp 1644969367
transform 1 0 24118 0 1 400
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_33
timestamp 1644969367
transform 1 0 23340 0 1 400
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_34
timestamp 1644969367
transform 1 0 22562 0 1 400
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_35
timestamp 1644969367
transform 1 0 21784 0 1 400
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_36
timestamp 1644969367
transform 1 0 21006 0 1 400
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_37
timestamp 1644969367
transform 1 0 20228 0 1 400
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_38
timestamp 1644969367
transform 1 0 19450 0 1 400
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_39
timestamp 1644969367
transform 1 0 18672 0 1 400
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_40
timestamp 1644969367
transform 1 0 17894 0 1 400
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_41
timestamp 1644969367
transform 1 0 17116 0 1 400
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_42
timestamp 1644969367
transform 1 0 16338 0 1 400
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_43
timestamp 1644969367
transform 1 0 15560 0 1 400
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_44
timestamp 1644969367
transform 1 0 14782 0 1 400
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_45
timestamp 1644969367
transform 1 0 14004 0 1 400
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_46
timestamp 1644969367
transform 1 0 13226 0 1 400
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_47
timestamp 1644969367
transform 1 0 12448 0 1 400
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_48
timestamp 1644969367
transform 1 0 11670 0 1 400
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_49
timestamp 1644969367
transform 1 0 10892 0 1 400
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_50
timestamp 1644969367
transform 1 0 10114 0 1 400
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_51
timestamp 1644969367
transform 1 0 9336 0 1 400
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_52
timestamp 1644969367
transform 1 0 8558 0 1 400
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_53
timestamp 1644969367
transform 1 0 7780 0 1 400
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_54
timestamp 1644969367
transform 1 0 7002 0 1 400
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_55
timestamp 1644969367
transform 1 0 6224 0 1 400
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_56
timestamp 1644969367
transform 1 0 5446 0 1 400
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_57
timestamp 1644969367
transform 1 0 4668 0 1 400
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_58
timestamp 1644969367
transform 1 0 3890 0 1 400
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_59
timestamp 1644969367
transform 1 0 3112 0 1 400
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_60
timestamp 1644969367
transform 1 0 2334 0 1 400
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_61
timestamp 1644969367
transform 1 0 1556 0 1 400
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_62
timestamp 1644969367
transform 1 0 778 0 1 400
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_63
timestamp 1644969367
transform 1 0 0 0 1 400
box 49 0 844 1508
<< labels >>
rlabel metal1 s 0 240 49792 268 4 sel_0
rlabel metal1 s 0 320 49792 348 4 sel_1
rlabel metal2 s 84 160 112 400 4 rbl0_out_0
rlabel metal2 s 694 80 722 400 4 rbl1_out_0
rlabel metal2 s 1640 160 1668 400 4 rbl0_out_1
rlabel metal2 s 2250 80 2278 400 4 rbl1_out_1
rlabel metal2 s 3196 160 3224 400 4 rbl0_out_2
rlabel metal2 s 3806 80 3834 400 4 rbl1_out_2
rlabel metal2 s 4752 160 4780 400 4 rbl0_out_3
rlabel metal2 s 5362 80 5390 400 4 rbl1_out_3
rlabel metal2 s 6308 160 6336 400 4 rbl0_out_4
rlabel metal2 s 6918 80 6946 400 4 rbl1_out_4
rlabel metal2 s 7864 160 7892 400 4 rbl0_out_5
rlabel metal2 s 8474 80 8502 400 4 rbl1_out_5
rlabel metal2 s 9420 160 9448 400 4 rbl0_out_6
rlabel metal2 s 10030 80 10058 400 4 rbl1_out_6
rlabel metal2 s 10976 160 11004 400 4 rbl0_out_7
rlabel metal2 s 11586 80 11614 400 4 rbl1_out_7
rlabel metal2 s 12532 160 12560 400 4 rbl0_out_8
rlabel metal2 s 13142 80 13170 400 4 rbl1_out_8
rlabel metal2 s 14088 160 14116 400 4 rbl0_out_9
rlabel metal2 s 14698 80 14726 400 4 rbl1_out_9
rlabel metal2 s 15644 160 15672 400 4 rbl0_out_10
rlabel metal2 s 16254 80 16282 400 4 rbl1_out_10
rlabel metal2 s 17200 160 17228 400 4 rbl0_out_11
rlabel metal2 s 17810 80 17838 400 4 rbl1_out_11
rlabel metal2 s 18756 160 18784 400 4 rbl0_out_12
rlabel metal2 s 19366 80 19394 400 4 rbl1_out_12
rlabel metal2 s 20312 160 20340 400 4 rbl0_out_13
rlabel metal2 s 20922 80 20950 400 4 rbl1_out_13
rlabel metal2 s 21868 160 21896 400 4 rbl0_out_14
rlabel metal2 s 22478 80 22506 400 4 rbl1_out_14
rlabel metal2 s 23424 160 23452 400 4 rbl0_out_15
rlabel metal2 s 24034 80 24062 400 4 rbl1_out_15
rlabel metal2 s 24980 160 25008 400 4 rbl0_out_16
rlabel metal2 s 25590 80 25618 400 4 rbl1_out_16
rlabel metal2 s 26536 160 26564 400 4 rbl0_out_17
rlabel metal2 s 27146 80 27174 400 4 rbl1_out_17
rlabel metal2 s 28092 160 28120 400 4 rbl0_out_18
rlabel metal2 s 28702 80 28730 400 4 rbl1_out_18
rlabel metal2 s 29648 160 29676 400 4 rbl0_out_19
rlabel metal2 s 30258 80 30286 400 4 rbl1_out_19
rlabel metal2 s 31204 160 31232 400 4 rbl0_out_20
rlabel metal2 s 31814 80 31842 400 4 rbl1_out_20
rlabel metal2 s 32760 160 32788 400 4 rbl0_out_21
rlabel metal2 s 33370 80 33398 400 4 rbl1_out_21
rlabel metal2 s 34316 160 34344 400 4 rbl0_out_22
rlabel metal2 s 34926 80 34954 400 4 rbl1_out_22
rlabel metal2 s 35872 160 35900 400 4 rbl0_out_23
rlabel metal2 s 36482 80 36510 400 4 rbl1_out_23
rlabel metal2 s 37428 160 37456 400 4 rbl0_out_24
rlabel metal2 s 38038 80 38066 400 4 rbl1_out_24
rlabel metal2 s 38984 160 39012 400 4 rbl0_out_25
rlabel metal2 s 39594 80 39622 400 4 rbl1_out_25
rlabel metal2 s 40540 160 40568 400 4 rbl0_out_26
rlabel metal2 s 41150 80 41178 400 4 rbl1_out_26
rlabel metal2 s 42096 160 42124 400 4 rbl0_out_27
rlabel metal2 s 42706 80 42734 400 4 rbl1_out_27
rlabel metal2 s 43652 160 43680 400 4 rbl0_out_28
rlabel metal2 s 44262 80 44290 400 4 rbl1_out_28
rlabel metal2 s 45208 160 45236 400 4 rbl0_out_29
rlabel metal2 s 45818 80 45846 400 4 rbl1_out_29
rlabel metal2 s 46764 160 46792 400 4 rbl0_out_30
rlabel metal2 s 47374 80 47402 400 4 rbl1_out_30
rlabel metal2 s 48320 160 48348 400 4 rbl0_out_31
rlabel metal2 s 48930 80 48958 400 4 rbl1_out_31
rlabel metal2 s 84 1852 112 1908 4 rbl0_0
rlabel metal2 s 694 1852 722 1908 4 rbl1_0
rlabel metal2 s 862 1852 890 1908 4 rbl0_1
rlabel metal2 s 1472 1852 1500 1908 4 rbl1_1
rlabel metal2 s 1640 1852 1668 1908 4 rbl0_2
rlabel metal2 s 2250 1852 2278 1908 4 rbl1_2
rlabel metal2 s 2418 1852 2446 1908 4 rbl0_3
rlabel metal2 s 3028 1852 3056 1908 4 rbl1_3
rlabel metal2 s 3196 1852 3224 1908 4 rbl0_4
rlabel metal2 s 3806 1852 3834 1908 4 rbl1_4
rlabel metal2 s 3974 1852 4002 1908 4 rbl0_5
rlabel metal2 s 4584 1852 4612 1908 4 rbl1_5
rlabel metal2 s 4752 1852 4780 1908 4 rbl0_6
rlabel metal2 s 5362 1852 5390 1908 4 rbl1_6
rlabel metal2 s 5530 1852 5558 1908 4 rbl0_7
rlabel metal2 s 6140 1852 6168 1908 4 rbl1_7
rlabel metal2 s 6308 1852 6336 1908 4 rbl0_8
rlabel metal2 s 6918 1852 6946 1908 4 rbl1_8
rlabel metal2 s 7086 1852 7114 1908 4 rbl0_9
rlabel metal2 s 7696 1852 7724 1908 4 rbl1_9
rlabel metal2 s 7864 1852 7892 1908 4 rbl0_10
rlabel metal2 s 8474 1852 8502 1908 4 rbl1_10
rlabel metal2 s 8642 1852 8670 1908 4 rbl0_11
rlabel metal2 s 9252 1852 9280 1908 4 rbl1_11
rlabel metal2 s 9420 1852 9448 1908 4 rbl0_12
rlabel metal2 s 10030 1852 10058 1908 4 rbl1_12
rlabel metal2 s 10198 1852 10226 1908 4 rbl0_13
rlabel metal2 s 10808 1852 10836 1908 4 rbl1_13
rlabel metal2 s 10976 1852 11004 1908 4 rbl0_14
rlabel metal2 s 11586 1852 11614 1908 4 rbl1_14
rlabel metal2 s 11754 1852 11782 1908 4 rbl0_15
rlabel metal2 s 12364 1852 12392 1908 4 rbl1_15
rlabel metal2 s 12532 1852 12560 1908 4 rbl0_16
rlabel metal2 s 13142 1852 13170 1908 4 rbl1_16
rlabel metal2 s 13310 1852 13338 1908 4 rbl0_17
rlabel metal2 s 13920 1852 13948 1908 4 rbl1_17
rlabel metal2 s 14088 1852 14116 1908 4 rbl0_18
rlabel metal2 s 14698 1852 14726 1908 4 rbl1_18
rlabel metal2 s 14866 1852 14894 1908 4 rbl0_19
rlabel metal2 s 15476 1852 15504 1908 4 rbl1_19
rlabel metal2 s 15644 1852 15672 1908 4 rbl0_20
rlabel metal2 s 16254 1852 16282 1908 4 rbl1_20
rlabel metal2 s 16422 1852 16450 1908 4 rbl0_21
rlabel metal2 s 17032 1852 17060 1908 4 rbl1_21
rlabel metal2 s 17200 1852 17228 1908 4 rbl0_22
rlabel metal2 s 17810 1852 17838 1908 4 rbl1_22
rlabel metal2 s 17978 1852 18006 1908 4 rbl0_23
rlabel metal2 s 18588 1852 18616 1908 4 rbl1_23
rlabel metal2 s 18756 1852 18784 1908 4 rbl0_24
rlabel metal2 s 19366 1852 19394 1908 4 rbl1_24
rlabel metal2 s 19534 1852 19562 1908 4 rbl0_25
rlabel metal2 s 20144 1852 20172 1908 4 rbl1_25
rlabel metal2 s 20312 1852 20340 1908 4 rbl0_26
rlabel metal2 s 20922 1852 20950 1908 4 rbl1_26
rlabel metal2 s 21090 1852 21118 1908 4 rbl0_27
rlabel metal2 s 21700 1852 21728 1908 4 rbl1_27
rlabel metal2 s 21868 1852 21896 1908 4 rbl0_28
rlabel metal2 s 22478 1852 22506 1908 4 rbl1_28
rlabel metal2 s 22646 1852 22674 1908 4 rbl0_29
rlabel metal2 s 23256 1852 23284 1908 4 rbl1_29
rlabel metal2 s 23424 1852 23452 1908 4 rbl0_30
rlabel metal2 s 24034 1852 24062 1908 4 rbl1_30
rlabel metal2 s 24202 1852 24230 1908 4 rbl0_31
rlabel metal2 s 24812 1852 24840 1908 4 rbl1_31
rlabel metal2 s 24980 1852 25008 1908 4 rbl0_32
rlabel metal2 s 25590 1852 25618 1908 4 rbl1_32
rlabel metal2 s 25758 1852 25786 1908 4 rbl0_33
rlabel metal2 s 26368 1852 26396 1908 4 rbl1_33
rlabel metal2 s 26536 1852 26564 1908 4 rbl0_34
rlabel metal2 s 27146 1852 27174 1908 4 rbl1_34
rlabel metal2 s 27314 1852 27342 1908 4 rbl0_35
rlabel metal2 s 27924 1852 27952 1908 4 rbl1_35
rlabel metal2 s 28092 1852 28120 1908 4 rbl0_36
rlabel metal2 s 28702 1852 28730 1908 4 rbl1_36
rlabel metal2 s 28870 1852 28898 1908 4 rbl0_37
rlabel metal2 s 29480 1852 29508 1908 4 rbl1_37
rlabel metal2 s 29648 1852 29676 1908 4 rbl0_38
rlabel metal2 s 30258 1852 30286 1908 4 rbl1_38
rlabel metal2 s 30426 1852 30454 1908 4 rbl0_39
rlabel metal2 s 31036 1852 31064 1908 4 rbl1_39
rlabel metal2 s 31204 1852 31232 1908 4 rbl0_40
rlabel metal2 s 31814 1852 31842 1908 4 rbl1_40
rlabel metal2 s 31982 1852 32010 1908 4 rbl0_41
rlabel metal2 s 32592 1852 32620 1908 4 rbl1_41
rlabel metal2 s 32760 1852 32788 1908 4 rbl0_42
rlabel metal2 s 33370 1852 33398 1908 4 rbl1_42
rlabel metal2 s 33538 1852 33566 1908 4 rbl0_43
rlabel metal2 s 34148 1852 34176 1908 4 rbl1_43
rlabel metal2 s 34316 1852 34344 1908 4 rbl0_44
rlabel metal2 s 34926 1852 34954 1908 4 rbl1_44
rlabel metal2 s 35094 1852 35122 1908 4 rbl0_45
rlabel metal2 s 35704 1852 35732 1908 4 rbl1_45
rlabel metal2 s 35872 1852 35900 1908 4 rbl0_46
rlabel metal2 s 36482 1852 36510 1908 4 rbl1_46
rlabel metal2 s 36650 1852 36678 1908 4 rbl0_47
rlabel metal2 s 37260 1852 37288 1908 4 rbl1_47
rlabel metal2 s 37428 1852 37456 1908 4 rbl0_48
rlabel metal2 s 38038 1852 38066 1908 4 rbl1_48
rlabel metal2 s 38206 1852 38234 1908 4 rbl0_49
rlabel metal2 s 38816 1852 38844 1908 4 rbl1_49
rlabel metal2 s 38984 1852 39012 1908 4 rbl0_50
rlabel metal2 s 39594 1852 39622 1908 4 rbl1_50
rlabel metal2 s 39762 1852 39790 1908 4 rbl0_51
rlabel metal2 s 40372 1852 40400 1908 4 rbl1_51
rlabel metal2 s 40540 1852 40568 1908 4 rbl0_52
rlabel metal2 s 41150 1852 41178 1908 4 rbl1_52
rlabel metal2 s 41318 1852 41346 1908 4 rbl0_53
rlabel metal2 s 41928 1852 41956 1908 4 rbl1_53
rlabel metal2 s 42096 1852 42124 1908 4 rbl0_54
rlabel metal2 s 42706 1852 42734 1908 4 rbl1_54
rlabel metal2 s 42874 1852 42902 1908 4 rbl0_55
rlabel metal2 s 43484 1852 43512 1908 4 rbl1_55
rlabel metal2 s 43652 1852 43680 1908 4 rbl0_56
rlabel metal2 s 44262 1852 44290 1908 4 rbl1_56
rlabel metal2 s 44430 1852 44458 1908 4 rbl0_57
rlabel metal2 s 45040 1852 45068 1908 4 rbl1_57
rlabel metal2 s 45208 1852 45236 1908 4 rbl0_58
rlabel metal2 s 45818 1852 45846 1908 4 rbl1_58
rlabel metal2 s 45986 1852 46014 1908 4 rbl0_59
rlabel metal2 s 46596 1852 46624 1908 4 rbl1_59
rlabel metal2 s 46764 1852 46792 1908 4 rbl0_60
rlabel metal2 s 47374 1852 47402 1908 4 rbl1_60
rlabel metal2 s 47542 1852 47570 1908 4 rbl0_61
rlabel metal2 s 48152 1852 48180 1908 4 rbl1_61
rlabel metal2 s 48320 1852 48348 1908 4 rbl0_62
rlabel metal2 s 48930 1852 48958 1908 4 rbl1_62
rlabel metal2 s 49098 1852 49126 1908 4 rbl0_63
rlabel metal2 s 49708 1852 49736 1908 4 rbl1_63
rlabel metal3 s 44280 1122 44412 1196 4 gnd
rlabel metal3 s 31832 1122 31964 1196 4 gnd
rlabel metal3 s 17828 1122 17960 1196 4 gnd
rlabel metal3 s 10048 1122 10180 1196 4 gnd
rlabel metal3 s 13160 1122 13292 1196 4 gnd
rlabel metal3 s 41168 1122 41300 1196 4 gnd
rlabel metal3 s 24052 1122 24184 1196 4 gnd
rlabel metal3 s 35722 1122 35854 1196 4 gnd
rlabel metal3 s 49726 1122 49858 1196 4 gnd
rlabel metal3 s 22496 1122 22628 1196 4 gnd
rlabel metal3 s 41946 1122 42078 1196 4 gnd
rlabel metal3 s 47392 1122 47524 1196 4 gnd
rlabel metal3 s 13938 1122 14070 1196 4 gnd
rlabel metal3 s 5380 1122 5512 1196 4 gnd
rlabel metal3 s 8492 1122 8624 1196 4 gnd
rlabel metal3 s 27164 1122 27296 1196 4 gnd
rlabel metal3 s 48170 1122 48302 1196 4 gnd
rlabel metal3 s 21718 1122 21850 1196 4 gnd
rlabel metal3 s 43502 1122 43634 1196 4 gnd
rlabel metal3 s 46614 1122 46746 1196 4 gnd
rlabel metal3 s 6936 1122 7068 1196 4 gnd
rlabel metal3 s 6158 1122 6290 1196 4 gnd
rlabel metal3 s 1490 1122 1622 1196 4 gnd
rlabel metal3 s 24830 1122 24962 1196 4 gnd
rlabel metal3 s 31054 1122 31186 1196 4 gnd
rlabel metal3 s 39612 1122 39744 1196 4 gnd
rlabel metal3 s 9270 1122 9402 1196 4 gnd
rlabel metal3 s 26386 1122 26518 1196 4 gnd
rlabel metal3 s 19384 1122 19516 1196 4 gnd
rlabel metal3 s 40390 1122 40522 1196 4 gnd
rlabel metal3 s 25608 1122 25740 1196 4 gnd
rlabel metal3 s 27942 1122 28074 1196 4 gnd
rlabel metal3 s 23274 1122 23406 1196 4 gnd
rlabel metal3 s 38834 1122 38966 1196 4 gnd
rlabel metal3 s 4602 1122 4734 1196 4 gnd
rlabel metal3 s 11604 1122 11736 1196 4 gnd
rlabel metal3 s 34944 1122 35076 1196 4 gnd
rlabel metal3 s 28720 1122 28852 1196 4 gnd
rlabel metal3 s 33388 1122 33520 1196 4 gnd
rlabel metal3 s 30276 1122 30408 1196 4 gnd
rlabel metal3 s 712 1122 844 1196 4 gnd
rlabel metal3 s 3046 1122 3178 1196 4 gnd
rlabel metal3 s 36500 1122 36632 1196 4 gnd
rlabel metal3 s 3824 1122 3956 1196 4 gnd
rlabel metal3 s 34166 1122 34298 1196 4 gnd
rlabel metal3 s 37278 1122 37410 1196 4 gnd
rlabel metal3 s 32610 1122 32742 1196 4 gnd
rlabel metal3 s 14716 1122 14848 1196 4 gnd
rlabel metal3 s 45836 1122 45968 1196 4 gnd
rlabel metal3 s 2268 1122 2400 1196 4 gnd
rlabel metal3 s 20162 1122 20294 1196 4 gnd
rlabel metal3 s 18606 1122 18738 1196 4 gnd
rlabel metal3 s 7714 1122 7846 1196 4 gnd
rlabel metal3 s 48948 1122 49080 1196 4 gnd
rlabel metal3 s 15494 1122 15626 1196 4 gnd
rlabel metal3 s 16272 1122 16404 1196 4 gnd
rlabel metal3 s 17050 1122 17182 1196 4 gnd
rlabel metal3 s 38056 1122 38188 1196 4 gnd
rlabel metal3 s 42724 1122 42856 1196 4 gnd
rlabel metal3 s 10826 1122 10958 1196 4 gnd
rlabel metal3 s 45058 1122 45190 1196 4 gnd
rlabel metal3 s 12382 1122 12514 1196 4 gnd
rlabel metal3 s 20940 1122 21072 1196 4 gnd
rlabel metal3 s 29498 1122 29630 1196 4 gnd
<< properties >>
string FIXED_BBOX 0 0 49792 1908
string GDS_FILE sram_0rw2r1w_32_128_sky130A.gds
string GDS_END 2723038
string GDS_START 2648242
<< end >>
