magic
tech sky130A
magscale 1 2
timestamp 1643671299
<< checkpaint >>
rect -1260 -1284 26934 2264
<< metal1 >>
rect 0 -5 25674 23
<< metal2 >>
rect 54 0 82 990
rect 532 0 560 990
rect 832 0 860 990
rect 1310 0 1338 990
rect 1610 0 1638 990
rect 2088 0 2116 990
rect 2388 0 2416 990
rect 2866 0 2894 990
rect 3166 0 3194 990
rect 3644 0 3672 990
rect 3944 0 3972 990
rect 4422 0 4450 990
rect 4722 0 4750 990
rect 5200 0 5228 990
rect 5500 0 5528 990
rect 5978 0 6006 990
rect 6278 0 6306 990
rect 6756 0 6784 990
rect 7056 0 7084 990
rect 7534 0 7562 990
rect 7834 0 7862 990
rect 8312 0 8340 990
rect 8612 0 8640 990
rect 9090 0 9118 990
rect 9390 0 9418 990
rect 9868 0 9896 990
rect 10168 0 10196 990
rect 10646 0 10674 990
rect 10946 0 10974 990
rect 11424 0 11452 990
rect 11724 0 11752 990
rect 12202 0 12230 990
rect 12502 0 12530 990
rect 12980 0 13008 990
rect 13280 0 13308 990
rect 13758 0 13786 990
rect 14058 0 14086 990
rect 14536 0 14564 990
rect 14836 0 14864 990
rect 15314 0 15342 990
rect 15614 0 15642 990
rect 16092 0 16120 990
rect 16392 0 16420 990
rect 16870 0 16898 990
rect 17170 0 17198 990
rect 17648 0 17676 990
rect 17948 0 17976 990
rect 18426 0 18454 990
rect 18726 0 18754 990
rect 19204 0 19232 990
rect 19504 0 19532 990
rect 19982 0 20010 990
rect 20282 0 20310 990
rect 20760 0 20788 990
rect 21060 0 21088 990
rect 21538 0 21566 990
rect 21838 0 21866 990
rect 22316 0 22344 990
rect 22616 0 22644 990
rect 23094 0 23122 990
rect 23394 0 23422 990
rect 23872 0 23900 990
rect 24172 0 24200 990
rect 24650 0 24678 990
rect 24950 0 24978 990
rect 25428 0 25456 990
<< metal3 >>
rect 163 850 223 910
rect 941 850 1001 910
rect 1719 850 1779 910
rect 2497 850 2557 910
rect 3275 850 3335 910
rect 4053 850 4113 910
rect 4831 850 4891 910
rect 5609 850 5669 910
rect 6387 850 6447 910
rect 7165 850 7225 910
rect 7943 850 8003 910
rect 8721 850 8781 910
rect 9499 850 9559 910
rect 10277 850 10337 910
rect 11055 850 11115 910
rect 11833 850 11893 910
rect 12611 850 12671 910
rect 13389 850 13449 910
rect 14167 850 14227 910
rect 14945 850 15005 910
rect 15723 850 15783 910
rect 16501 850 16561 910
rect 17279 850 17339 910
rect 18057 850 18117 910
rect 18835 850 18895 910
rect 19613 850 19673 910
rect 20391 850 20451 910
rect 21169 850 21229 910
rect 21947 850 22007 910
rect 22725 850 22785 910
rect 23503 850 23563 910
rect 24281 850 24341 910
rect 25059 850 25119 910
use precharge_multiport_0  precharge_multiport_0_0
timestamp 1643671299
transform 1 0 24896 0 1 0
box 0 -24 778 1004
use precharge_multiport_0  precharge_multiport_0_1
timestamp 1643671299
transform 1 0 24118 0 1 0
box 0 -24 778 1004
use precharge_multiport_0  precharge_multiport_0_2
timestamp 1643671299
transform 1 0 23340 0 1 0
box 0 -24 778 1004
use precharge_multiport_0  precharge_multiport_0_3
timestamp 1643671299
transform 1 0 22562 0 1 0
box 0 -24 778 1004
use precharge_multiport_0  precharge_multiport_0_4
timestamp 1643671299
transform 1 0 21784 0 1 0
box 0 -24 778 1004
use precharge_multiport_0  precharge_multiport_0_5
timestamp 1643671299
transform 1 0 21006 0 1 0
box 0 -24 778 1004
use precharge_multiport_0  precharge_multiport_0_6
timestamp 1643671299
transform 1 0 20228 0 1 0
box 0 -24 778 1004
use precharge_multiport_0  precharge_multiport_0_7
timestamp 1643671299
transform 1 0 19450 0 1 0
box 0 -24 778 1004
use precharge_multiport_0  precharge_multiport_0_8
timestamp 1643671299
transform 1 0 18672 0 1 0
box 0 -24 778 1004
use precharge_multiport_0  precharge_multiport_0_9
timestamp 1643671299
transform 1 0 17894 0 1 0
box 0 -24 778 1004
use precharge_multiport_0  precharge_multiport_0_10
timestamp 1643671299
transform 1 0 17116 0 1 0
box 0 -24 778 1004
use precharge_multiport_0  precharge_multiport_0_11
timestamp 1643671299
transform 1 0 16338 0 1 0
box 0 -24 778 1004
use precharge_multiport_0  precharge_multiport_0_12
timestamp 1643671299
transform 1 0 15560 0 1 0
box 0 -24 778 1004
use precharge_multiport_0  precharge_multiport_0_13
timestamp 1643671299
transform 1 0 14782 0 1 0
box 0 -24 778 1004
use precharge_multiport_0  precharge_multiport_0_14
timestamp 1643671299
transform 1 0 14004 0 1 0
box 0 -24 778 1004
use precharge_multiport_0  precharge_multiport_0_15
timestamp 1643671299
transform 1 0 13226 0 1 0
box 0 -24 778 1004
use precharge_multiport_0  precharge_multiport_0_16
timestamp 1643671299
transform 1 0 12448 0 1 0
box 0 -24 778 1004
use precharge_multiport_0  precharge_multiport_0_17
timestamp 1643671299
transform 1 0 11670 0 1 0
box 0 -24 778 1004
use precharge_multiport_0  precharge_multiport_0_18
timestamp 1643671299
transform 1 0 10892 0 1 0
box 0 -24 778 1004
use precharge_multiport_0  precharge_multiport_0_19
timestamp 1643671299
transform 1 0 10114 0 1 0
box 0 -24 778 1004
use precharge_multiport_0  precharge_multiport_0_20
timestamp 1643671299
transform 1 0 9336 0 1 0
box 0 -24 778 1004
use precharge_multiport_0  precharge_multiport_0_21
timestamp 1643671299
transform 1 0 8558 0 1 0
box 0 -24 778 1004
use precharge_multiport_0  precharge_multiport_0_22
timestamp 1643671299
transform 1 0 7780 0 1 0
box 0 -24 778 1004
use precharge_multiport_0  precharge_multiport_0_23
timestamp 1643671299
transform 1 0 7002 0 1 0
box 0 -24 778 1004
use precharge_multiport_0  precharge_multiport_0_24
timestamp 1643671299
transform 1 0 6224 0 1 0
box 0 -24 778 1004
use precharge_multiport_0  precharge_multiport_0_25
timestamp 1643671299
transform 1 0 5446 0 1 0
box 0 -24 778 1004
use precharge_multiport_0  precharge_multiport_0_26
timestamp 1643671299
transform 1 0 4668 0 1 0
box 0 -24 778 1004
use precharge_multiport_0  precharge_multiport_0_27
timestamp 1643671299
transform 1 0 3890 0 1 0
box 0 -24 778 1004
use precharge_multiport_0  precharge_multiport_0_28
timestamp 1643671299
transform 1 0 3112 0 1 0
box 0 -24 778 1004
use precharge_multiport_0  precharge_multiport_0_29
timestamp 1643671299
transform 1 0 2334 0 1 0
box 0 -24 778 1004
use precharge_multiport_0  precharge_multiport_0_30
timestamp 1643671299
transform 1 0 1556 0 1 0
box 0 -24 778 1004
use precharge_multiport_0  precharge_multiport_0_31
timestamp 1643671299
transform 1 0 778 0 1 0
box 0 -24 778 1004
use precharge_multiport_0  precharge_multiport_0_32
timestamp 1643671299
transform 1 0 0 0 1 0
box 0 -24 778 1004
<< labels >>
rlabel metal1 s 0 -4 25674 22 4 en_bar
rlabel metal3 s 22724 850 22784 910 4 vdd
rlabel metal3 s 2496 850 2556 910 4 vdd
rlabel metal3 s 5608 850 5668 910 4 vdd
rlabel metal3 s 6386 850 6446 910 4 vdd
rlabel metal3 s 15722 850 15782 910 4 vdd
rlabel metal3 s 18834 850 18894 910 4 vdd
rlabel metal3 s 18056 850 18116 910 4 vdd
rlabel metal3 s 8720 850 8780 910 4 vdd
rlabel metal3 s 11832 850 11892 910 4 vdd
rlabel metal3 s 162 850 222 910 4 vdd
rlabel metal3 s 4052 850 4112 910 4 vdd
rlabel metal3 s 14944 850 15004 910 4 vdd
rlabel metal3 s 10276 850 10336 910 4 vdd
rlabel metal3 s 7164 850 7224 910 4 vdd
rlabel metal3 s 940 850 1000 910 4 vdd
rlabel metal3 s 12610 850 12670 910 4 vdd
rlabel metal3 s 17278 850 17338 910 4 vdd
rlabel metal3 s 16500 850 16560 910 4 vdd
rlabel metal3 s 24280 850 24340 910 4 vdd
rlabel metal3 s 21946 850 22006 910 4 vdd
rlabel metal3 s 23502 850 23562 910 4 vdd
rlabel metal3 s 11054 850 11114 910 4 vdd
rlabel metal3 s 4830 850 4890 910 4 vdd
rlabel metal3 s 7942 850 8002 910 4 vdd
rlabel metal3 s 13388 850 13448 910 4 vdd
rlabel metal3 s 21168 850 21228 910 4 vdd
rlabel metal3 s 20390 850 20450 910 4 vdd
rlabel metal3 s 3274 850 3334 910 4 vdd
rlabel metal3 s 19612 850 19672 910 4 vdd
rlabel metal3 s 9498 850 9558 910 4 vdd
rlabel metal3 s 25058 850 25118 910 4 vdd
rlabel metal3 s 1718 850 1778 910 4 vdd
rlabel metal3 s 14166 850 14226 910 4 vdd
rlabel metal2 s 54 0 82 990 4 rbl0_0
rlabel metal2 s 532 0 560 990 4 rbl1_0
rlabel metal2 s 832 0 860 990 4 rbl0_1
rlabel metal2 s 1310 0 1338 990 4 rbl1_1
rlabel metal2 s 1610 0 1638 990 4 rbl0_2
rlabel metal2 s 2088 0 2116 990 4 rbl1_2
rlabel metal2 s 2388 0 2416 990 4 rbl0_3
rlabel metal2 s 2866 0 2894 990 4 rbl1_3
rlabel metal2 s 3166 0 3194 990 4 rbl0_4
rlabel metal2 s 3644 0 3672 990 4 rbl1_4
rlabel metal2 s 3944 0 3972 990 4 rbl0_5
rlabel metal2 s 4422 0 4450 990 4 rbl1_5
rlabel metal2 s 4722 0 4750 990 4 rbl0_6
rlabel metal2 s 5200 0 5228 990 4 rbl1_6
rlabel metal2 s 5500 0 5528 990 4 rbl0_7
rlabel metal2 s 5978 0 6006 990 4 rbl1_7
rlabel metal2 s 6278 0 6306 990 4 rbl0_8
rlabel metal2 s 6756 0 6784 990 4 rbl1_8
rlabel metal2 s 7056 0 7084 990 4 rbl0_9
rlabel metal2 s 7534 0 7562 990 4 rbl1_9
rlabel metal2 s 7834 0 7862 990 4 rbl0_10
rlabel metal2 s 8312 0 8340 990 4 rbl1_10
rlabel metal2 s 8612 0 8640 990 4 rbl0_11
rlabel metal2 s 9090 0 9118 990 4 rbl1_11
rlabel metal2 s 9390 0 9418 990 4 rbl0_12
rlabel metal2 s 9868 0 9896 990 4 rbl1_12
rlabel metal2 s 10168 0 10196 990 4 rbl0_13
rlabel metal2 s 10646 0 10674 990 4 rbl1_13
rlabel metal2 s 10946 0 10974 990 4 rbl0_14
rlabel metal2 s 11424 0 11452 990 4 rbl1_14
rlabel metal2 s 11724 0 11752 990 4 rbl0_15
rlabel metal2 s 12202 0 12230 990 4 rbl1_15
rlabel metal2 s 12502 0 12530 990 4 rbl0_16
rlabel metal2 s 12980 0 13008 990 4 rbl1_16
rlabel metal2 s 13280 0 13308 990 4 rbl0_17
rlabel metal2 s 13758 0 13786 990 4 rbl1_17
rlabel metal2 s 14058 0 14086 990 4 rbl0_18
rlabel metal2 s 14536 0 14564 990 4 rbl1_18
rlabel metal2 s 14836 0 14864 990 4 rbl0_19
rlabel metal2 s 15314 0 15342 990 4 rbl1_19
rlabel metal2 s 15614 0 15642 990 4 rbl0_20
rlabel metal2 s 16092 0 16120 990 4 rbl1_20
rlabel metal2 s 16392 0 16420 990 4 rbl0_21
rlabel metal2 s 16870 0 16898 990 4 rbl1_21
rlabel metal2 s 17170 0 17198 990 4 rbl0_22
rlabel metal2 s 17648 0 17676 990 4 rbl1_22
rlabel metal2 s 17948 0 17976 990 4 rbl0_23
rlabel metal2 s 18426 0 18454 990 4 rbl1_23
rlabel metal2 s 18726 0 18754 990 4 rbl0_24
rlabel metal2 s 19204 0 19232 990 4 rbl1_24
rlabel metal2 s 19504 0 19532 990 4 rbl0_25
rlabel metal2 s 19982 0 20010 990 4 rbl1_25
rlabel metal2 s 20282 0 20310 990 4 rbl0_26
rlabel metal2 s 20760 0 20788 990 4 rbl1_26
rlabel metal2 s 21060 0 21088 990 4 rbl0_27
rlabel metal2 s 21538 0 21566 990 4 rbl1_27
rlabel metal2 s 21838 0 21866 990 4 rbl0_28
rlabel metal2 s 22316 0 22344 990 4 rbl1_28
rlabel metal2 s 22616 0 22644 990 4 rbl0_29
rlabel metal2 s 23094 0 23122 990 4 rbl1_29
rlabel metal2 s 23394 0 23422 990 4 rbl0_30
rlabel metal2 s 23872 0 23900 990 4 rbl1_30
rlabel metal2 s 24172 0 24200 990 4 rbl0_31
rlabel metal2 s 24650 0 24678 990 4 rbl1_31
rlabel metal2 s 24950 0 24978 990 4 rbl0_32
rlabel metal2 s 25428 0 25456 990 4 rbl1_32
<< properties >>
string FIXED_BBOX 0 0 25674 990
string GDS_FILE sram_0rw2r1w_16_32_sky130A.gds
string GDS_END 772798
string GDS_START 750012
<< end >>
