magic
tech sky130A
magscale 1 2
timestamp 1643678851
<< checkpaint >>
rect -1235 -1176 1385 1345
<< labels >>
rlabel mvvaractor s 75 84 75 84 4 G
rlabel mvpsubdiff s 25 84 25 84 4 S
rlabel mvpsubdiff s 125 84 125 84 4 D
<< properties >>
string GDS_FILE sram_0rw2r1w_16_128_sky130A.gds
string GDS_END 1882938
string GDS_START 1882254
<< end >>
