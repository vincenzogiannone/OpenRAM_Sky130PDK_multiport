magic
tech sky130A
magscale 1 2
timestamp 1643593061
<< checkpaint >>
rect -1260 -1302 7690 25922
<< metal1 >>
rect 5331 23998 5744 24026
rect 5331 23906 5359 23998
rect 6370 23928 6398 23956
rect 5240 23878 5442 23906
rect 5240 23760 5268 23878
rect 5187 23732 5268 23760
rect 5187 23644 5215 23732
rect 5240 23644 5268 23732
rect 5331 23644 5359 23878
rect 6370 23802 6398 23830
rect 5166 23616 5359 23644
rect 5187 23522 5215 23616
rect 5166 23494 5215 23522
rect 5240 23376 5268 23616
rect 6370 23576 6398 23604
rect 5166 23348 5268 23376
rect 6370 22536 6398 22564
rect 5187 22380 5264 22408
rect 5187 22072 5215 22380
rect 6370 22310 6398 22338
rect 5240 22234 5442 22262
rect 5240 22072 5268 22234
rect 6370 22184 6398 22212
rect 5166 22044 5268 22072
rect 5331 22114 5744 22142
rect 5187 21926 5215 22044
rect 5166 21898 5215 21926
rect 5331 21804 5359 22114
rect 5166 21776 5359 21804
rect 5331 20922 5744 20950
rect 5331 20830 5359 20922
rect 6370 20852 6398 20880
rect 5240 20802 5442 20830
rect 5240 20684 5268 20802
rect 5187 20656 5268 20684
rect 5187 20616 5215 20656
rect 5240 20616 5268 20656
rect 5331 20616 5359 20802
rect 6370 20726 6398 20754
rect 5166 20588 5359 20616
rect 5187 20494 5215 20588
rect 5166 20466 5215 20494
rect 5240 20348 5268 20588
rect 6370 20500 6398 20528
rect 5166 20320 5268 20348
rect 6370 19460 6398 19488
rect 5187 19304 5264 19332
rect 5187 19044 5215 19304
rect 6370 19234 6398 19262
rect 5240 19158 5442 19186
rect 5240 19044 5268 19158
rect 6370 19108 6398 19136
rect 5166 19016 5268 19044
rect 5331 19038 5744 19066
rect 5187 18898 5215 19016
rect 5166 18870 5215 18898
rect 5331 18776 5359 19038
rect 5166 18748 5359 18776
rect 5331 17846 5744 17874
rect 5331 17754 5359 17846
rect 6370 17776 6398 17804
rect 5240 17726 5442 17754
rect 5240 17608 5268 17726
rect 5187 17588 5268 17608
rect 5331 17588 5359 17726
rect 6370 17650 6398 17678
rect 5166 17560 5359 17588
rect 5187 17466 5215 17560
rect 5166 17438 5215 17466
rect 5240 17320 5268 17560
rect 6370 17424 6398 17452
rect 5166 17292 5268 17320
rect 6370 16384 6398 16412
rect 5187 16228 5264 16256
rect 5187 16016 5215 16228
rect 6370 16158 6398 16186
rect 5240 16082 5442 16110
rect 5240 16016 5268 16082
rect 6370 16032 6398 16060
rect 5166 15988 5268 16016
rect 5187 15870 5215 15988
rect 5166 15842 5215 15870
rect 5331 15962 5744 15990
rect 5331 15748 5359 15962
rect 5166 15720 5359 15748
rect 5331 14770 5744 14798
rect 5331 14678 5359 14770
rect 6370 14700 6398 14728
rect 5240 14650 5442 14678
rect 5240 14560 5268 14650
rect 5331 14560 5359 14650
rect 6370 14574 6398 14602
rect 5166 14532 5359 14560
rect 5187 14504 5268 14532
rect 5187 14438 5215 14504
rect 5166 14410 5215 14438
rect 5240 14292 5268 14504
rect 6370 14348 6398 14376
rect 5166 14264 5268 14292
rect 6370 13308 6398 13336
rect 5187 13152 5264 13180
rect 5187 12988 5215 13152
rect 6370 13082 6398 13110
rect 5240 13006 5442 13034
rect 5240 12988 5268 13006
rect 5166 12960 5268 12988
rect 5187 12842 5215 12960
rect 6370 12956 6398 12984
rect 5166 12814 5215 12842
rect 5331 12886 5744 12914
rect 5331 12720 5359 12886
rect 5166 12692 5359 12720
rect 5331 11694 5744 11722
rect 5331 11602 5359 11694
rect 6370 11624 6398 11652
rect 5240 11574 5442 11602
rect 5240 11532 5268 11574
rect 5331 11532 5359 11574
rect 5166 11504 5359 11532
rect 5240 11456 5268 11504
rect 6370 11498 6398 11526
rect 5187 11428 5268 11456
rect 5187 11410 5215 11428
rect 5166 11382 5215 11410
rect 5240 11264 5268 11428
rect 6370 11272 6398 11300
rect 5166 11236 5268 11264
rect 6370 10232 6398 10260
rect 5187 10076 5264 10104
rect 5187 9960 5215 10076
rect 6370 10006 6398 10034
rect 5166 9958 5268 9960
rect 5166 9932 5442 9958
rect 5187 9814 5215 9932
rect 5240 9930 5442 9932
rect 6370 9880 6398 9908
rect 5166 9786 5215 9814
rect 5331 9810 5744 9838
rect 5331 9692 5359 9810
rect 5166 9664 5359 9692
rect 5331 8618 5744 8646
rect 5331 8526 5359 8618
rect 6370 8548 6398 8576
rect 5240 8504 5442 8526
rect 5166 8498 5442 8504
rect 5166 8476 5359 8498
rect 5166 8380 5215 8382
rect 5240 8380 5268 8476
rect 6370 8422 6398 8450
rect 5166 8354 5268 8380
rect 5187 8352 5268 8354
rect 5240 8236 5268 8352
rect 5166 8208 5268 8236
rect 6370 8196 6398 8224
rect 6370 7156 6398 7184
rect 5187 7000 5264 7028
rect 5187 6932 5215 7000
rect 5166 6904 5268 6932
rect 6370 6930 6398 6958
rect 5187 6786 5215 6904
rect 5240 6882 5268 6904
rect 5240 6854 5442 6882
rect 6370 6804 6398 6832
rect 5166 6758 5215 6786
rect 5331 6734 5744 6762
rect 5331 6664 5359 6734
rect 5166 6636 5359 6664
rect 5331 5542 5744 5570
rect 5331 5476 5359 5542
rect 5166 5450 5359 5476
rect 6370 5472 6398 5500
rect 5166 5448 5442 5450
rect 5240 5422 5442 5448
rect 5166 5326 5215 5354
rect 5187 5304 5215 5326
rect 5240 5304 5268 5422
rect 6370 5346 6398 5374
rect 5187 5276 5268 5304
rect 5240 5208 5268 5276
rect 5166 5180 5268 5208
rect 6370 5120 6398 5148
rect 6370 4080 6398 4108
rect 5187 3924 5264 3952
rect 5187 3904 5215 3924
rect 5166 3876 5268 3904
rect 5187 3758 5215 3876
rect 5240 3806 5268 3876
rect 6370 3854 6398 3882
rect 5240 3778 5442 3806
rect 5166 3730 5215 3758
rect 6370 3728 6398 3756
rect 5331 3658 5744 3686
rect 5331 3636 5359 3658
rect 5166 3608 5359 3636
rect 5331 2466 5744 2494
rect 5331 2448 5359 2466
rect 5166 2420 5359 2448
rect 6370 2396 6398 2424
rect 5240 2346 5442 2374
rect 5166 2298 5215 2326
rect 5187 2228 5215 2298
rect 5240 2228 5268 2346
rect 6370 2270 6398 2298
rect 5187 2200 5268 2228
rect 5240 2180 5268 2200
rect 5166 2152 5268 2180
rect 6370 2044 6398 2072
rect 6370 1004 6398 1032
rect 5166 848 5268 876
rect 5187 730 5215 848
rect 5166 702 5215 730
rect 5240 730 5268 848
rect 6370 778 6398 806
rect 5240 702 5442 730
rect 6370 652 6398 680
rect 5331 608 5744 610
rect 5166 582 5744 608
rect 5166 580 5359 582
<< metal2 >>
rect 18 0 46 24632
rect 102 0 130 24632
rect 186 0 214 24632
rect 270 0 298 24632
rect 354 0 382 24632
rect 438 0 466 24632
rect 5008 24594 5222 24622
<< metal3 >>
rect 828 24602 888 24662
rect 1700 24602 1760 24662
rect 6368 24578 6428 24638
rect 5164 24194 5224 24254
rect 828 23062 888 23122
rect 1700 23062 1760 23122
rect 6368 23040 6428 23100
rect 5164 22680 5224 22740
rect 828 21522 888 21582
rect 1700 21522 1760 21582
rect 6368 21502 6428 21562
rect 5164 21166 5224 21226
rect 828 19982 888 20042
rect 1700 19982 1760 20042
rect 6368 19964 6428 20024
rect 5164 19652 5224 19712
rect 828 18442 888 18502
rect 1700 18442 1760 18502
rect 6368 18426 6428 18486
rect 5164 18138 5224 18198
rect 6368 16888 6428 16948
rect 5164 16624 5224 16684
rect 828 15366 888 15426
rect 1700 15366 1760 15426
rect 6368 15350 6428 15410
rect 5164 15110 5224 15170
rect 828 13826 888 13886
rect 1700 13826 1760 13886
rect 6368 13812 6428 13872
rect 5164 13596 5224 13656
rect 828 12286 888 12346
rect 1700 12286 1760 12346
rect 6368 12274 6428 12334
rect 5164 12082 5224 12142
rect 828 10746 888 10806
rect 1700 10746 1760 10806
rect 6368 10736 6428 10796
rect 5164 10568 5224 10628
rect 828 9206 888 9266
rect 1700 9206 1760 9266
rect 6368 9198 6428 9258
rect 5164 9054 5224 9114
rect 6368 7660 6428 7720
rect 5164 7540 5224 7600
rect 828 6130 888 6190
rect 1700 6130 1760 6190
rect 6368 6122 6428 6182
rect 5164 6026 5224 6086
rect 828 4590 888 4650
rect 1700 4590 1760 4650
rect 6368 4584 6428 4644
rect 5164 4512 5224 4572
rect 828 3050 888 3110
rect 1700 3050 1760 3110
rect 5164 2998 5224 3058
rect 6368 3046 6428 3106
rect 828 1510 888 1570
rect 1700 1510 1760 1570
rect 5164 1484 5224 1544
rect 6368 1508 6428 1568
rect 828 -30 888 30
rect 1700 -30 1760 30
rect 5164 -30 5224 30
rect 6368 -30 6428 30
use wordline_driver_array  wordline_driver_array_0
timestamp 1643593061
transform 1 0 5194 0 1 0
box 0 -42 1236 24650
use hierarchical_decoder  hierarchical_decoder_0
timestamp 1643593061
transform 1 0 0 0 1 0
box 0 -42 5226 24662
<< labels >>
rlabel metal2 s 18 0 46 24632 4 addr0
rlabel metal2 s 102 0 130 24632 4 addr1
rlabel metal2 s 186 0 214 24632 4 addr2
rlabel metal2 s 270 0 298 24632 4 addr3
rlabel metal2 s 354 0 382 24632 4 addr4
rlabel metal2 s 438 0 466 24632 4 addr5
rlabel metal1 s 6370 778 6398 806 4 rwl0_0
rlabel metal1 s 6370 1004 6398 1032 4 rwl1_0
rlabel metal1 s 6370 652 6398 680 4 wwl0_0
rlabel metal1 s 6370 2270 6398 2298 4 rwl0_1
rlabel metal1 s 6370 2044 6398 2072 4 rwl1_1
rlabel metal1 s 6370 2396 6398 2424 4 wwl0_1
rlabel metal1 s 6370 3854 6398 3882 4 rwl0_2
rlabel metal1 s 6370 4080 6398 4108 4 rwl1_2
rlabel metal1 s 6370 3728 6398 3756 4 wwl0_2
rlabel metal1 s 6370 5346 6398 5374 4 rwl0_3
rlabel metal1 s 6370 5120 6398 5148 4 rwl1_3
rlabel metal1 s 6370 5472 6398 5500 4 wwl0_3
rlabel metal1 s 6370 6930 6398 6958 4 rwl0_4
rlabel metal1 s 6370 7156 6398 7184 4 rwl1_4
rlabel metal1 s 6370 6804 6398 6832 4 wwl0_4
rlabel metal1 s 6370 8422 6398 8450 4 rwl0_5
rlabel metal1 s 6370 8196 6398 8224 4 rwl1_5
rlabel metal1 s 6370 8548 6398 8576 4 wwl0_5
rlabel metal1 s 6370 10006 6398 10034 4 rwl0_6
rlabel metal1 s 6370 10232 6398 10260 4 rwl1_6
rlabel metal1 s 6370 9880 6398 9908 4 wwl0_6
rlabel metal1 s 6370 11498 6398 11526 4 rwl0_7
rlabel metal1 s 6370 11272 6398 11300 4 rwl1_7
rlabel metal1 s 6370 11624 6398 11652 4 wwl0_7
rlabel metal1 s 6370 13082 6398 13110 4 rwl0_8
rlabel metal1 s 6370 13308 6398 13336 4 rwl1_8
rlabel metal1 s 6370 12956 6398 12984 4 wwl0_8
rlabel metal1 s 6370 14574 6398 14602 4 rwl0_9
rlabel metal1 s 6370 14348 6398 14376 4 rwl1_9
rlabel metal1 s 6370 14700 6398 14728 4 wwl0_9
rlabel metal1 s 6370 16158 6398 16186 4 rwl0_10
rlabel metal1 s 6370 16384 6398 16412 4 rwl1_10
rlabel metal1 s 6370 16032 6398 16060 4 wwl0_10
rlabel metal1 s 6370 17650 6398 17678 4 rwl0_11
rlabel metal1 s 6370 17424 6398 17452 4 rwl1_11
rlabel metal1 s 6370 17776 6398 17804 4 wwl0_11
rlabel metal1 s 6370 19234 6398 19262 4 rwl0_12
rlabel metal1 s 6370 19460 6398 19488 4 rwl1_12
rlabel metal1 s 6370 19108 6398 19136 4 wwl0_12
rlabel metal1 s 6370 20726 6398 20754 4 rwl0_13
rlabel metal1 s 6370 20500 6398 20528 4 rwl1_13
rlabel metal1 s 6370 20852 6398 20880 4 wwl0_13
rlabel metal1 s 6370 22310 6398 22338 4 rwl0_14
rlabel metal1 s 6370 22536 6398 22564 4 rwl1_14
rlabel metal1 s 6370 22184 6398 22212 4 wwl0_14
rlabel metal1 s 6370 23802 6398 23830 4 rwl0_15
rlabel metal1 s 6370 23576 6398 23604 4 rwl1_15
rlabel metal1 s 6370 23928 6398 23956 4 wwl0_15
rlabel metal2 s 5194 24594 5222 24622 4 wl_en
rlabel metal3 s 1700 19982 1760 20042 4 vdd
rlabel metal3 s 5164 7540 5224 7600 4 vdd
rlabel metal3 s 828 23062 888 23122 4 vdd
rlabel metal3 s 1700 13826 1760 13886 4 vdd
rlabel metal3 s 5164 13596 5224 13656 4 vdd
rlabel metal3 s 828 19982 888 20042 4 vdd
rlabel metal3 s 5164 10568 5224 10628 4 vdd
rlabel metal3 s 828 1510 888 1570 4 vdd
rlabel metal3 s 6368 1508 6428 1568 4 vdd
rlabel metal3 s 6368 19964 6428 20024 4 vdd
rlabel metal3 s 828 10746 888 10806 4 vdd
rlabel metal3 s 5164 19652 5224 19712 4 vdd
rlabel metal3 s 1700 1510 1760 1570 4 vdd
rlabel metal3 s 5164 16624 5224 16684 4 vdd
rlabel metal3 s 6368 13812 6428 13872 4 vdd
rlabel metal3 s 6368 10736 6428 10796 4 vdd
rlabel metal3 s 828 13826 888 13886 4 vdd
rlabel metal3 s 6368 23040 6428 23100 4 vdd
rlabel metal3 s 5164 22680 5224 22740 4 vdd
rlabel metal3 s 1700 4590 1760 4650 4 vdd
rlabel metal3 s 6368 16888 6428 16948 4 vdd
rlabel metal3 s 5164 1484 5224 1544 4 vdd
rlabel metal3 s 5164 4512 5224 4572 4 vdd
rlabel metal3 s 1700 23062 1760 23122 4 vdd
rlabel metal3 s 1700 10746 1760 10806 4 vdd
rlabel metal3 s 828 4590 888 4650 4 vdd
rlabel metal3 s 6368 7660 6428 7720 4 vdd
rlabel metal3 s 6368 4584 6428 4644 4 vdd
rlabel metal3 s 5164 6026 5224 6086 4 gnd
rlabel metal3 s 1700 -30 1760 30 4 gnd
rlabel metal3 s 1700 24602 1760 24662 4 gnd
rlabel metal3 s 828 21522 888 21582 4 gnd
rlabel metal3 s 828 3050 888 3110 4 gnd
rlabel metal3 s 5164 18138 5224 18198 4 gnd
rlabel metal3 s 5164 2998 5224 3058 4 gnd
rlabel metal3 s 828 15366 888 15426 4 gnd
rlabel metal3 s 828 6130 888 6190 4 gnd
rlabel metal3 s 5164 15110 5224 15170 4 gnd
rlabel metal3 s 5164 9054 5224 9114 4 gnd
rlabel metal3 s 5164 -30 5224 30 4 gnd
rlabel metal3 s 6368 24578 6428 24638 4 gnd
rlabel metal3 s 1700 9206 1760 9266 4 gnd
rlabel metal3 s 828 9206 888 9266 4 gnd
rlabel metal3 s 828 12286 888 12346 4 gnd
rlabel metal3 s 5164 12082 5224 12142 4 gnd
rlabel metal3 s 1700 6130 1760 6190 4 gnd
rlabel metal3 s 828 -30 888 30 4 gnd
rlabel metal3 s 6368 18426 6428 18486 4 gnd
rlabel metal3 s 5164 24194 5224 24254 4 gnd
rlabel metal3 s 6368 15350 6428 15410 4 gnd
rlabel metal3 s 5164 21166 5224 21226 4 gnd
rlabel metal3 s 6368 -30 6428 30 4 gnd
rlabel metal3 s 1700 12286 1760 12346 4 gnd
rlabel metal3 s 1700 3050 1760 3110 4 gnd
rlabel metal3 s 6368 9198 6428 9258 4 gnd
rlabel metal3 s 6368 12274 6428 12334 4 gnd
rlabel metal3 s 6368 21502 6428 21562 4 gnd
rlabel metal3 s 1700 15366 1760 15426 4 gnd
rlabel metal3 s 6368 3046 6428 3106 4 gnd
rlabel metal3 s 828 24602 888 24662 4 gnd
rlabel metal3 s 1700 21522 1760 21582 4 gnd
rlabel metal3 s 6368 6122 6428 6182 4 gnd
rlabel metal3 s 1700 18442 1760 18502 4 gnd
rlabel metal3 s 828 18442 888 18502 4 gnd
<< properties >>
string FIXED_BBOX 0 0 6434 24660
string GDS_FILE sram_0rw2r1w_2_16_sky130A.gds
string GDS_END 318098
string GDS_START 274016
<< end >>
