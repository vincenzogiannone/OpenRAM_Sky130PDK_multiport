magic
tech sky130A
magscale 1 2
timestamp 1644951705
<< checkpaint >>
rect -1296 -1277 2744 2155
<< nwell >>
rect -36 402 1484 895
<< locali >>
rect 0 821 1448 855
rect 48 340 114 406
rect 721 356 755 390
rect 0 -17 1448 17
use pinv_4  pinv_4_0
timestamp 1644951705
transform 1 0 0 0 1 0
box -36 -17 1484 895
<< labels >>
rlabel locali s 738 373 738 373 4 Z
rlabel locali s 81 373 81 373 4 A
rlabel locali s 724 0 724 0 4 gnd
rlabel locali s 724 838 724 838 4 vdd
<< properties >>
string FIXED_BBOX 0 0 1448 838
string GDS_FILE sram_0rw2r1w_16_128_sky130A.gds
string GDS_END 2021828
string GDS_START 2020984
<< end >>
