magic
tech sky130A
magscale 1 2
timestamp 1644949024
<< checkpaint >>
rect -1260 -1263 4138 2310
<< metal1 >>
rect 104 954 110 1006
rect 162 954 168 1006
rect 376 954 382 1006
rect 434 954 440 1006
rect 882 954 888 1006
rect 940 954 946 1006
rect 1154 954 1160 1006
rect 1212 954 1218 1006
rect 1660 954 1666 1006
rect 1718 954 1724 1006
rect 1932 954 1938 1006
rect 1990 954 1996 1006
rect 2438 954 2444 1006
rect 2496 954 2502 1006
rect 2710 954 2716 1006
rect 2768 954 2774 1006
rect 104 8 110 60
rect 162 8 168 60
rect 376 8 382 60
rect 434 8 440 60
rect 882 8 888 60
rect 940 8 946 60
rect 1154 8 1160 60
rect 1212 8 1218 60
rect 1660 8 1666 60
rect 1718 8 1724 60
rect 1932 8 1938 60
rect 1990 8 1996 60
rect 2438 8 2444 60
rect 2496 8 2502 60
rect 2710 8 2716 60
rect 2768 8 2774 60
<< via1 >>
rect 110 954 162 1006
rect 382 954 434 1006
rect 888 954 940 1006
rect 1160 954 1212 1006
rect 1666 954 1718 1006
rect 1938 954 1990 1006
rect 2444 954 2496 1006
rect 2716 954 2768 1006
rect 110 8 162 60
rect 382 8 434 60
rect 888 8 940 60
rect 1160 8 1212 60
rect 1666 8 1718 60
rect 1938 8 1990 60
rect 2444 8 2496 60
rect 2716 8 2768 60
<< metal2 >>
rect 108 1008 164 1017
rect 108 943 164 952
rect 380 1008 436 1017
rect 380 943 436 952
rect 886 1008 942 1017
rect 886 943 942 952
rect 1158 1008 1214 1017
rect 1158 943 1214 952
rect 1664 1008 1720 1017
rect 1664 943 1720 952
rect 1936 1008 1992 1017
rect 1936 943 1992 952
rect 2442 1008 2498 1017
rect 2442 943 2498 952
rect 2714 1008 2770 1017
rect 2714 943 2770 952
rect 14 0 42 240
rect 108 62 164 71
rect 108 -3 164 6
rect 202 0 230 240
rect 286 0 314 240
rect 380 62 436 71
rect 380 -3 436 6
rect 474 0 502 240
rect 792 0 820 240
rect 886 62 942 71
rect 886 -3 942 6
rect 980 0 1008 240
rect 1064 0 1092 240
rect 1158 62 1214 71
rect 1158 -3 1214 6
rect 1252 0 1280 240
rect 1570 0 1598 240
rect 1664 62 1720 71
rect 1664 -3 1720 6
rect 1758 0 1786 240
rect 1842 0 1870 240
rect 1936 62 1992 71
rect 1936 -3 1992 6
rect 2030 0 2058 240
rect 2348 0 2376 240
rect 2442 62 2498 71
rect 2442 -3 2498 6
rect 2536 0 2564 240
rect 2620 0 2648 240
rect 2714 62 2770 71
rect 2714 -3 2770 6
rect 2808 0 2836 240
<< via2 >>
rect 108 1006 164 1008
rect 108 954 110 1006
rect 110 954 162 1006
rect 162 954 164 1006
rect 108 952 164 954
rect 380 1006 436 1008
rect 380 954 382 1006
rect 382 954 434 1006
rect 434 954 436 1006
rect 380 952 436 954
rect 886 1006 942 1008
rect 886 954 888 1006
rect 888 954 940 1006
rect 940 954 942 1006
rect 886 952 942 954
rect 1158 1006 1214 1008
rect 1158 954 1160 1006
rect 1160 954 1212 1006
rect 1212 954 1214 1006
rect 1158 952 1214 954
rect 1664 1006 1720 1008
rect 1664 954 1666 1006
rect 1666 954 1718 1006
rect 1718 954 1720 1006
rect 1664 952 1720 954
rect 1936 1006 1992 1008
rect 1936 954 1938 1006
rect 1938 954 1990 1006
rect 1990 954 1992 1006
rect 1936 952 1992 954
rect 2442 1006 2498 1008
rect 2442 954 2444 1006
rect 2444 954 2496 1006
rect 2496 954 2498 1006
rect 2442 952 2498 954
rect 2714 1006 2770 1008
rect 2714 954 2716 1006
rect 2716 954 2768 1006
rect 2768 954 2770 1006
rect 2714 952 2770 954
rect 108 60 164 62
rect 108 8 110 60
rect 110 8 162 60
rect 162 8 164 60
rect 108 6 164 8
rect 380 60 436 62
rect 380 8 382 60
rect 382 8 434 60
rect 434 8 436 60
rect 380 6 436 8
rect 886 60 942 62
rect 886 8 888 60
rect 888 8 940 60
rect 940 8 942 60
rect 886 6 942 8
rect 1158 60 1214 62
rect 1158 8 1160 60
rect 1160 8 1212 60
rect 1212 8 1214 60
rect 1158 6 1214 8
rect 1664 60 1720 62
rect 1664 8 1666 60
rect 1666 8 1718 60
rect 1718 8 1720 60
rect 1664 6 1720 8
rect 1936 60 1992 62
rect 1936 8 1938 60
rect 1938 8 1990 60
rect 1990 8 1992 60
rect 1936 6 1992 8
rect 2442 60 2498 62
rect 2442 8 2444 60
rect 2444 8 2496 60
rect 2496 8 2498 60
rect 2442 6 2498 8
rect 2714 60 2770 62
rect 2714 8 2716 60
rect 2716 8 2768 60
rect 2768 8 2770 60
rect 2714 6 2770 8
<< metal3 >>
rect 70 1008 202 1017
rect 70 952 108 1008
rect 164 952 202 1008
rect 70 943 202 952
rect 342 1008 474 1017
rect 342 952 380 1008
rect 436 952 474 1008
rect 342 943 474 952
rect 848 1008 980 1017
rect 848 952 886 1008
rect 942 952 980 1008
rect 848 943 980 952
rect 1120 1008 1252 1017
rect 1120 952 1158 1008
rect 1214 952 1252 1008
rect 1120 943 1252 952
rect 1626 1008 1758 1017
rect 1626 952 1664 1008
rect 1720 952 1758 1008
rect 1626 943 1758 952
rect 1898 1008 2030 1017
rect 1898 952 1936 1008
rect 1992 952 2030 1008
rect 1898 943 2030 952
rect 2404 1008 2536 1017
rect 2404 952 2442 1008
rect 2498 952 2536 1008
rect 2404 943 2536 952
rect 2676 1008 2808 1017
rect 2676 952 2714 1008
rect 2770 952 2808 1008
rect 2676 943 2808 952
rect 70 62 202 71
rect 70 6 108 62
rect 164 6 202 62
rect 70 -3 202 6
rect 342 62 474 71
rect 342 6 380 62
rect 436 6 474 62
rect 342 -3 474 6
rect 848 62 980 71
rect 848 6 886 62
rect 942 6 980 62
rect 848 -3 980 6
rect 1120 62 1252 71
rect 1120 6 1158 62
rect 1214 6 1252 62
rect 1120 -3 1252 6
rect 1626 62 1758 71
rect 1626 6 1664 62
rect 1720 6 1758 62
rect 1626 -3 1758 6
rect 1898 62 2030 71
rect 1898 6 1936 62
rect 1992 6 2030 62
rect 1898 -3 2030 6
rect 2404 62 2536 71
rect 2404 6 2442 62
rect 2498 6 2536 62
rect 2404 -3 2536 6
rect 2676 62 2808 71
rect 2676 6 2714 62
rect 2770 6 2808 62
rect 2676 -3 2808 6
use contact_18  contact_18_0
timestamp 1644949024
transform 1 0 2676 0 1 943
box 0 0 1 1
use contact_17  contact_17_0
timestamp 1644949024
transform 1 0 2710 0 1 948
box 0 0 1 1
use contact_18  contact_18_1
timestamp 1644949024
transform 1 0 2676 0 1 -3
box 0 0 1 1
use contact_17  contact_17_1
timestamp 1644949024
transform 1 0 2710 0 1 2
box 0 0 1 1
use contact_18  contact_18_2
timestamp 1644949024
transform 1 0 2404 0 1 943
box 0 0 1 1
use contact_17  contact_17_2
timestamp 1644949024
transform 1 0 2438 0 1 948
box 0 0 1 1
use contact_18  contact_18_3
timestamp 1644949024
transform 1 0 2404 0 1 -3
box 0 0 1 1
use contact_17  contact_17_3
timestamp 1644949024
transform 1 0 2438 0 1 2
box 0 0 1 1
use contact_18  contact_18_4
timestamp 1644949024
transform 1 0 1898 0 1 943
box 0 0 1 1
use contact_17  contact_17_4
timestamp 1644949024
transform 1 0 1932 0 1 948
box 0 0 1 1
use contact_18  contact_18_5
timestamp 1644949024
transform 1 0 1898 0 1 -3
box 0 0 1 1
use contact_17  contact_17_5
timestamp 1644949024
transform 1 0 1932 0 1 2
box 0 0 1 1
use contact_18  contact_18_6
timestamp 1644949024
transform 1 0 1626 0 1 943
box 0 0 1 1
use contact_17  contact_17_6
timestamp 1644949024
transform 1 0 1660 0 1 948
box 0 0 1 1
use contact_18  contact_18_7
timestamp 1644949024
transform 1 0 1626 0 1 -3
box 0 0 1 1
use contact_17  contact_17_7
timestamp 1644949024
transform 1 0 1660 0 1 2
box 0 0 1 1
use contact_18  contact_18_8
timestamp 1644949024
transform 1 0 1120 0 1 943
box 0 0 1 1
use contact_17  contact_17_8
timestamp 1644949024
transform 1 0 1154 0 1 948
box 0 0 1 1
use contact_18  contact_18_9
timestamp 1644949024
transform 1 0 1120 0 1 -3
box 0 0 1 1
use contact_17  contact_17_9
timestamp 1644949024
transform 1 0 1154 0 1 2
box 0 0 1 1
use contact_18  contact_18_10
timestamp 1644949024
transform 1 0 848 0 1 943
box 0 0 1 1
use contact_17  contact_17_10
timestamp 1644949024
transform 1 0 882 0 1 948
box 0 0 1 1
use contact_18  contact_18_11
timestamp 1644949024
transform 1 0 848 0 1 -3
box 0 0 1 1
use contact_17  contact_17_11
timestamp 1644949024
transform 1 0 882 0 1 2
box 0 0 1 1
use contact_18  contact_18_12
timestamp 1644949024
transform 1 0 342 0 1 943
box 0 0 1 1
use contact_17  contact_17_12
timestamp 1644949024
transform 1 0 376 0 1 948
box 0 0 1 1
use contact_18  contact_18_13
timestamp 1644949024
transform 1 0 342 0 1 -3
box 0 0 1 1
use contact_17  contact_17_13
timestamp 1644949024
transform 1 0 376 0 1 2
box 0 0 1 1
use contact_18  contact_18_14
timestamp 1644949024
transform 1 0 70 0 1 943
box 0 0 1 1
use contact_17  contact_17_14
timestamp 1644949024
transform 1 0 104 0 1 948
box 0 0 1 1
use contact_18  contact_18_15
timestamp 1644949024
transform 1 0 70 0 1 -3
box 0 0 1 1
use contact_17  contact_17_15
timestamp 1644949024
transform 1 0 104 0 1 2
box 0 0 1 1
use sense_amp_multiport  sense_amp_multiport_0
timestamp 1644949024
transform 1 0 2606 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_1
timestamp 1644949024
transform 1 0 2334 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_2
timestamp 1644949024
transform 1 0 1828 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_3
timestamp 1644949024
transform 1 0 1556 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_4
timestamp 1644949024
transform 1 0 1050 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_5
timestamp 1644949024
transform 1 0 778 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_6
timestamp 1644949024
transform 1 0 272 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_7
timestamp 1644949024
transform 1 0 0 0 1 0
box 0 0 272 1050
<< labels >>
rlabel metal3 s 1120 -3 1252 71 4 gnd
rlabel metal3 s 2404 -3 2536 71 4 gnd
rlabel metal3 s 342 -3 474 71 4 gnd
rlabel metal3 s 848 -3 980 71 4 gnd
rlabel metal3 s 70 -3 202 71 4 gnd
rlabel metal3 s 1626 -3 1758 71 4 gnd
rlabel metal3 s 2676 -3 2808 71 4 gnd
rlabel metal3 s 1898 -3 2030 71 4 gnd
rlabel metal3 s 2404 943 2536 1017 4 vdd
rlabel metal3 s 1626 943 1758 1017 4 vdd
rlabel metal3 s 1898 943 2030 1017 4 vdd
rlabel metal3 s 342 943 474 1017 4 vdd
rlabel metal3 s 1120 943 1252 1017 4 vdd
rlabel metal3 s 70 943 202 1017 4 vdd
rlabel metal3 s 2676 943 2808 1017 4 vdd
rlabel metal3 s 848 943 980 1017 4 vdd
rlabel metal2 s 14 0 42 240 4 rbl_0
rlabel metal2 s 202 0 230 240 4 data_0
rlabel metal2 s 286 0 314 240 4 rbl_1
rlabel metal2 s 474 0 502 240 4 data_1
rlabel metal2 s 792 0 820 240 4 rbl_2
rlabel metal2 s 980 0 1008 240 4 data_2
rlabel metal2 s 1064 0 1092 240 4 rbl_3
rlabel metal2 s 1252 0 1280 240 4 data_3
rlabel metal2 s 1570 0 1598 240 4 rbl_4
rlabel metal2 s 1758 0 1786 240 4 data_4
rlabel metal2 s 1842 0 1870 240 4 rbl_5
rlabel metal2 s 2030 0 2058 240 4 data_5
rlabel metal2 s 2348 0 2376 240 4 rbl_6
rlabel metal2 s 2536 0 2564 240 4 data_6
rlabel metal2 s 2620 0 2648 240 4 rbl_7
rlabel metal2 s 2808 0 2836 240 4 data_7
<< properties >>
string FIXED_BBOX 2676 -3 2808 0
string GDS_FILE sram_0rw2r1w_4_16_sky130A.gds
string GDS_END 210086
string GDS_START 201266
<< end >>
