magic
tech sky130A
magscale 1 2
timestamp 1644969367
<< checkpaint >>
rect -1260 -1302 2530 99734
<< metal1 >>
rect 1172 98406 1178 98458
rect 1230 98406 1236 98458
rect 536 97822 618 97850
rect 1176 97752 1204 97780
rect 234 97702 318 97730
rect 1176 97626 1204 97654
rect 56 97556 126 97584
rect 1176 97400 1204 97428
rect 1172 96868 1178 96920
rect 1230 96868 1236 96920
rect 1176 96360 1204 96388
rect 56 96204 126 96232
rect 1176 96134 1204 96162
rect 234 96058 318 96086
rect 1176 96008 1204 96036
rect 536 95938 618 95966
rect 1172 95330 1178 95382
rect 1230 95330 1236 95382
rect 536 94746 618 94774
rect 1176 94676 1204 94704
rect 234 94626 318 94654
rect 1176 94550 1204 94578
rect 56 94480 126 94508
rect 1176 94324 1204 94352
rect 1172 93792 1178 93844
rect 1230 93792 1236 93844
rect 1176 93284 1204 93312
rect 56 93128 126 93156
rect 1176 93058 1204 93086
rect 234 92982 318 93010
rect 1176 92932 1204 92960
rect 536 92862 618 92890
rect 1172 92254 1178 92306
rect 1230 92254 1236 92306
rect 536 91670 618 91698
rect 1176 91600 1204 91628
rect 234 91550 318 91578
rect 1176 91474 1204 91502
rect 56 91404 126 91432
rect 1176 91248 1204 91276
rect 1172 90716 1178 90768
rect 1230 90716 1236 90768
rect 1176 90208 1204 90236
rect 56 90052 126 90080
rect 1176 89982 1204 90010
rect 234 89906 318 89934
rect 1176 89856 1204 89884
rect 536 89786 618 89814
rect 1172 89178 1178 89230
rect 1230 89178 1236 89230
rect 536 88594 618 88622
rect 1176 88524 1204 88552
rect 234 88474 318 88502
rect 1176 88398 1204 88426
rect 56 88328 126 88356
rect 1176 88172 1204 88200
rect 1172 87640 1178 87692
rect 1230 87640 1236 87692
rect 1176 87132 1204 87160
rect 56 86976 126 87004
rect 1176 86906 1204 86934
rect 234 86830 318 86858
rect 1176 86780 1204 86808
rect 536 86710 618 86738
rect 1172 86102 1178 86154
rect 1230 86102 1236 86154
rect 536 85518 618 85546
rect 1176 85448 1204 85476
rect 234 85398 318 85426
rect 1176 85322 1204 85350
rect 56 85252 126 85280
rect 1176 85096 1204 85124
rect 1172 84564 1178 84616
rect 1230 84564 1236 84616
rect 1176 84056 1204 84084
rect 56 83900 126 83928
rect 1176 83830 1204 83858
rect 234 83754 318 83782
rect 1176 83704 1204 83732
rect 536 83634 618 83662
rect 1172 83026 1178 83078
rect 1230 83026 1236 83078
rect 536 82442 618 82470
rect 1176 82372 1204 82400
rect 234 82322 318 82350
rect 1176 82246 1204 82274
rect 56 82176 126 82204
rect 1176 82020 1204 82048
rect 1172 81488 1178 81540
rect 1230 81488 1236 81540
rect 1176 80980 1204 81008
rect 56 80824 126 80852
rect 1176 80754 1204 80782
rect 234 80678 318 80706
rect 1176 80628 1204 80656
rect 536 80558 618 80586
rect 1172 79950 1178 80002
rect 1230 79950 1236 80002
rect 536 79366 618 79394
rect 1176 79296 1204 79324
rect 234 79246 318 79274
rect 1176 79170 1204 79198
rect 56 79100 126 79128
rect 1176 78944 1204 78972
rect 1172 78412 1178 78464
rect 1230 78412 1236 78464
rect 1176 77904 1204 77932
rect 56 77748 126 77776
rect 1176 77678 1204 77706
rect 234 77602 318 77630
rect 1176 77552 1204 77580
rect 536 77482 618 77510
rect 1172 76874 1178 76926
rect 1230 76874 1236 76926
rect 536 76290 618 76318
rect 1176 76220 1204 76248
rect 234 76170 318 76198
rect 1176 76094 1204 76122
rect 56 76024 126 76052
rect 1176 75868 1204 75896
rect 1172 75336 1178 75388
rect 1230 75336 1236 75388
rect 1176 74828 1204 74856
rect 56 74672 126 74700
rect 1176 74602 1204 74630
rect 234 74526 318 74554
rect 1176 74476 1204 74504
rect 536 74406 618 74434
rect 1172 73798 1178 73850
rect 1230 73798 1236 73850
rect 536 73214 618 73242
rect 1176 73144 1204 73172
rect 234 73094 318 73122
rect 1176 73018 1204 73046
rect 56 72948 126 72976
rect 1176 72792 1204 72820
rect 1172 72260 1178 72312
rect 1230 72260 1236 72312
rect 1176 71752 1204 71780
rect 56 71596 126 71624
rect 1176 71526 1204 71554
rect 234 71450 318 71478
rect 1176 71400 1204 71428
rect 536 71330 618 71358
rect 1172 70722 1178 70774
rect 1230 70722 1236 70774
rect 536 70138 618 70166
rect 1176 70068 1204 70096
rect 234 70018 318 70046
rect 1176 69942 1204 69970
rect 56 69872 126 69900
rect 1176 69716 1204 69744
rect 1172 69184 1178 69236
rect 1230 69184 1236 69236
rect 1176 68676 1204 68704
rect 56 68520 126 68548
rect 1176 68450 1204 68478
rect 234 68374 318 68402
rect 1176 68324 1204 68352
rect 536 68254 618 68282
rect 1172 67646 1178 67698
rect 1230 67646 1236 67698
rect 536 67062 618 67090
rect 1176 66992 1204 67020
rect 234 66942 318 66970
rect 1176 66866 1204 66894
rect 56 66796 126 66824
rect 1176 66640 1204 66668
rect 1172 66108 1178 66160
rect 1230 66108 1236 66160
rect 1176 65600 1204 65628
rect 56 65444 126 65472
rect 1176 65374 1204 65402
rect 234 65298 318 65326
rect 1176 65248 1204 65276
rect 536 65178 618 65206
rect 1172 64570 1178 64622
rect 1230 64570 1236 64622
rect 536 63986 618 64014
rect 1176 63916 1204 63944
rect 234 63866 318 63894
rect 1176 63790 1204 63818
rect 56 63720 126 63748
rect 1176 63564 1204 63592
rect 1172 63032 1178 63084
rect 1230 63032 1236 63084
rect 1176 62524 1204 62552
rect 56 62368 126 62396
rect 1176 62298 1204 62326
rect 234 62222 318 62250
rect 1176 62172 1204 62200
rect 536 62102 618 62130
rect 1172 61494 1178 61546
rect 1230 61494 1236 61546
rect 536 60910 618 60938
rect 1176 60840 1204 60868
rect 234 60790 318 60818
rect 1176 60714 1204 60742
rect 56 60644 126 60672
rect 1176 60488 1204 60516
rect 1172 59956 1178 60008
rect 1230 59956 1236 60008
rect 1176 59448 1204 59476
rect 56 59292 126 59320
rect 1176 59222 1204 59250
rect 234 59146 318 59174
rect 1176 59096 1204 59124
rect 536 59026 618 59054
rect 1172 58418 1178 58470
rect 1230 58418 1236 58470
rect 536 57834 618 57862
rect 1176 57764 1204 57792
rect 234 57714 318 57742
rect 1176 57638 1204 57666
rect 56 57568 126 57596
rect 1176 57412 1204 57440
rect 1172 56880 1178 56932
rect 1230 56880 1236 56932
rect 1176 56372 1204 56400
rect 56 56216 126 56244
rect 1176 56146 1204 56174
rect 234 56070 318 56098
rect 1176 56020 1204 56048
rect 536 55950 618 55978
rect 1172 55342 1178 55394
rect 1230 55342 1236 55394
rect 536 54758 618 54786
rect 1176 54688 1204 54716
rect 234 54638 318 54666
rect 1176 54562 1204 54590
rect 56 54492 126 54520
rect 1176 54336 1204 54364
rect 1172 53804 1178 53856
rect 1230 53804 1236 53856
rect 1176 53296 1204 53324
rect 56 53140 126 53168
rect 1176 53070 1204 53098
rect 234 52994 318 53022
rect 1176 52944 1204 52972
rect 536 52874 618 52902
rect 1172 52266 1178 52318
rect 1230 52266 1236 52318
rect 536 51682 618 51710
rect 1176 51612 1204 51640
rect 234 51562 318 51590
rect 1176 51486 1204 51514
rect 56 51416 126 51444
rect 1176 51260 1204 51288
rect 1172 50728 1178 50780
rect 1230 50728 1236 50780
rect 1176 50220 1204 50248
rect 56 50064 126 50092
rect 1176 49994 1204 50022
rect 234 49918 318 49946
rect 1176 49868 1204 49896
rect 536 49798 618 49826
rect 1172 49190 1178 49242
rect 1230 49190 1236 49242
rect 536 48606 618 48634
rect 1176 48536 1204 48564
rect 234 48486 318 48514
rect 1176 48410 1204 48438
rect 56 48340 126 48368
rect 1176 48184 1204 48212
rect 1172 47652 1178 47704
rect 1230 47652 1236 47704
rect 1176 47144 1204 47172
rect 56 46988 126 47016
rect 1176 46918 1204 46946
rect 234 46842 318 46870
rect 1176 46792 1204 46820
rect 536 46722 618 46750
rect 1172 46114 1178 46166
rect 1230 46114 1236 46166
rect 536 45530 618 45558
rect 1176 45460 1204 45488
rect 234 45410 318 45438
rect 1176 45334 1204 45362
rect 56 45264 126 45292
rect 1176 45108 1204 45136
rect 1172 44576 1178 44628
rect 1230 44576 1236 44628
rect 1176 44068 1204 44096
rect 56 43912 126 43940
rect 1176 43842 1204 43870
rect 234 43766 318 43794
rect 1176 43716 1204 43744
rect 536 43646 618 43674
rect 1172 43038 1178 43090
rect 1230 43038 1236 43090
rect 536 42454 618 42482
rect 1176 42384 1204 42412
rect 234 42334 318 42362
rect 1176 42258 1204 42286
rect 56 42188 126 42216
rect 1176 42032 1204 42060
rect 1172 41500 1178 41552
rect 1230 41500 1236 41552
rect 1176 40992 1204 41020
rect 56 40836 126 40864
rect 1176 40766 1204 40794
rect 234 40690 318 40718
rect 1176 40640 1204 40668
rect 536 40570 618 40598
rect 1172 39962 1178 40014
rect 1230 39962 1236 40014
rect 536 39378 618 39406
rect 1176 39308 1204 39336
rect 234 39258 318 39286
rect 1176 39182 1204 39210
rect 56 39112 126 39140
rect 1176 38956 1204 38984
rect 1172 38424 1178 38476
rect 1230 38424 1236 38476
rect 1176 37916 1204 37944
rect 56 37760 126 37788
rect 1176 37690 1204 37718
rect 234 37614 318 37642
rect 1176 37564 1204 37592
rect 536 37494 618 37522
rect 1172 36886 1178 36938
rect 1230 36886 1236 36938
rect 536 36302 618 36330
rect 1176 36232 1204 36260
rect 234 36182 318 36210
rect 1176 36106 1204 36134
rect 56 36036 126 36064
rect 1176 35880 1204 35908
rect 1172 35348 1178 35400
rect 1230 35348 1236 35400
rect 1176 34840 1204 34868
rect 56 34684 126 34712
rect 1176 34614 1204 34642
rect 234 34538 318 34566
rect 1176 34488 1204 34516
rect 536 34418 618 34446
rect 1172 33810 1178 33862
rect 1230 33810 1236 33862
rect 536 33226 618 33254
rect 1176 33156 1204 33184
rect 234 33106 318 33134
rect 1176 33030 1204 33058
rect 56 32960 126 32988
rect 1176 32804 1204 32832
rect 1172 32272 1178 32324
rect 1230 32272 1236 32324
rect 1176 31764 1204 31792
rect 56 31608 126 31636
rect 1176 31538 1204 31566
rect 234 31462 318 31490
rect 1176 31412 1204 31440
rect 536 31342 618 31370
rect 1172 30734 1178 30786
rect 1230 30734 1236 30786
rect 536 30150 618 30178
rect 1176 30080 1204 30108
rect 234 30030 318 30058
rect 1176 29954 1204 29982
rect 56 29884 126 29912
rect 1176 29728 1204 29756
rect 1172 29196 1178 29248
rect 1230 29196 1236 29248
rect 1176 28688 1204 28716
rect 56 28532 126 28560
rect 1176 28462 1204 28490
rect 234 28386 318 28414
rect 1176 28336 1204 28364
rect 536 28266 618 28294
rect 1172 27658 1178 27710
rect 1230 27658 1236 27710
rect 536 27074 618 27102
rect 1176 27004 1204 27032
rect 234 26954 318 26982
rect 1176 26878 1204 26906
rect 56 26808 126 26836
rect 1176 26652 1204 26680
rect 1172 26120 1178 26172
rect 1230 26120 1236 26172
rect 1176 25612 1204 25640
rect 56 25456 126 25484
rect 1176 25386 1204 25414
rect 234 25310 318 25338
rect 1176 25260 1204 25288
rect 536 25190 618 25218
rect 1172 24582 1178 24634
rect 1230 24582 1236 24634
rect 536 23998 618 24026
rect 1176 23928 1204 23956
rect 234 23878 318 23906
rect 1176 23802 1204 23830
rect 56 23732 126 23760
rect 1176 23576 1204 23604
rect 1172 23044 1178 23096
rect 1230 23044 1236 23096
rect 1176 22536 1204 22564
rect 56 22380 126 22408
rect 1176 22310 1204 22338
rect 234 22234 318 22262
rect 1176 22184 1204 22212
rect 536 22114 618 22142
rect 1172 21506 1178 21558
rect 1230 21506 1236 21558
rect 536 20922 618 20950
rect 1176 20852 1204 20880
rect 234 20802 318 20830
rect 1176 20726 1204 20754
rect 56 20656 126 20684
rect 1176 20500 1204 20528
rect 1172 19968 1178 20020
rect 1230 19968 1236 20020
rect 1176 19460 1204 19488
rect 56 19304 126 19332
rect 1176 19234 1204 19262
rect 234 19158 318 19186
rect 1176 19108 1204 19136
rect 536 19038 618 19066
rect 1172 18430 1178 18482
rect 1230 18430 1236 18482
rect 536 17846 618 17874
rect 1176 17776 1204 17804
rect 234 17726 318 17754
rect 1176 17650 1204 17678
rect 56 17580 126 17608
rect 1176 17424 1204 17452
rect 1172 16892 1178 16944
rect 1230 16892 1236 16944
rect 1176 16384 1204 16412
rect 56 16228 126 16256
rect 1176 16158 1204 16186
rect 234 16082 318 16110
rect 1176 16032 1204 16060
rect 536 15962 618 15990
rect 1172 15354 1178 15406
rect 1230 15354 1236 15406
rect 536 14770 618 14798
rect 1176 14700 1204 14728
rect 234 14650 318 14678
rect 1176 14574 1204 14602
rect 56 14504 126 14532
rect 1176 14348 1204 14376
rect 1172 13816 1178 13868
rect 1230 13816 1236 13868
rect 1176 13308 1204 13336
rect 56 13152 126 13180
rect 1176 13082 1204 13110
rect 234 13006 318 13034
rect 1176 12956 1204 12984
rect 536 12886 618 12914
rect 1172 12278 1178 12330
rect 1230 12278 1236 12330
rect 536 11694 618 11722
rect 1176 11624 1204 11652
rect 234 11574 318 11602
rect 1176 11498 1204 11526
rect 56 11428 126 11456
rect 1176 11272 1204 11300
rect 1172 10740 1178 10792
rect 1230 10740 1236 10792
rect 1176 10232 1204 10260
rect 56 10076 126 10104
rect 1176 10006 1204 10034
rect 234 9930 318 9958
rect 1176 9880 1204 9908
rect 536 9810 618 9838
rect 1172 9202 1178 9254
rect 1230 9202 1236 9254
rect 536 8618 618 8646
rect 1176 8548 1204 8576
rect 234 8498 318 8526
rect 1176 8422 1204 8450
rect 56 8352 126 8380
rect 1176 8196 1204 8224
rect 1172 7664 1178 7716
rect 1230 7664 1236 7716
rect 1176 7156 1204 7184
rect 56 7000 126 7028
rect 1176 6930 1204 6958
rect 234 6854 318 6882
rect 1176 6804 1204 6832
rect 536 6734 618 6762
rect 1172 6126 1178 6178
rect 1230 6126 1236 6178
rect 536 5542 618 5570
rect 1176 5472 1204 5500
rect 234 5422 318 5450
rect 1176 5346 1204 5374
rect 56 5276 126 5304
rect 1176 5120 1204 5148
rect 1172 4588 1178 4640
rect 1230 4588 1236 4640
rect 1176 4080 1204 4108
rect 56 3924 126 3952
rect 1176 3854 1204 3882
rect 234 3778 318 3806
rect 1176 3728 1204 3756
rect 536 3658 618 3686
rect 1172 3050 1178 3102
rect 1230 3050 1236 3102
rect 536 2466 618 2494
rect 1176 2396 1204 2424
rect 234 2346 318 2374
rect 1176 2270 1204 2298
rect 56 2200 126 2228
rect 1176 2044 1204 2072
rect 1172 1512 1178 1564
rect 1230 1512 1236 1564
rect 1176 1004 1204 1032
rect 56 848 126 876
rect 1176 778 1204 806
rect 234 702 318 730
rect 1176 652 1204 680
rect 536 582 618 610
rect 1172 -26 1178 26
rect 1230 -26 1236 26
<< via1 >>
rect 1178 98406 1230 98458
rect 1178 96868 1230 96920
rect 1178 95330 1230 95382
rect 1178 93792 1230 93844
rect 1178 92254 1230 92306
rect 1178 90716 1230 90768
rect 1178 89178 1230 89230
rect 1178 87640 1230 87692
rect 1178 86102 1230 86154
rect 1178 84564 1230 84616
rect 1178 83026 1230 83078
rect 1178 81488 1230 81540
rect 1178 79950 1230 80002
rect 1178 78412 1230 78464
rect 1178 76874 1230 76926
rect 1178 75336 1230 75388
rect 1178 73798 1230 73850
rect 1178 72260 1230 72312
rect 1178 70722 1230 70774
rect 1178 69184 1230 69236
rect 1178 67646 1230 67698
rect 1178 66108 1230 66160
rect 1178 64570 1230 64622
rect 1178 63032 1230 63084
rect 1178 61494 1230 61546
rect 1178 59956 1230 60008
rect 1178 58418 1230 58470
rect 1178 56880 1230 56932
rect 1178 55342 1230 55394
rect 1178 53804 1230 53856
rect 1178 52266 1230 52318
rect 1178 50728 1230 50780
rect 1178 49190 1230 49242
rect 1178 47652 1230 47704
rect 1178 46114 1230 46166
rect 1178 44576 1230 44628
rect 1178 43038 1230 43090
rect 1178 41500 1230 41552
rect 1178 39962 1230 40014
rect 1178 38424 1230 38476
rect 1178 36886 1230 36938
rect 1178 35348 1230 35400
rect 1178 33810 1230 33862
rect 1178 32272 1230 32324
rect 1178 30734 1230 30786
rect 1178 29196 1230 29248
rect 1178 27658 1230 27710
rect 1178 26120 1230 26172
rect 1178 24582 1230 24634
rect 1178 23044 1230 23096
rect 1178 21506 1230 21558
rect 1178 19968 1230 20020
rect 1178 18430 1230 18482
rect 1178 16892 1230 16944
rect 1178 15354 1230 15406
rect 1178 13816 1230 13868
rect 1178 12278 1230 12330
rect 1178 10740 1230 10792
rect 1178 9202 1230 9254
rect 1178 7664 1230 7716
rect 1178 6126 1230 6178
rect 1178 4588 1230 4640
rect 1178 3050 1230 3102
rect 1178 1512 1230 1564
rect 1178 -26 1230 26
<< metal2 >>
rect 1176 98460 1232 98469
rect 0 0 28 98432
rect 1176 98395 1232 98404
rect 192 97724 220 97752
rect 1176 96922 1232 96931
rect 1176 96857 1232 96866
rect 192 96036 220 96064
rect 1176 95384 1232 95393
rect 1176 95319 1232 95328
rect 192 94648 220 94676
rect 1176 93846 1232 93855
rect 1176 93781 1232 93790
rect 192 92960 220 92988
rect 1176 92308 1232 92317
rect 1176 92243 1232 92252
rect 192 91572 220 91600
rect 1176 90770 1232 90779
rect 1176 90705 1232 90714
rect 192 89884 220 89912
rect 1176 89232 1232 89241
rect 1176 89167 1232 89176
rect 192 88496 220 88524
rect 1176 87694 1232 87703
rect 1176 87629 1232 87638
rect 192 86808 220 86836
rect 1176 86156 1232 86165
rect 1176 86091 1232 86100
rect 192 85420 220 85448
rect 1176 84618 1232 84627
rect 1176 84553 1232 84562
rect 192 83732 220 83760
rect 1176 83080 1232 83089
rect 1176 83015 1232 83024
rect 192 82344 220 82372
rect 1176 81542 1232 81551
rect 1176 81477 1232 81486
rect 192 80656 220 80684
rect 1176 80004 1232 80013
rect 1176 79939 1232 79948
rect 192 79268 220 79296
rect 1176 78466 1232 78475
rect 1176 78401 1232 78410
rect 192 77580 220 77608
rect 1176 76928 1232 76937
rect 1176 76863 1232 76872
rect 192 76192 220 76220
rect 1176 75390 1232 75399
rect 1176 75325 1232 75334
rect 192 74504 220 74532
rect 1176 73852 1232 73861
rect 1176 73787 1232 73796
rect 192 73116 220 73144
rect 1176 72314 1232 72323
rect 1176 72249 1232 72258
rect 192 71428 220 71456
rect 1176 70776 1232 70785
rect 1176 70711 1232 70720
rect 192 70040 220 70068
rect 1176 69238 1232 69247
rect 1176 69173 1232 69182
rect 192 68352 220 68380
rect 1176 67700 1232 67709
rect 1176 67635 1232 67644
rect 192 66964 220 66992
rect 1176 66162 1232 66171
rect 1176 66097 1232 66106
rect 192 65276 220 65304
rect 1176 64624 1232 64633
rect 1176 64559 1232 64568
rect 192 63888 220 63916
rect 1176 63086 1232 63095
rect 1176 63021 1232 63030
rect 192 62200 220 62228
rect 1176 61548 1232 61557
rect 1176 61483 1232 61492
rect 192 60812 220 60840
rect 1176 60010 1232 60019
rect 1176 59945 1232 59954
rect 192 59124 220 59152
rect 1176 58472 1232 58481
rect 1176 58407 1232 58416
rect 192 57736 220 57764
rect 1176 56934 1232 56943
rect 1176 56869 1232 56878
rect 192 56048 220 56076
rect 1176 55396 1232 55405
rect 1176 55331 1232 55340
rect 192 54660 220 54688
rect 1176 53858 1232 53867
rect 1176 53793 1232 53802
rect 192 52972 220 53000
rect 1176 52320 1232 52329
rect 1176 52255 1232 52264
rect 192 51584 220 51612
rect 1176 50782 1232 50791
rect 1176 50717 1232 50726
rect 192 49896 220 49924
rect 1176 49244 1232 49253
rect 1176 49179 1232 49188
rect 192 48508 220 48536
rect 1176 47706 1232 47715
rect 1176 47641 1232 47650
rect 192 46820 220 46848
rect 1176 46168 1232 46177
rect 1176 46103 1232 46112
rect 192 45432 220 45460
rect 1176 44630 1232 44639
rect 1176 44565 1232 44574
rect 192 43744 220 43772
rect 1176 43092 1232 43101
rect 1176 43027 1232 43036
rect 192 42356 220 42384
rect 1176 41554 1232 41563
rect 1176 41489 1232 41498
rect 192 40668 220 40696
rect 1176 40016 1232 40025
rect 1176 39951 1232 39960
rect 192 39280 220 39308
rect 1176 38478 1232 38487
rect 1176 38413 1232 38422
rect 192 37592 220 37620
rect 1176 36940 1232 36949
rect 1176 36875 1232 36884
rect 192 36204 220 36232
rect 1176 35402 1232 35411
rect 1176 35337 1232 35346
rect 192 34516 220 34544
rect 1176 33864 1232 33873
rect 1176 33799 1232 33808
rect 192 33128 220 33156
rect 1176 32326 1232 32335
rect 1176 32261 1232 32270
rect 192 31440 220 31468
rect 1176 30788 1232 30797
rect 1176 30723 1232 30732
rect 192 30052 220 30080
rect 1176 29250 1232 29259
rect 1176 29185 1232 29194
rect 192 28364 220 28392
rect 1176 27712 1232 27721
rect 1176 27647 1232 27656
rect 192 26976 220 27004
rect 1176 26174 1232 26183
rect 1176 26109 1232 26118
rect 192 25288 220 25316
rect 1176 24636 1232 24645
rect 1176 24571 1232 24580
rect 192 23900 220 23928
rect 1176 23098 1232 23107
rect 1176 23033 1232 23042
rect 192 22212 220 22240
rect 1176 21560 1232 21569
rect 1176 21495 1232 21504
rect 192 20824 220 20852
rect 1176 20022 1232 20031
rect 1176 19957 1232 19966
rect 192 19136 220 19164
rect 1176 18484 1232 18493
rect 1176 18419 1232 18428
rect 192 17748 220 17776
rect 1176 16946 1232 16955
rect 1176 16881 1232 16890
rect 192 16060 220 16088
rect 1176 15408 1232 15417
rect 1176 15343 1232 15352
rect 192 14672 220 14700
rect 1176 13870 1232 13879
rect 1176 13805 1232 13814
rect 192 12984 220 13012
rect 1176 12332 1232 12341
rect 1176 12267 1232 12276
rect 192 11596 220 11624
rect 1176 10794 1232 10803
rect 1176 10729 1232 10738
rect 192 9908 220 9936
rect 1176 9256 1232 9265
rect 1176 9191 1232 9200
rect 192 8520 220 8548
rect 1176 7718 1232 7727
rect 1176 7653 1232 7662
rect 192 6832 220 6860
rect 1176 6180 1232 6189
rect 1176 6115 1232 6124
rect 192 5444 220 5472
rect 1176 4642 1232 4651
rect 1176 4577 1232 4586
rect 192 3756 220 3784
rect 1176 3104 1232 3113
rect 1176 3039 1232 3048
rect 192 2368 220 2396
rect 1176 1566 1232 1575
rect 1176 1501 1232 1510
rect 192 680 220 708
rect 1176 28 1232 37
rect 1176 -37 1232 -28
<< via2 >>
rect 1176 98458 1232 98460
rect 1176 98406 1178 98458
rect 1178 98406 1230 98458
rect 1230 98406 1232 98458
rect 1176 98404 1232 98406
rect 1176 96920 1232 96922
rect 1176 96868 1178 96920
rect 1178 96868 1230 96920
rect 1230 96868 1232 96920
rect 1176 96866 1232 96868
rect 1176 95382 1232 95384
rect 1176 95330 1178 95382
rect 1178 95330 1230 95382
rect 1230 95330 1232 95382
rect 1176 95328 1232 95330
rect 1176 93844 1232 93846
rect 1176 93792 1178 93844
rect 1178 93792 1230 93844
rect 1230 93792 1232 93844
rect 1176 93790 1232 93792
rect 1176 92306 1232 92308
rect 1176 92254 1178 92306
rect 1178 92254 1230 92306
rect 1230 92254 1232 92306
rect 1176 92252 1232 92254
rect 1176 90768 1232 90770
rect 1176 90716 1178 90768
rect 1178 90716 1230 90768
rect 1230 90716 1232 90768
rect 1176 90714 1232 90716
rect 1176 89230 1232 89232
rect 1176 89178 1178 89230
rect 1178 89178 1230 89230
rect 1230 89178 1232 89230
rect 1176 89176 1232 89178
rect 1176 87692 1232 87694
rect 1176 87640 1178 87692
rect 1178 87640 1230 87692
rect 1230 87640 1232 87692
rect 1176 87638 1232 87640
rect 1176 86154 1232 86156
rect 1176 86102 1178 86154
rect 1178 86102 1230 86154
rect 1230 86102 1232 86154
rect 1176 86100 1232 86102
rect 1176 84616 1232 84618
rect 1176 84564 1178 84616
rect 1178 84564 1230 84616
rect 1230 84564 1232 84616
rect 1176 84562 1232 84564
rect 1176 83078 1232 83080
rect 1176 83026 1178 83078
rect 1178 83026 1230 83078
rect 1230 83026 1232 83078
rect 1176 83024 1232 83026
rect 1176 81540 1232 81542
rect 1176 81488 1178 81540
rect 1178 81488 1230 81540
rect 1230 81488 1232 81540
rect 1176 81486 1232 81488
rect 1176 80002 1232 80004
rect 1176 79950 1178 80002
rect 1178 79950 1230 80002
rect 1230 79950 1232 80002
rect 1176 79948 1232 79950
rect 1176 78464 1232 78466
rect 1176 78412 1178 78464
rect 1178 78412 1230 78464
rect 1230 78412 1232 78464
rect 1176 78410 1232 78412
rect 1176 76926 1232 76928
rect 1176 76874 1178 76926
rect 1178 76874 1230 76926
rect 1230 76874 1232 76926
rect 1176 76872 1232 76874
rect 1176 75388 1232 75390
rect 1176 75336 1178 75388
rect 1178 75336 1230 75388
rect 1230 75336 1232 75388
rect 1176 75334 1232 75336
rect 1176 73850 1232 73852
rect 1176 73798 1178 73850
rect 1178 73798 1230 73850
rect 1230 73798 1232 73850
rect 1176 73796 1232 73798
rect 1176 72312 1232 72314
rect 1176 72260 1178 72312
rect 1178 72260 1230 72312
rect 1230 72260 1232 72312
rect 1176 72258 1232 72260
rect 1176 70774 1232 70776
rect 1176 70722 1178 70774
rect 1178 70722 1230 70774
rect 1230 70722 1232 70774
rect 1176 70720 1232 70722
rect 1176 69236 1232 69238
rect 1176 69184 1178 69236
rect 1178 69184 1230 69236
rect 1230 69184 1232 69236
rect 1176 69182 1232 69184
rect 1176 67698 1232 67700
rect 1176 67646 1178 67698
rect 1178 67646 1230 67698
rect 1230 67646 1232 67698
rect 1176 67644 1232 67646
rect 1176 66160 1232 66162
rect 1176 66108 1178 66160
rect 1178 66108 1230 66160
rect 1230 66108 1232 66160
rect 1176 66106 1232 66108
rect 1176 64622 1232 64624
rect 1176 64570 1178 64622
rect 1178 64570 1230 64622
rect 1230 64570 1232 64622
rect 1176 64568 1232 64570
rect 1176 63084 1232 63086
rect 1176 63032 1178 63084
rect 1178 63032 1230 63084
rect 1230 63032 1232 63084
rect 1176 63030 1232 63032
rect 1176 61546 1232 61548
rect 1176 61494 1178 61546
rect 1178 61494 1230 61546
rect 1230 61494 1232 61546
rect 1176 61492 1232 61494
rect 1176 60008 1232 60010
rect 1176 59956 1178 60008
rect 1178 59956 1230 60008
rect 1230 59956 1232 60008
rect 1176 59954 1232 59956
rect 1176 58470 1232 58472
rect 1176 58418 1178 58470
rect 1178 58418 1230 58470
rect 1230 58418 1232 58470
rect 1176 58416 1232 58418
rect 1176 56932 1232 56934
rect 1176 56880 1178 56932
rect 1178 56880 1230 56932
rect 1230 56880 1232 56932
rect 1176 56878 1232 56880
rect 1176 55394 1232 55396
rect 1176 55342 1178 55394
rect 1178 55342 1230 55394
rect 1230 55342 1232 55394
rect 1176 55340 1232 55342
rect 1176 53856 1232 53858
rect 1176 53804 1178 53856
rect 1178 53804 1230 53856
rect 1230 53804 1232 53856
rect 1176 53802 1232 53804
rect 1176 52318 1232 52320
rect 1176 52266 1178 52318
rect 1178 52266 1230 52318
rect 1230 52266 1232 52318
rect 1176 52264 1232 52266
rect 1176 50780 1232 50782
rect 1176 50728 1178 50780
rect 1178 50728 1230 50780
rect 1230 50728 1232 50780
rect 1176 50726 1232 50728
rect 1176 49242 1232 49244
rect 1176 49190 1178 49242
rect 1178 49190 1230 49242
rect 1230 49190 1232 49242
rect 1176 49188 1232 49190
rect 1176 47704 1232 47706
rect 1176 47652 1178 47704
rect 1178 47652 1230 47704
rect 1230 47652 1232 47704
rect 1176 47650 1232 47652
rect 1176 46166 1232 46168
rect 1176 46114 1178 46166
rect 1178 46114 1230 46166
rect 1230 46114 1232 46166
rect 1176 46112 1232 46114
rect 1176 44628 1232 44630
rect 1176 44576 1178 44628
rect 1178 44576 1230 44628
rect 1230 44576 1232 44628
rect 1176 44574 1232 44576
rect 1176 43090 1232 43092
rect 1176 43038 1178 43090
rect 1178 43038 1230 43090
rect 1230 43038 1232 43090
rect 1176 43036 1232 43038
rect 1176 41552 1232 41554
rect 1176 41500 1178 41552
rect 1178 41500 1230 41552
rect 1230 41500 1232 41552
rect 1176 41498 1232 41500
rect 1176 40014 1232 40016
rect 1176 39962 1178 40014
rect 1178 39962 1230 40014
rect 1230 39962 1232 40014
rect 1176 39960 1232 39962
rect 1176 38476 1232 38478
rect 1176 38424 1178 38476
rect 1178 38424 1230 38476
rect 1230 38424 1232 38476
rect 1176 38422 1232 38424
rect 1176 36938 1232 36940
rect 1176 36886 1178 36938
rect 1178 36886 1230 36938
rect 1230 36886 1232 36938
rect 1176 36884 1232 36886
rect 1176 35400 1232 35402
rect 1176 35348 1178 35400
rect 1178 35348 1230 35400
rect 1230 35348 1232 35400
rect 1176 35346 1232 35348
rect 1176 33862 1232 33864
rect 1176 33810 1178 33862
rect 1178 33810 1230 33862
rect 1230 33810 1232 33862
rect 1176 33808 1232 33810
rect 1176 32324 1232 32326
rect 1176 32272 1178 32324
rect 1178 32272 1230 32324
rect 1230 32272 1232 32324
rect 1176 32270 1232 32272
rect 1176 30786 1232 30788
rect 1176 30734 1178 30786
rect 1178 30734 1230 30786
rect 1230 30734 1232 30786
rect 1176 30732 1232 30734
rect 1176 29248 1232 29250
rect 1176 29196 1178 29248
rect 1178 29196 1230 29248
rect 1230 29196 1232 29248
rect 1176 29194 1232 29196
rect 1176 27710 1232 27712
rect 1176 27658 1178 27710
rect 1178 27658 1230 27710
rect 1230 27658 1232 27710
rect 1176 27656 1232 27658
rect 1176 26172 1232 26174
rect 1176 26120 1178 26172
rect 1178 26120 1230 26172
rect 1230 26120 1232 26172
rect 1176 26118 1232 26120
rect 1176 24634 1232 24636
rect 1176 24582 1178 24634
rect 1178 24582 1230 24634
rect 1230 24582 1232 24634
rect 1176 24580 1232 24582
rect 1176 23096 1232 23098
rect 1176 23044 1178 23096
rect 1178 23044 1230 23096
rect 1230 23044 1232 23096
rect 1176 23042 1232 23044
rect 1176 21558 1232 21560
rect 1176 21506 1178 21558
rect 1178 21506 1230 21558
rect 1230 21506 1232 21558
rect 1176 21504 1232 21506
rect 1176 20020 1232 20022
rect 1176 19968 1178 20020
rect 1178 19968 1230 20020
rect 1230 19968 1232 20020
rect 1176 19966 1232 19968
rect 1176 18482 1232 18484
rect 1176 18430 1178 18482
rect 1178 18430 1230 18482
rect 1230 18430 1232 18482
rect 1176 18428 1232 18430
rect 1176 16944 1232 16946
rect 1176 16892 1178 16944
rect 1178 16892 1230 16944
rect 1230 16892 1232 16944
rect 1176 16890 1232 16892
rect 1176 15406 1232 15408
rect 1176 15354 1178 15406
rect 1178 15354 1230 15406
rect 1230 15354 1232 15406
rect 1176 15352 1232 15354
rect 1176 13868 1232 13870
rect 1176 13816 1178 13868
rect 1178 13816 1230 13868
rect 1230 13816 1232 13868
rect 1176 13814 1232 13816
rect 1176 12330 1232 12332
rect 1176 12278 1178 12330
rect 1178 12278 1230 12330
rect 1230 12278 1232 12330
rect 1176 12276 1232 12278
rect 1176 10792 1232 10794
rect 1176 10740 1178 10792
rect 1178 10740 1230 10792
rect 1230 10740 1232 10792
rect 1176 10738 1232 10740
rect 1176 9254 1232 9256
rect 1176 9202 1178 9254
rect 1178 9202 1230 9254
rect 1230 9202 1232 9254
rect 1176 9200 1232 9202
rect 1176 7716 1232 7718
rect 1176 7664 1178 7716
rect 1178 7664 1230 7716
rect 1230 7664 1232 7716
rect 1176 7662 1232 7664
rect 1176 6178 1232 6180
rect 1176 6126 1178 6178
rect 1178 6126 1230 6178
rect 1230 6126 1232 6178
rect 1176 6124 1232 6126
rect 1176 4640 1232 4642
rect 1176 4588 1178 4640
rect 1178 4588 1230 4640
rect 1230 4588 1232 4640
rect 1176 4586 1232 4588
rect 1176 3102 1232 3104
rect 1176 3050 1178 3102
rect 1178 3050 1230 3102
rect 1230 3050 1232 3102
rect 1176 3048 1232 3050
rect 1176 1564 1232 1566
rect 1176 1512 1178 1564
rect 1178 1512 1230 1564
rect 1230 1512 1232 1564
rect 1176 1510 1232 1512
rect 1176 26 1232 28
rect 1176 -26 1178 26
rect 1178 -26 1230 26
rect 1230 -26 1232 26
rect 1176 -28 1232 -26
<< metal3 >>
rect 1138 98460 1270 98469
rect 1138 98404 1176 98460
rect 1232 98404 1270 98460
rect 1138 98395 1270 98404
rect 1138 96922 1270 96931
rect 1138 96866 1176 96922
rect 1232 96866 1270 96922
rect 1138 96857 1270 96866
rect 1138 95384 1270 95393
rect 1138 95328 1176 95384
rect 1232 95328 1270 95384
rect 1138 95319 1270 95328
rect 1138 93846 1270 93855
rect 1138 93790 1176 93846
rect 1232 93790 1270 93846
rect 1138 93781 1270 93790
rect 1138 92308 1270 92317
rect 1138 92252 1176 92308
rect 1232 92252 1270 92308
rect 1138 92243 1270 92252
rect 1138 90770 1270 90779
rect 1138 90714 1176 90770
rect 1232 90714 1270 90770
rect 1138 90705 1270 90714
rect 1138 89232 1270 89241
rect 1138 89176 1176 89232
rect 1232 89176 1270 89232
rect 1138 89167 1270 89176
rect 1138 87694 1270 87703
rect 1138 87638 1176 87694
rect 1232 87638 1270 87694
rect 1138 87629 1270 87638
rect 1138 86156 1270 86165
rect 1138 86100 1176 86156
rect 1232 86100 1270 86156
rect 1138 86091 1270 86100
rect 1138 84618 1270 84627
rect 1138 84562 1176 84618
rect 1232 84562 1270 84618
rect 1138 84553 1270 84562
rect 1138 83080 1270 83089
rect 1138 83024 1176 83080
rect 1232 83024 1270 83080
rect 1138 83015 1270 83024
rect 1138 81542 1270 81551
rect 1138 81486 1176 81542
rect 1232 81486 1270 81542
rect 1138 81477 1270 81486
rect 1138 80004 1270 80013
rect 1138 79948 1176 80004
rect 1232 79948 1270 80004
rect 1138 79939 1270 79948
rect 1138 78466 1270 78475
rect 1138 78410 1176 78466
rect 1232 78410 1270 78466
rect 1138 78401 1270 78410
rect 1138 76928 1270 76937
rect 1138 76872 1176 76928
rect 1232 76872 1270 76928
rect 1138 76863 1270 76872
rect 1138 75390 1270 75399
rect 1138 75334 1176 75390
rect 1232 75334 1270 75390
rect 1138 75325 1270 75334
rect 1138 73852 1270 73861
rect 1138 73796 1176 73852
rect 1232 73796 1270 73852
rect 1138 73787 1270 73796
rect 1138 72314 1270 72323
rect 1138 72258 1176 72314
rect 1232 72258 1270 72314
rect 1138 72249 1270 72258
rect 1138 70776 1270 70785
rect 1138 70720 1176 70776
rect 1232 70720 1270 70776
rect 1138 70711 1270 70720
rect 1138 69238 1270 69247
rect 1138 69182 1176 69238
rect 1232 69182 1270 69238
rect 1138 69173 1270 69182
rect 1138 67700 1270 67709
rect 1138 67644 1176 67700
rect 1232 67644 1270 67700
rect 1138 67635 1270 67644
rect 1138 66162 1270 66171
rect 1138 66106 1176 66162
rect 1232 66106 1270 66162
rect 1138 66097 1270 66106
rect 1138 64624 1270 64633
rect 1138 64568 1176 64624
rect 1232 64568 1270 64624
rect 1138 64559 1270 64568
rect 1138 63086 1270 63095
rect 1138 63030 1176 63086
rect 1232 63030 1270 63086
rect 1138 63021 1270 63030
rect 1138 61548 1270 61557
rect 1138 61492 1176 61548
rect 1232 61492 1270 61548
rect 1138 61483 1270 61492
rect 1138 60010 1270 60019
rect 1138 59954 1176 60010
rect 1232 59954 1270 60010
rect 1138 59945 1270 59954
rect 1138 58472 1270 58481
rect 1138 58416 1176 58472
rect 1232 58416 1270 58472
rect 1138 58407 1270 58416
rect 1138 56934 1270 56943
rect 1138 56878 1176 56934
rect 1232 56878 1270 56934
rect 1138 56869 1270 56878
rect 1138 55396 1270 55405
rect 1138 55340 1176 55396
rect 1232 55340 1270 55396
rect 1138 55331 1270 55340
rect 1138 53858 1270 53867
rect 1138 53802 1176 53858
rect 1232 53802 1270 53858
rect 1138 53793 1270 53802
rect 1138 52320 1270 52329
rect 1138 52264 1176 52320
rect 1232 52264 1270 52320
rect 1138 52255 1270 52264
rect 1138 50782 1270 50791
rect 1138 50726 1176 50782
rect 1232 50726 1270 50782
rect 1138 50717 1270 50726
rect 1138 49244 1270 49253
rect 1138 49188 1176 49244
rect 1232 49188 1270 49244
rect 1138 49179 1270 49188
rect 1138 47706 1270 47715
rect 1138 47650 1176 47706
rect 1232 47650 1270 47706
rect 1138 47641 1270 47650
rect 1138 46168 1270 46177
rect 1138 46112 1176 46168
rect 1232 46112 1270 46168
rect 1138 46103 1270 46112
rect 1138 44630 1270 44639
rect 1138 44574 1176 44630
rect 1232 44574 1270 44630
rect 1138 44565 1270 44574
rect 1138 43092 1270 43101
rect 1138 43036 1176 43092
rect 1232 43036 1270 43092
rect 1138 43027 1270 43036
rect 1138 41554 1270 41563
rect 1138 41498 1176 41554
rect 1232 41498 1270 41554
rect 1138 41489 1270 41498
rect 1138 40016 1270 40025
rect 1138 39960 1176 40016
rect 1232 39960 1270 40016
rect 1138 39951 1270 39960
rect 1138 38478 1270 38487
rect 1138 38422 1176 38478
rect 1232 38422 1270 38478
rect 1138 38413 1270 38422
rect 1138 36940 1270 36949
rect 1138 36884 1176 36940
rect 1232 36884 1270 36940
rect 1138 36875 1270 36884
rect 1138 35402 1270 35411
rect 1138 35346 1176 35402
rect 1232 35346 1270 35402
rect 1138 35337 1270 35346
rect 1138 33864 1270 33873
rect 1138 33808 1176 33864
rect 1232 33808 1270 33864
rect 1138 33799 1270 33808
rect 1138 32326 1270 32335
rect 1138 32270 1176 32326
rect 1232 32270 1270 32326
rect 1138 32261 1270 32270
rect 1138 30788 1270 30797
rect 1138 30732 1176 30788
rect 1232 30732 1270 30788
rect 1138 30723 1270 30732
rect 1138 29250 1270 29259
rect 1138 29194 1176 29250
rect 1232 29194 1270 29250
rect 1138 29185 1270 29194
rect 1138 27712 1270 27721
rect 1138 27656 1176 27712
rect 1232 27656 1270 27712
rect 1138 27647 1270 27656
rect 1138 26174 1270 26183
rect 1138 26118 1176 26174
rect 1232 26118 1270 26174
rect 1138 26109 1270 26118
rect 1138 24636 1270 24645
rect 1138 24580 1176 24636
rect 1232 24580 1270 24636
rect 1138 24571 1270 24580
rect 1138 23098 1270 23107
rect 1138 23042 1176 23098
rect 1232 23042 1270 23098
rect 1138 23033 1270 23042
rect 1138 21560 1270 21569
rect 1138 21504 1176 21560
rect 1232 21504 1270 21560
rect 1138 21495 1270 21504
rect 1138 20022 1270 20031
rect 1138 19966 1176 20022
rect 1232 19966 1270 20022
rect 1138 19957 1270 19966
rect 1138 18484 1270 18493
rect 1138 18428 1176 18484
rect 1232 18428 1270 18484
rect 1138 18419 1270 18428
rect 1138 16946 1270 16955
rect 1138 16890 1176 16946
rect 1232 16890 1270 16946
rect 1138 16881 1270 16890
rect 1138 15408 1270 15417
rect 1138 15352 1176 15408
rect 1232 15352 1270 15408
rect 1138 15343 1270 15352
rect 1138 13870 1270 13879
rect 1138 13814 1176 13870
rect 1232 13814 1270 13870
rect 1138 13805 1270 13814
rect 1138 12332 1270 12341
rect 1138 12276 1176 12332
rect 1232 12276 1270 12332
rect 1138 12267 1270 12276
rect 1138 10794 1270 10803
rect 1138 10738 1176 10794
rect 1232 10738 1270 10794
rect 1138 10729 1270 10738
rect 1138 9256 1270 9265
rect 1138 9200 1176 9256
rect 1232 9200 1270 9256
rect 1138 9191 1270 9200
rect 1138 7718 1270 7727
rect 1138 7662 1176 7718
rect 1232 7662 1270 7718
rect 1138 7653 1270 7662
rect 1138 6180 1270 6189
rect 1138 6124 1176 6180
rect 1232 6124 1270 6180
rect 1138 6115 1270 6124
rect 1138 4642 1270 4651
rect 1138 4586 1176 4642
rect 1232 4586 1270 4642
rect 1138 4577 1270 4586
rect 1138 3104 1270 3113
rect 1138 3048 1176 3104
rect 1232 3048 1270 3104
rect 1138 3039 1270 3048
rect 1138 1566 1270 1575
rect 1138 1510 1176 1566
rect 1232 1510 1270 1566
rect 1138 1501 1270 1510
rect 1138 28 1270 37
rect 1138 -28 1176 28
rect 1232 -28 1270 28
rect 1138 -37 1270 -28
use contact_18  contact_18_0
timestamp 1644969367
transform 1 0 1138 0 1 98395
box 0 0 1 1
use contact_17  contact_17_0
timestamp 1644969367
transform 1 0 1172 0 1 98400
box 0 0 1 1
use contact_18  contact_18_1
timestamp 1644969367
transform 1 0 1138 0 1 96857
box 0 0 1 1
use contact_17  contact_17_1
timestamp 1644969367
transform 1 0 1172 0 1 96862
box 0 0 1 1
use contact_18  contact_18_2
timestamp 1644969367
transform 1 0 1138 0 1 95319
box 0 0 1 1
use contact_17  contact_17_2
timestamp 1644969367
transform 1 0 1172 0 1 95324
box 0 0 1 1
use contact_18  contact_18_3
timestamp 1644969367
transform 1 0 1138 0 1 96857
box 0 0 1 1
use contact_17  contact_17_3
timestamp 1644969367
transform 1 0 1172 0 1 96862
box 0 0 1 1
use contact_18  contact_18_4
timestamp 1644969367
transform 1 0 1138 0 1 95319
box 0 0 1 1
use contact_17  contact_17_4
timestamp 1644969367
transform 1 0 1172 0 1 95324
box 0 0 1 1
use contact_18  contact_18_5
timestamp 1644969367
transform 1 0 1138 0 1 93781
box 0 0 1 1
use contact_17  contact_17_5
timestamp 1644969367
transform 1 0 1172 0 1 93786
box 0 0 1 1
use contact_18  contact_18_6
timestamp 1644969367
transform 1 0 1138 0 1 92243
box 0 0 1 1
use contact_17  contact_17_6
timestamp 1644969367
transform 1 0 1172 0 1 92248
box 0 0 1 1
use contact_18  contact_18_7
timestamp 1644969367
transform 1 0 1138 0 1 93781
box 0 0 1 1
use contact_17  contact_17_7
timestamp 1644969367
transform 1 0 1172 0 1 93786
box 0 0 1 1
use contact_18  contact_18_8
timestamp 1644969367
transform 1 0 1138 0 1 92243
box 0 0 1 1
use contact_17  contact_17_8
timestamp 1644969367
transform 1 0 1172 0 1 92248
box 0 0 1 1
use contact_18  contact_18_9
timestamp 1644969367
transform 1 0 1138 0 1 90705
box 0 0 1 1
use contact_17  contact_17_9
timestamp 1644969367
transform 1 0 1172 0 1 90710
box 0 0 1 1
use contact_18  contact_18_10
timestamp 1644969367
transform 1 0 1138 0 1 89167
box 0 0 1 1
use contact_17  contact_17_10
timestamp 1644969367
transform 1 0 1172 0 1 89172
box 0 0 1 1
use contact_18  contact_18_11
timestamp 1644969367
transform 1 0 1138 0 1 90705
box 0 0 1 1
use contact_17  contact_17_11
timestamp 1644969367
transform 1 0 1172 0 1 90710
box 0 0 1 1
use contact_18  contact_18_12
timestamp 1644969367
transform 1 0 1138 0 1 89167
box 0 0 1 1
use contact_17  contact_17_12
timestamp 1644969367
transform 1 0 1172 0 1 89172
box 0 0 1 1
use contact_18  contact_18_13
timestamp 1644969367
transform 1 0 1138 0 1 87629
box 0 0 1 1
use contact_17  contact_17_13
timestamp 1644969367
transform 1 0 1172 0 1 87634
box 0 0 1 1
use contact_18  contact_18_14
timestamp 1644969367
transform 1 0 1138 0 1 86091
box 0 0 1 1
use contact_17  contact_17_14
timestamp 1644969367
transform 1 0 1172 0 1 86096
box 0 0 1 1
use contact_18  contact_18_15
timestamp 1644969367
transform 1 0 1138 0 1 87629
box 0 0 1 1
use contact_17  contact_17_15
timestamp 1644969367
transform 1 0 1172 0 1 87634
box 0 0 1 1
use contact_18  contact_18_16
timestamp 1644969367
transform 1 0 1138 0 1 86091
box 0 0 1 1
use contact_17  contact_17_16
timestamp 1644969367
transform 1 0 1172 0 1 86096
box 0 0 1 1
use contact_18  contact_18_17
timestamp 1644969367
transform 1 0 1138 0 1 84553
box 0 0 1 1
use contact_17  contact_17_17
timestamp 1644969367
transform 1 0 1172 0 1 84558
box 0 0 1 1
use contact_18  contact_18_18
timestamp 1644969367
transform 1 0 1138 0 1 83015
box 0 0 1 1
use contact_17  contact_17_18
timestamp 1644969367
transform 1 0 1172 0 1 83020
box 0 0 1 1
use contact_18  contact_18_19
timestamp 1644969367
transform 1 0 1138 0 1 84553
box 0 0 1 1
use contact_17  contact_17_19
timestamp 1644969367
transform 1 0 1172 0 1 84558
box 0 0 1 1
use contact_18  contact_18_20
timestamp 1644969367
transform 1 0 1138 0 1 83015
box 0 0 1 1
use contact_17  contact_17_20
timestamp 1644969367
transform 1 0 1172 0 1 83020
box 0 0 1 1
use contact_18  contact_18_21
timestamp 1644969367
transform 1 0 1138 0 1 81477
box 0 0 1 1
use contact_17  contact_17_21
timestamp 1644969367
transform 1 0 1172 0 1 81482
box 0 0 1 1
use contact_18  contact_18_22
timestamp 1644969367
transform 1 0 1138 0 1 79939
box 0 0 1 1
use contact_17  contact_17_22
timestamp 1644969367
transform 1 0 1172 0 1 79944
box 0 0 1 1
use contact_18  contact_18_23
timestamp 1644969367
transform 1 0 1138 0 1 81477
box 0 0 1 1
use contact_17  contact_17_23
timestamp 1644969367
transform 1 0 1172 0 1 81482
box 0 0 1 1
use contact_18  contact_18_24
timestamp 1644969367
transform 1 0 1138 0 1 79939
box 0 0 1 1
use contact_17  contact_17_24
timestamp 1644969367
transform 1 0 1172 0 1 79944
box 0 0 1 1
use contact_18  contact_18_25
timestamp 1644969367
transform 1 0 1138 0 1 78401
box 0 0 1 1
use contact_17  contact_17_25
timestamp 1644969367
transform 1 0 1172 0 1 78406
box 0 0 1 1
use contact_18  contact_18_26
timestamp 1644969367
transform 1 0 1138 0 1 76863
box 0 0 1 1
use contact_17  contact_17_26
timestamp 1644969367
transform 1 0 1172 0 1 76868
box 0 0 1 1
use contact_18  contact_18_27
timestamp 1644969367
transform 1 0 1138 0 1 78401
box 0 0 1 1
use contact_17  contact_17_27
timestamp 1644969367
transform 1 0 1172 0 1 78406
box 0 0 1 1
use contact_18  contact_18_28
timestamp 1644969367
transform 1 0 1138 0 1 76863
box 0 0 1 1
use contact_17  contact_17_28
timestamp 1644969367
transform 1 0 1172 0 1 76868
box 0 0 1 1
use contact_18  contact_18_29
timestamp 1644969367
transform 1 0 1138 0 1 75325
box 0 0 1 1
use contact_17  contact_17_29
timestamp 1644969367
transform 1 0 1172 0 1 75330
box 0 0 1 1
use contact_18  contact_18_30
timestamp 1644969367
transform 1 0 1138 0 1 73787
box 0 0 1 1
use contact_17  contact_17_30
timestamp 1644969367
transform 1 0 1172 0 1 73792
box 0 0 1 1
use contact_18  contact_18_31
timestamp 1644969367
transform 1 0 1138 0 1 75325
box 0 0 1 1
use contact_17  contact_17_31
timestamp 1644969367
transform 1 0 1172 0 1 75330
box 0 0 1 1
use contact_18  contact_18_32
timestamp 1644969367
transform 1 0 1138 0 1 73787
box 0 0 1 1
use contact_17  contact_17_32
timestamp 1644969367
transform 1 0 1172 0 1 73792
box 0 0 1 1
use contact_18  contact_18_33
timestamp 1644969367
transform 1 0 1138 0 1 72249
box 0 0 1 1
use contact_17  contact_17_33
timestamp 1644969367
transform 1 0 1172 0 1 72254
box 0 0 1 1
use contact_18  contact_18_34
timestamp 1644969367
transform 1 0 1138 0 1 70711
box 0 0 1 1
use contact_17  contact_17_34
timestamp 1644969367
transform 1 0 1172 0 1 70716
box 0 0 1 1
use contact_18  contact_18_35
timestamp 1644969367
transform 1 0 1138 0 1 72249
box 0 0 1 1
use contact_17  contact_17_35
timestamp 1644969367
transform 1 0 1172 0 1 72254
box 0 0 1 1
use contact_18  contact_18_36
timestamp 1644969367
transform 1 0 1138 0 1 70711
box 0 0 1 1
use contact_17  contact_17_36
timestamp 1644969367
transform 1 0 1172 0 1 70716
box 0 0 1 1
use contact_18  contact_18_37
timestamp 1644969367
transform 1 0 1138 0 1 69173
box 0 0 1 1
use contact_17  contact_17_37
timestamp 1644969367
transform 1 0 1172 0 1 69178
box 0 0 1 1
use contact_18  contact_18_38
timestamp 1644969367
transform 1 0 1138 0 1 67635
box 0 0 1 1
use contact_17  contact_17_38
timestamp 1644969367
transform 1 0 1172 0 1 67640
box 0 0 1 1
use contact_18  contact_18_39
timestamp 1644969367
transform 1 0 1138 0 1 69173
box 0 0 1 1
use contact_17  contact_17_39
timestamp 1644969367
transform 1 0 1172 0 1 69178
box 0 0 1 1
use contact_18  contact_18_40
timestamp 1644969367
transform 1 0 1138 0 1 67635
box 0 0 1 1
use contact_17  contact_17_40
timestamp 1644969367
transform 1 0 1172 0 1 67640
box 0 0 1 1
use contact_18  contact_18_41
timestamp 1644969367
transform 1 0 1138 0 1 66097
box 0 0 1 1
use contact_17  contact_17_41
timestamp 1644969367
transform 1 0 1172 0 1 66102
box 0 0 1 1
use contact_18  contact_18_42
timestamp 1644969367
transform 1 0 1138 0 1 64559
box 0 0 1 1
use contact_17  contact_17_42
timestamp 1644969367
transform 1 0 1172 0 1 64564
box 0 0 1 1
use contact_18  contact_18_43
timestamp 1644969367
transform 1 0 1138 0 1 66097
box 0 0 1 1
use contact_17  contact_17_43
timestamp 1644969367
transform 1 0 1172 0 1 66102
box 0 0 1 1
use contact_18  contact_18_44
timestamp 1644969367
transform 1 0 1138 0 1 64559
box 0 0 1 1
use contact_17  contact_17_44
timestamp 1644969367
transform 1 0 1172 0 1 64564
box 0 0 1 1
use contact_18  contact_18_45
timestamp 1644969367
transform 1 0 1138 0 1 63021
box 0 0 1 1
use contact_17  contact_17_45
timestamp 1644969367
transform 1 0 1172 0 1 63026
box 0 0 1 1
use contact_18  contact_18_46
timestamp 1644969367
transform 1 0 1138 0 1 61483
box 0 0 1 1
use contact_17  contact_17_46
timestamp 1644969367
transform 1 0 1172 0 1 61488
box 0 0 1 1
use contact_18  contact_18_47
timestamp 1644969367
transform 1 0 1138 0 1 63021
box 0 0 1 1
use contact_17  contact_17_47
timestamp 1644969367
transform 1 0 1172 0 1 63026
box 0 0 1 1
use contact_18  contact_18_48
timestamp 1644969367
transform 1 0 1138 0 1 61483
box 0 0 1 1
use contact_17  contact_17_48
timestamp 1644969367
transform 1 0 1172 0 1 61488
box 0 0 1 1
use contact_18  contact_18_49
timestamp 1644969367
transform 1 0 1138 0 1 59945
box 0 0 1 1
use contact_17  contact_17_49
timestamp 1644969367
transform 1 0 1172 0 1 59950
box 0 0 1 1
use contact_18  contact_18_50
timestamp 1644969367
transform 1 0 1138 0 1 58407
box 0 0 1 1
use contact_17  contact_17_50
timestamp 1644969367
transform 1 0 1172 0 1 58412
box 0 0 1 1
use contact_18  contact_18_51
timestamp 1644969367
transform 1 0 1138 0 1 59945
box 0 0 1 1
use contact_17  contact_17_51
timestamp 1644969367
transform 1 0 1172 0 1 59950
box 0 0 1 1
use contact_18  contact_18_52
timestamp 1644969367
transform 1 0 1138 0 1 58407
box 0 0 1 1
use contact_17  contact_17_52
timestamp 1644969367
transform 1 0 1172 0 1 58412
box 0 0 1 1
use contact_18  contact_18_53
timestamp 1644969367
transform 1 0 1138 0 1 56869
box 0 0 1 1
use contact_17  contact_17_53
timestamp 1644969367
transform 1 0 1172 0 1 56874
box 0 0 1 1
use contact_18  contact_18_54
timestamp 1644969367
transform 1 0 1138 0 1 55331
box 0 0 1 1
use contact_17  contact_17_54
timestamp 1644969367
transform 1 0 1172 0 1 55336
box 0 0 1 1
use contact_18  contact_18_55
timestamp 1644969367
transform 1 0 1138 0 1 56869
box 0 0 1 1
use contact_17  contact_17_55
timestamp 1644969367
transform 1 0 1172 0 1 56874
box 0 0 1 1
use contact_18  contact_18_56
timestamp 1644969367
transform 1 0 1138 0 1 55331
box 0 0 1 1
use contact_17  contact_17_56
timestamp 1644969367
transform 1 0 1172 0 1 55336
box 0 0 1 1
use contact_18  contact_18_57
timestamp 1644969367
transform 1 0 1138 0 1 53793
box 0 0 1 1
use contact_17  contact_17_57
timestamp 1644969367
transform 1 0 1172 0 1 53798
box 0 0 1 1
use contact_18  contact_18_58
timestamp 1644969367
transform 1 0 1138 0 1 52255
box 0 0 1 1
use contact_17  contact_17_58
timestamp 1644969367
transform 1 0 1172 0 1 52260
box 0 0 1 1
use contact_18  contact_18_59
timestamp 1644969367
transform 1 0 1138 0 1 53793
box 0 0 1 1
use contact_17  contact_17_59
timestamp 1644969367
transform 1 0 1172 0 1 53798
box 0 0 1 1
use contact_18  contact_18_60
timestamp 1644969367
transform 1 0 1138 0 1 52255
box 0 0 1 1
use contact_17  contact_17_60
timestamp 1644969367
transform 1 0 1172 0 1 52260
box 0 0 1 1
use contact_18  contact_18_61
timestamp 1644969367
transform 1 0 1138 0 1 50717
box 0 0 1 1
use contact_17  contact_17_61
timestamp 1644969367
transform 1 0 1172 0 1 50722
box 0 0 1 1
use contact_18  contact_18_62
timestamp 1644969367
transform 1 0 1138 0 1 49179
box 0 0 1 1
use contact_17  contact_17_62
timestamp 1644969367
transform 1 0 1172 0 1 49184
box 0 0 1 1
use contact_18  contact_18_63
timestamp 1644969367
transform 1 0 1138 0 1 50717
box 0 0 1 1
use contact_17  contact_17_63
timestamp 1644969367
transform 1 0 1172 0 1 50722
box 0 0 1 1
use contact_18  contact_18_64
timestamp 1644969367
transform 1 0 1138 0 1 49179
box 0 0 1 1
use contact_17  contact_17_64
timestamp 1644969367
transform 1 0 1172 0 1 49184
box 0 0 1 1
use contact_18  contact_18_65
timestamp 1644969367
transform 1 0 1138 0 1 47641
box 0 0 1 1
use contact_17  contact_17_65
timestamp 1644969367
transform 1 0 1172 0 1 47646
box 0 0 1 1
use contact_18  contact_18_66
timestamp 1644969367
transform 1 0 1138 0 1 46103
box 0 0 1 1
use contact_17  contact_17_66
timestamp 1644969367
transform 1 0 1172 0 1 46108
box 0 0 1 1
use contact_18  contact_18_67
timestamp 1644969367
transform 1 0 1138 0 1 47641
box 0 0 1 1
use contact_17  contact_17_67
timestamp 1644969367
transform 1 0 1172 0 1 47646
box 0 0 1 1
use contact_18  contact_18_68
timestamp 1644969367
transform 1 0 1138 0 1 46103
box 0 0 1 1
use contact_17  contact_17_68
timestamp 1644969367
transform 1 0 1172 0 1 46108
box 0 0 1 1
use contact_18  contact_18_69
timestamp 1644969367
transform 1 0 1138 0 1 44565
box 0 0 1 1
use contact_17  contact_17_69
timestamp 1644969367
transform 1 0 1172 0 1 44570
box 0 0 1 1
use contact_18  contact_18_70
timestamp 1644969367
transform 1 0 1138 0 1 43027
box 0 0 1 1
use contact_17  contact_17_70
timestamp 1644969367
transform 1 0 1172 0 1 43032
box 0 0 1 1
use contact_18  contact_18_71
timestamp 1644969367
transform 1 0 1138 0 1 44565
box 0 0 1 1
use contact_17  contact_17_71
timestamp 1644969367
transform 1 0 1172 0 1 44570
box 0 0 1 1
use contact_18  contact_18_72
timestamp 1644969367
transform 1 0 1138 0 1 43027
box 0 0 1 1
use contact_17  contact_17_72
timestamp 1644969367
transform 1 0 1172 0 1 43032
box 0 0 1 1
use contact_18  contact_18_73
timestamp 1644969367
transform 1 0 1138 0 1 41489
box 0 0 1 1
use contact_17  contact_17_73
timestamp 1644969367
transform 1 0 1172 0 1 41494
box 0 0 1 1
use contact_18  contact_18_74
timestamp 1644969367
transform 1 0 1138 0 1 39951
box 0 0 1 1
use contact_17  contact_17_74
timestamp 1644969367
transform 1 0 1172 0 1 39956
box 0 0 1 1
use contact_18  contact_18_75
timestamp 1644969367
transform 1 0 1138 0 1 41489
box 0 0 1 1
use contact_17  contact_17_75
timestamp 1644969367
transform 1 0 1172 0 1 41494
box 0 0 1 1
use contact_18  contact_18_76
timestamp 1644969367
transform 1 0 1138 0 1 39951
box 0 0 1 1
use contact_17  contact_17_76
timestamp 1644969367
transform 1 0 1172 0 1 39956
box 0 0 1 1
use contact_18  contact_18_77
timestamp 1644969367
transform 1 0 1138 0 1 38413
box 0 0 1 1
use contact_17  contact_17_77
timestamp 1644969367
transform 1 0 1172 0 1 38418
box 0 0 1 1
use contact_18  contact_18_78
timestamp 1644969367
transform 1 0 1138 0 1 36875
box 0 0 1 1
use contact_17  contact_17_78
timestamp 1644969367
transform 1 0 1172 0 1 36880
box 0 0 1 1
use contact_18  contact_18_79
timestamp 1644969367
transform 1 0 1138 0 1 38413
box 0 0 1 1
use contact_17  contact_17_79
timestamp 1644969367
transform 1 0 1172 0 1 38418
box 0 0 1 1
use contact_18  contact_18_80
timestamp 1644969367
transform 1 0 1138 0 1 36875
box 0 0 1 1
use contact_17  contact_17_80
timestamp 1644969367
transform 1 0 1172 0 1 36880
box 0 0 1 1
use contact_18  contact_18_81
timestamp 1644969367
transform 1 0 1138 0 1 35337
box 0 0 1 1
use contact_17  contact_17_81
timestamp 1644969367
transform 1 0 1172 0 1 35342
box 0 0 1 1
use contact_18  contact_18_82
timestamp 1644969367
transform 1 0 1138 0 1 33799
box 0 0 1 1
use contact_17  contact_17_82
timestamp 1644969367
transform 1 0 1172 0 1 33804
box 0 0 1 1
use contact_18  contact_18_83
timestamp 1644969367
transform 1 0 1138 0 1 35337
box 0 0 1 1
use contact_17  contact_17_83
timestamp 1644969367
transform 1 0 1172 0 1 35342
box 0 0 1 1
use contact_18  contact_18_84
timestamp 1644969367
transform 1 0 1138 0 1 33799
box 0 0 1 1
use contact_17  contact_17_84
timestamp 1644969367
transform 1 0 1172 0 1 33804
box 0 0 1 1
use contact_18  contact_18_85
timestamp 1644969367
transform 1 0 1138 0 1 32261
box 0 0 1 1
use contact_17  contact_17_85
timestamp 1644969367
transform 1 0 1172 0 1 32266
box 0 0 1 1
use contact_18  contact_18_86
timestamp 1644969367
transform 1 0 1138 0 1 30723
box 0 0 1 1
use contact_17  contact_17_86
timestamp 1644969367
transform 1 0 1172 0 1 30728
box 0 0 1 1
use contact_18  contact_18_87
timestamp 1644969367
transform 1 0 1138 0 1 32261
box 0 0 1 1
use contact_17  contact_17_87
timestamp 1644969367
transform 1 0 1172 0 1 32266
box 0 0 1 1
use contact_18  contact_18_88
timestamp 1644969367
transform 1 0 1138 0 1 30723
box 0 0 1 1
use contact_17  contact_17_88
timestamp 1644969367
transform 1 0 1172 0 1 30728
box 0 0 1 1
use contact_18  contact_18_89
timestamp 1644969367
transform 1 0 1138 0 1 29185
box 0 0 1 1
use contact_17  contact_17_89
timestamp 1644969367
transform 1 0 1172 0 1 29190
box 0 0 1 1
use contact_18  contact_18_90
timestamp 1644969367
transform 1 0 1138 0 1 27647
box 0 0 1 1
use contact_17  contact_17_90
timestamp 1644969367
transform 1 0 1172 0 1 27652
box 0 0 1 1
use contact_18  contact_18_91
timestamp 1644969367
transform 1 0 1138 0 1 29185
box 0 0 1 1
use contact_17  contact_17_91
timestamp 1644969367
transform 1 0 1172 0 1 29190
box 0 0 1 1
use contact_18  contact_18_92
timestamp 1644969367
transform 1 0 1138 0 1 27647
box 0 0 1 1
use contact_17  contact_17_92
timestamp 1644969367
transform 1 0 1172 0 1 27652
box 0 0 1 1
use contact_18  contact_18_93
timestamp 1644969367
transform 1 0 1138 0 1 26109
box 0 0 1 1
use contact_17  contact_17_93
timestamp 1644969367
transform 1 0 1172 0 1 26114
box 0 0 1 1
use contact_18  contact_18_94
timestamp 1644969367
transform 1 0 1138 0 1 24571
box 0 0 1 1
use contact_17  contact_17_94
timestamp 1644969367
transform 1 0 1172 0 1 24576
box 0 0 1 1
use contact_18  contact_18_95
timestamp 1644969367
transform 1 0 1138 0 1 26109
box 0 0 1 1
use contact_17  contact_17_95
timestamp 1644969367
transform 1 0 1172 0 1 26114
box 0 0 1 1
use contact_18  contact_18_96
timestamp 1644969367
transform 1 0 1138 0 1 24571
box 0 0 1 1
use contact_17  contact_17_96
timestamp 1644969367
transform 1 0 1172 0 1 24576
box 0 0 1 1
use contact_18  contact_18_97
timestamp 1644969367
transform 1 0 1138 0 1 23033
box 0 0 1 1
use contact_17  contact_17_97
timestamp 1644969367
transform 1 0 1172 0 1 23038
box 0 0 1 1
use contact_18  contact_18_98
timestamp 1644969367
transform 1 0 1138 0 1 21495
box 0 0 1 1
use contact_17  contact_17_98
timestamp 1644969367
transform 1 0 1172 0 1 21500
box 0 0 1 1
use contact_18  contact_18_99
timestamp 1644969367
transform 1 0 1138 0 1 23033
box 0 0 1 1
use contact_17  contact_17_99
timestamp 1644969367
transform 1 0 1172 0 1 23038
box 0 0 1 1
use contact_18  contact_18_100
timestamp 1644969367
transform 1 0 1138 0 1 21495
box 0 0 1 1
use contact_17  contact_17_100
timestamp 1644969367
transform 1 0 1172 0 1 21500
box 0 0 1 1
use contact_18  contact_18_101
timestamp 1644969367
transform 1 0 1138 0 1 19957
box 0 0 1 1
use contact_17  contact_17_101
timestamp 1644969367
transform 1 0 1172 0 1 19962
box 0 0 1 1
use contact_18  contact_18_102
timestamp 1644969367
transform 1 0 1138 0 1 18419
box 0 0 1 1
use contact_17  contact_17_102
timestamp 1644969367
transform 1 0 1172 0 1 18424
box 0 0 1 1
use contact_18  contact_18_103
timestamp 1644969367
transform 1 0 1138 0 1 19957
box 0 0 1 1
use contact_17  contact_17_103
timestamp 1644969367
transform 1 0 1172 0 1 19962
box 0 0 1 1
use contact_18  contact_18_104
timestamp 1644969367
transform 1 0 1138 0 1 18419
box 0 0 1 1
use contact_17  contact_17_104
timestamp 1644969367
transform 1 0 1172 0 1 18424
box 0 0 1 1
use contact_18  contact_18_105
timestamp 1644969367
transform 1 0 1138 0 1 16881
box 0 0 1 1
use contact_17  contact_17_105
timestamp 1644969367
transform 1 0 1172 0 1 16886
box 0 0 1 1
use contact_18  contact_18_106
timestamp 1644969367
transform 1 0 1138 0 1 15343
box 0 0 1 1
use contact_17  contact_17_106
timestamp 1644969367
transform 1 0 1172 0 1 15348
box 0 0 1 1
use contact_18  contact_18_107
timestamp 1644969367
transform 1 0 1138 0 1 16881
box 0 0 1 1
use contact_17  contact_17_107
timestamp 1644969367
transform 1 0 1172 0 1 16886
box 0 0 1 1
use contact_18  contact_18_108
timestamp 1644969367
transform 1 0 1138 0 1 15343
box 0 0 1 1
use contact_17  contact_17_108
timestamp 1644969367
transform 1 0 1172 0 1 15348
box 0 0 1 1
use contact_18  contact_18_109
timestamp 1644969367
transform 1 0 1138 0 1 13805
box 0 0 1 1
use contact_17  contact_17_109
timestamp 1644969367
transform 1 0 1172 0 1 13810
box 0 0 1 1
use contact_18  contact_18_110
timestamp 1644969367
transform 1 0 1138 0 1 12267
box 0 0 1 1
use contact_17  contact_17_110
timestamp 1644969367
transform 1 0 1172 0 1 12272
box 0 0 1 1
use contact_18  contact_18_111
timestamp 1644969367
transform 1 0 1138 0 1 13805
box 0 0 1 1
use contact_17  contact_17_111
timestamp 1644969367
transform 1 0 1172 0 1 13810
box 0 0 1 1
use contact_18  contact_18_112
timestamp 1644969367
transform 1 0 1138 0 1 12267
box 0 0 1 1
use contact_17  contact_17_112
timestamp 1644969367
transform 1 0 1172 0 1 12272
box 0 0 1 1
use contact_18  contact_18_113
timestamp 1644969367
transform 1 0 1138 0 1 10729
box 0 0 1 1
use contact_17  contact_17_113
timestamp 1644969367
transform 1 0 1172 0 1 10734
box 0 0 1 1
use contact_18  contact_18_114
timestamp 1644969367
transform 1 0 1138 0 1 9191
box 0 0 1 1
use contact_17  contact_17_114
timestamp 1644969367
transform 1 0 1172 0 1 9196
box 0 0 1 1
use contact_18  contact_18_115
timestamp 1644969367
transform 1 0 1138 0 1 10729
box 0 0 1 1
use contact_17  contact_17_115
timestamp 1644969367
transform 1 0 1172 0 1 10734
box 0 0 1 1
use contact_18  contact_18_116
timestamp 1644969367
transform 1 0 1138 0 1 9191
box 0 0 1 1
use contact_17  contact_17_116
timestamp 1644969367
transform 1 0 1172 0 1 9196
box 0 0 1 1
use contact_18  contact_18_117
timestamp 1644969367
transform 1 0 1138 0 1 7653
box 0 0 1 1
use contact_17  contact_17_117
timestamp 1644969367
transform 1 0 1172 0 1 7658
box 0 0 1 1
use contact_18  contact_18_118
timestamp 1644969367
transform 1 0 1138 0 1 6115
box 0 0 1 1
use contact_17  contact_17_118
timestamp 1644969367
transform 1 0 1172 0 1 6120
box 0 0 1 1
use contact_18  contact_18_119
timestamp 1644969367
transform 1 0 1138 0 1 7653
box 0 0 1 1
use contact_17  contact_17_119
timestamp 1644969367
transform 1 0 1172 0 1 7658
box 0 0 1 1
use contact_18  contact_18_120
timestamp 1644969367
transform 1 0 1138 0 1 6115
box 0 0 1 1
use contact_17  contact_17_120
timestamp 1644969367
transform 1 0 1172 0 1 6120
box 0 0 1 1
use contact_18  contact_18_121
timestamp 1644969367
transform 1 0 1138 0 1 4577
box 0 0 1 1
use contact_17  contact_17_121
timestamp 1644969367
transform 1 0 1172 0 1 4582
box 0 0 1 1
use contact_18  contact_18_122
timestamp 1644969367
transform 1 0 1138 0 1 3039
box 0 0 1 1
use contact_17  contact_17_122
timestamp 1644969367
transform 1 0 1172 0 1 3044
box 0 0 1 1
use contact_18  contact_18_123
timestamp 1644969367
transform 1 0 1138 0 1 4577
box 0 0 1 1
use contact_17  contact_17_123
timestamp 1644969367
transform 1 0 1172 0 1 4582
box 0 0 1 1
use contact_18  contact_18_124
timestamp 1644969367
transform 1 0 1138 0 1 3039
box 0 0 1 1
use contact_17  contact_17_124
timestamp 1644969367
transform 1 0 1172 0 1 3044
box 0 0 1 1
use contact_18  contact_18_125
timestamp 1644969367
transform 1 0 1138 0 1 1501
box 0 0 1 1
use contact_17  contact_17_125
timestamp 1644969367
transform 1 0 1172 0 1 1506
box 0 0 1 1
use contact_18  contact_18_126
timestamp 1644969367
transform 1 0 1138 0 1 -37
box 0 0 1 1
use contact_17  contact_17_126
timestamp 1644969367
transform 1 0 1172 0 1 -32
box 0 0 1 1
use contact_18  contact_18_127
timestamp 1644969367
transform 1 0 1138 0 1 1501
box 0 0 1 1
use contact_17  contact_17_127
timestamp 1644969367
transform 1 0 1172 0 1 1506
box 0 0 1 1
use wordline_driver_cell  wordline_driver_cell_0
timestamp 1644969367
transform 1 0 0 0 -1 98432
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_1
timestamp 1644969367
transform 1 0 0 0 1 95356
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_2
timestamp 1644969367
transform 1 0 0 0 -1 95356
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_3
timestamp 1644969367
transform 1 0 0 0 1 92280
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_4
timestamp 1644969367
transform 1 0 0 0 -1 92280
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_5
timestamp 1644969367
transform 1 0 0 0 1 89204
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_6
timestamp 1644969367
transform 1 0 0 0 -1 89204
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_7
timestamp 1644969367
transform 1 0 0 0 1 86128
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_8
timestamp 1644969367
transform 1 0 0 0 -1 86128
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_9
timestamp 1644969367
transform 1 0 0 0 1 83052
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_10
timestamp 1644969367
transform 1 0 0 0 -1 83052
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_11
timestamp 1644969367
transform 1 0 0 0 1 79976
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_12
timestamp 1644969367
transform 1 0 0 0 -1 79976
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_13
timestamp 1644969367
transform 1 0 0 0 1 76900
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_14
timestamp 1644969367
transform 1 0 0 0 -1 76900
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_15
timestamp 1644969367
transform 1 0 0 0 1 73824
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_16
timestamp 1644969367
transform 1 0 0 0 -1 73824
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_17
timestamp 1644969367
transform 1 0 0 0 1 70748
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_18
timestamp 1644969367
transform 1 0 0 0 -1 70748
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_19
timestamp 1644969367
transform 1 0 0 0 1 67672
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_20
timestamp 1644969367
transform 1 0 0 0 -1 67672
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_21
timestamp 1644969367
transform 1 0 0 0 1 64596
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_22
timestamp 1644969367
transform 1 0 0 0 -1 64596
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_23
timestamp 1644969367
transform 1 0 0 0 1 61520
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_24
timestamp 1644969367
transform 1 0 0 0 -1 61520
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_25
timestamp 1644969367
transform 1 0 0 0 1 58444
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_26
timestamp 1644969367
transform 1 0 0 0 -1 58444
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_27
timestamp 1644969367
transform 1 0 0 0 1 55368
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_28
timestamp 1644969367
transform 1 0 0 0 -1 55368
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_29
timestamp 1644969367
transform 1 0 0 0 1 52292
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_30
timestamp 1644969367
transform 1 0 0 0 -1 52292
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_31
timestamp 1644969367
transform 1 0 0 0 1 49216
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_32
timestamp 1644969367
transform 1 0 0 0 -1 49216
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_33
timestamp 1644969367
transform 1 0 0 0 1 46140
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_34
timestamp 1644969367
transform 1 0 0 0 -1 46140
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_35
timestamp 1644969367
transform 1 0 0 0 1 43064
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_36
timestamp 1644969367
transform 1 0 0 0 -1 43064
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_37
timestamp 1644969367
transform 1 0 0 0 1 39988
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_38
timestamp 1644969367
transform 1 0 0 0 -1 39988
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_39
timestamp 1644969367
transform 1 0 0 0 1 36912
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_40
timestamp 1644969367
transform 1 0 0 0 -1 36912
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_41
timestamp 1644969367
transform 1 0 0 0 1 33836
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_42
timestamp 1644969367
transform 1 0 0 0 -1 33836
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_43
timestamp 1644969367
transform 1 0 0 0 1 30760
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_44
timestamp 1644969367
transform 1 0 0 0 -1 30760
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_45
timestamp 1644969367
transform 1 0 0 0 1 27684
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_46
timestamp 1644969367
transform 1 0 0 0 -1 27684
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_47
timestamp 1644969367
transform 1 0 0 0 1 24608
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_48
timestamp 1644969367
transform 1 0 0 0 -1 24608
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_49
timestamp 1644969367
transform 1 0 0 0 1 21532
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_50
timestamp 1644969367
transform 1 0 0 0 -1 21532
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_51
timestamp 1644969367
transform 1 0 0 0 1 18456
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_52
timestamp 1644969367
transform 1 0 0 0 -1 18456
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_53
timestamp 1644969367
transform 1 0 0 0 1 15380
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_54
timestamp 1644969367
transform 1 0 0 0 -1 15380
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_55
timestamp 1644969367
transform 1 0 0 0 1 12304
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_56
timestamp 1644969367
transform 1 0 0 0 -1 12304
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_57
timestamp 1644969367
transform 1 0 0 0 1 9228
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_58
timestamp 1644969367
transform 1 0 0 0 -1 9228
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_59
timestamp 1644969367
transform 1 0 0 0 1 6152
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_60
timestamp 1644969367
transform 1 0 0 0 -1 6152
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_61
timestamp 1644969367
transform 1 0 0 0 1 3076
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_62
timestamp 1644969367
transform 1 0 0 0 -1 3076
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_63
timestamp 1644969367
transform 1 0 0 0 1 0
box 0 -42 1204 1616
<< labels >>
rlabel metal2 s 0 0 28 98432 4 wl_en
rlabel metal1 s 56 848 126 876 4 in0_0
rlabel metal1 s 234 702 318 730 4 in1_0
rlabel metal1 s 536 582 618 610 4 in2_0
rlabel metal1 s 1176 778 1204 806 4 rwl0_0
rlabel metal1 s 1176 1004 1204 1032 4 rwl1_0
rlabel metal1 s 1176 652 1204 680 4 wwl0_0
rlabel metal1 s 56 2200 126 2228 4 in0_1
rlabel metal1 s 234 2346 318 2374 4 in1_1
rlabel metal1 s 536 2466 618 2494 4 in2_1
rlabel metal1 s 1176 2270 1204 2298 4 rwl0_1
rlabel metal1 s 1176 2044 1204 2072 4 rwl1_1
rlabel metal1 s 1176 2396 1204 2424 4 wwl0_1
rlabel metal1 s 56 3924 126 3952 4 in0_2
rlabel metal1 s 234 3778 318 3806 4 in1_2
rlabel metal1 s 536 3658 618 3686 4 in2_2
rlabel metal1 s 1176 3854 1204 3882 4 rwl0_2
rlabel metal1 s 1176 4080 1204 4108 4 rwl1_2
rlabel metal1 s 1176 3728 1204 3756 4 wwl0_2
rlabel metal1 s 56 5276 126 5304 4 in0_3
rlabel metal1 s 234 5422 318 5450 4 in1_3
rlabel metal1 s 536 5542 618 5570 4 in2_3
rlabel metal1 s 1176 5346 1204 5374 4 rwl0_3
rlabel metal1 s 1176 5120 1204 5148 4 rwl1_3
rlabel metal1 s 1176 5472 1204 5500 4 wwl0_3
rlabel metal1 s 56 7000 126 7028 4 in0_4
rlabel metal1 s 234 6854 318 6882 4 in1_4
rlabel metal1 s 536 6734 618 6762 4 in2_4
rlabel metal1 s 1176 6930 1204 6958 4 rwl0_4
rlabel metal1 s 1176 7156 1204 7184 4 rwl1_4
rlabel metal1 s 1176 6804 1204 6832 4 wwl0_4
rlabel metal1 s 56 8352 126 8380 4 in0_5
rlabel metal1 s 234 8498 318 8526 4 in1_5
rlabel metal1 s 536 8618 618 8646 4 in2_5
rlabel metal1 s 1176 8422 1204 8450 4 rwl0_5
rlabel metal1 s 1176 8196 1204 8224 4 rwl1_5
rlabel metal1 s 1176 8548 1204 8576 4 wwl0_5
rlabel metal1 s 56 10076 126 10104 4 in0_6
rlabel metal1 s 234 9930 318 9958 4 in1_6
rlabel metal1 s 536 9810 618 9838 4 in2_6
rlabel metal1 s 1176 10006 1204 10034 4 rwl0_6
rlabel metal1 s 1176 10232 1204 10260 4 rwl1_6
rlabel metal1 s 1176 9880 1204 9908 4 wwl0_6
rlabel metal1 s 56 11428 126 11456 4 in0_7
rlabel metal1 s 234 11574 318 11602 4 in1_7
rlabel metal1 s 536 11694 618 11722 4 in2_7
rlabel metal1 s 1176 11498 1204 11526 4 rwl0_7
rlabel metal1 s 1176 11272 1204 11300 4 rwl1_7
rlabel metal1 s 1176 11624 1204 11652 4 wwl0_7
rlabel metal1 s 56 13152 126 13180 4 in0_8
rlabel metal1 s 234 13006 318 13034 4 in1_8
rlabel metal1 s 536 12886 618 12914 4 in2_8
rlabel metal1 s 1176 13082 1204 13110 4 rwl0_8
rlabel metal1 s 1176 13308 1204 13336 4 rwl1_8
rlabel metal1 s 1176 12956 1204 12984 4 wwl0_8
rlabel metal1 s 56 14504 126 14532 4 in0_9
rlabel metal1 s 234 14650 318 14678 4 in1_9
rlabel metal1 s 536 14770 618 14798 4 in2_9
rlabel metal1 s 1176 14574 1204 14602 4 rwl0_9
rlabel metal1 s 1176 14348 1204 14376 4 rwl1_9
rlabel metal1 s 1176 14700 1204 14728 4 wwl0_9
rlabel metal1 s 56 16228 126 16256 4 in0_10
rlabel metal1 s 234 16082 318 16110 4 in1_10
rlabel metal1 s 536 15962 618 15990 4 in2_10
rlabel metal1 s 1176 16158 1204 16186 4 rwl0_10
rlabel metal1 s 1176 16384 1204 16412 4 rwl1_10
rlabel metal1 s 1176 16032 1204 16060 4 wwl0_10
rlabel metal1 s 56 17580 126 17608 4 in0_11
rlabel metal1 s 234 17726 318 17754 4 in1_11
rlabel metal1 s 536 17846 618 17874 4 in2_11
rlabel metal1 s 1176 17650 1204 17678 4 rwl0_11
rlabel metal1 s 1176 17424 1204 17452 4 rwl1_11
rlabel metal1 s 1176 17776 1204 17804 4 wwl0_11
rlabel metal1 s 56 19304 126 19332 4 in0_12
rlabel metal1 s 234 19158 318 19186 4 in1_12
rlabel metal1 s 536 19038 618 19066 4 in2_12
rlabel metal1 s 1176 19234 1204 19262 4 rwl0_12
rlabel metal1 s 1176 19460 1204 19488 4 rwl1_12
rlabel metal1 s 1176 19108 1204 19136 4 wwl0_12
rlabel metal1 s 56 20656 126 20684 4 in0_13
rlabel metal1 s 234 20802 318 20830 4 in1_13
rlabel metal1 s 536 20922 618 20950 4 in2_13
rlabel metal1 s 1176 20726 1204 20754 4 rwl0_13
rlabel metal1 s 1176 20500 1204 20528 4 rwl1_13
rlabel metal1 s 1176 20852 1204 20880 4 wwl0_13
rlabel metal1 s 56 22380 126 22408 4 in0_14
rlabel metal1 s 234 22234 318 22262 4 in1_14
rlabel metal1 s 536 22114 618 22142 4 in2_14
rlabel metal1 s 1176 22310 1204 22338 4 rwl0_14
rlabel metal1 s 1176 22536 1204 22564 4 rwl1_14
rlabel metal1 s 1176 22184 1204 22212 4 wwl0_14
rlabel metal1 s 56 23732 126 23760 4 in0_15
rlabel metal1 s 234 23878 318 23906 4 in1_15
rlabel metal1 s 536 23998 618 24026 4 in2_15
rlabel metal1 s 1176 23802 1204 23830 4 rwl0_15
rlabel metal1 s 1176 23576 1204 23604 4 rwl1_15
rlabel metal1 s 1176 23928 1204 23956 4 wwl0_15
rlabel metal1 s 56 25456 126 25484 4 in0_16
rlabel metal1 s 234 25310 318 25338 4 in1_16
rlabel metal1 s 536 25190 618 25218 4 in2_16
rlabel metal1 s 1176 25386 1204 25414 4 rwl0_16
rlabel metal1 s 1176 25612 1204 25640 4 rwl1_16
rlabel metal1 s 1176 25260 1204 25288 4 wwl0_16
rlabel metal1 s 56 26808 126 26836 4 in0_17
rlabel metal1 s 234 26954 318 26982 4 in1_17
rlabel metal1 s 536 27074 618 27102 4 in2_17
rlabel metal1 s 1176 26878 1204 26906 4 rwl0_17
rlabel metal1 s 1176 26652 1204 26680 4 rwl1_17
rlabel metal1 s 1176 27004 1204 27032 4 wwl0_17
rlabel metal1 s 56 28532 126 28560 4 in0_18
rlabel metal1 s 234 28386 318 28414 4 in1_18
rlabel metal1 s 536 28266 618 28294 4 in2_18
rlabel metal1 s 1176 28462 1204 28490 4 rwl0_18
rlabel metal1 s 1176 28688 1204 28716 4 rwl1_18
rlabel metal1 s 1176 28336 1204 28364 4 wwl0_18
rlabel metal1 s 56 29884 126 29912 4 in0_19
rlabel metal1 s 234 30030 318 30058 4 in1_19
rlabel metal1 s 536 30150 618 30178 4 in2_19
rlabel metal1 s 1176 29954 1204 29982 4 rwl0_19
rlabel metal1 s 1176 29728 1204 29756 4 rwl1_19
rlabel metal1 s 1176 30080 1204 30108 4 wwl0_19
rlabel metal1 s 56 31608 126 31636 4 in0_20
rlabel metal1 s 234 31462 318 31490 4 in1_20
rlabel metal1 s 536 31342 618 31370 4 in2_20
rlabel metal1 s 1176 31538 1204 31566 4 rwl0_20
rlabel metal1 s 1176 31764 1204 31792 4 rwl1_20
rlabel metal1 s 1176 31412 1204 31440 4 wwl0_20
rlabel metal1 s 56 32960 126 32988 4 in0_21
rlabel metal1 s 234 33106 318 33134 4 in1_21
rlabel metal1 s 536 33226 618 33254 4 in2_21
rlabel metal1 s 1176 33030 1204 33058 4 rwl0_21
rlabel metal1 s 1176 32804 1204 32832 4 rwl1_21
rlabel metal1 s 1176 33156 1204 33184 4 wwl0_21
rlabel metal1 s 56 34684 126 34712 4 in0_22
rlabel metal1 s 234 34538 318 34566 4 in1_22
rlabel metal1 s 536 34418 618 34446 4 in2_22
rlabel metal1 s 1176 34614 1204 34642 4 rwl0_22
rlabel metal1 s 1176 34840 1204 34868 4 rwl1_22
rlabel metal1 s 1176 34488 1204 34516 4 wwl0_22
rlabel metal1 s 56 36036 126 36064 4 in0_23
rlabel metal1 s 234 36182 318 36210 4 in1_23
rlabel metal1 s 536 36302 618 36330 4 in2_23
rlabel metal1 s 1176 36106 1204 36134 4 rwl0_23
rlabel metal1 s 1176 35880 1204 35908 4 rwl1_23
rlabel metal1 s 1176 36232 1204 36260 4 wwl0_23
rlabel metal1 s 56 37760 126 37788 4 in0_24
rlabel metal1 s 234 37614 318 37642 4 in1_24
rlabel metal1 s 536 37494 618 37522 4 in2_24
rlabel metal1 s 1176 37690 1204 37718 4 rwl0_24
rlabel metal1 s 1176 37916 1204 37944 4 rwl1_24
rlabel metal1 s 1176 37564 1204 37592 4 wwl0_24
rlabel metal1 s 56 39112 126 39140 4 in0_25
rlabel metal1 s 234 39258 318 39286 4 in1_25
rlabel metal1 s 536 39378 618 39406 4 in2_25
rlabel metal1 s 1176 39182 1204 39210 4 rwl0_25
rlabel metal1 s 1176 38956 1204 38984 4 rwl1_25
rlabel metal1 s 1176 39308 1204 39336 4 wwl0_25
rlabel metal1 s 56 40836 126 40864 4 in0_26
rlabel metal1 s 234 40690 318 40718 4 in1_26
rlabel metal1 s 536 40570 618 40598 4 in2_26
rlabel metal1 s 1176 40766 1204 40794 4 rwl0_26
rlabel metal1 s 1176 40992 1204 41020 4 rwl1_26
rlabel metal1 s 1176 40640 1204 40668 4 wwl0_26
rlabel metal1 s 56 42188 126 42216 4 in0_27
rlabel metal1 s 234 42334 318 42362 4 in1_27
rlabel metal1 s 536 42454 618 42482 4 in2_27
rlabel metal1 s 1176 42258 1204 42286 4 rwl0_27
rlabel metal1 s 1176 42032 1204 42060 4 rwl1_27
rlabel metal1 s 1176 42384 1204 42412 4 wwl0_27
rlabel metal1 s 56 43912 126 43940 4 in0_28
rlabel metal1 s 234 43766 318 43794 4 in1_28
rlabel metal1 s 536 43646 618 43674 4 in2_28
rlabel metal1 s 1176 43842 1204 43870 4 rwl0_28
rlabel metal1 s 1176 44068 1204 44096 4 rwl1_28
rlabel metal1 s 1176 43716 1204 43744 4 wwl0_28
rlabel metal1 s 56 45264 126 45292 4 in0_29
rlabel metal1 s 234 45410 318 45438 4 in1_29
rlabel metal1 s 536 45530 618 45558 4 in2_29
rlabel metal1 s 1176 45334 1204 45362 4 rwl0_29
rlabel metal1 s 1176 45108 1204 45136 4 rwl1_29
rlabel metal1 s 1176 45460 1204 45488 4 wwl0_29
rlabel metal1 s 56 46988 126 47016 4 in0_30
rlabel metal1 s 234 46842 318 46870 4 in1_30
rlabel metal1 s 536 46722 618 46750 4 in2_30
rlabel metal1 s 1176 46918 1204 46946 4 rwl0_30
rlabel metal1 s 1176 47144 1204 47172 4 rwl1_30
rlabel metal1 s 1176 46792 1204 46820 4 wwl0_30
rlabel metal1 s 56 48340 126 48368 4 in0_31
rlabel metal1 s 234 48486 318 48514 4 in1_31
rlabel metal1 s 536 48606 618 48634 4 in2_31
rlabel metal1 s 1176 48410 1204 48438 4 rwl0_31
rlabel metal1 s 1176 48184 1204 48212 4 rwl1_31
rlabel metal1 s 1176 48536 1204 48564 4 wwl0_31
rlabel metal1 s 56 50064 126 50092 4 in0_32
rlabel metal1 s 234 49918 318 49946 4 in1_32
rlabel metal1 s 536 49798 618 49826 4 in2_32
rlabel metal1 s 1176 49994 1204 50022 4 rwl0_32
rlabel metal1 s 1176 50220 1204 50248 4 rwl1_32
rlabel metal1 s 1176 49868 1204 49896 4 wwl0_32
rlabel metal1 s 56 51416 126 51444 4 in0_33
rlabel metal1 s 234 51562 318 51590 4 in1_33
rlabel metal1 s 536 51682 618 51710 4 in2_33
rlabel metal1 s 1176 51486 1204 51514 4 rwl0_33
rlabel metal1 s 1176 51260 1204 51288 4 rwl1_33
rlabel metal1 s 1176 51612 1204 51640 4 wwl0_33
rlabel metal1 s 56 53140 126 53168 4 in0_34
rlabel metal1 s 234 52994 318 53022 4 in1_34
rlabel metal1 s 536 52874 618 52902 4 in2_34
rlabel metal1 s 1176 53070 1204 53098 4 rwl0_34
rlabel metal1 s 1176 53296 1204 53324 4 rwl1_34
rlabel metal1 s 1176 52944 1204 52972 4 wwl0_34
rlabel metal1 s 56 54492 126 54520 4 in0_35
rlabel metal1 s 234 54638 318 54666 4 in1_35
rlabel metal1 s 536 54758 618 54786 4 in2_35
rlabel metal1 s 1176 54562 1204 54590 4 rwl0_35
rlabel metal1 s 1176 54336 1204 54364 4 rwl1_35
rlabel metal1 s 1176 54688 1204 54716 4 wwl0_35
rlabel metal1 s 56 56216 126 56244 4 in0_36
rlabel metal1 s 234 56070 318 56098 4 in1_36
rlabel metal1 s 536 55950 618 55978 4 in2_36
rlabel metal1 s 1176 56146 1204 56174 4 rwl0_36
rlabel metal1 s 1176 56372 1204 56400 4 rwl1_36
rlabel metal1 s 1176 56020 1204 56048 4 wwl0_36
rlabel metal1 s 56 57568 126 57596 4 in0_37
rlabel metal1 s 234 57714 318 57742 4 in1_37
rlabel metal1 s 536 57834 618 57862 4 in2_37
rlabel metal1 s 1176 57638 1204 57666 4 rwl0_37
rlabel metal1 s 1176 57412 1204 57440 4 rwl1_37
rlabel metal1 s 1176 57764 1204 57792 4 wwl0_37
rlabel metal1 s 56 59292 126 59320 4 in0_38
rlabel metal1 s 234 59146 318 59174 4 in1_38
rlabel metal1 s 536 59026 618 59054 4 in2_38
rlabel metal1 s 1176 59222 1204 59250 4 rwl0_38
rlabel metal1 s 1176 59448 1204 59476 4 rwl1_38
rlabel metal1 s 1176 59096 1204 59124 4 wwl0_38
rlabel metal1 s 56 60644 126 60672 4 in0_39
rlabel metal1 s 234 60790 318 60818 4 in1_39
rlabel metal1 s 536 60910 618 60938 4 in2_39
rlabel metal1 s 1176 60714 1204 60742 4 rwl0_39
rlabel metal1 s 1176 60488 1204 60516 4 rwl1_39
rlabel metal1 s 1176 60840 1204 60868 4 wwl0_39
rlabel metal1 s 56 62368 126 62396 4 in0_40
rlabel metal1 s 234 62222 318 62250 4 in1_40
rlabel metal1 s 536 62102 618 62130 4 in2_40
rlabel metal1 s 1176 62298 1204 62326 4 rwl0_40
rlabel metal1 s 1176 62524 1204 62552 4 rwl1_40
rlabel metal1 s 1176 62172 1204 62200 4 wwl0_40
rlabel metal1 s 56 63720 126 63748 4 in0_41
rlabel metal1 s 234 63866 318 63894 4 in1_41
rlabel metal1 s 536 63986 618 64014 4 in2_41
rlabel metal1 s 1176 63790 1204 63818 4 rwl0_41
rlabel metal1 s 1176 63564 1204 63592 4 rwl1_41
rlabel metal1 s 1176 63916 1204 63944 4 wwl0_41
rlabel metal1 s 56 65444 126 65472 4 in0_42
rlabel metal1 s 234 65298 318 65326 4 in1_42
rlabel metal1 s 536 65178 618 65206 4 in2_42
rlabel metal1 s 1176 65374 1204 65402 4 rwl0_42
rlabel metal1 s 1176 65600 1204 65628 4 rwl1_42
rlabel metal1 s 1176 65248 1204 65276 4 wwl0_42
rlabel metal1 s 56 66796 126 66824 4 in0_43
rlabel metal1 s 234 66942 318 66970 4 in1_43
rlabel metal1 s 536 67062 618 67090 4 in2_43
rlabel metal1 s 1176 66866 1204 66894 4 rwl0_43
rlabel metal1 s 1176 66640 1204 66668 4 rwl1_43
rlabel metal1 s 1176 66992 1204 67020 4 wwl0_43
rlabel metal1 s 56 68520 126 68548 4 in0_44
rlabel metal1 s 234 68374 318 68402 4 in1_44
rlabel metal1 s 536 68254 618 68282 4 in2_44
rlabel metal1 s 1176 68450 1204 68478 4 rwl0_44
rlabel metal1 s 1176 68676 1204 68704 4 rwl1_44
rlabel metal1 s 1176 68324 1204 68352 4 wwl0_44
rlabel metal1 s 56 69872 126 69900 4 in0_45
rlabel metal1 s 234 70018 318 70046 4 in1_45
rlabel metal1 s 536 70138 618 70166 4 in2_45
rlabel metal1 s 1176 69942 1204 69970 4 rwl0_45
rlabel metal1 s 1176 69716 1204 69744 4 rwl1_45
rlabel metal1 s 1176 70068 1204 70096 4 wwl0_45
rlabel metal1 s 56 71596 126 71624 4 in0_46
rlabel metal1 s 234 71450 318 71478 4 in1_46
rlabel metal1 s 536 71330 618 71358 4 in2_46
rlabel metal1 s 1176 71526 1204 71554 4 rwl0_46
rlabel metal1 s 1176 71752 1204 71780 4 rwl1_46
rlabel metal1 s 1176 71400 1204 71428 4 wwl0_46
rlabel metal1 s 56 72948 126 72976 4 in0_47
rlabel metal1 s 234 73094 318 73122 4 in1_47
rlabel metal1 s 536 73214 618 73242 4 in2_47
rlabel metal1 s 1176 73018 1204 73046 4 rwl0_47
rlabel metal1 s 1176 72792 1204 72820 4 rwl1_47
rlabel metal1 s 1176 73144 1204 73172 4 wwl0_47
rlabel metal1 s 56 74672 126 74700 4 in0_48
rlabel metal1 s 234 74526 318 74554 4 in1_48
rlabel metal1 s 536 74406 618 74434 4 in2_48
rlabel metal1 s 1176 74602 1204 74630 4 rwl0_48
rlabel metal1 s 1176 74828 1204 74856 4 rwl1_48
rlabel metal1 s 1176 74476 1204 74504 4 wwl0_48
rlabel metal1 s 56 76024 126 76052 4 in0_49
rlabel metal1 s 234 76170 318 76198 4 in1_49
rlabel metal1 s 536 76290 618 76318 4 in2_49
rlabel metal1 s 1176 76094 1204 76122 4 rwl0_49
rlabel metal1 s 1176 75868 1204 75896 4 rwl1_49
rlabel metal1 s 1176 76220 1204 76248 4 wwl0_49
rlabel metal1 s 56 77748 126 77776 4 in0_50
rlabel metal1 s 234 77602 318 77630 4 in1_50
rlabel metal1 s 536 77482 618 77510 4 in2_50
rlabel metal1 s 1176 77678 1204 77706 4 rwl0_50
rlabel metal1 s 1176 77904 1204 77932 4 rwl1_50
rlabel metal1 s 1176 77552 1204 77580 4 wwl0_50
rlabel metal1 s 56 79100 126 79128 4 in0_51
rlabel metal1 s 234 79246 318 79274 4 in1_51
rlabel metal1 s 536 79366 618 79394 4 in2_51
rlabel metal1 s 1176 79170 1204 79198 4 rwl0_51
rlabel metal1 s 1176 78944 1204 78972 4 rwl1_51
rlabel metal1 s 1176 79296 1204 79324 4 wwl0_51
rlabel metal1 s 56 80824 126 80852 4 in0_52
rlabel metal1 s 234 80678 318 80706 4 in1_52
rlabel metal1 s 536 80558 618 80586 4 in2_52
rlabel metal1 s 1176 80754 1204 80782 4 rwl0_52
rlabel metal1 s 1176 80980 1204 81008 4 rwl1_52
rlabel metal1 s 1176 80628 1204 80656 4 wwl0_52
rlabel metal1 s 56 82176 126 82204 4 in0_53
rlabel metal1 s 234 82322 318 82350 4 in1_53
rlabel metal1 s 536 82442 618 82470 4 in2_53
rlabel metal1 s 1176 82246 1204 82274 4 rwl0_53
rlabel metal1 s 1176 82020 1204 82048 4 rwl1_53
rlabel metal1 s 1176 82372 1204 82400 4 wwl0_53
rlabel metal1 s 56 83900 126 83928 4 in0_54
rlabel metal1 s 234 83754 318 83782 4 in1_54
rlabel metal1 s 536 83634 618 83662 4 in2_54
rlabel metal1 s 1176 83830 1204 83858 4 rwl0_54
rlabel metal1 s 1176 84056 1204 84084 4 rwl1_54
rlabel metal1 s 1176 83704 1204 83732 4 wwl0_54
rlabel metal1 s 56 85252 126 85280 4 in0_55
rlabel metal1 s 234 85398 318 85426 4 in1_55
rlabel metal1 s 536 85518 618 85546 4 in2_55
rlabel metal1 s 1176 85322 1204 85350 4 rwl0_55
rlabel metal1 s 1176 85096 1204 85124 4 rwl1_55
rlabel metal1 s 1176 85448 1204 85476 4 wwl0_55
rlabel metal1 s 56 86976 126 87004 4 in0_56
rlabel metal1 s 234 86830 318 86858 4 in1_56
rlabel metal1 s 536 86710 618 86738 4 in2_56
rlabel metal1 s 1176 86906 1204 86934 4 rwl0_56
rlabel metal1 s 1176 87132 1204 87160 4 rwl1_56
rlabel metal1 s 1176 86780 1204 86808 4 wwl0_56
rlabel metal1 s 56 88328 126 88356 4 in0_57
rlabel metal1 s 234 88474 318 88502 4 in1_57
rlabel metal1 s 536 88594 618 88622 4 in2_57
rlabel metal1 s 1176 88398 1204 88426 4 rwl0_57
rlabel metal1 s 1176 88172 1204 88200 4 rwl1_57
rlabel metal1 s 1176 88524 1204 88552 4 wwl0_57
rlabel metal1 s 56 90052 126 90080 4 in0_58
rlabel metal1 s 234 89906 318 89934 4 in1_58
rlabel metal1 s 536 89786 618 89814 4 in2_58
rlabel metal1 s 1176 89982 1204 90010 4 rwl0_58
rlabel metal1 s 1176 90208 1204 90236 4 rwl1_58
rlabel metal1 s 1176 89856 1204 89884 4 wwl0_58
rlabel metal1 s 56 91404 126 91432 4 in0_59
rlabel metal1 s 234 91550 318 91578 4 in1_59
rlabel metal1 s 536 91670 618 91698 4 in2_59
rlabel metal1 s 1176 91474 1204 91502 4 rwl0_59
rlabel metal1 s 1176 91248 1204 91276 4 rwl1_59
rlabel metal1 s 1176 91600 1204 91628 4 wwl0_59
rlabel metal1 s 56 93128 126 93156 4 in0_60
rlabel metal1 s 234 92982 318 93010 4 in1_60
rlabel metal1 s 536 92862 618 92890 4 in2_60
rlabel metal1 s 1176 93058 1204 93086 4 rwl0_60
rlabel metal1 s 1176 93284 1204 93312 4 rwl1_60
rlabel metal1 s 1176 92932 1204 92960 4 wwl0_60
rlabel metal1 s 56 94480 126 94508 4 in0_61
rlabel metal1 s 234 94626 318 94654 4 in1_61
rlabel metal1 s 536 94746 618 94774 4 in2_61
rlabel metal1 s 1176 94550 1204 94578 4 rwl0_61
rlabel metal1 s 1176 94324 1204 94352 4 rwl1_61
rlabel metal1 s 1176 94676 1204 94704 4 wwl0_61
rlabel metal1 s 56 96204 126 96232 4 in0_62
rlabel metal1 s 234 96058 318 96086 4 in1_62
rlabel metal1 s 536 95938 618 95966 4 in2_62
rlabel metal1 s 1176 96134 1204 96162 4 rwl0_62
rlabel metal1 s 1176 96360 1204 96388 4 rwl1_62
rlabel metal1 s 1176 96008 1204 96036 4 wwl0_62
rlabel metal1 s 56 97556 126 97584 4 in0_63
rlabel metal1 s 234 97702 318 97730 4 in1_63
rlabel metal1 s 536 97822 618 97850 4 in2_63
rlabel metal1 s 1176 97626 1204 97654 4 rwl0_63
rlabel metal1 s 1176 97400 1204 97428 4 rwl1_63
rlabel metal1 s 1176 97752 1204 97780 4 wwl0_63
rlabel metal3 s 1138 10729 1270 10803 4 vdd
rlabel metal3 s 1138 69173 1270 69247 4 vdd
rlabel metal3 s 1138 41489 1270 41563 4 vdd
rlabel metal3 s 1138 90705 1270 90779 4 vdd
rlabel metal3 s 1138 16881 1270 16955 4 vdd
rlabel metal3 s 1138 56869 1270 56943 4 vdd
rlabel metal3 s 1204 90742 1204 90742 4 vdd
rlabel metal3 s 1138 93781 1270 93855 4 vdd
rlabel metal3 s 1138 38413 1270 38487 4 vdd
rlabel metal3 s 1138 35337 1270 35411 4 vdd
rlabel metal3 s 1138 44565 1270 44639 4 vdd
rlabel metal3 s 1204 44602 1204 44602 4 vdd
rlabel metal3 s 1138 26109 1270 26183 4 vdd
rlabel metal3 s 1138 4577 1270 4651 4 vdd
rlabel metal3 s 1138 84553 1270 84627 4 vdd
rlabel metal3 s 1138 75325 1270 75399 4 vdd
rlabel metal3 s 1138 23033 1270 23107 4 vdd
rlabel metal3 s 1138 47641 1270 47715 4 vdd
rlabel metal3 s 1138 13805 1270 13879 4 vdd
rlabel metal3 s 1138 72249 1270 72323 4 vdd
rlabel metal3 s 1138 7653 1270 7727 4 vdd
rlabel metal3 s 1138 50717 1270 50791 4 vdd
rlabel metal3 s 1204 50754 1204 50754 4 vdd
rlabel metal3 s 1138 63021 1270 63095 4 vdd
rlabel metal3 s 1138 29185 1270 29259 4 vdd
rlabel metal3 s 1138 19957 1270 20031 4 vdd
rlabel metal3 s 1138 32261 1270 32335 4 vdd
rlabel metal3 s 1138 1501 1270 1575 4 vdd
rlabel metal3 s 1204 1538 1204 1538 4 vdd
rlabel metal3 s 1138 96857 1270 96931 4 vdd
rlabel metal3 s 1138 87629 1270 87703 4 vdd
rlabel metal3 s 1138 53793 1270 53867 4 vdd
rlabel metal3 s 1204 53830 1204 53830 4 vdd
rlabel metal3 s 1138 66097 1270 66171 4 vdd
rlabel metal3 s 1138 59945 1270 60019 4 vdd
rlabel metal3 s 1138 81477 1270 81551 4 vdd
rlabel metal3 s 1138 78401 1270 78475 4 vdd
rlabel metal3 s 1204 10766 1204 10766 4 vdd
rlabel metal3 s 1138 33799 1270 33873 4 gnd
rlabel metal3 s 1138 52255 1270 52329 4 gnd
rlabel metal3 s 1138 70711 1270 70785 4 gnd
rlabel metal3 s 1138 21495 1270 21569 4 gnd
rlabel metal3 s 1138 49179 1270 49253 4 gnd
rlabel metal3 s 1138 79939 1270 80013 4 gnd
rlabel metal3 s 1138 58407 1270 58481 4 gnd
rlabel metal3 s 1138 76863 1270 76937 4 gnd
rlabel metal3 s 1138 86091 1270 86165 4 gnd
rlabel metal3 s 1138 27647 1270 27721 4 gnd
rlabel metal3 s 1138 67635 1270 67709 4 gnd
rlabel metal3 s 1138 46103 1270 46177 4 gnd
rlabel metal3 s 1138 83015 1270 83089 4 gnd
rlabel metal3 s 1138 6115 1270 6189 4 gnd
rlabel metal3 s 1138 89167 1270 89241 4 gnd
rlabel metal3 s 1138 55331 1270 55405 4 gnd
rlabel metal3 s 1138 36875 1270 36949 4 gnd
rlabel metal3 s 1138 3039 1270 3113 4 gnd
rlabel metal3 s 1138 30723 1270 30797 4 gnd
rlabel metal3 s 1138 92243 1270 92317 4 gnd
rlabel metal3 s 1138 9191 1270 9265 4 gnd
rlabel metal3 s 1138 95319 1270 95393 4 gnd
rlabel metal3 s 1138 15343 1270 15417 4 gnd
rlabel metal3 s 1138 39951 1270 40025 4 gnd
rlabel metal3 s 1138 12267 1270 12341 4 gnd
rlabel metal3 s 1138 98395 1270 98469 4 gnd
rlabel metal3 s 1138 -37 1270 37 4 gnd
rlabel metal3 s 1138 73787 1270 73861 4 gnd
rlabel metal3 s 1138 24571 1270 24645 4 gnd
rlabel metal3 s 1138 43027 1270 43101 4 gnd
rlabel metal3 s 1138 18419 1270 18493 4 gnd
rlabel metal3 s 1138 64559 1270 64633 4 gnd
rlabel metal3 s 1138 61483 1270 61557 4 gnd
<< properties >>
string FIXED_BBOX 1138 -37 1270 0
string GDS_FILE sram_0rw2r1w_32_128_sky130A.gds
string GDS_END 3236724
string GDS_START 3124954
<< end >>
