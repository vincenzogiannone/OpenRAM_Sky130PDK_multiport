magic
tech sky130A
timestamp 1642866255
<< nwell >>
rect 0 488 747 808
<< nmos >>
rect 47 115 62 215
rect 95 115 110 215
rect 143 115 158 215
rect 191 115 206 215
rect 239 115 254 215
rect 287 115 302 215
rect 389 115 404 215
rect 437 115 452 215
rect 485 115 500 215
rect 537 115 552 157
rect 637 115 652 157
rect 685 115 700 157
<< pmos >>
rect 47 506 62 548
rect 95 506 110 548
rect 143 506 158 548
rect 191 506 206 548
rect 239 506 254 548
rect 287 506 302 548
rect 389 506 404 548
rect 437 506 452 548
rect 485 506 500 548
rect 537 506 552 641
rect 637 506 652 641
rect 685 506 700 641
<< ndiff >>
rect 18 198 47 215
rect 18 181 22 198
rect 39 181 47 198
rect 18 149 47 181
rect 18 132 22 149
rect 39 132 47 149
rect 18 115 47 132
rect 62 115 95 215
rect 110 115 143 215
rect 158 198 191 215
rect 158 181 166 198
rect 183 181 191 198
rect 158 149 191 181
rect 158 132 166 149
rect 183 132 191 149
rect 158 115 191 132
rect 206 115 239 215
rect 254 115 287 215
rect 302 198 331 215
rect 302 181 310 198
rect 327 181 331 198
rect 302 149 331 181
rect 302 132 310 149
rect 327 132 331 149
rect 302 115 331 132
rect 360 198 389 215
rect 360 181 364 198
rect 381 181 389 198
rect 360 149 389 181
rect 360 132 364 149
rect 381 132 389 149
rect 360 115 389 132
rect 404 115 437 215
rect 452 115 485 215
rect 500 198 529 215
rect 500 181 508 198
rect 525 181 529 198
rect 500 157 529 181
rect 500 149 537 157
rect 500 132 508 149
rect 525 132 537 149
rect 500 115 537 132
rect 552 144 581 157
rect 552 127 560 144
rect 577 127 581 144
rect 552 115 581 127
rect 608 144 637 157
rect 608 127 612 144
rect 629 127 637 144
rect 608 115 637 127
rect 652 144 685 157
rect 652 127 660 144
rect 677 127 685 144
rect 652 115 685 127
rect 700 144 729 157
rect 700 127 708 144
rect 725 127 729 144
rect 700 115 729 127
<< pdiff >>
rect 508 624 537 641
rect 508 607 512 624
rect 529 607 537 624
rect 508 582 537 607
rect 508 565 512 582
rect 529 565 537 582
rect 508 548 537 565
rect 18 535 47 548
rect 18 518 22 535
rect 39 518 47 535
rect 18 506 47 518
rect 62 535 95 548
rect 62 518 70 535
rect 87 518 95 535
rect 62 506 95 518
rect 110 535 143 548
rect 110 518 118 535
rect 135 518 143 535
rect 110 506 143 518
rect 158 535 191 548
rect 158 518 166 535
rect 183 518 191 535
rect 158 506 191 518
rect 206 535 239 548
rect 206 518 214 535
rect 231 518 239 535
rect 206 506 239 518
rect 254 535 287 548
rect 254 518 262 535
rect 279 518 287 535
rect 254 506 287 518
rect 302 535 331 548
rect 302 518 310 535
rect 327 518 331 535
rect 302 506 331 518
rect 360 535 389 548
rect 360 518 364 535
rect 381 518 389 535
rect 360 506 389 518
rect 404 535 437 548
rect 404 518 412 535
rect 429 518 437 535
rect 404 506 437 518
rect 452 535 485 548
rect 452 518 460 535
rect 477 518 485 535
rect 452 506 485 518
rect 500 540 537 548
rect 500 523 512 540
rect 529 523 537 540
rect 500 506 537 523
rect 552 624 581 641
rect 552 607 560 624
rect 577 607 581 624
rect 552 582 581 607
rect 552 565 560 582
rect 577 565 581 582
rect 552 540 581 565
rect 552 523 560 540
rect 577 523 581 540
rect 552 506 581 523
rect 608 624 637 641
rect 608 607 612 624
rect 629 607 637 624
rect 608 582 637 607
rect 608 565 612 582
rect 629 565 637 582
rect 608 540 637 565
rect 608 523 612 540
rect 629 523 637 540
rect 608 506 637 523
rect 652 624 685 641
rect 652 607 660 624
rect 677 607 685 624
rect 652 582 685 607
rect 652 565 660 582
rect 677 565 685 582
rect 652 540 685 565
rect 652 523 660 540
rect 677 523 685 540
rect 652 506 685 523
rect 700 624 729 641
rect 700 607 708 624
rect 725 607 729 624
rect 700 582 729 607
rect 700 565 708 582
rect 725 565 729 582
rect 700 540 729 565
rect 700 523 708 540
rect 725 523 729 540
rect 700 506 729 523
<< ndiffc >>
rect 22 181 39 198
rect 22 132 39 149
rect 166 181 183 198
rect 166 132 183 149
rect 310 181 327 198
rect 310 132 327 149
rect 364 181 381 198
rect 364 132 381 149
rect 508 181 525 198
rect 508 132 525 149
rect 560 127 577 144
rect 612 127 629 144
rect 660 127 677 144
rect 708 127 725 144
<< pdiffc >>
rect 512 607 529 624
rect 512 565 529 582
rect 22 518 39 535
rect 70 518 87 535
rect 118 518 135 535
rect 166 518 183 535
rect 214 518 231 535
rect 262 518 279 535
rect 310 518 327 535
rect 364 518 381 535
rect 412 518 429 535
rect 460 518 477 535
rect 512 523 529 540
rect 560 607 577 624
rect 560 565 577 582
rect 560 523 577 540
rect 612 607 629 624
rect 612 565 629 582
rect 612 523 629 540
rect 660 607 677 624
rect 660 565 677 582
rect 660 523 677 540
rect 708 607 725 624
rect 708 565 725 582
rect 708 523 725 540
<< psubdiff >>
rect 120 9 156 21
rect 120 -9 129 9
rect 147 -9 156 9
rect 120 -21 156 -9
rect 277 9 313 21
rect 277 -9 286 9
rect 304 -9 313 9
rect 277 -21 313 -9
rect 434 9 470 21
rect 434 -9 443 9
rect 461 -9 470 9
rect 434 -21 470 -9
rect 591 9 627 21
rect 591 -9 600 9
rect 618 -9 627 9
rect 591 -21 627 -9
<< nsubdiff >>
rect 120 766 156 778
rect 120 748 129 766
rect 147 748 156 766
rect 120 736 156 748
rect 277 766 313 778
rect 277 748 286 766
rect 304 748 313 766
rect 277 736 313 748
rect 434 766 470 778
rect 434 748 443 766
rect 461 748 470 766
rect 434 736 470 748
rect 591 766 627 778
rect 591 748 600 766
rect 618 748 627 766
rect 591 736 627 748
<< psubdiffcont >>
rect 129 -9 147 9
rect 286 -9 304 9
rect 443 -9 461 9
rect 600 -9 618 9
<< nsubdiffcont >>
rect 129 748 147 766
rect 286 748 304 766
rect 443 748 461 766
rect 600 748 618 766
<< poly >>
rect 537 641 552 654
rect 637 641 652 654
rect 685 641 700 654
rect 47 548 62 561
rect 95 548 110 561
rect 143 548 158 561
rect 191 548 206 561
rect 239 548 254 561
rect 287 548 302 561
rect 389 548 404 561
rect 437 548 452 561
rect 485 548 500 561
rect 47 489 62 506
rect 35 481 62 489
rect 35 464 40 481
rect 57 464 62 481
rect 35 456 62 464
rect 95 461 110 506
rect 47 215 62 456
rect 83 453 110 461
rect 83 436 88 453
rect 105 436 110 453
rect 83 428 110 436
rect 143 433 158 506
rect 95 215 110 428
rect 131 425 158 433
rect 131 408 136 425
rect 153 408 158 425
rect 131 400 158 408
rect 191 405 206 506
rect 143 215 158 400
rect 179 397 206 405
rect 179 380 184 397
rect 201 380 206 397
rect 179 372 206 380
rect 239 377 254 506
rect 191 215 206 372
rect 227 369 254 377
rect 227 352 232 369
rect 249 352 254 369
rect 227 344 254 352
rect 287 349 302 506
rect 239 215 254 344
rect 275 341 302 349
rect 275 324 280 341
rect 297 324 302 341
rect 275 316 302 324
rect 389 321 404 506
rect 287 215 302 316
rect 377 313 404 321
rect 377 296 382 313
rect 399 296 404 313
rect 377 288 404 296
rect 437 293 452 506
rect 389 215 404 288
rect 425 285 452 293
rect 425 268 430 285
rect 447 268 452 285
rect 425 260 452 268
rect 485 265 500 506
rect 537 319 552 506
rect 525 311 552 319
rect 525 294 530 311
rect 547 294 552 311
rect 525 286 552 294
rect 437 215 452 260
rect 473 257 500 265
rect 473 240 478 257
rect 495 240 500 257
rect 473 232 500 240
rect 485 215 500 232
rect 537 157 552 286
rect 637 420 652 506
rect 685 489 700 506
rect 673 481 700 489
rect 673 464 678 481
rect 695 464 700 481
rect 673 456 700 464
rect 637 412 664 420
rect 637 395 642 412
rect 659 395 664 412
rect 637 387 664 395
rect 637 157 652 387
rect 685 157 700 456
rect 47 102 62 115
rect 95 102 110 115
rect 143 102 158 115
rect 191 102 206 115
rect 239 102 254 115
rect 287 102 302 115
rect 389 102 404 115
rect 437 102 452 115
rect 485 102 500 115
rect 537 102 552 115
rect 637 102 652 115
rect 685 102 700 115
<< polycont >>
rect 40 464 57 481
rect 88 436 105 453
rect 136 408 153 425
rect 184 380 201 397
rect 232 352 249 369
rect 280 324 297 341
rect 382 296 399 313
rect 430 268 447 285
rect 530 294 547 311
rect 478 240 495 257
rect 678 464 695 481
rect 642 395 659 412
<< locali >>
rect 129 766 147 774
rect 286 766 304 774
rect 443 766 461 774
rect 600 766 618 774
rect 70 748 129 766
rect 147 748 286 766
rect 304 748 443 766
rect 461 748 600 766
rect 618 748 677 766
rect 70 548 87 748
rect 129 740 147 748
rect 166 548 183 748
rect 262 740 304 748
rect 412 740 461 748
rect 262 548 279 740
rect 412 548 429 740
rect 512 641 529 748
rect 600 740 618 748
rect 660 641 677 748
rect 508 624 532 641
rect 508 607 512 624
rect 529 607 532 624
rect 508 582 532 607
rect 508 565 512 582
rect 529 565 532 582
rect 18 535 42 548
rect 18 518 22 535
rect 39 518 42 535
rect 18 506 42 518
rect 67 535 90 548
rect 67 518 70 535
rect 87 518 90 535
rect 67 506 90 518
rect 115 535 138 548
rect 115 518 118 535
rect 135 518 138 535
rect 115 506 138 518
rect 163 535 186 548
rect 163 518 166 535
rect 183 518 186 535
rect 163 506 186 518
rect 211 535 234 548
rect 211 518 214 535
rect 231 518 234 535
rect 211 506 234 518
rect 259 535 282 548
rect 259 518 262 535
rect 279 518 282 535
rect 259 506 282 518
rect 307 535 331 548
rect 307 518 310 535
rect 327 518 331 535
rect 307 506 331 518
rect 360 535 384 548
rect 360 518 364 535
rect 381 518 384 535
rect 360 506 384 518
rect 409 535 432 548
rect 409 518 412 535
rect 429 518 432 535
rect 409 506 432 518
rect 457 535 480 548
rect 457 518 460 535
rect 477 518 480 535
rect 457 506 480 518
rect 508 540 532 565
rect 508 523 512 540
rect 529 523 532 540
rect 508 506 532 523
rect 557 624 581 641
rect 557 607 560 624
rect 577 607 581 624
rect 557 582 581 607
rect 557 565 560 582
rect 577 565 581 582
rect 557 540 581 565
rect 557 523 560 540
rect 577 523 581 540
rect 557 506 581 523
rect 40 481 57 489
rect 40 456 57 464
rect 348 467 364 484
rect 88 453 105 461
rect 88 428 105 436
rect 136 425 153 433
rect 136 400 153 408
rect 184 397 201 405
rect 307 388 331 405
rect 184 372 201 380
rect 232 369 249 377
rect 232 344 249 352
rect 280 341 297 349
rect 280 316 297 324
rect 314 299 331 388
rect 22 282 331 299
rect 22 215 39 282
rect 348 265 365 467
rect 463 327 480 506
rect 382 313 399 321
rect 463 311 547 327
rect 463 310 530 311
rect 382 288 399 296
rect 310 248 365 265
rect 430 285 447 293
rect 530 286 547 294
rect 564 304 581 506
rect 608 624 632 641
rect 608 607 612 624
rect 629 607 632 624
rect 608 582 632 607
rect 608 565 612 582
rect 629 565 632 582
rect 608 540 632 565
rect 608 523 612 540
rect 629 523 632 540
rect 608 506 632 523
rect 657 624 680 641
rect 657 607 660 624
rect 677 607 680 624
rect 657 582 680 607
rect 657 565 660 582
rect 677 565 680 582
rect 657 540 680 565
rect 657 523 660 540
rect 677 523 680 540
rect 657 506 680 523
rect 705 624 729 641
rect 705 607 708 624
rect 725 607 729 624
rect 705 582 729 607
rect 705 565 708 582
rect 725 565 729 582
rect 705 540 729 565
rect 705 523 708 540
rect 725 523 729 540
rect 705 506 729 523
rect 608 365 625 506
rect 678 481 695 489
rect 678 456 695 464
rect 712 438 729 506
rect 642 412 659 420
rect 642 387 659 395
rect 564 287 567 304
rect 430 260 447 268
rect 478 257 495 265
rect 310 215 327 248
rect 478 232 495 240
rect 18 198 42 215
rect 18 181 22 198
rect 39 181 42 198
rect 18 149 42 181
rect 18 132 22 149
rect 39 132 42 149
rect 18 115 42 132
rect 163 198 186 215
rect 163 181 166 198
rect 183 181 186 198
rect 163 149 186 181
rect 163 132 166 149
rect 183 132 186 149
rect 163 115 186 132
rect 307 198 331 215
rect 307 181 310 198
rect 327 181 331 198
rect 307 149 331 181
rect 307 132 310 149
rect 327 132 331 149
rect 307 115 331 132
rect 360 198 384 215
rect 360 181 364 198
rect 381 181 384 198
rect 360 149 384 181
rect 360 132 364 149
rect 381 132 384 149
rect 360 115 384 132
rect 505 198 529 215
rect 505 181 508 198
rect 525 181 529 198
rect 505 149 529 181
rect 564 157 581 287
rect 505 132 508 149
rect 525 132 529 149
rect 505 115 529 132
rect 557 144 581 157
rect 557 127 560 144
rect 577 127 581 144
rect 557 115 581 127
rect 608 157 625 348
rect 712 157 729 421
rect 608 144 632 157
rect 608 127 612 144
rect 629 127 632 144
rect 608 115 632 127
rect 657 144 680 157
rect 657 127 660 144
rect 677 127 680 144
rect 657 115 680 127
rect 705 144 729 157
rect 705 127 708 144
rect 725 127 729 144
rect 705 115 729 127
rect 129 9 147 21
rect 166 9 183 115
rect 286 9 304 21
rect 443 9 461 21
rect 508 9 525 115
rect 600 9 618 21
rect 660 9 677 115
rect 70 -9 129 9
rect 147 -9 286 9
rect 304 -9 443 9
rect 461 -9 600 9
rect 618 -9 677 9
rect 129 -21 147 -9
rect 286 -21 304 -9
rect 443 -21 461 -9
rect 600 -21 618 -9
<< viali >>
rect 129 748 147 766
rect 286 748 304 766
rect 443 748 461 766
rect 600 748 618 766
rect 22 518 39 535
rect 118 518 135 535
rect 214 518 231 535
rect 310 518 327 535
rect 364 518 381 535
rect 460 518 477 535
rect 40 464 57 481
rect 364 467 381 484
rect 88 436 105 453
rect 136 408 153 425
rect 184 380 201 397
rect 290 388 307 405
rect 232 352 249 369
rect 280 324 297 341
rect 382 296 399 313
rect 530 294 547 311
rect 678 464 695 481
rect 712 421 729 438
rect 642 395 659 412
rect 608 348 625 365
rect 567 287 584 304
rect 430 268 447 285
rect 478 240 495 257
rect 364 132 381 149
rect 129 -9 147 9
rect 286 -9 304 9
rect 443 -9 461 9
rect 600 -9 618 9
<< metal1 >>
rect 0 766 747 772
rect 0 748 129 766
rect 147 748 286 766
rect 304 748 443 766
rect 461 748 600 766
rect 618 748 747 766
rect 0 742 747 748
rect 19 535 138 541
rect 19 518 22 535
rect 39 527 118 535
rect 39 518 42 527
rect 19 512 42 518
rect 115 518 118 527
rect 135 518 138 535
rect 115 512 138 518
rect 211 535 330 541
rect 211 518 214 535
rect 231 527 310 535
rect 231 518 234 527
rect 211 512 234 518
rect 307 518 310 527
rect 327 518 330 535
rect 307 512 330 518
rect 361 535 480 541
rect 361 518 364 535
rect 381 527 460 535
rect 381 518 384 527
rect 361 512 384 518
rect 457 518 460 527
rect 477 518 480 535
rect 457 512 480 518
rect 124 494 138 512
rect 36 481 63 488
rect 36 471 40 481
rect 35 464 40 471
rect 57 464 63 481
rect 124 480 253 494
rect 35 457 63 464
rect 84 453 111 460
rect 84 443 88 453
rect 83 436 88 443
rect 105 436 111 453
rect 83 429 111 436
rect 132 425 159 432
rect 132 415 136 425
rect 131 408 136 415
rect 153 408 159 425
rect 131 401 159 408
rect 239 418 253 480
rect 316 490 330 512
rect 316 487 384 490
rect 316 484 698 487
rect 316 476 364 484
rect 361 467 364 476
rect 381 481 698 484
rect 381 473 678 481
rect 381 467 384 473
rect 361 461 384 467
rect 675 464 678 473
rect 695 464 698 481
rect 675 458 698 464
rect 709 438 732 444
rect 709 421 712 438
rect 729 424 747 438
rect 729 421 732 424
rect 239 412 662 418
rect 709 415 732 421
rect 239 405 642 412
rect 239 404 290 405
rect 180 397 207 404
rect 180 387 184 397
rect 179 380 184 387
rect 201 380 207 397
rect 287 388 290 404
rect 307 404 642 405
rect 307 388 310 404
rect 639 395 642 404
rect 659 395 662 412
rect 639 389 662 395
rect 287 382 310 388
rect 179 373 207 380
rect 228 369 255 376
rect 228 359 232 369
rect 227 352 232 359
rect 249 352 255 369
rect 227 345 255 352
rect 605 365 628 371
rect 605 348 608 365
rect 625 351 747 365
rect 625 348 628 351
rect 276 341 303 348
rect 605 342 628 348
rect 276 331 280 341
rect 275 324 280 331
rect 297 324 303 341
rect 275 317 303 324
rect 378 313 405 320
rect 378 303 382 313
rect 377 296 382 303
rect 399 296 405 313
rect 377 289 405 296
rect 527 311 550 317
rect 527 294 530 311
rect 547 294 550 311
rect 426 285 453 292
rect 527 288 550 294
rect 426 275 430 285
rect 425 268 430 275
rect 447 268 453 285
rect 425 261 453 268
rect 474 257 501 264
rect 474 247 478 257
rect 473 240 478 247
rect 495 240 501 257
rect 473 233 501 240
rect 536 155 550 288
rect 564 304 587 310
rect 564 287 567 304
rect 584 290 747 304
rect 584 287 587 290
rect 564 281 587 287
rect 361 149 550 155
rect 361 132 364 149
rect 381 141 550 149
rect 381 132 384 141
rect 361 126 384 132
rect 0 9 747 15
rect 0 -9 129 9
rect 147 -9 286 9
rect 304 -9 443 9
rect 461 -9 600 9
rect 618 -9 747 9
rect 0 -15 747 -9
<< labels >>
flabel metal1 35 464 35 464 0 FreeSans 80 0 0 0 A0
port 0 nsew
flabel metal1 83 435 83 435 0 FreeSans 80 0 0 0 B0
port 1 nsew
flabel metal1 131 405 131 405 0 FreeSans 80 0 0 0 C0
port 2 nsew
flabel metal1 179 378 179 378 0 FreeSans 80 0 0 0 A1
port 3 nsew
flabel metal1 227 350 227 350 0 FreeSans 80 0 0 0 B1
port 4 nsew
flabel metal1 275 322 275 322 0 FreeSans 80 0 0 0 C1
port 5 nsew
flabel metal1 377 296 377 296 0 FreeSans 80 0 0 0 A2
port 6 nsew
flabel metal1 425 268 425 268 0 FreeSans 80 0 0 0 B2
port 7 nsew
flabel metal1 473 239 473 239 0 FreeSans 80 0 0 0 C2
port 8 nsew
flabel metal1 738 431 738 431 0 FreeSans 80 0 0 0 OUT1
port 9 nsew
flabel metal1 737 357 737 357 0 FreeSans 80 0 0 0 OUT0
port 10 nsew
flabel metal1 736 296 736 296 0 FreeSans 80 0 0 0 OUT2
port 11 nsew
flabel metal1 355 756 355 756 0 FreeSans 80 0 0 0 vdd
port 12 nsew
flabel metal1 348 0 348 0 0 FreeSans 80 0 0 0 gnd
port 13 nsew
flabel metal1 179 482 179 482 0 FreeSans 80 0 0 0 net3
flabel ndiff 217 158 217 158 0 FreeSans 80 0 0 0 net4
flabel ndiff 266 157 266 157 0 FreeSans 80 0 0 0 net5
flabel metal1 326 480 326 480 0 FreeSans 80 0 0 0 net6
flabel ndiff 126 157 126 157 0 FreeSans 80 0 0 0 net1
flabel ndiff 79 153 79 153 0 FreeSans 80 0 0 0 net2
flabel ndiff 466 170 466 170 0 FreeSans 80 0 0 0 net7
flabel ndiff 420 168 420 168 0 FreeSans 80 0 0 0 net8
flabel locali 475 375 475 375 0 FreeSans 80 0 0 0 net9
<< properties >>
string FIXED_BBOX 0 0 747 757
<< end >>
