magic
tech sky130A
magscale 1 2
timestamp 1643671299
<< checkpaint >>
rect -1263 -1302 2742 2176
<< via1 >>
rect 715 812 767 864
rect 715 -26 767 26
<< metal2 >>
rect 721 866 761 872
rect 0 328 28 838
rect 721 804 761 810
rect 0 0 28 272
rect 180 232 234 260
rect 1260 228 1314 256
rect 721 28 761 34
rect 721 -34 761 -28
<< via2 >>
rect 713 864 769 866
rect 713 812 715 864
rect 715 812 767 864
rect 767 812 769 864
rect 713 810 769 812
rect -1 272 55 328
rect 713 26 769 28
rect 713 -26 715 26
rect 715 -26 767 26
rect 767 -26 769 26
rect 713 -28 769 -26
<< metal3 >>
rect 711 866 771 868
rect 711 810 713 866
rect 769 810 771 866
rect 711 808 771 810
rect -3 328 1482 330
rect -3 272 -1 328
rect 55 272 1482 328
rect -3 270 1482 272
rect 711 28 771 30
rect 711 -28 713 28
rect 769 -28 771 28
rect 711 -30 771 -28
use contact_18  contact_18_0
timestamp 1643671299
transform 1 0 -3 0 1 270
box 0 0 1 1
use contact_18  contact_18_1
timestamp 1643671299
transform 1 0 711 0 1 -30
box 0 0 1 1
use contact_17  contact_17_0
timestamp 1643671299
transform 1 0 726 0 1 -15
box 0 0 1 1
use contact_18  contact_18_2
timestamp 1643671299
transform 1 0 711 0 1 808
box 0 0 1 1
use contact_17  contact_17_1
timestamp 1643671299
transform 1 0 726 0 1 823
box 0 0 1 1
use dff  dff_0
timestamp 1643671299
transform 1 0 0 0 1 0
box 0 -42 1482 916
<< labels >>
rlabel metal3 s 711 808 771 868 4 vdd
rlabel metal3 s 711 -30 771 30 4 gnd
rlabel metal2 s 180 232 234 260 4 din_0
rlabel metal2 s 1260 228 1314 256 4 dout_0
rlabel metal3 s 0 270 1482 330 4 clk
<< properties >>
string FIXED_BBOX 711 -30 771 0
string GDS_FILE sram_0rw2r1w_16_32_sky130A.gds
string GDS_END 1233572
string GDS_START 1232080
<< end >>
