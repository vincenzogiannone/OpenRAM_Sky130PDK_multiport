magic
tech sky130A
magscale 1 2
timestamp 1643671299
<< checkpaint >>
rect -1271 -1302 5952 25926
<< viali >>
rect 2115 23887 2149 23921
rect 2115 22263 2149 22297
rect 2115 20807 2149 20841
rect 2115 19183 2149 19217
rect 2115 14651 2149 14685
rect 2115 13027 2149 13061
rect 2115 11571 2149 11605
rect 2115 9947 2149 9981
rect 2115 5415 2149 5449
rect 2115 3791 2149 3825
rect 2115 2335 2149 2369
rect 2115 711 2149 745
<< metal1 >>
rect 2103 23919 2106 23927
rect 2077 23889 2106 23919
rect 2103 23881 2106 23889
rect 2158 23919 2161 23927
rect 2158 23889 2188 23919
rect 2158 23881 2161 23889
rect 3058 23730 4142 23758
rect 2854 23674 4046 23702
rect 2514 23618 3950 23646
rect 4282 23616 4648 23644
rect 3058 23562 3746 23590
rect 2854 23506 3650 23534
rect 4364 23494 4648 23522
rect 2446 23450 3554 23478
rect 3058 23394 3458 23422
rect 2854 23338 3362 23366
rect 4572 23348 4648 23376
rect 2378 23282 3266 23310
rect 2103 22295 2106 22303
rect 2077 22265 2106 22295
rect 2103 22257 2106 22265
rect 2158 22295 2161 22303
rect 2158 22265 2188 22295
rect 2158 22257 2161 22265
rect 2446 22110 3266 22138
rect 2786 22054 3362 22082
rect 4572 22044 4648 22072
rect 3058 21998 3458 22026
rect 2514 21942 3554 21970
rect 2786 21886 3650 21914
rect 4364 21898 4648 21926
rect 3058 21830 3746 21858
rect 2582 21774 3950 21802
rect 4282 21776 4648 21804
rect 2786 21718 4046 21746
rect 3058 21662 4142 21690
rect 381 20810 561 20838
rect 2103 20839 2106 20847
rect 2077 20809 2106 20839
rect 2103 20801 2106 20809
rect 2158 20839 2161 20847
rect 2158 20809 2188 20839
rect 2158 20801 2161 20809
rect 3058 20702 4142 20730
rect 2786 20646 4046 20674
rect 2378 20590 3950 20618
rect 4282 20588 4648 20616
rect 3058 20534 3746 20562
rect 2718 20478 3650 20506
rect 4364 20466 4648 20494
rect 2582 20422 3554 20450
rect 3058 20366 3458 20394
rect 2718 20310 3362 20338
rect 4572 20320 4648 20348
rect 2514 20254 3266 20282
rect 313 19186 493 19214
rect 2103 19215 2106 19223
rect 2077 19185 2106 19215
rect 2103 19177 2106 19185
rect 2158 19215 2161 19223
rect 2158 19185 2188 19215
rect 2158 19177 2161 19185
rect 2582 19082 3266 19110
rect 2650 19026 3362 19054
rect 4572 19016 4648 19044
rect 3058 18970 3458 18998
rect 2378 18914 3554 18942
rect 2718 18858 3650 18886
rect 4364 18870 4648 18898
rect 3058 18802 3746 18830
rect 2446 18746 3950 18774
rect 4282 18748 4648 18776
rect 2718 18690 4046 18718
rect 3058 18634 4142 18662
rect 3058 17674 4142 17702
rect 2650 17618 4046 17646
rect 2514 17562 3950 17590
rect 4282 17560 4648 17588
rect 3058 17506 3746 17534
rect 2650 17450 3650 17478
rect 4364 17438 4648 17466
rect 2446 17394 3554 17422
rect 3058 17338 3458 17366
rect 2650 17282 3362 17310
rect 4572 17292 4648 17320
rect 2378 17226 3266 17254
rect 2446 16054 3266 16082
rect 2854 15998 3362 16026
rect 4572 15988 4648 16016
rect 2990 15942 3458 15970
rect 2514 15886 3554 15914
rect 2854 15830 3650 15858
rect 4364 15842 4648 15870
rect 2990 15774 3746 15802
rect 2582 15718 3950 15746
rect 4282 15720 4648 15748
rect 2854 15662 4046 15690
rect 2990 15606 4142 15634
rect 2103 14683 2106 14691
rect 2077 14653 2106 14683
rect 2103 14645 2106 14653
rect 2158 14683 2161 14691
rect 2158 14653 2188 14683
rect 2158 14645 2161 14653
rect 2990 14646 4142 14674
rect 2854 14590 4046 14618
rect 2378 14534 3950 14562
rect 4282 14532 4648 14560
rect 2990 14478 3746 14506
rect 2786 14422 3650 14450
rect 4364 14410 4648 14438
rect 2582 14366 3554 14394
rect 2990 14310 3458 14338
rect 2786 14254 3362 14282
rect 4572 14264 4648 14292
rect 2514 14198 3266 14226
rect 2103 13059 2106 13067
rect 2077 13029 2106 13059
rect 2103 13021 2106 13029
rect 2158 13059 2161 13067
rect 2158 13029 2188 13059
rect 2158 13021 2161 13029
rect 2582 13026 3266 13054
rect 2718 12970 3362 12998
rect 4572 12960 4648 12988
rect 2990 12914 3458 12942
rect 2378 12858 3554 12886
rect 2786 12802 3650 12830
rect 4364 12814 4648 12842
rect 2990 12746 3746 12774
rect 2446 12690 3950 12718
rect 4282 12692 4648 12720
rect 2786 12634 4046 12662
rect 2990 12578 4142 12606
rect 245 11574 561 11602
rect 2103 11603 2106 11611
rect 2077 11573 2106 11603
rect 2103 11565 2106 11573
rect 2158 11603 2161 11611
rect 2990 11618 4142 11646
rect 2158 11573 2188 11603
rect 2158 11565 2161 11573
rect 2718 11562 4046 11590
rect 2514 11506 3950 11534
rect 4282 11504 4648 11532
rect 2990 11450 3746 11478
rect 2718 11394 3650 11422
rect 4364 11382 4648 11410
rect 2446 11338 3554 11366
rect 2990 11282 3458 11310
rect 2718 11226 3362 11254
rect 4572 11236 4648 11264
rect 2378 11170 3266 11198
rect 177 9950 493 9978
rect 2103 9979 2106 9987
rect 2077 9949 2106 9979
rect 2103 9941 2106 9949
rect 2158 9979 2161 9987
rect 2446 9998 3266 10026
rect 2158 9949 2188 9979
rect 2158 9941 2161 9949
rect 2650 9942 3362 9970
rect 4572 9932 4648 9960
rect 2990 9886 3458 9914
rect 2514 9830 3554 9858
rect 2650 9774 3650 9802
rect 4364 9786 4648 9814
rect 2990 9718 3746 9746
rect 2582 9662 3950 9690
rect 4282 9664 4648 9692
rect 2650 9606 4046 9634
rect 2990 9550 4142 9578
rect 2990 8590 4142 8618
rect 2650 8534 4046 8562
rect 2378 8478 3950 8506
rect 4282 8476 4648 8504
rect 2922 8422 3746 8450
rect 2854 8366 3650 8394
rect 4364 8354 4648 8382
rect 2582 8310 3554 8338
rect 2922 8254 3458 8282
rect 2854 8198 3362 8226
rect 4572 8208 4648 8236
rect 2514 8142 3266 8170
rect 2582 6970 3266 6998
rect 2786 6914 3362 6942
rect 4572 6904 4648 6932
rect 2922 6858 3458 6886
rect 2378 6802 3554 6830
rect 2854 6746 3650 6774
rect 4364 6758 4648 6786
rect 2922 6690 3746 6718
rect 2446 6634 3950 6662
rect 4282 6636 4648 6664
rect 2854 6578 4046 6606
rect 2922 6522 4142 6550
rect 2922 5562 4142 5590
rect 2786 5506 4046 5534
rect 2103 5447 2106 5455
rect 2077 5417 2106 5447
rect 2103 5409 2106 5417
rect 2158 5447 2161 5455
rect 2158 5417 2188 5447
rect 2514 5450 3950 5478
rect 4282 5448 4648 5476
rect 2158 5409 2161 5417
rect 2922 5394 3746 5422
rect 2786 5338 3650 5366
rect 4364 5326 4648 5354
rect 2446 5282 3554 5310
rect 2922 5226 3458 5254
rect 2786 5170 3362 5198
rect 4572 5180 4648 5208
rect 2378 5114 3266 5142
rect 2446 3942 3266 3970
rect 2718 3886 3362 3914
rect 4572 3876 4648 3904
rect 2103 3823 2106 3831
rect 2077 3793 2106 3823
rect 2103 3785 2106 3793
rect 2158 3823 2161 3831
rect 2158 3793 2188 3823
rect 2922 3830 3458 3858
rect 2158 3785 2161 3793
rect 2514 3774 3554 3802
rect 2718 3718 3650 3746
rect 4364 3730 4648 3758
rect 2922 3662 3746 3690
rect 2582 3606 3950 3634
rect 4282 3608 4648 3636
rect 2718 3550 4046 3578
rect 2922 3494 4142 3522
rect 2922 2534 4142 2562
rect 2718 2478 4046 2506
rect 2378 2422 3950 2450
rect 4282 2420 4648 2448
rect 109 2338 561 2366
rect 2103 2367 2106 2375
rect 2077 2337 2106 2367
rect 2103 2329 2106 2337
rect 2158 2367 2161 2375
rect 2158 2337 2188 2367
rect 2922 2366 3746 2394
rect 2158 2329 2161 2337
rect 2650 2310 3650 2338
rect 4364 2298 4648 2326
rect 2582 2254 3554 2282
rect 2922 2198 3458 2226
rect 2650 2142 3362 2170
rect 4572 2152 4648 2180
rect 2514 2086 3266 2114
rect 2354 914 2530 942
rect 2450 858 2802 886
rect 4572 848 4648 876
rect 2546 802 3006 830
rect 41 714 493 742
rect 2103 743 2106 751
rect 2077 713 2106 743
rect 2103 705 2106 713
rect 2158 743 2161 751
rect 2158 713 2188 743
rect 2378 746 3554 774
rect 2158 705 2161 713
rect 2650 690 3650 718
rect 4364 702 4648 730
rect 2922 634 3746 662
rect 2446 578 3950 606
rect 4282 580 4648 608
rect 2650 522 4046 550
rect 2922 466 4142 494
<< via1 >>
rect 4636 24198 4688 24250
rect 2106 23921 2158 23930
rect 2106 23887 2115 23921
rect 2115 23887 2149 23921
rect 2149 23887 2158 23921
rect 2106 23878 2158 23887
rect 3006 23718 3058 23770
rect 2802 23662 2854 23714
rect 2462 23606 2514 23658
rect 3006 23550 3058 23602
rect 2802 23494 2854 23546
rect 2394 23438 2446 23490
rect 3006 23382 3058 23434
rect 2802 23326 2854 23378
rect 2326 23270 2378 23322
rect 4636 22684 4688 22736
rect 2106 22297 2158 22306
rect 2106 22263 2115 22297
rect 2115 22263 2149 22297
rect 2149 22263 2158 22297
rect 2106 22254 2158 22263
rect 2394 22098 2446 22150
rect 2734 22042 2786 22094
rect 3006 21986 3058 22038
rect 2462 21930 2514 21982
rect 2734 21874 2786 21926
rect 3006 21818 3058 21870
rect 2530 21762 2582 21814
rect 2734 21706 2786 21758
rect 3006 21650 3058 21702
rect 4636 21170 4688 21222
rect 329 20798 381 20850
rect 561 20798 613 20850
rect 2106 20841 2158 20850
rect 2106 20807 2115 20841
rect 2115 20807 2149 20841
rect 2149 20807 2158 20841
rect 2106 20798 2158 20807
rect 3006 20690 3058 20742
rect 2734 20634 2786 20686
rect 2326 20578 2378 20630
rect 3006 20522 3058 20574
rect 2666 20466 2718 20518
rect 2530 20410 2582 20462
rect 3006 20354 3058 20406
rect 2666 20298 2718 20350
rect 2462 20242 2514 20294
rect 4636 19656 4688 19708
rect 261 19174 313 19226
rect 493 19174 545 19226
rect 2106 19217 2158 19226
rect 2106 19183 2115 19217
rect 2115 19183 2149 19217
rect 2149 19183 2158 19217
rect 2106 19174 2158 19183
rect 2530 19070 2582 19122
rect 2598 19014 2650 19066
rect 3006 18958 3058 19010
rect 2326 18902 2378 18954
rect 2666 18846 2718 18898
rect 3006 18790 3058 18842
rect 2394 18734 2446 18786
rect 2666 18678 2718 18730
rect 3006 18622 3058 18674
rect 4636 18142 4688 18194
rect 3006 17662 3058 17714
rect 2598 17606 2650 17658
rect 2462 17550 2514 17602
rect 3006 17494 3058 17546
rect 2598 17438 2650 17490
rect 2394 17382 2446 17434
rect 3006 17326 3058 17378
rect 2598 17270 2650 17322
rect 2326 17214 2378 17266
rect 4636 16628 4688 16680
rect 2394 16042 2446 16094
rect 2802 15986 2854 16038
rect 2938 15930 2990 15982
rect 2462 15874 2514 15926
rect 2802 15818 2854 15870
rect 2938 15762 2990 15814
rect 2530 15706 2582 15758
rect 2802 15650 2854 15702
rect 2938 15594 2990 15646
rect 4636 15114 4688 15166
rect 2106 14685 2158 14694
rect 2106 14651 2115 14685
rect 2115 14651 2149 14685
rect 2149 14651 2158 14685
rect 2106 14642 2158 14651
rect 2938 14634 2990 14686
rect 2802 14578 2854 14630
rect 2326 14522 2378 14574
rect 2938 14466 2990 14518
rect 2734 14410 2786 14462
rect 2530 14354 2582 14406
rect 2938 14298 2990 14350
rect 2734 14242 2786 14294
rect 2462 14186 2514 14238
rect 4636 13600 4688 13652
rect 2106 13061 2158 13070
rect 2106 13027 2115 13061
rect 2115 13027 2149 13061
rect 2149 13027 2158 13061
rect 2106 13018 2158 13027
rect 2530 13014 2582 13066
rect 2666 12958 2718 13010
rect 2938 12902 2990 12954
rect 2326 12846 2378 12898
rect 2734 12790 2786 12842
rect 2938 12734 2990 12786
rect 2394 12678 2446 12730
rect 2734 12622 2786 12674
rect 2938 12566 2990 12618
rect 4636 12086 4688 12138
rect 193 11562 245 11614
rect 561 11562 613 11614
rect 2106 11605 2158 11614
rect 2106 11571 2115 11605
rect 2115 11571 2149 11605
rect 2149 11571 2158 11605
rect 2938 11606 2990 11658
rect 2106 11562 2158 11571
rect 2666 11550 2718 11602
rect 2462 11494 2514 11546
rect 2938 11438 2990 11490
rect 2666 11382 2718 11434
rect 2394 11326 2446 11378
rect 2938 11270 2990 11322
rect 2666 11214 2718 11266
rect 2326 11158 2378 11210
rect 4636 10572 4688 10624
rect 125 9938 177 9990
rect 493 9938 545 9990
rect 2106 9981 2158 9990
rect 2106 9947 2115 9981
rect 2115 9947 2149 9981
rect 2149 9947 2158 9981
rect 2394 9986 2446 10038
rect 2106 9938 2158 9947
rect 2598 9930 2650 9982
rect 2938 9874 2990 9926
rect 2462 9818 2514 9870
rect 2598 9762 2650 9814
rect 2938 9706 2990 9758
rect 2530 9650 2582 9702
rect 2598 9594 2650 9646
rect 2938 9538 2990 9590
rect 4636 9058 4688 9110
rect 2938 8578 2990 8630
rect 2598 8522 2650 8574
rect 2326 8466 2378 8518
rect 2870 8410 2922 8462
rect 2802 8354 2854 8406
rect 2530 8298 2582 8350
rect 2870 8242 2922 8294
rect 2802 8186 2854 8238
rect 2462 8130 2514 8182
rect 4636 7544 4688 7596
rect 2530 6958 2582 7010
rect 2734 6902 2786 6954
rect 2870 6846 2922 6898
rect 2326 6790 2378 6842
rect 2802 6734 2854 6786
rect 2870 6678 2922 6730
rect 2394 6622 2446 6674
rect 2802 6566 2854 6618
rect 2870 6510 2922 6562
rect 4636 6030 4688 6082
rect 2870 5550 2922 5602
rect 2734 5494 2786 5546
rect 2106 5449 2158 5458
rect 2106 5415 2115 5449
rect 2115 5415 2149 5449
rect 2149 5415 2158 5449
rect 2462 5438 2514 5490
rect 2106 5406 2158 5415
rect 2870 5382 2922 5434
rect 2734 5326 2786 5378
rect 2394 5270 2446 5322
rect 2870 5214 2922 5266
rect 2734 5158 2786 5210
rect 2326 5102 2378 5154
rect 4636 4516 4688 4568
rect 2394 3930 2446 3982
rect 2666 3874 2718 3926
rect 2106 3825 2158 3834
rect 2106 3791 2115 3825
rect 2115 3791 2149 3825
rect 2149 3791 2158 3825
rect 2870 3818 2922 3870
rect 2106 3782 2158 3791
rect 2462 3762 2514 3814
rect 2666 3706 2718 3758
rect 2870 3650 2922 3702
rect 2530 3594 2582 3646
rect 2666 3538 2718 3590
rect 2870 3482 2922 3534
rect 4636 3002 4688 3054
rect 2870 2522 2922 2574
rect 2666 2466 2718 2518
rect 2326 2410 2378 2462
rect 57 2326 109 2378
rect 561 2326 613 2378
rect 2106 2369 2158 2378
rect 2106 2335 2115 2369
rect 2115 2335 2149 2369
rect 2149 2335 2158 2369
rect 2870 2354 2922 2406
rect 2106 2326 2158 2335
rect 2598 2298 2650 2350
rect 2530 2242 2582 2294
rect 2870 2186 2922 2238
rect 2598 2130 2650 2182
rect 2462 2074 2514 2126
rect 4636 1488 4688 1540
rect 2530 902 2582 954
rect 2802 846 2854 898
rect 3006 790 3058 842
rect -11 702 41 754
rect 493 702 545 754
rect 2106 745 2158 754
rect 2106 711 2115 745
rect 2115 711 2149 745
rect 2149 711 2158 745
rect 2326 734 2378 786
rect 2106 702 2158 711
rect 2598 678 2650 730
rect 2870 622 2922 674
rect 2394 566 2446 618
rect 2598 510 2650 562
rect 2870 454 2922 506
rect 4636 -26 4688 26
<< metal2 >>
rect 1 754 29 24632
rect 69 2378 97 24632
rect 137 9990 165 24632
rect 205 11614 233 24632
rect 273 19226 301 24632
rect 341 20850 369 24632
rect 2112 23932 2152 23938
rect 2112 23870 2152 23876
rect 2338 23322 2366 24660
rect 2406 23490 2434 24660
rect 2474 23658 2502 24660
rect 2112 22308 2152 22314
rect 2112 22246 2152 22252
rect 2112 20852 2152 20858
rect 1 0 29 702
rect 69 0 97 2326
rect 137 0 165 9938
rect 205 0 233 11562
rect 273 0 301 19174
rect 341 0 369 20798
rect 2112 20790 2152 20796
rect 2338 20630 2366 23270
rect 2406 22150 2434 23438
rect 2112 19228 2152 19234
rect 2112 19166 2152 19172
rect 2338 18954 2366 20578
rect 2338 17266 2366 18902
rect 2406 18786 2434 22098
rect 2474 21982 2502 23606
rect 2474 20294 2502 21930
rect 2542 21814 2570 24660
rect 2542 20462 2570 21762
rect 2406 17434 2434 18734
rect 2474 17602 2502 20242
rect 2542 19122 2570 20410
rect 2112 14696 2152 14702
rect 2112 14634 2152 14640
rect 2338 14574 2366 17214
rect 2406 16094 2434 17382
rect 2112 13072 2152 13078
rect 2112 13010 2152 13016
rect 2338 12898 2366 14522
rect 2112 11616 2152 11622
rect 2112 11554 2152 11560
rect 2338 11210 2366 12846
rect 2406 12730 2434 16042
rect 2474 15926 2502 17550
rect 2474 14238 2502 15874
rect 2542 15758 2570 19070
rect 2610 19066 2638 24660
rect 2678 20518 2706 24660
rect 2746 22094 2774 24660
rect 2814 23714 2842 24660
rect 2814 23546 2842 23662
rect 2814 23378 2842 23494
rect 2746 21926 2774 22042
rect 2746 21758 2774 21874
rect 2746 20686 2774 21706
rect 2678 20350 2706 20466
rect 2610 17658 2638 19014
rect 2678 18898 2706 20298
rect 2678 18730 2706 18846
rect 2610 17490 2638 17606
rect 2610 17322 2638 17438
rect 2542 14406 2570 15706
rect 2406 11378 2434 12678
rect 2474 11546 2502 14186
rect 2542 13066 2570 14354
rect 2112 9992 2152 9998
rect 2112 9930 2152 9936
rect 2338 8518 2366 11158
rect 2406 10038 2434 11326
rect 2338 6842 2366 8466
rect 2112 5460 2152 5466
rect 2112 5398 2152 5404
rect 2338 5154 2366 6790
rect 2406 6674 2434 9986
rect 2474 9870 2502 11494
rect 2474 8182 2502 9818
rect 2542 9702 2570 13014
rect 2610 9982 2638 17270
rect 2678 13010 2706 18678
rect 2746 14462 2774 20634
rect 2814 16038 2842 23326
rect 2882 18500 2910 24660
rect 2950 20040 2978 24660
rect 3018 23770 3046 24660
rect 3018 23602 3046 23718
rect 3018 23434 3046 23550
rect 3018 22038 3046 23382
rect 3086 23120 3114 24660
rect 4642 24252 4682 24258
rect 4642 24190 4682 24196
rect 3018 21870 3046 21986
rect 3018 21702 3046 21818
rect 3018 21580 3046 21650
rect 3018 20742 3046 21524
rect 3018 20574 3046 20690
rect 3018 20406 3046 20522
rect 2814 15870 2842 15986
rect 2814 15702 2842 15818
rect 2814 14630 2842 15650
rect 2746 14294 2774 14410
rect 2678 11602 2706 12958
rect 2746 12842 2774 14242
rect 2814 13884 2842 14578
rect 2746 12674 2774 12790
rect 2746 12344 2774 12622
rect 2678 11434 2706 11550
rect 2678 11266 2706 11382
rect 2678 10804 2706 11214
rect 2610 9814 2638 9930
rect 2542 8350 2570 9650
rect 2610 9646 2638 9762
rect 2610 9264 2638 9594
rect 2610 8574 2638 9208
rect 2406 5322 2434 6622
rect 2474 5490 2502 8130
rect 2542 7010 2570 8298
rect 2112 3836 2152 3842
rect 2112 3774 2152 3780
rect 2338 2462 2366 5102
rect 2406 3982 2434 5270
rect 2112 2380 2152 2386
rect 2112 2318 2152 2324
rect 2338 786 2366 2410
rect 2406 1568 2434 3930
rect 2474 3814 2502 5438
rect 2542 4648 2570 6958
rect 2474 3108 2502 3762
rect 2542 3646 2570 4592
rect 2474 2126 2502 3052
rect 2542 2294 2570 3594
rect 2610 2350 2638 8522
rect 2678 3926 2706 10748
rect 2746 6954 2774 12288
rect 2814 8406 2842 13828
rect 2882 8462 2910 18444
rect 2950 15982 2978 19984
rect 3018 19010 3046 20354
rect 3018 18842 3046 18958
rect 3018 18674 3046 18790
rect 3018 17714 3046 18622
rect 3018 17546 3046 17662
rect 3018 17378 3046 17494
rect 2950 15814 2978 15930
rect 2950 15646 2978 15762
rect 2950 14686 2978 15594
rect 2950 14518 2978 14634
rect 2950 14350 2978 14466
rect 2950 12954 2978 14298
rect 2950 12786 2978 12902
rect 2950 12618 2978 12734
rect 2950 11658 2978 12566
rect 2950 11490 2978 11606
rect 2950 11322 2978 11438
rect 2950 9926 2978 11270
rect 2950 9758 2978 9874
rect 2950 9590 2978 9706
rect 2950 8630 2978 9538
rect 2814 8238 2842 8354
rect 2882 8294 2910 8410
rect 2746 5546 2774 6902
rect 2814 6786 2842 8186
rect 2882 6898 2910 8242
rect 2814 6618 2842 6734
rect 2882 6730 2910 6846
rect 2746 5378 2774 5494
rect 2746 5210 2774 5326
rect 2678 3758 2706 3874
rect 2678 3590 2706 3706
rect 2678 2518 2706 3538
rect 2112 756 2152 762
rect 2112 694 2152 700
rect 2338 28 2366 734
rect 2406 618 2434 1512
rect 2406 0 2434 566
rect 2474 0 2502 2074
rect 2542 954 2570 2242
rect 2610 2182 2638 2298
rect 2542 0 2570 902
rect 2610 730 2638 2130
rect 2610 562 2638 678
rect 2610 0 2638 510
rect 2678 0 2706 2466
rect 2746 0 2774 5158
rect 2814 898 2842 6566
rect 2882 6562 2910 6678
rect 2882 5602 2910 6510
rect 2882 5434 2910 5550
rect 2882 5266 2910 5382
rect 2882 3870 2910 5214
rect 2882 3702 2910 3818
rect 2882 3534 2910 3650
rect 2882 2574 2910 3482
rect 2882 2406 2910 2522
rect 2882 2238 2910 2354
rect 2814 0 2842 846
rect 2882 674 2910 2186
rect 2882 506 2910 622
rect 2882 0 2910 454
rect 2950 0 2978 8578
rect 3018 842 3046 17326
rect 3018 0 3046 790
rect 3086 0 3114 23064
rect 4642 22738 4682 22744
rect 4642 22676 4682 22682
rect 4642 21224 4682 21230
rect 4642 21162 4682 21168
rect 4642 19710 4682 19716
rect 4642 19648 4682 19654
rect 4642 18196 4682 18202
rect 4642 18134 4682 18140
rect 4642 16682 4682 16688
rect 4642 16620 4682 16626
rect 4642 15168 4682 15174
rect 4642 15106 4682 15112
rect 4642 13654 4682 13660
rect 4642 13592 4682 13598
rect 4642 12140 4682 12146
rect 4642 12078 4682 12084
rect 4642 10626 4682 10632
rect 4642 10564 4682 10570
rect 4642 9112 4682 9118
rect 4642 9050 4682 9056
rect 4642 7598 4682 7604
rect 4642 7536 4682 7542
rect 4642 6084 4682 6090
rect 4642 6022 4682 6028
rect 4642 4570 4682 4576
rect 4642 4508 4682 4514
rect 4642 3056 4682 3062
rect 4642 2994 4682 3000
rect 4642 1542 4682 1548
rect 4642 1480 4682 1486
rect 4642 28 4682 34
rect 4642 -34 4682 -28
<< via2 >>
rect 2104 23930 2160 23932
rect 2104 23878 2106 23930
rect 2106 23878 2158 23930
rect 2158 23878 2160 23930
rect 2104 23876 2160 23878
rect 2104 22306 2160 22308
rect 2104 22254 2106 22306
rect 2106 22254 2158 22306
rect 2158 22254 2160 22306
rect 2104 22252 2160 22254
rect 2104 20850 2160 20852
rect 2104 20798 2106 20850
rect 2106 20798 2158 20850
rect 2158 20798 2160 20850
rect 2104 20796 2160 20798
rect 2104 19226 2160 19228
rect 2104 19174 2106 19226
rect 2106 19174 2158 19226
rect 2158 19174 2160 19226
rect 2104 19172 2160 19174
rect 2104 14694 2160 14696
rect 2104 14642 2106 14694
rect 2106 14642 2158 14694
rect 2158 14642 2160 14694
rect 2104 14640 2160 14642
rect 2104 13070 2160 13072
rect 2104 13018 2106 13070
rect 2106 13018 2158 13070
rect 2158 13018 2160 13070
rect 2104 13016 2160 13018
rect 2104 11614 2160 11616
rect 2104 11562 2106 11614
rect 2106 11562 2158 11614
rect 2158 11562 2160 11614
rect 2104 11560 2160 11562
rect 2104 9990 2160 9992
rect 2104 9938 2106 9990
rect 2106 9938 2158 9990
rect 2158 9938 2160 9990
rect 2104 9936 2160 9938
rect 2104 5458 2160 5460
rect 2104 5406 2106 5458
rect 2106 5406 2158 5458
rect 2158 5406 2160 5458
rect 2104 5404 2160 5406
rect 4634 24250 4690 24252
rect 4634 24198 4636 24250
rect 4636 24198 4688 24250
rect 4688 24198 4690 24250
rect 4634 24196 4690 24198
rect 3072 23064 3128 23120
rect 3004 21524 3060 21580
rect 2936 19984 2992 20040
rect 2868 18444 2924 18500
rect 2800 13828 2856 13884
rect 2732 12288 2788 12344
rect 2664 10748 2720 10804
rect 2596 9208 2652 9264
rect 2104 3834 2160 3836
rect 2104 3782 2106 3834
rect 2106 3782 2158 3834
rect 2158 3782 2160 3834
rect 2104 3780 2160 3782
rect 2104 2378 2160 2380
rect 2104 2326 2106 2378
rect 2106 2326 2158 2378
rect 2158 2326 2160 2378
rect 2104 2324 2160 2326
rect 2528 4592 2584 4648
rect 2460 3052 2516 3108
rect 2392 1512 2448 1568
rect 2104 754 2160 756
rect 2104 702 2106 754
rect 2106 702 2158 754
rect 2158 702 2160 754
rect 2104 700 2160 702
rect 2324 -28 2380 28
rect 4634 22736 4690 22738
rect 4634 22684 4636 22736
rect 4636 22684 4688 22736
rect 4688 22684 4690 22736
rect 4634 22682 4690 22684
rect 4634 21222 4690 21224
rect 4634 21170 4636 21222
rect 4636 21170 4688 21222
rect 4688 21170 4690 21222
rect 4634 21168 4690 21170
rect 4634 19708 4690 19710
rect 4634 19656 4636 19708
rect 4636 19656 4688 19708
rect 4688 19656 4690 19708
rect 4634 19654 4690 19656
rect 4634 18194 4690 18196
rect 4634 18142 4636 18194
rect 4636 18142 4688 18194
rect 4688 18142 4690 18194
rect 4634 18140 4690 18142
rect 4634 16680 4690 16682
rect 4634 16628 4636 16680
rect 4636 16628 4688 16680
rect 4688 16628 4690 16680
rect 4634 16626 4690 16628
rect 4634 15166 4690 15168
rect 4634 15114 4636 15166
rect 4636 15114 4688 15166
rect 4688 15114 4690 15166
rect 4634 15112 4690 15114
rect 4634 13652 4690 13654
rect 4634 13600 4636 13652
rect 4636 13600 4688 13652
rect 4688 13600 4690 13652
rect 4634 13598 4690 13600
rect 4634 12138 4690 12140
rect 4634 12086 4636 12138
rect 4636 12086 4688 12138
rect 4688 12086 4690 12138
rect 4634 12084 4690 12086
rect 4634 10624 4690 10626
rect 4634 10572 4636 10624
rect 4636 10572 4688 10624
rect 4688 10572 4690 10624
rect 4634 10570 4690 10572
rect 4634 9110 4690 9112
rect 4634 9058 4636 9110
rect 4636 9058 4688 9110
rect 4688 9058 4690 9110
rect 4634 9056 4690 9058
rect 4634 7596 4690 7598
rect 4634 7544 4636 7596
rect 4636 7544 4688 7596
rect 4688 7544 4690 7596
rect 4634 7542 4690 7544
rect 4634 6082 4690 6084
rect 4634 6030 4636 6082
rect 4636 6030 4688 6082
rect 4688 6030 4690 6082
rect 4634 6028 4690 6030
rect 4634 4568 4690 4570
rect 4634 4516 4636 4568
rect 4636 4516 4688 4568
rect 4688 4516 4690 4568
rect 4634 4514 4690 4516
rect 4634 3054 4690 3056
rect 4634 3002 4636 3054
rect 4636 3002 4688 3054
rect 4688 3002 4690 3054
rect 4634 3000 4690 3002
rect 4634 1540 4690 1542
rect 4634 1488 4636 1540
rect 4636 1488 4688 1540
rect 4688 1488 4690 1540
rect 4634 1486 4690 1488
rect 4634 26 4690 28
rect 4634 -26 4636 26
rect 4636 -26 4688 26
rect 4688 -26 4690 26
rect 4634 -28 4690 -26
<< metal3 >>
rect 651 24602 711 24662
rect 1410 24602 1470 24662
rect 4632 24252 4692 24254
rect 4632 24196 4634 24252
rect 4690 24196 4692 24252
rect 4632 24194 4692 24196
rect 2102 23932 2162 23934
rect 2102 23876 2104 23932
rect 2160 23876 2162 23932
rect 2102 23122 2162 23876
rect 651 23062 711 23122
rect 1410 23062 1470 23122
rect 2102 23120 3130 23122
rect 2102 23064 3072 23120
rect 3128 23064 3130 23120
rect 2102 23062 3130 23064
rect 4632 22738 4692 22740
rect 4632 22682 4634 22738
rect 4690 22682 4692 22738
rect 4632 22680 4692 22682
rect 2102 22308 2162 22310
rect 2102 22252 2104 22308
rect 2160 22252 2162 22308
rect 2102 21582 2162 22252
rect 651 21522 711 21582
rect 1410 21522 1470 21582
rect 2102 21580 3062 21582
rect 2102 21524 3004 21580
rect 3060 21524 3062 21580
rect 2102 21522 3062 21524
rect 4632 21224 4692 21226
rect 4632 21168 4634 21224
rect 4690 21168 4692 21224
rect 4632 21166 4692 21168
rect 2102 20852 2162 20854
rect 2102 20796 2104 20852
rect 2160 20796 2162 20852
rect 2102 20042 2162 20796
rect 651 19982 711 20042
rect 1410 19982 1470 20042
rect 2102 20040 2994 20042
rect 2102 19984 2936 20040
rect 2992 19984 2994 20040
rect 2102 19982 2994 19984
rect 4632 19710 4692 19712
rect 4632 19654 4634 19710
rect 4690 19654 4692 19710
rect 4632 19652 4692 19654
rect 2102 19228 2162 19230
rect 2102 19172 2104 19228
rect 2160 19172 2162 19228
rect 2102 18502 2162 19172
rect 651 18442 711 18502
rect 1410 18442 1470 18502
rect 2102 18500 2926 18502
rect 2102 18444 2868 18500
rect 2924 18444 2926 18500
rect 2102 18442 2926 18444
rect 4632 18196 4692 18198
rect 4632 18140 4634 18196
rect 4690 18140 4692 18196
rect 4632 18138 4692 18140
rect 4632 16682 4692 16684
rect 4632 16626 4634 16682
rect 4690 16626 4692 16682
rect 4632 16624 4692 16626
rect 651 15366 711 15426
rect 1410 15366 1470 15426
rect 4632 15168 4692 15170
rect 4632 15112 4634 15168
rect 4690 15112 4692 15168
rect 4632 15110 4692 15112
rect 2102 14696 2162 14698
rect 2102 14640 2104 14696
rect 2160 14640 2162 14696
rect 2102 13886 2162 14640
rect 651 13826 711 13886
rect 1410 13826 1470 13886
rect 2102 13884 2858 13886
rect 2102 13828 2800 13884
rect 2856 13828 2858 13884
rect 2102 13826 2858 13828
rect 4632 13654 4692 13656
rect 4632 13598 4634 13654
rect 4690 13598 4692 13654
rect 4632 13596 4692 13598
rect 2102 13072 2162 13074
rect 2102 13016 2104 13072
rect 2160 13016 2162 13072
rect 2102 12346 2162 13016
rect 651 12286 711 12346
rect 1410 12286 1470 12346
rect 2102 12344 2790 12346
rect 2102 12288 2732 12344
rect 2788 12288 2790 12344
rect 2102 12286 2790 12288
rect 4632 12140 4692 12142
rect 4632 12084 4634 12140
rect 4690 12084 4692 12140
rect 4632 12082 4692 12084
rect 2102 11616 2162 11618
rect 2102 11560 2104 11616
rect 2160 11560 2162 11616
rect 2102 10806 2162 11560
rect 651 10746 711 10806
rect 1410 10746 1470 10806
rect 2102 10804 2722 10806
rect 2102 10748 2664 10804
rect 2720 10748 2722 10804
rect 2102 10746 2722 10748
rect 4632 10626 4692 10628
rect 4632 10570 4634 10626
rect 4690 10570 4692 10626
rect 4632 10568 4692 10570
rect 2102 9992 2162 9994
rect 2102 9936 2104 9992
rect 2160 9936 2162 9992
rect 2102 9266 2162 9936
rect 651 9206 711 9266
rect 1410 9206 1470 9266
rect 2102 9264 2654 9266
rect 2102 9208 2596 9264
rect 2652 9208 2654 9264
rect 2102 9206 2654 9208
rect 4632 9112 4692 9114
rect 4632 9056 4634 9112
rect 4690 9056 4692 9112
rect 4632 9054 4692 9056
rect 4632 7598 4692 7600
rect 4632 7542 4634 7598
rect 4690 7542 4692 7598
rect 4632 7540 4692 7542
rect 651 6130 711 6190
rect 1410 6130 1470 6190
rect 4632 6084 4692 6086
rect 4632 6028 4634 6084
rect 4690 6028 4692 6084
rect 4632 6026 4692 6028
rect 2102 5460 2162 5462
rect 2102 5404 2104 5460
rect 2160 5404 2162 5460
rect 2102 4650 2162 5404
rect 651 4590 711 4650
rect 1410 4590 1470 4650
rect 2102 4648 2586 4650
rect 2102 4592 2528 4648
rect 2584 4592 2586 4648
rect 2102 4590 2586 4592
rect 4632 4570 4692 4572
rect 4632 4514 4634 4570
rect 4690 4514 4692 4570
rect 4632 4512 4692 4514
rect 2102 3836 2162 3838
rect 2102 3780 2104 3836
rect 2160 3780 2162 3836
rect 2102 3110 2162 3780
rect 651 3050 711 3110
rect 1410 3050 1470 3110
rect 2102 3108 2518 3110
rect 2102 3052 2460 3108
rect 2516 3052 2518 3108
rect 2102 3050 2518 3052
rect 4632 3056 4692 3058
rect 4632 3000 4634 3056
rect 4690 3000 4692 3056
rect 4632 2998 4692 3000
rect 2102 2380 2162 2382
rect 2102 2324 2104 2380
rect 2160 2324 2162 2380
rect 2102 1570 2162 2324
rect 651 1510 711 1570
rect 1410 1510 1470 1570
rect 2102 1568 2450 1570
rect 2102 1512 2392 1568
rect 2448 1512 2450 1568
rect 2102 1510 2450 1512
rect 4632 1542 4692 1544
rect 4632 1486 4634 1542
rect 4690 1486 4692 1542
rect 4632 1484 4692 1486
rect 2102 756 2162 758
rect 2102 700 2104 756
rect 2160 700 2162 756
rect 2102 30 2162 700
rect 651 -30 711 30
rect 1410 -30 1470 30
rect 2102 28 2382 30
rect 2102 -28 2324 28
rect 2380 -28 2382 28
rect 2102 -30 2382 -28
rect 4632 28 4692 30
rect 4632 -28 4634 28
rect 4690 -28 4692 28
rect 4632 -30 4692 -28
use contact_18  contact_18_0
timestamp 1643671299
transform 1 0 4632 0 1 -30
box 0 0 1 1
use contact_17  contact_17_0
timestamp 1643671299
transform 1 0 4647 0 1 -15
box 0 0 1 1
use contact_18  contact_18_1
timestamp 1643671299
transform 1 0 4632 0 1 1484
box 0 0 1 1
use contact_17  contact_17_1
timestamp 1643671299
transform 1 0 4647 0 1 1499
box 0 0 1 1
use contact_18  contact_18_2
timestamp 1643671299
transform 1 0 4632 0 1 -30
box 0 0 1 1
use contact_17  contact_17_2
timestamp 1643671299
transform 1 0 4647 0 1 -15
box 0 0 1 1
use contact_18  contact_18_3
timestamp 1643671299
transform 1 0 4632 0 1 1484
box 0 0 1 1
use contact_17  contact_17_3
timestamp 1643671299
transform 1 0 4647 0 1 1499
box 0 0 1 1
use contact_18  contact_18_4
timestamp 1643671299
transform 1 0 4632 0 1 -30
box 0 0 1 1
use contact_17  contact_17_4
timestamp 1643671299
transform 1 0 4647 0 1 -15
box 0 0 1 1
use contact_18  contact_18_5
timestamp 1643671299
transform 1 0 4632 0 1 1484
box 0 0 1 1
use contact_17  contact_17_5
timestamp 1643671299
transform 1 0 4647 0 1 1499
box 0 0 1 1
use contact_18  contact_18_6
timestamp 1643671299
transform 1 0 4632 0 1 -30
box 0 0 1 1
use contact_17  contact_17_6
timestamp 1643671299
transform 1 0 4647 0 1 -15
box 0 0 1 1
use contact_18  contact_18_7
timestamp 1643671299
transform 1 0 4632 0 1 1484
box 0 0 1 1
use contact_17  contact_17_7
timestamp 1643671299
transform 1 0 4647 0 1 1499
box 0 0 1 1
use contact_18  contact_18_8
timestamp 1643671299
transform 1 0 4632 0 1 -30
box 0 0 1 1
use contact_17  contact_17_8
timestamp 1643671299
transform 1 0 4647 0 1 -15
box 0 0 1 1
use contact_18  contact_18_9
timestamp 1643671299
transform 1 0 4632 0 1 1484
box 0 0 1 1
use contact_17  contact_17_9
timestamp 1643671299
transform 1 0 4647 0 1 1499
box 0 0 1 1
use contact_18  contact_18_10
timestamp 1643671299
transform 1 0 4632 0 1 -30
box 0 0 1 1
use contact_17  contact_17_10
timestamp 1643671299
transform 1 0 4647 0 1 -15
box 0 0 1 1
use contact_18  contact_18_11
timestamp 1643671299
transform 1 0 4632 0 1 1484
box 0 0 1 1
use contact_17  contact_17_11
timestamp 1643671299
transform 1 0 4647 0 1 1499
box 0 0 1 1
use contact_18  contact_18_12
timestamp 1643671299
transform 1 0 4632 0 1 -30
box 0 0 1 1
use contact_17  contact_17_12
timestamp 1643671299
transform 1 0 4647 0 1 -15
box 0 0 1 1
use contact_18  contact_18_13
timestamp 1643671299
transform 1 0 4632 0 1 1484
box 0 0 1 1
use contact_17  contact_17_13
timestamp 1643671299
transform 1 0 4647 0 1 1499
box 0 0 1 1
use contact_18  contact_18_14
timestamp 1643671299
transform 1 0 4632 0 1 -30
box 0 0 1 1
use contact_17  contact_17_14
timestamp 1643671299
transform 1 0 4647 0 1 -15
box 0 0 1 1
use contact_18  contact_18_15
timestamp 1643671299
transform 1 0 4632 0 1 1484
box 0 0 1 1
use contact_17  contact_17_15
timestamp 1643671299
transform 1 0 4647 0 1 1499
box 0 0 1 1
use contact_18  contact_18_16
timestamp 1643671299
transform 1 0 4632 0 1 -30
box 0 0 1 1
use contact_17  contact_17_16
timestamp 1643671299
transform 1 0 4647 0 1 -15
box 0 0 1 1
use contact_18  contact_18_17
timestamp 1643671299
transform 1 0 4632 0 1 1484
box 0 0 1 1
use contact_17  contact_17_17
timestamp 1643671299
transform 1 0 4647 0 1 1499
box 0 0 1 1
use contact_18  contact_18_18
timestamp 1643671299
transform 1 0 4632 0 1 -30
box 0 0 1 1
use contact_17  contact_17_18
timestamp 1643671299
transform 1 0 4647 0 1 -15
box 0 0 1 1
use contact_18  contact_18_19
timestamp 1643671299
transform 1 0 4632 0 1 1484
box 0 0 1 1
use contact_17  contact_17_19
timestamp 1643671299
transform 1 0 4647 0 1 1499
box 0 0 1 1
use contact_18  contact_18_20
timestamp 1643671299
transform 1 0 4632 0 1 -30
box 0 0 1 1
use contact_17  contact_17_20
timestamp 1643671299
transform 1 0 4647 0 1 -15
box 0 0 1 1
use contact_18  contact_18_21
timestamp 1643671299
transform 1 0 4632 0 1 1484
box 0 0 1 1
use contact_17  contact_17_21
timestamp 1643671299
transform 1 0 4647 0 1 1499
box 0 0 1 1
use contact_18  contact_18_22
timestamp 1643671299
transform 1 0 4632 0 1 -30
box 0 0 1 1
use contact_17  contact_17_22
timestamp 1643671299
transform 1 0 4647 0 1 -15
box 0 0 1 1
use contact_18  contact_18_23
timestamp 1643671299
transform 1 0 4632 0 1 1484
box 0 0 1 1
use contact_17  contact_17_23
timestamp 1643671299
transform 1 0 4647 0 1 1499
box 0 0 1 1
use contact_18  contact_18_24
timestamp 1643671299
transform 1 0 4632 0 1 -30
box 0 0 1 1
use contact_17  contact_17_24
timestamp 1643671299
transform 1 0 4647 0 1 -15
box 0 0 1 1
use contact_18  contact_18_25
timestamp 1643671299
transform 1 0 4632 0 1 1484
box 0 0 1 1
use contact_17  contact_17_25
timestamp 1643671299
transform 1 0 4647 0 1 1499
box 0 0 1 1
use contact_18  contact_18_26
timestamp 1643671299
transform 1 0 4632 0 1 -30
box 0 0 1 1
use contact_17  contact_17_26
timestamp 1643671299
transform 1 0 4647 0 1 -15
box 0 0 1 1
use contact_18  contact_18_27
timestamp 1643671299
transform 1 0 4632 0 1 1484
box 0 0 1 1
use contact_17  contact_17_27
timestamp 1643671299
transform 1 0 4647 0 1 1499
box 0 0 1 1
use contact_18  contact_18_28
timestamp 1643671299
transform 1 0 4632 0 1 -30
box 0 0 1 1
use contact_17  contact_17_28
timestamp 1643671299
transform 1 0 4647 0 1 -15
box 0 0 1 1
use contact_18  contact_18_29
timestamp 1643671299
transform 1 0 4632 0 1 1484
box 0 0 1 1
use contact_17  contact_17_29
timestamp 1643671299
transform 1 0 4647 0 1 1499
box 0 0 1 1
use contact_18  contact_18_30
timestamp 1643671299
transform 1 0 4632 0 1 -30
box 0 0 1 1
use contact_17  contact_17_30
timestamp 1643671299
transform 1 0 4647 0 1 -15
box 0 0 1 1
use contact_18  contact_18_31
timestamp 1643671299
transform 1 0 4632 0 1 1484
box 0 0 1 1
use contact_17  contact_17_31
timestamp 1643671299
transform 1 0 4647 0 1 1499
box 0 0 1 1
use contact_18  contact_18_32
timestamp 1643671299
transform 1 0 4632 0 1 -30
box 0 0 1 1
use contact_17  contact_17_32
timestamp 1643671299
transform 1 0 4647 0 1 -15
box 0 0 1 1
use contact_18  contact_18_33
timestamp 1643671299
transform 1 0 4632 0 1 1484
box 0 0 1 1
use contact_17  contact_17_33
timestamp 1643671299
transform 1 0 4647 0 1 1499
box 0 0 1 1
use contact_18  contact_18_34
timestamp 1643671299
transform 1 0 4632 0 1 -30
box 0 0 1 1
use contact_17  contact_17_34
timestamp 1643671299
transform 1 0 4647 0 1 -15
box 0 0 1 1
use contact_18  contact_18_35
timestamp 1643671299
transform 1 0 4632 0 1 1484
box 0 0 1 1
use contact_17  contact_17_35
timestamp 1643671299
transform 1 0 4647 0 1 1499
box 0 0 1 1
use contact_18  contact_18_36
timestamp 1643671299
transform 1 0 4632 0 1 -30
box 0 0 1 1
use contact_17  contact_17_36
timestamp 1643671299
transform 1 0 4647 0 1 -15
box 0 0 1 1
use contact_18  contact_18_37
timestamp 1643671299
transform 1 0 4632 0 1 1484
box 0 0 1 1
use contact_17  contact_17_37
timestamp 1643671299
transform 1 0 4647 0 1 1499
box 0 0 1 1
use contact_18  contact_18_38
timestamp 1643671299
transform 1 0 4632 0 1 -30
box 0 0 1 1
use contact_17  contact_17_38
timestamp 1643671299
transform 1 0 4647 0 1 -15
box 0 0 1 1
use contact_18  contact_18_39
timestamp 1643671299
transform 1 0 4632 0 1 1484
box 0 0 1 1
use contact_17  contact_17_39
timestamp 1643671299
transform 1 0 4647 0 1 1499
box 0 0 1 1
use contact_18  contact_18_40
timestamp 1643671299
transform 1 0 4632 0 1 -30
box 0 0 1 1
use contact_17  contact_17_40
timestamp 1643671299
transform 1 0 4647 0 1 -15
box 0 0 1 1
use contact_18  contact_18_41
timestamp 1643671299
transform 1 0 4632 0 1 1484
box 0 0 1 1
use contact_17  contact_17_41
timestamp 1643671299
transform 1 0 4647 0 1 1499
box 0 0 1 1
use contact_18  contact_18_42
timestamp 1643671299
transform 1 0 4632 0 1 -30
box 0 0 1 1
use contact_17  contact_17_42
timestamp 1643671299
transform 1 0 4647 0 1 -15
box 0 0 1 1
use contact_18  contact_18_43
timestamp 1643671299
transform 1 0 4632 0 1 1484
box 0 0 1 1
use contact_17  contact_17_43
timestamp 1643671299
transform 1 0 4647 0 1 1499
box 0 0 1 1
use contact_18  contact_18_44
timestamp 1643671299
transform 1 0 4632 0 1 -30
box 0 0 1 1
use contact_17  contact_17_44
timestamp 1643671299
transform 1 0 4647 0 1 -15
box 0 0 1 1
use contact_18  contact_18_45
timestamp 1643671299
transform 1 0 4632 0 1 1484
box 0 0 1 1
use contact_17  contact_17_45
timestamp 1643671299
transform 1 0 4647 0 1 1499
box 0 0 1 1
use contact_18  contact_18_46
timestamp 1643671299
transform 1 0 4632 0 1 -30
box 0 0 1 1
use contact_17  contact_17_46
timestamp 1643671299
transform 1 0 4647 0 1 -15
box 0 0 1 1
use contact_18  contact_18_47
timestamp 1643671299
transform 1 0 4632 0 1 1484
box 0 0 1 1
use contact_17  contact_17_47
timestamp 1643671299
transform 1 0 4647 0 1 1499
box 0 0 1 1
use contact_18  contact_18_48
timestamp 1643671299
transform 1 0 4632 0 1 -30
box 0 0 1 1
use contact_17  contact_17_48
timestamp 1643671299
transform 1 0 4647 0 1 -15
box 0 0 1 1
use contact_18  contact_18_49
timestamp 1643671299
transform 1 0 4632 0 1 1484
box 0 0 1 1
use contact_17  contact_17_49
timestamp 1643671299
transform 1 0 4647 0 1 1499
box 0 0 1 1
use contact_18  contact_18_50
timestamp 1643671299
transform 1 0 4632 0 1 -30
box 0 0 1 1
use contact_17  contact_17_50
timestamp 1643671299
transform 1 0 4647 0 1 -15
box 0 0 1 1
use contact_18  contact_18_51
timestamp 1643671299
transform 1 0 4632 0 1 1484
box 0 0 1 1
use contact_17  contact_17_51
timestamp 1643671299
transform 1 0 4647 0 1 1499
box 0 0 1 1
use contact_18  contact_18_52
timestamp 1643671299
transform 1 0 4632 0 1 -30
box 0 0 1 1
use contact_17  contact_17_52
timestamp 1643671299
transform 1 0 4647 0 1 -15
box 0 0 1 1
use contact_18  contact_18_53
timestamp 1643671299
transform 1 0 4632 0 1 1484
box 0 0 1 1
use contact_17  contact_17_53
timestamp 1643671299
transform 1 0 4647 0 1 1499
box 0 0 1 1
use contact_18  contact_18_54
timestamp 1643671299
transform 1 0 4632 0 1 -30
box 0 0 1 1
use contact_17  contact_17_54
timestamp 1643671299
transform 1 0 4647 0 1 -15
box 0 0 1 1
use contact_18  contact_18_55
timestamp 1643671299
transform 1 0 4632 0 1 1484
box 0 0 1 1
use contact_17  contact_17_55
timestamp 1643671299
transform 1 0 4647 0 1 1499
box 0 0 1 1
use contact_18  contact_18_56
timestamp 1643671299
transform 1 0 4632 0 1 -30
box 0 0 1 1
use contact_17  contact_17_56
timestamp 1643671299
transform 1 0 4647 0 1 -15
box 0 0 1 1
use contact_18  contact_18_57
timestamp 1643671299
transform 1 0 4632 0 1 1484
box 0 0 1 1
use contact_17  contact_17_57
timestamp 1643671299
transform 1 0 4647 0 1 1499
box 0 0 1 1
use contact_18  contact_18_58
timestamp 1643671299
transform 1 0 4632 0 1 -30
box 0 0 1 1
use contact_17  contact_17_58
timestamp 1643671299
transform 1 0 4647 0 1 -15
box 0 0 1 1
use contact_18  contact_18_59
timestamp 1643671299
transform 1 0 4632 0 1 1484
box 0 0 1 1
use contact_17  contact_17_59
timestamp 1643671299
transform 1 0 4647 0 1 1499
box 0 0 1 1
use contact_18  contact_18_60
timestamp 1643671299
transform 1 0 4632 0 1 -30
box 0 0 1 1
use contact_17  contact_17_60
timestamp 1643671299
transform 1 0 4647 0 1 -15
box 0 0 1 1
use contact_18  contact_18_61
timestamp 1643671299
transform 1 0 4632 0 1 1484
box 0 0 1 1
use contact_17  contact_17_61
timestamp 1643671299
transform 1 0 4647 0 1 1499
box 0 0 1 1
use contact_18  contact_18_62
timestamp 1643671299
transform 1 0 4632 0 1 -30
box 0 0 1 1
use contact_17  contact_17_62
timestamp 1643671299
transform 1 0 4647 0 1 -15
box 0 0 1 1
use contact_18  contact_18_63
timestamp 1643671299
transform 1 0 4632 0 1 1484
box 0 0 1 1
use contact_17  contact_17_63
timestamp 1643671299
transform 1 0 4647 0 1 1499
box 0 0 1 1
use contact_18  contact_18_64
timestamp 1643671299
transform 1 0 4632 0 1 24194
box 0 0 1 1
use contact_17  contact_17_64
timestamp 1643671299
transform 1 0 4647 0 1 24209
box 0 0 1 1
use contact_18  contact_18_65
timestamp 1643671299
transform 1 0 4632 0 1 22680
box 0 0 1 1
use contact_17  contact_17_65
timestamp 1643671299
transform 1 0 4647 0 1 22695
box 0 0 1 1
use contact_18  contact_18_66
timestamp 1643671299
transform 1 0 4632 0 1 21166
box 0 0 1 1
use contact_17  contact_17_66
timestamp 1643671299
transform 1 0 4647 0 1 21181
box 0 0 1 1
use contact_18  contact_18_67
timestamp 1643671299
transform 1 0 4632 0 1 22680
box 0 0 1 1
use contact_17  contact_17_67
timestamp 1643671299
transform 1 0 4647 0 1 22695
box 0 0 1 1
use contact_18  contact_18_68
timestamp 1643671299
transform 1 0 4632 0 1 21166
box 0 0 1 1
use contact_17  contact_17_68
timestamp 1643671299
transform 1 0 4647 0 1 21181
box 0 0 1 1
use contact_18  contact_18_69
timestamp 1643671299
transform 1 0 4632 0 1 19652
box 0 0 1 1
use contact_17  contact_17_69
timestamp 1643671299
transform 1 0 4647 0 1 19667
box 0 0 1 1
use contact_18  contact_18_70
timestamp 1643671299
transform 1 0 4632 0 1 18138
box 0 0 1 1
use contact_17  contact_17_70
timestamp 1643671299
transform 1 0 4647 0 1 18153
box 0 0 1 1
use contact_18  contact_18_71
timestamp 1643671299
transform 1 0 4632 0 1 19652
box 0 0 1 1
use contact_17  contact_17_71
timestamp 1643671299
transform 1 0 4647 0 1 19667
box 0 0 1 1
use contact_18  contact_18_72
timestamp 1643671299
transform 1 0 4632 0 1 18138
box 0 0 1 1
use contact_17  contact_17_72
timestamp 1643671299
transform 1 0 4647 0 1 18153
box 0 0 1 1
use contact_18  contact_18_73
timestamp 1643671299
transform 1 0 4632 0 1 16624
box 0 0 1 1
use contact_17  contact_17_73
timestamp 1643671299
transform 1 0 4647 0 1 16639
box 0 0 1 1
use contact_18  contact_18_74
timestamp 1643671299
transform 1 0 4632 0 1 15110
box 0 0 1 1
use contact_17  contact_17_74
timestamp 1643671299
transform 1 0 4647 0 1 15125
box 0 0 1 1
use contact_18  contact_18_75
timestamp 1643671299
transform 1 0 4632 0 1 16624
box 0 0 1 1
use contact_17  contact_17_75
timestamp 1643671299
transform 1 0 4647 0 1 16639
box 0 0 1 1
use contact_18  contact_18_76
timestamp 1643671299
transform 1 0 4632 0 1 15110
box 0 0 1 1
use contact_17  contact_17_76
timestamp 1643671299
transform 1 0 4647 0 1 15125
box 0 0 1 1
use contact_18  contact_18_77
timestamp 1643671299
transform 1 0 4632 0 1 13596
box 0 0 1 1
use contact_17  contact_17_77
timestamp 1643671299
transform 1 0 4647 0 1 13611
box 0 0 1 1
use contact_18  contact_18_78
timestamp 1643671299
transform 1 0 4632 0 1 12082
box 0 0 1 1
use contact_17  contact_17_78
timestamp 1643671299
transform 1 0 4647 0 1 12097
box 0 0 1 1
use contact_18  contact_18_79
timestamp 1643671299
transform 1 0 4632 0 1 13596
box 0 0 1 1
use contact_17  contact_17_79
timestamp 1643671299
transform 1 0 4647 0 1 13611
box 0 0 1 1
use contact_18  contact_18_80
timestamp 1643671299
transform 1 0 4632 0 1 12082
box 0 0 1 1
use contact_17  contact_17_80
timestamp 1643671299
transform 1 0 4647 0 1 12097
box 0 0 1 1
use contact_18  contact_18_81
timestamp 1643671299
transform 1 0 4632 0 1 10568
box 0 0 1 1
use contact_17  contact_17_81
timestamp 1643671299
transform 1 0 4647 0 1 10583
box 0 0 1 1
use contact_18  contact_18_82
timestamp 1643671299
transform 1 0 4632 0 1 9054
box 0 0 1 1
use contact_17  contact_17_82
timestamp 1643671299
transform 1 0 4647 0 1 9069
box 0 0 1 1
use contact_18  contact_18_83
timestamp 1643671299
transform 1 0 4632 0 1 10568
box 0 0 1 1
use contact_17  contact_17_83
timestamp 1643671299
transform 1 0 4647 0 1 10583
box 0 0 1 1
use contact_18  contact_18_84
timestamp 1643671299
transform 1 0 4632 0 1 9054
box 0 0 1 1
use contact_17  contact_17_84
timestamp 1643671299
transform 1 0 4647 0 1 9069
box 0 0 1 1
use contact_18  contact_18_85
timestamp 1643671299
transform 1 0 4632 0 1 7540
box 0 0 1 1
use contact_17  contact_17_85
timestamp 1643671299
transform 1 0 4647 0 1 7555
box 0 0 1 1
use contact_18  contact_18_86
timestamp 1643671299
transform 1 0 4632 0 1 6026
box 0 0 1 1
use contact_17  contact_17_86
timestamp 1643671299
transform 1 0 4647 0 1 6041
box 0 0 1 1
use contact_18  contact_18_87
timestamp 1643671299
transform 1 0 4632 0 1 7540
box 0 0 1 1
use contact_17  contact_17_87
timestamp 1643671299
transform 1 0 4647 0 1 7555
box 0 0 1 1
use contact_18  contact_18_88
timestamp 1643671299
transform 1 0 4632 0 1 6026
box 0 0 1 1
use contact_17  contact_17_88
timestamp 1643671299
transform 1 0 4647 0 1 6041
box 0 0 1 1
use contact_18  contact_18_89
timestamp 1643671299
transform 1 0 4632 0 1 4512
box 0 0 1 1
use contact_17  contact_17_89
timestamp 1643671299
transform 1 0 4647 0 1 4527
box 0 0 1 1
use contact_18  contact_18_90
timestamp 1643671299
transform 1 0 4632 0 1 2998
box 0 0 1 1
use contact_17  contact_17_90
timestamp 1643671299
transform 1 0 4647 0 1 3013
box 0 0 1 1
use contact_18  contact_18_91
timestamp 1643671299
transform 1 0 4632 0 1 4512
box 0 0 1 1
use contact_17  contact_17_91
timestamp 1643671299
transform 1 0 4647 0 1 4527
box 0 0 1 1
use contact_18  contact_18_92
timestamp 1643671299
transform 1 0 4632 0 1 2998
box 0 0 1 1
use contact_17  contact_17_92
timestamp 1643671299
transform 1 0 4647 0 1 3013
box 0 0 1 1
use contact_18  contact_18_93
timestamp 1643671299
transform 1 0 4632 0 1 1484
box 0 0 1 1
use contact_17  contact_17_93
timestamp 1643671299
transform 1 0 4647 0 1 1499
box 0 0 1 1
use contact_18  contact_18_94
timestamp 1643671299
transform 1 0 4632 0 1 -30
box 0 0 1 1
use contact_17  contact_17_94
timestamp 1643671299
transform 1 0 4647 0 1 -15
box 0 0 1 1
use contact_18  contact_18_95
timestamp 1643671299
transform 1 0 4632 0 1 1484
box 0 0 1 1
use contact_17  contact_17_95
timestamp 1643671299
transform 1 0 4647 0 1 1499
box 0 0 1 1
use contact_20  contact_20_0
timestamp 1643671299
transform 1 0 3070 0 1 23062
box 0 0 1 1
use contact_18  contact_18_96
timestamp 1643671299
transform 1 0 2102 0 1 23874
box 0 0 1 1
use contact_17  contact_17_96
timestamp 1643671299
transform 1 0 2117 0 1 23889
box 0 0 1 1
use contact_13  contact_13_0
timestamp 1643671299
transform 1 0 2103 0 1 23881
box 0 0 1 1
use contact_20  contact_20_1
timestamp 1643671299
transform 1 0 3002 0 1 21522
box 0 0 1 1
use contact_18  contact_18_97
timestamp 1643671299
transform 1 0 2102 0 1 22250
box 0 0 1 1
use contact_17  contact_17_97
timestamp 1643671299
transform 1 0 2117 0 1 22265
box 0 0 1 1
use contact_13  contact_13_1
timestamp 1643671299
transform 1 0 2103 0 1 22257
box 0 0 1 1
use contact_20  contact_20_2
timestamp 1643671299
transform 1 0 2934 0 1 19982
box 0 0 1 1
use contact_18  contact_18_98
timestamp 1643671299
transform 1 0 2102 0 1 20794
box 0 0 1 1
use contact_17  contact_17_98
timestamp 1643671299
transform 1 0 2117 0 1 20809
box 0 0 1 1
use contact_13  contact_13_2
timestamp 1643671299
transform 1 0 2103 0 1 20801
box 0 0 1 1
use contact_20  contact_20_3
timestamp 1643671299
transform 1 0 2866 0 1 18442
box 0 0 1 1
use contact_18  contact_18_99
timestamp 1643671299
transform 1 0 2102 0 1 19170
box 0 0 1 1
use contact_17  contact_17_99
timestamp 1643671299
transform 1 0 2117 0 1 19185
box 0 0 1 1
use contact_13  contact_13_3
timestamp 1643671299
transform 1 0 2103 0 1 19177
box 0 0 1 1
use contact_20  contact_20_4
timestamp 1643671299
transform 1 0 2798 0 1 13826
box 0 0 1 1
use contact_18  contact_18_100
timestamp 1643671299
transform 1 0 2102 0 1 14638
box 0 0 1 1
use contact_17  contact_17_100
timestamp 1643671299
transform 1 0 2117 0 1 14653
box 0 0 1 1
use contact_13  contact_13_4
timestamp 1643671299
transform 1 0 2103 0 1 14645
box 0 0 1 1
use contact_20  contact_20_5
timestamp 1643671299
transform 1 0 2730 0 1 12286
box 0 0 1 1
use contact_18  contact_18_101
timestamp 1643671299
transform 1 0 2102 0 1 13014
box 0 0 1 1
use contact_17  contact_17_101
timestamp 1643671299
transform 1 0 2117 0 1 13029
box 0 0 1 1
use contact_13  contact_13_5
timestamp 1643671299
transform 1 0 2103 0 1 13021
box 0 0 1 1
use contact_20  contact_20_6
timestamp 1643671299
transform 1 0 2662 0 1 10746
box 0 0 1 1
use contact_18  contact_18_102
timestamp 1643671299
transform 1 0 2102 0 1 11558
box 0 0 1 1
use contact_17  contact_17_102
timestamp 1643671299
transform 1 0 2117 0 1 11573
box 0 0 1 1
use contact_13  contact_13_6
timestamp 1643671299
transform 1 0 2103 0 1 11565
box 0 0 1 1
use contact_20  contact_20_7
timestamp 1643671299
transform 1 0 2594 0 1 9206
box 0 0 1 1
use contact_18  contact_18_103
timestamp 1643671299
transform 1 0 2102 0 1 9934
box 0 0 1 1
use contact_17  contact_17_103
timestamp 1643671299
transform 1 0 2117 0 1 9949
box 0 0 1 1
use contact_13  contact_13_7
timestamp 1643671299
transform 1 0 2103 0 1 9941
box 0 0 1 1
use contact_20  contact_20_8
timestamp 1643671299
transform 1 0 2526 0 1 4590
box 0 0 1 1
use contact_18  contact_18_104
timestamp 1643671299
transform 1 0 2102 0 1 5402
box 0 0 1 1
use contact_17  contact_17_104
timestamp 1643671299
transform 1 0 2117 0 1 5417
box 0 0 1 1
use contact_13  contact_13_8
timestamp 1643671299
transform 1 0 2103 0 1 5409
box 0 0 1 1
use contact_20  contact_20_9
timestamp 1643671299
transform 1 0 2458 0 1 3050
box 0 0 1 1
use contact_18  contact_18_105
timestamp 1643671299
transform 1 0 2102 0 1 3778
box 0 0 1 1
use contact_17  contact_17_105
timestamp 1643671299
transform 1 0 2117 0 1 3793
box 0 0 1 1
use contact_13  contact_13_9
timestamp 1643671299
transform 1 0 2103 0 1 3785
box 0 0 1 1
use contact_20  contact_20_10
timestamp 1643671299
transform 1 0 2390 0 1 1510
box 0 0 1 1
use contact_18  contact_18_106
timestamp 1643671299
transform 1 0 2102 0 1 2322
box 0 0 1 1
use contact_17  contact_17_106
timestamp 1643671299
transform 1 0 2117 0 1 2337
box 0 0 1 1
use contact_13  contact_13_10
timestamp 1643671299
transform 1 0 2103 0 1 2329
box 0 0 1 1
use contact_20  contact_20_11
timestamp 1643671299
transform 1 0 2322 0 1 -30
box 0 0 1 1
use contact_18  contact_18_107
timestamp 1643671299
transform 1 0 2102 0 1 698
box 0 0 1 1
use contact_17  contact_17_107
timestamp 1643671299
transform 1 0 2117 0 1 713
box 0 0 1 1
use contact_13  contact_13_11
timestamp 1643671299
transform 1 0 2103 0 1 705
box 0 0 1 1
use contact_14  contact_14_0
timestamp 1643671299
transform 1 0 3017 0 1 801
box 0 0 1 1
use contact_14  contact_14_1
timestamp 1643671299
transform 1 0 2813 0 1 857
box 0 0 1 1
use contact_14  contact_14_2
timestamp 1643671299
transform 1 0 2541 0 1 913
box 0 0 1 1
use contact_14  contact_14_3
timestamp 1643671299
transform 1 0 3017 0 1 23729
box 0 0 1 1
use contact_14  contact_14_4
timestamp 1643671299
transform 1 0 2813 0 1 23673
box 0 0 1 1
use contact_14  contact_14_5
timestamp 1643671299
transform 1 0 2473 0 1 23617
box 0 0 1 1
use contact_14  contact_14_6
timestamp 1643671299
transform 1 0 3017 0 1 23561
box 0 0 1 1
use contact_14  contact_14_7
timestamp 1643671299
transform 1 0 2813 0 1 23505
box 0 0 1 1
use contact_14  contact_14_8
timestamp 1643671299
transform 1 0 2405 0 1 23449
box 0 0 1 1
use contact_14  contact_14_9
timestamp 1643671299
transform 1 0 3017 0 1 23393
box 0 0 1 1
use contact_14  contact_14_10
timestamp 1643671299
transform 1 0 2813 0 1 23337
box 0 0 1 1
use contact_14  contact_14_11
timestamp 1643671299
transform 1 0 2337 0 1 23281
box 0 0 1 1
use contact_14  contact_14_12
timestamp 1643671299
transform 1 0 3017 0 1 21661
box 0 0 1 1
use contact_14  contact_14_13
timestamp 1643671299
transform 1 0 2745 0 1 21717
box 0 0 1 1
use contact_14  contact_14_14
timestamp 1643671299
transform 1 0 2541 0 1 21773
box 0 0 1 1
use contact_14  contact_14_15
timestamp 1643671299
transform 1 0 3017 0 1 21829
box 0 0 1 1
use contact_14  contact_14_16
timestamp 1643671299
transform 1 0 2745 0 1 21885
box 0 0 1 1
use contact_14  contact_14_17
timestamp 1643671299
transform 1 0 2473 0 1 21941
box 0 0 1 1
use contact_14  contact_14_18
timestamp 1643671299
transform 1 0 3017 0 1 21997
box 0 0 1 1
use contact_14  contact_14_19
timestamp 1643671299
transform 1 0 2745 0 1 22053
box 0 0 1 1
use contact_14  contact_14_20
timestamp 1643671299
transform 1 0 2405 0 1 22109
box 0 0 1 1
use contact_14  contact_14_21
timestamp 1643671299
transform 1 0 3017 0 1 20701
box 0 0 1 1
use contact_14  contact_14_22
timestamp 1643671299
transform 1 0 2745 0 1 20645
box 0 0 1 1
use contact_14  contact_14_23
timestamp 1643671299
transform 1 0 2337 0 1 20589
box 0 0 1 1
use contact_14  contact_14_24
timestamp 1643671299
transform 1 0 3017 0 1 20533
box 0 0 1 1
use contact_14  contact_14_25
timestamp 1643671299
transform 1 0 2677 0 1 20477
box 0 0 1 1
use contact_14  contact_14_26
timestamp 1643671299
transform 1 0 2541 0 1 20421
box 0 0 1 1
use contact_14  contact_14_27
timestamp 1643671299
transform 1 0 3017 0 1 20365
box 0 0 1 1
use contact_14  contact_14_28
timestamp 1643671299
transform 1 0 2677 0 1 20309
box 0 0 1 1
use contact_14  contact_14_29
timestamp 1643671299
transform 1 0 2473 0 1 20253
box 0 0 1 1
use contact_14  contact_14_30
timestamp 1643671299
transform 1 0 3017 0 1 18633
box 0 0 1 1
use contact_14  contact_14_31
timestamp 1643671299
transform 1 0 2677 0 1 18689
box 0 0 1 1
use contact_14  contact_14_32
timestamp 1643671299
transform 1 0 2405 0 1 18745
box 0 0 1 1
use contact_14  contact_14_33
timestamp 1643671299
transform 1 0 3017 0 1 18801
box 0 0 1 1
use contact_14  contact_14_34
timestamp 1643671299
transform 1 0 2677 0 1 18857
box 0 0 1 1
use contact_14  contact_14_35
timestamp 1643671299
transform 1 0 2337 0 1 18913
box 0 0 1 1
use contact_14  contact_14_36
timestamp 1643671299
transform 1 0 3017 0 1 18969
box 0 0 1 1
use contact_14  contact_14_37
timestamp 1643671299
transform 1 0 2609 0 1 19025
box 0 0 1 1
use contact_14  contact_14_38
timestamp 1643671299
transform 1 0 2541 0 1 19081
box 0 0 1 1
use contact_14  contact_14_39
timestamp 1643671299
transform 1 0 3017 0 1 17673
box 0 0 1 1
use contact_14  contact_14_40
timestamp 1643671299
transform 1 0 2609 0 1 17617
box 0 0 1 1
use contact_14  contact_14_41
timestamp 1643671299
transform 1 0 2473 0 1 17561
box 0 0 1 1
use contact_14  contact_14_42
timestamp 1643671299
transform 1 0 3017 0 1 17505
box 0 0 1 1
use contact_14  contact_14_43
timestamp 1643671299
transform 1 0 2609 0 1 17449
box 0 0 1 1
use contact_14  contact_14_44
timestamp 1643671299
transform 1 0 2405 0 1 17393
box 0 0 1 1
use contact_14  contact_14_45
timestamp 1643671299
transform 1 0 3017 0 1 17337
box 0 0 1 1
use contact_14  contact_14_46
timestamp 1643671299
transform 1 0 2609 0 1 17281
box 0 0 1 1
use contact_14  contact_14_47
timestamp 1643671299
transform 1 0 2337 0 1 17225
box 0 0 1 1
use contact_14  contact_14_48
timestamp 1643671299
transform 1 0 2949 0 1 15605
box 0 0 1 1
use contact_14  contact_14_49
timestamp 1643671299
transform 1 0 2813 0 1 15661
box 0 0 1 1
use contact_14  contact_14_50
timestamp 1643671299
transform 1 0 2541 0 1 15717
box 0 0 1 1
use contact_14  contact_14_51
timestamp 1643671299
transform 1 0 2949 0 1 15773
box 0 0 1 1
use contact_14  contact_14_52
timestamp 1643671299
transform 1 0 2813 0 1 15829
box 0 0 1 1
use contact_14  contact_14_53
timestamp 1643671299
transform 1 0 2473 0 1 15885
box 0 0 1 1
use contact_14  contact_14_54
timestamp 1643671299
transform 1 0 2949 0 1 15941
box 0 0 1 1
use contact_14  contact_14_55
timestamp 1643671299
transform 1 0 2813 0 1 15997
box 0 0 1 1
use contact_14  contact_14_56
timestamp 1643671299
transform 1 0 2405 0 1 16053
box 0 0 1 1
use contact_14  contact_14_57
timestamp 1643671299
transform 1 0 2949 0 1 14645
box 0 0 1 1
use contact_14  contact_14_58
timestamp 1643671299
transform 1 0 2813 0 1 14589
box 0 0 1 1
use contact_14  contact_14_59
timestamp 1643671299
transform 1 0 2337 0 1 14533
box 0 0 1 1
use contact_14  contact_14_60
timestamp 1643671299
transform 1 0 2949 0 1 14477
box 0 0 1 1
use contact_14  contact_14_61
timestamp 1643671299
transform 1 0 2745 0 1 14421
box 0 0 1 1
use contact_14  contact_14_62
timestamp 1643671299
transform 1 0 2541 0 1 14365
box 0 0 1 1
use contact_14  contact_14_63
timestamp 1643671299
transform 1 0 2949 0 1 14309
box 0 0 1 1
use contact_14  contact_14_64
timestamp 1643671299
transform 1 0 2745 0 1 14253
box 0 0 1 1
use contact_14  contact_14_65
timestamp 1643671299
transform 1 0 2473 0 1 14197
box 0 0 1 1
use contact_14  contact_14_66
timestamp 1643671299
transform 1 0 2949 0 1 12577
box 0 0 1 1
use contact_14  contact_14_67
timestamp 1643671299
transform 1 0 2745 0 1 12633
box 0 0 1 1
use contact_14  contact_14_68
timestamp 1643671299
transform 1 0 2405 0 1 12689
box 0 0 1 1
use contact_14  contact_14_69
timestamp 1643671299
transform 1 0 2949 0 1 12745
box 0 0 1 1
use contact_14  contact_14_70
timestamp 1643671299
transform 1 0 2745 0 1 12801
box 0 0 1 1
use contact_14  contact_14_71
timestamp 1643671299
transform 1 0 2337 0 1 12857
box 0 0 1 1
use contact_14  contact_14_72
timestamp 1643671299
transform 1 0 2949 0 1 12913
box 0 0 1 1
use contact_14  contact_14_73
timestamp 1643671299
transform 1 0 2677 0 1 12969
box 0 0 1 1
use contact_14  contact_14_74
timestamp 1643671299
transform 1 0 2541 0 1 13025
box 0 0 1 1
use contact_14  contact_14_75
timestamp 1643671299
transform 1 0 2949 0 1 11617
box 0 0 1 1
use contact_14  contact_14_76
timestamp 1643671299
transform 1 0 2677 0 1 11561
box 0 0 1 1
use contact_14  contact_14_77
timestamp 1643671299
transform 1 0 2473 0 1 11505
box 0 0 1 1
use contact_14  contact_14_78
timestamp 1643671299
transform 1 0 2949 0 1 11449
box 0 0 1 1
use contact_14  contact_14_79
timestamp 1643671299
transform 1 0 2677 0 1 11393
box 0 0 1 1
use contact_14  contact_14_80
timestamp 1643671299
transform 1 0 2405 0 1 11337
box 0 0 1 1
use contact_14  contact_14_81
timestamp 1643671299
transform 1 0 2949 0 1 11281
box 0 0 1 1
use contact_14  contact_14_82
timestamp 1643671299
transform 1 0 2677 0 1 11225
box 0 0 1 1
use contact_14  contact_14_83
timestamp 1643671299
transform 1 0 2337 0 1 11169
box 0 0 1 1
use contact_14  contact_14_84
timestamp 1643671299
transform 1 0 2949 0 1 9549
box 0 0 1 1
use contact_14  contact_14_85
timestamp 1643671299
transform 1 0 2609 0 1 9605
box 0 0 1 1
use contact_14  contact_14_86
timestamp 1643671299
transform 1 0 2541 0 1 9661
box 0 0 1 1
use contact_14  contact_14_87
timestamp 1643671299
transform 1 0 2949 0 1 9717
box 0 0 1 1
use contact_14  contact_14_88
timestamp 1643671299
transform 1 0 2609 0 1 9773
box 0 0 1 1
use contact_14  contact_14_89
timestamp 1643671299
transform 1 0 2473 0 1 9829
box 0 0 1 1
use contact_14  contact_14_90
timestamp 1643671299
transform 1 0 2949 0 1 9885
box 0 0 1 1
use contact_14  contact_14_91
timestamp 1643671299
transform 1 0 2609 0 1 9941
box 0 0 1 1
use contact_14  contact_14_92
timestamp 1643671299
transform 1 0 2405 0 1 9997
box 0 0 1 1
use contact_14  contact_14_93
timestamp 1643671299
transform 1 0 2949 0 1 8589
box 0 0 1 1
use contact_14  contact_14_94
timestamp 1643671299
transform 1 0 2609 0 1 8533
box 0 0 1 1
use contact_14  contact_14_95
timestamp 1643671299
transform 1 0 2337 0 1 8477
box 0 0 1 1
use contact_14  contact_14_96
timestamp 1643671299
transform 1 0 2881 0 1 8421
box 0 0 1 1
use contact_14  contact_14_97
timestamp 1643671299
transform 1 0 2813 0 1 8365
box 0 0 1 1
use contact_14  contact_14_98
timestamp 1643671299
transform 1 0 2541 0 1 8309
box 0 0 1 1
use contact_14  contact_14_99
timestamp 1643671299
transform 1 0 2881 0 1 8253
box 0 0 1 1
use contact_14  contact_14_100
timestamp 1643671299
transform 1 0 2813 0 1 8197
box 0 0 1 1
use contact_14  contact_14_101
timestamp 1643671299
transform 1 0 2473 0 1 8141
box 0 0 1 1
use contact_14  contact_14_102
timestamp 1643671299
transform 1 0 2881 0 1 6521
box 0 0 1 1
use contact_14  contact_14_103
timestamp 1643671299
transform 1 0 2813 0 1 6577
box 0 0 1 1
use contact_14  contact_14_104
timestamp 1643671299
transform 1 0 2405 0 1 6633
box 0 0 1 1
use contact_14  contact_14_105
timestamp 1643671299
transform 1 0 2881 0 1 6689
box 0 0 1 1
use contact_14  contact_14_106
timestamp 1643671299
transform 1 0 2813 0 1 6745
box 0 0 1 1
use contact_14  contact_14_107
timestamp 1643671299
transform 1 0 2337 0 1 6801
box 0 0 1 1
use contact_14  contact_14_108
timestamp 1643671299
transform 1 0 2881 0 1 6857
box 0 0 1 1
use contact_14  contact_14_109
timestamp 1643671299
transform 1 0 2745 0 1 6913
box 0 0 1 1
use contact_14  contact_14_110
timestamp 1643671299
transform 1 0 2541 0 1 6969
box 0 0 1 1
use contact_14  contact_14_111
timestamp 1643671299
transform 1 0 2881 0 1 5561
box 0 0 1 1
use contact_14  contact_14_112
timestamp 1643671299
transform 1 0 2745 0 1 5505
box 0 0 1 1
use contact_14  contact_14_113
timestamp 1643671299
transform 1 0 2473 0 1 5449
box 0 0 1 1
use contact_14  contact_14_114
timestamp 1643671299
transform 1 0 2881 0 1 5393
box 0 0 1 1
use contact_14  contact_14_115
timestamp 1643671299
transform 1 0 2745 0 1 5337
box 0 0 1 1
use contact_14  contact_14_116
timestamp 1643671299
transform 1 0 2405 0 1 5281
box 0 0 1 1
use contact_14  contact_14_117
timestamp 1643671299
transform 1 0 2881 0 1 5225
box 0 0 1 1
use contact_14  contact_14_118
timestamp 1643671299
transform 1 0 2745 0 1 5169
box 0 0 1 1
use contact_14  contact_14_119
timestamp 1643671299
transform 1 0 2337 0 1 5113
box 0 0 1 1
use contact_14  contact_14_120
timestamp 1643671299
transform 1 0 2881 0 1 3493
box 0 0 1 1
use contact_14  contact_14_121
timestamp 1643671299
transform 1 0 2677 0 1 3549
box 0 0 1 1
use contact_14  contact_14_122
timestamp 1643671299
transform 1 0 2541 0 1 3605
box 0 0 1 1
use contact_14  contact_14_123
timestamp 1643671299
transform 1 0 2881 0 1 3661
box 0 0 1 1
use contact_14  contact_14_124
timestamp 1643671299
transform 1 0 2677 0 1 3717
box 0 0 1 1
use contact_14  contact_14_125
timestamp 1643671299
transform 1 0 2473 0 1 3773
box 0 0 1 1
use contact_14  contact_14_126
timestamp 1643671299
transform 1 0 2881 0 1 3829
box 0 0 1 1
use contact_14  contact_14_127
timestamp 1643671299
transform 1 0 2677 0 1 3885
box 0 0 1 1
use contact_14  contact_14_128
timestamp 1643671299
transform 1 0 2405 0 1 3941
box 0 0 1 1
use contact_14  contact_14_129
timestamp 1643671299
transform 1 0 2881 0 1 2533
box 0 0 1 1
use contact_14  contact_14_130
timestamp 1643671299
transform 1 0 2677 0 1 2477
box 0 0 1 1
use contact_14  contact_14_131
timestamp 1643671299
transform 1 0 2337 0 1 2421
box 0 0 1 1
use contact_14  contact_14_132
timestamp 1643671299
transform 1 0 2881 0 1 2365
box 0 0 1 1
use contact_14  contact_14_133
timestamp 1643671299
transform 1 0 2609 0 1 2309
box 0 0 1 1
use contact_14  contact_14_134
timestamp 1643671299
transform 1 0 2541 0 1 2253
box 0 0 1 1
use contact_14  contact_14_135
timestamp 1643671299
transform 1 0 2881 0 1 2197
box 0 0 1 1
use contact_14  contact_14_136
timestamp 1643671299
transform 1 0 2609 0 1 2141
box 0 0 1 1
use contact_14  contact_14_137
timestamp 1643671299
transform 1 0 2473 0 1 2085
box 0 0 1 1
use contact_14  contact_14_138
timestamp 1643671299
transform 1 0 2881 0 1 465
box 0 0 1 1
use contact_14  contact_14_139
timestamp 1643671299
transform 1 0 2609 0 1 521
box 0 0 1 1
use contact_14  contact_14_140
timestamp 1643671299
transform 1 0 2405 0 1 577
box 0 0 1 1
use contact_14  contact_14_141
timestamp 1643671299
transform 1 0 2881 0 1 633
box 0 0 1 1
use contact_14  contact_14_142
timestamp 1643671299
transform 1 0 2609 0 1 689
box 0 0 1 1
use contact_14  contact_14_143
timestamp 1643671299
transform 1 0 2337 0 1 745
box 0 0 1 1
use contact_14  contact_14_144
timestamp 1643671299
transform 1 0 340 0 1 20809
box 0 0 1 1
use contact_17  contact_17_108
timestamp 1643671299
transform 1 0 572 0 1 20809
box 0 0 1 1
use contact_14  contact_14_145
timestamp 1643671299
transform 1 0 272 0 1 19185
box 0 0 1 1
use contact_17  contact_17_109
timestamp 1643671299
transform 1 0 504 0 1 19185
box 0 0 1 1
use contact_14  contact_14_146
timestamp 1643671299
transform 1 0 204 0 1 11573
box 0 0 1 1
use contact_17  contact_17_110
timestamp 1643671299
transform 1 0 572 0 1 11573
box 0 0 1 1
use contact_14  contact_14_147
timestamp 1643671299
transform 1 0 136 0 1 9949
box 0 0 1 1
use contact_17  contact_17_111
timestamp 1643671299
transform 1 0 504 0 1 9949
box 0 0 1 1
use contact_14  contact_14_148
timestamp 1643671299
transform 1 0 68 0 1 2337
box 0 0 1 1
use contact_17  contact_17_112
timestamp 1643671299
transform 1 0 572 0 1 2337
box 0 0 1 1
use contact_14  contact_14_149
timestamp 1643671299
transform 1 0 0 0 1 713
box 0 0 1 1
use contact_17  contact_17_113
timestamp 1643671299
transform 1 0 504 0 1 713
box 0 0 1 1
use dec_cell3_2r1w  dec_cell3_2r1w_0
timestamp 1643671299
transform 1 0 2270 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_1
timestamp 1643671299
transform 1 0 2270 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_2
timestamp 1643671299
transform 1 0 2270 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_3
timestamp 1643671299
transform 1 0 2270 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_4
timestamp 1643671299
transform 1 0 2270 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_5
timestamp 1643671299
transform 1 0 2270 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_6
timestamp 1643671299
transform 1 0 2270 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_7
timestamp 1643671299
transform 1 0 2270 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_8
timestamp 1643671299
transform 1 0 2270 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_9
timestamp 1643671299
transform 1 0 2270 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_10
timestamp 1643671299
transform 1 0 2270 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_11
timestamp 1643671299
transform 1 0 2270 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_12
timestamp 1643671299
transform 1 0 2270 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_13
timestamp 1643671299
transform 1 0 2270 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_14
timestamp 1643671299
transform 1 0 2270 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_15
timestamp 1643671299
transform 1 0 2270 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_16
timestamp 1643671299
transform 1 0 2270 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_17
timestamp 1643671299
transform 1 0 2270 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_18
timestamp 1643671299
transform 1 0 2270 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_19
timestamp 1643671299
transform 1 0 2270 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_20
timestamp 1643671299
transform 1 0 2270 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_21
timestamp 1643671299
transform 1 0 2270 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_22
timestamp 1643671299
transform 1 0 2270 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_23
timestamp 1643671299
transform 1 0 2270 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_24
timestamp 1643671299
transform 1 0 2270 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_25
timestamp 1643671299
transform 1 0 2270 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_26
timestamp 1643671299
transform 1 0 2270 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_27
timestamp 1643671299
transform 1 0 2270 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_28
timestamp 1643671299
transform 1 0 2270 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_29
timestamp 1643671299
transform 1 0 2270 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_30
timestamp 1643671299
transform 1 0 2270 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_31
timestamp 1643671299
transform 1 0 2270 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_32
timestamp 1643671299
transform 1 0 3154 0 -1 24224
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_33
timestamp 1643671299
transform 1 0 3154 0 1 21196
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_34
timestamp 1643671299
transform 1 0 3154 0 -1 21196
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_35
timestamp 1643671299
transform 1 0 3154 0 1 18168
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_36
timestamp 1643671299
transform 1 0 3154 0 -1 18168
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_37
timestamp 1643671299
transform 1 0 3154 0 1 15140
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_38
timestamp 1643671299
transform 1 0 3154 0 -1 15140
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_39
timestamp 1643671299
transform 1 0 3154 0 1 12112
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_40
timestamp 1643671299
transform 1 0 3154 0 -1 12112
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_41
timestamp 1643671299
transform 1 0 3154 0 1 9084
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_42
timestamp 1643671299
transform 1 0 3154 0 -1 9084
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_43
timestamp 1643671299
transform 1 0 3154 0 1 6056
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_44
timestamp 1643671299
transform 1 0 3154 0 -1 6056
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_45
timestamp 1643671299
transform 1 0 3154 0 1 3028
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_46
timestamp 1643671299
transform 1 0 3154 0 -1 3028
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_47
timestamp 1643671299
transform 1 0 3154 0 1 0
box 0 -42 1494 1616
use hierarchical_predecode2x4  hierarchical_predecode2x4_0
timestamp 1643671299
transform 1 0 437 0 1 18472
box 0 -34 1869 6194
use hierarchical_predecode2x4  hierarchical_predecode2x4_1
timestamp 1643671299
transform 1 0 437 0 1 9236
box 0 -34 1869 6194
use hierarchical_predecode2x4  hierarchical_predecode2x4_2
timestamp 1643671299
transform 1 0 437 0 1 0
box 0 -34 1869 6194
<< labels >>
rlabel metal2 s 1 0 29 24632 4 addr_0
rlabel metal2 s 69 0 97 24632 4 addr_1
rlabel metal2 s 137 0 165 24632 4 addr_2
rlabel metal2 s 205 0 233 24632 4 addr_3
rlabel metal2 s 273 0 301 24632 4 addr_4
rlabel metal2 s 341 0 369 24632 4 addr_5
rlabel metal1 s 4364 702 4648 730 4 decode0_0
rlabel metal1 s 4572 848 4648 876 4 decode1_0
rlabel metal1 s 4282 580 4648 608 4 decode2_0
rlabel metal1 s 4364 2298 4648 2326 4 decode0_1
rlabel metal1 s 4572 2152 4648 2180 4 decode1_1
rlabel metal1 s 4282 2420 4648 2448 4 decode2_1
rlabel metal1 s 4364 3730 4648 3758 4 decode0_2
rlabel metal1 s 4572 3876 4648 3904 4 decode1_2
rlabel metal1 s 4282 3608 4648 3636 4 decode2_2
rlabel metal1 s 4364 5326 4648 5354 4 decode0_3
rlabel metal1 s 4572 5180 4648 5208 4 decode1_3
rlabel metal1 s 4282 5448 4648 5476 4 decode2_3
rlabel metal1 s 4364 6758 4648 6786 4 decode0_4
rlabel metal1 s 4572 6904 4648 6932 4 decode1_4
rlabel metal1 s 4282 6636 4648 6664 4 decode2_4
rlabel metal1 s 4364 8354 4648 8382 4 decode0_5
rlabel metal1 s 4572 8208 4648 8236 4 decode1_5
rlabel metal1 s 4282 8476 4648 8504 4 decode2_5
rlabel metal1 s 4364 9786 4648 9814 4 decode0_6
rlabel metal1 s 4572 9932 4648 9960 4 decode1_6
rlabel metal1 s 4282 9664 4648 9692 4 decode2_6
rlabel metal1 s 4364 11382 4648 11410 4 decode0_7
rlabel metal1 s 4572 11236 4648 11264 4 decode1_7
rlabel metal1 s 4282 11504 4648 11532 4 decode2_7
rlabel metal1 s 4364 12814 4648 12842 4 decode0_8
rlabel metal1 s 4572 12960 4648 12988 4 decode1_8
rlabel metal1 s 4282 12692 4648 12720 4 decode2_8
rlabel metal1 s 4364 14410 4648 14438 4 decode0_9
rlabel metal1 s 4572 14264 4648 14292 4 decode1_9
rlabel metal1 s 4282 14532 4648 14560 4 decode2_9
rlabel metal1 s 4364 15842 4648 15870 4 decode0_10
rlabel metal1 s 4572 15988 4648 16016 4 decode1_10
rlabel metal1 s 4282 15720 4648 15748 4 decode2_10
rlabel metal1 s 4364 17438 4648 17466 4 decode0_11
rlabel metal1 s 4572 17292 4648 17320 4 decode1_11
rlabel metal1 s 4282 17560 4648 17588 4 decode2_11
rlabel metal1 s 4364 18870 4648 18898 4 decode0_12
rlabel metal1 s 4572 19016 4648 19044 4 decode1_12
rlabel metal1 s 4282 18748 4648 18776 4 decode2_12
rlabel metal1 s 4364 20466 4648 20494 4 decode0_13
rlabel metal1 s 4572 20320 4648 20348 4 decode1_13
rlabel metal1 s 4282 20588 4648 20616 4 decode2_13
rlabel metal1 s 4364 21898 4648 21926 4 decode0_14
rlabel metal1 s 4572 22044 4648 22072 4 decode1_14
rlabel metal1 s 4282 21776 4648 21804 4 decode2_14
rlabel metal1 s 4364 23494 4648 23522 4 decode0_15
rlabel metal1 s 4572 23348 4648 23376 4 decode1_15
rlabel metal1 s 4282 23616 4648 23644 4 decode2_15
rlabel metal2 s 2338 0 2366 24660 4 predecode_0
rlabel metal2 s 2406 0 2434 24660 4 predecode_1
rlabel metal2 s 2474 0 2502 24660 4 predecode_2
rlabel metal2 s 2542 0 2570 24660 4 predecode_3
rlabel metal2 s 2610 0 2638 24660 4 predecode_4
rlabel metal2 s 2678 0 2706 24660 4 predecode_5
rlabel metal2 s 2746 0 2774 24660 4 predecode_6
rlabel metal2 s 2814 0 2842 24660 4 predecode_7
rlabel metal2 s 2882 0 2910 24660 4 predecode_8
rlabel metal2 s 2950 0 2978 24660 4 predecode_9
rlabel metal2 s 3018 0 3046 24660 4 predecode_10
rlabel metal2 s 3086 0 3114 24660 4 predecode_11
rlabel metal3 s 651 23062 711 23122 4 vdd
rlabel metal3 s 1410 1510 1470 1570 4 vdd
rlabel metal3 s 4632 4512 4692 4572 4 vdd
rlabel metal3 s 651 4590 711 4650 4 vdd
rlabel metal3 s 1410 13826 1470 13886 4 vdd
rlabel metal3 s 4632 16624 4692 16684 4 vdd
rlabel metal3 s 1410 10746 1470 10806 4 vdd
rlabel metal3 s 1410 19982 1470 20042 4 vdd
rlabel metal3 s 4632 1484 4692 1544 4 vdd
rlabel metal3 s 4632 22680 4692 22740 4 vdd
rlabel metal3 s 651 13826 711 13886 4 vdd
rlabel metal3 s 4632 13596 4692 13656 4 vdd
rlabel metal3 s 4632 7540 4692 7600 4 vdd
rlabel metal3 s 4632 10568 4692 10628 4 vdd
rlabel metal3 s 1410 23062 1470 23122 4 vdd
rlabel metal3 s 651 10746 711 10806 4 vdd
rlabel metal3 s 4632 19652 4692 19712 4 vdd
rlabel metal3 s 1410 4590 1470 4650 4 vdd
rlabel metal3 s 651 19982 711 20042 4 vdd
rlabel metal3 s 651 1510 711 1570 4 vdd
rlabel metal3 s 1410 18442 1470 18502 4 gnd
rlabel metal3 s 4632 -30 4692 30 4 gnd
rlabel metal3 s 651 15366 711 15426 4 gnd
rlabel metal3 s 651 12286 711 12346 4 gnd
rlabel metal3 s 1410 15366 1470 15426 4 gnd
rlabel metal3 s 651 -30 711 30 4 gnd
rlabel metal3 s 651 3050 711 3110 4 gnd
rlabel metal3 s 1410 21522 1470 21582 4 gnd
rlabel metal3 s 4632 6026 4692 6086 4 gnd
rlabel metal3 s 651 21522 711 21582 4 gnd
rlabel metal3 s 651 24602 711 24662 4 gnd
rlabel metal3 s 1410 -30 1470 30 4 gnd
rlabel metal3 s 4632 21166 4692 21226 4 gnd
rlabel metal3 s 1410 6130 1470 6190 4 gnd
rlabel metal3 s 4632 9054 4692 9114 4 gnd
rlabel metal3 s 4632 18138 4692 18198 4 gnd
rlabel metal3 s 1410 12286 1470 12346 4 gnd
rlabel metal3 s 4632 15110 4692 15170 4 gnd
rlabel metal3 s 1410 3050 1470 3110 4 gnd
rlabel metal3 s 1410 24602 1470 24662 4 gnd
rlabel metal3 s 1410 9206 1470 9266 4 gnd
rlabel metal3 s 4632 12082 4692 12142 4 gnd
rlabel metal3 s 4632 2998 4692 3058 4 gnd
rlabel metal3 s 4632 24194 4692 24254 4 gnd
rlabel metal3 s 651 18442 711 18502 4 gnd
rlabel metal3 s 651 6130 711 6190 4 gnd
rlabel metal3 s 651 9206 711 9266 4 gnd
<< properties >>
string FIXED_BBOX 4632 -30 4692 0
string GDS_FILE sram_0rw2r1w_16_32_sky130A.gds
string GDS_END 1004136
string GDS_START 935670
<< end >>
