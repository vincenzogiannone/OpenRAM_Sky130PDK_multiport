magic
tech sky130A
magscale 1 2
timestamp 1644951705
<< checkpaint >>
rect -1296 -1277 5876 2155
<< nwell >>
rect -36 402 4616 895
<< pwell >>
rect 4470 51 4520 133
<< psubdiff >>
rect 4470 109 4520 133
rect 4470 75 4478 109
rect 4512 75 4520 109
rect 4470 51 4520 75
<< nsubdiff >>
rect 4470 763 4520 787
rect 4470 729 4478 763
rect 4512 729 4520 763
rect 4470 705 4520 729
<< psubdiffcont >>
rect 4478 75 4512 109
<< nsubdiffcont >>
rect 4478 729 4512 763
<< poly >>
rect 114 402 144 435
rect 48 386 144 402
rect 48 352 64 386
rect 98 352 144 386
rect 48 336 144 352
rect 114 206 144 336
<< polycont >>
rect 64 352 98 386
<< locali >>
rect 0 821 4580 855
rect 62 606 96 821
rect 274 606 308 821
rect 490 606 524 821
rect 706 606 740 821
rect 922 606 956 821
rect 1138 606 1172 821
rect 1354 606 1388 821
rect 1570 606 1604 821
rect 1786 606 1820 821
rect 2002 606 2036 821
rect 2218 606 2252 821
rect 2434 606 2468 821
rect 2650 606 2684 821
rect 2866 606 2900 821
rect 3082 606 3116 821
rect 3298 606 3332 821
rect 3514 606 3548 821
rect 3730 606 3764 821
rect 3946 606 3980 821
rect 4162 606 4196 821
rect 4374 606 4408 821
rect 4478 763 4512 821
rect 4478 713 4512 729
rect 48 386 114 402
rect 48 352 64 386
rect 98 352 114 386
rect 48 336 114 352
rect 2218 386 2252 572
rect 2218 352 2269 386
rect 2218 167 2252 352
rect 4478 109 4512 125
rect 62 17 96 67
rect 274 17 308 67
rect 490 17 524 67
rect 706 17 740 67
rect 922 17 956 67
rect 1138 17 1172 67
rect 1354 17 1388 67
rect 1570 17 1604 67
rect 1786 17 1820 67
rect 2002 17 2036 67
rect 2218 17 2252 67
rect 2434 17 2468 67
rect 2650 17 2684 67
rect 2866 17 2900 67
rect 3082 17 3116 67
rect 3298 17 3332 67
rect 3514 17 3548 67
rect 3730 17 3764 67
rect 3946 17 3980 67
rect 4162 17 4196 67
rect 4374 17 4408 67
rect 4478 17 4512 75
rect 0 -17 4580 17
use contact_12  contact_12_0
timestamp 1644951705
transform 1 0 48 0 1 336
box 0 0 1 1
use contact_11  contact_11_0
timestamp 1644951705
transform 1 0 4470 0 1 51
box 0 0 1 1
use contact_10  contact_10_0
timestamp 1644951705
transform 1 0 4470 0 1 705
box 0 0 1 1
use nmos_m40_w0_495_sli_dli_da_p  nmos_m40_w0_495_sli_dli_da_p_0
timestamp 1644951705
transform 1 0 54 0 1 51
box 0 -26 4362 155
use pmos_m40_w1_480_sli_dli_da_p  pmos_m40_w1_480_sli_dli_da_p_0
timestamp 1644951705
transform 1 0 54 0 1 491
box -59 -56 4421 350
<< labels >>
rlabel locali s 81 369 81 369 4 A
rlabel locali s 2252 369 2252 369 4 Z
rlabel locali s 2290 0 2290 0 4 gnd
rlabel locali s 2290 838 2290 838 4 vdd
<< properties >>
string FIXED_BBOX 0 0 4580 838
string GDS_FILE sram_0rw2r1w_16_128_sky130A.gds
string GDS_END 2002584
string GDS_START 1998532
<< end >>
