magic
tech sky130A
magscale 1 2
timestamp 1643593061
<< checkpaint >>
rect -1296 -1277 2528 2155
<< nwell >>
rect -36 402 1268 895
<< locali >>
rect 0 821 1232 855
rect 48 340 114 406
rect 613 356 647 390
rect 0 -17 1232 17
use pinv_9  pinv_9_0
timestamp 1643593061
transform 1 0 0 0 1 0
box -36 -17 1268 895
<< labels >>
rlabel locali s 630 373 630 373 4 Z
rlabel locali s 81 373 81 373 4 A
rlabel locali s 616 0 616 0 4 gnd
rlabel locali s 616 838 616 838 4 vdd
<< properties >>
string FIXED_BBOX 0 0 1232 838
string GDS_FILE sram_0rw2r1w_2_16_sky130A.gds
string GDS_END 560084
string GDS_START 559240
<< end >>
