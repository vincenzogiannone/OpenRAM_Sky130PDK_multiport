* NGSPICE file created from sram_0rw2r1w_4_16_sky130A.ext - technology: sky130A

.subckt dff clk vdd gnd D Q
X0 net3 net2 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.35e+06u l=150000u
X1 gnd net7 a_922_96# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 vdd clk clkb vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.35e+06u l=150000u
X3 net3 net2 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 vdd net3 net4 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.35e+06u l=150000u
X5 gnd net3 a_474_96# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 gnd clk clkb gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_922_96# clkb net6 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_474_96# clk net2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 net4 clkb net2 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.35e+06u l=150000u
X10 net6 clk net3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 net2 clkb net1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 net7 net6 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.35e+06u l=150000u
X13 net8 clk net6 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.35e+06u l=150000u
X14 net2 clk net1 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.35e+06u l=150000u
X15 net1 D gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 vdd net7 net8 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.35e+06u l=150000u
X17 net1 D vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.35e+06u l=150000u
X18 net6 clkb net3 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.35e+06u l=150000u
X19 Q net7 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.35e+06u l=150000u
X20 net7 net6 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 Q net7 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt nmos_m4_w0_420_sli_dli_da_p S S_uq0 S_uq1 gnd D G
X0 D G S_uq1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 D G S gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 S G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 S_uq0 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt pmos_m4_w1_260_sli_dli_da_p w_n59_42# S S_uq0 S_uq1 gnd D G
X0 D G S w_n59_42# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.26e+06u l=150000u
X1 S G D w_n59_42# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.26e+06u l=150000u
X2 S_uq0 G D w_n59_42# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.26e+06u l=150000u
X3 D G S_uq1 w_n59_42# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.26e+06u l=150000u
.ends

.subckt pinv_1 Z gnd vdd A
Xnmos_m4_w0_420_sli_dli_da_p_0 gnd gnd gnd gnd Z A nmos_m4_w0_420_sli_dli_da_p
Xpmos_m4_w1_260_sli_dli_da_p_0 vdd vdd vdd vdd gnd Z A pmos_m4_w1_260_sli_dli_da_p
.ends

.subckt nmos_m2_w0_420_sli_dli_da_p S S_uq0 gnd D G
X0 D G S gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 S_uq0 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt pmos_m2_w1_260_sli_dli_da_p w_n59_42# S S_uq0 gnd D G
X0 S_uq0 G D w_n59_42# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.26e+06u l=150000u
X1 D G S w_n59_42# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.26e+06u l=150000u
.ends

.subckt pinv_0 Z gnd vdd A
Xnmos_m2_w0_420_sli_dli_da_p_0 gnd gnd gnd Z A nmos_m2_w0_420_sli_dli_da_p
Xpmos_m2_w1_260_sli_dli_da_p_0 vdd vdd vdd gnd Z A pmos_m2_w1_260_sli_dli_da_p
.ends

.subckt dff_buf_0 pinv_1_0/vdd clk Q D Qb gnd vdd
Xdff_0 clk vdd gnd D dff_0/Q dff
Xpinv_1_0 Q gnd pinv_1_0/vdd Qb pinv_1
Xpinv_0_0 Qb gnd pinv_1_0/vdd dff_0/Q pinv_0
.ends

.subckt dff_buf_array vdd dout_0 dout_1 din_1 dout_bar_0 dout_bar_1 din_0
Xdff_buf_0_1 dff_buf_0_1/pinv_1_0/vdd vdd dout_0 din_0 dout_bar_0 vdd vdd dff_buf_0
Xdff_buf_0_0 dff_buf_0_1/pinv_1_0/vdd vdd dout_1 din_1 dout_bar_1 vdd vdd dff_buf_0
.ends

.subckt nmos_m1_w0_420_sli_dli_da_p S gnd D G
X0 D G S gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt pmos_m1_w1_260_sli_dli_da_p w_n59_42# S gnd D G
X0 D G S w_n59_42# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.26e+06u l=150000u
.ends

.subckt pinv_3 A Z gnd vdd
Xnmos_m1_w0_420_sli_dli_da_p_0 gnd gnd Z A nmos_m1_w0_420_sli_dli_da_p
Xpmos_m1_w1_260_sli_dli_da_p_0 vdd vdd gnd Z A pmos_m1_w1_260_sli_dli_da_p
.ends

.subckt nmos_m5_w0_420_sli_dli_da_p S S_uq0 S_uq1 gnd D G
X0 D G S_uq1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 D G S gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 S G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 D G S_uq0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 S_uq0 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt pmos_m5_w1_260_sli_dli_da_p w_n59_42# S S_uq0 S_uq1 gnd D G
X0 D G S w_n59_42# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.26e+06u l=150000u
X1 S G D w_n59_42# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.26e+06u l=150000u
X2 D G S_uq0 w_n59_42# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.26e+06u l=150000u
X3 S_uq0 G D w_n59_42# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.26e+06u l=150000u
X4 D G S_uq1 w_n59_42# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.26e+06u l=150000u
.ends

.subckt pinv_9 Z gnd vdd A
Xnmos_m5_w0_420_sli_dli_da_p_0 gnd gnd gnd gnd Z A nmos_m5_w0_420_sli_dli_da_p
Xpmos_m5_w1_260_sli_dli_da_p_0 vdd vdd vdd vdd gnd Z A pmos_m5_w1_260_sli_dli_da_p
.ends

.subckt pinv_5 Z A gnd vdd
Xnmos_m1_w0_420_sli_dli_da_p_0 gnd gnd Z A nmos_m1_w0_420_sli_dli_da_p
Xpmos_m1_w1_260_sli_dli_da_p_0 vdd vdd gnd Z A pmos_m1_w1_260_sli_dli_da_p
.ends

.subckt pinv_6 vdd Z gnd A
Xnmos_m2_w0_420_sli_dli_da_p_0 gnd gnd gnd Z A nmos_m2_w0_420_sli_dli_da_p
Xpmos_m2_w1_260_sli_dli_da_p_0 vdd vdd vdd gnd Z A pmos_m2_w1_260_sli_dli_da_p
.ends

.subckt pdriver_1 vdd Z gnd A
Xpinv_9_0 Z gnd vdd pinv_9_0/A pinv_9
Xpinv_5_0 pinv_6_0/A pinv_5_1/Z gnd vdd pinv_5
Xpinv_5_1 pinv_5_1/Z A gnd vdd pinv_5
Xpinv_6_0 vdd pinv_9_0/A gnd pinv_6_0/A pinv_6
.ends

.subckt pmos_m1_w1_260_sli_dli w_n59_42# S gnd D G
X0 D G S w_n59_42# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.26e+06u l=150000u
.ends

.subckt nmos_m1_w0_840_sli_dactive S gnd G a_90_0#
X0 a_90_0# G S gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
.ends

.subckt nmos_m1_w0_840_sactive_dli a_0_0# gnd D G
X0 D G a_0_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
.ends

.subckt pnand2_0 w_n36_402# Z gnd A vdd B
Xpmos_m1_w1_260_sli_dli_0 w_n36_402# Z gnd vdd B pmos_m1_w1_260_sli_dli
Xpmos_m1_w1_260_sli_dli_1 w_n36_402# vdd gnd Z A pmos_m1_w1_260_sli_dli
Xnmos_m1_w0_840_sli_dactive_0 gnd gnd A nmos_m1_w0_840_sactive_dli_0/a_0_0# nmos_m1_w0_840_sli_dactive
Xnmos_m1_w0_840_sactive_dli_0 nmos_m1_w0_840_sactive_dli_0/a_0_0# gnd Z B nmos_m1_w0_840_sactive_dli
.ends

.subckt pmos_m11_w1_375_sli_dli_da_p S S_uq0 S_uq1 S_uq3 S_uq2 S_uq4 gnd w_n59_53#
+ D G
X0 D G S_uq3 w_n59_53# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=150000u
X1 D G S w_n59_53# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=150000u
X2 S_uq3 G D w_n59_53# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=150000u
X3 D G S_uq0 w_n59_53# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=150000u
X4 S G D w_n59_53# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=150000u
X5 S_uq0 G D w_n59_53# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=150000u
X6 D G S_uq2 w_n59_53# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=150000u
X7 D G S_uq1 w_n59_53# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=150000u
X8 S_uq2 G D w_n59_53# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=150000u
X9 S_uq1 G D w_n59_53# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=150000u
X10 D G S_uq4 w_n59_53# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=150000u
.ends

.subckt nmos_m11_w0_460_sli_dli_da_p S S_uq0 S_uq1 S_uq3 S_uq2 S_uq4 gnd D G
X0 S_uq1 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=460000u l=150000u
X1 D G S_uq4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=460000u l=150000u
X2 D G S_uq3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=460000u l=150000u
X3 D G S gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=460000u l=150000u
X4 S_uq3 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=460000u l=150000u
X5 D G S_uq0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=460000u l=150000u
X6 S G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=460000u l=150000u
X7 S_uq0 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=460000u l=150000u
X8 D G S_uq2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=460000u l=150000u
X9 D G S_uq1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=460000u l=150000u
X10 S_uq2 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=460000u l=150000u
.ends

.subckt pinv_2 gnd vdd Z A
Xpmos_m11_w1_375_sli_dli_da_p_0 vdd vdd vdd vdd vdd vdd gnd vdd Z A pmos_m11_w1_375_sli_dli_da_p
Xnmos_m11_w0_460_sli_dli_da_p_0 gnd gnd gnd gnd gnd gnd gnd Z A nmos_m11_w0_460_sli_dli_da_p
.ends

.subckt pdriver vdd gnd Z A
Xpinv_2_0 gnd vdd Z A pinv_2
.ends

.subckt pand2 vdd gnd Z A B
Xpnand2_0_0 vdd pdriver_0/A gnd A vdd B pnand2_0
Xpdriver_0 vdd gnd Z pdriver_0/A pdriver
.ends

.subckt pnand2_1 Z gnd vdd A
Xpmos_m1_w1_260_sli_dli_0 vdd Z gnd vdd B pmos_m1_w1_260_sli_dli
Xpmos_m1_w1_260_sli_dli_1 vdd vdd gnd Z A pmos_m1_w1_260_sli_dli
Xnmos_m1_w0_840_sli_dactive_0 gnd gnd A nmos_m1_w0_840_sactive_dli_0/a_0_0# nmos_m1_w0_840_sli_dactive
Xnmos_m1_w0_840_sactive_dli_0 nmos_m1_w0_840_sactive_dli_0/a_0_0# gnd Z B nmos_m1_w0_840_sactive_dli
.ends

.subckt pdriver_2 Z gnd vdd A
Xpinv_5_0 Z pinv_5_1/Z gnd vdd pinv_5
Xpinv_5_1 pinv_5_1/Z A gnd vdd pinv_5
.ends

.subckt pmos_m6_w1_260_sli_dli_da_p w_n59_42# S S_uq0 S_uq1 S_uq2 gnd D G
X0 D G S_uq1 w_n59_42# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.26e+06u l=150000u
X1 S_uq1 G D w_n59_42# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.26e+06u l=150000u
X2 D G S w_n59_42# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.26e+06u l=150000u
X3 S G D w_n59_42# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.26e+06u l=150000u
X4 S_uq0 G D w_n59_42# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.26e+06u l=150000u
X5 D G S_uq2 w_n59_42# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.26e+06u l=150000u
.ends

.subckt nmos_m6_w0_420_sli_dli_da_p S S_uq0 S_uq1 S_uq2 gnd D G
X0 S_uq0 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 D G S_uq2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 D G S_uq1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 S_uq1 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 D G S gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 S G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt pinv_7 Z gnd vdd A
Xpmos_m6_w1_260_sli_dli_da_p_0 vdd vdd vdd vdd vdd gnd Z A pmos_m6_w1_260_sli_dli_da_p
Xnmos_m6_w0_420_sli_dli_da_p_0 gnd gnd gnd gnd gnd Z A nmos_m6_w0_420_sli_dli_da_p
.ends

.subckt nmos_m16_w0_470_sli_dli_da_p S S_uq0 S_uq1 S_uq3 S_uq2 S_uq4 S_uq5 S_uq6 S_uq7
+ gnd D G
X0 S_uq4 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=470000u l=150000u
X1 D G S_uq7 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=470000u l=150000u
X2 S_uq1 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=470000u l=150000u
X3 S_uq0 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=470000u l=150000u
X4 D G S_uq6 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=470000u l=150000u
X5 D G S_uq3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=470000u l=150000u
X6 S_uq6 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=470000u l=150000u
X7 D G S_uq2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=470000u l=150000u
X8 D G S gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=470000u l=150000u
X9 S_uq3 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=470000u l=150000u
X10 S_uq2 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=470000u l=150000u
X11 S G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=470000u l=150000u
X12 D G S_uq5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=470000u l=150000u
X13 D G S_uq4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=470000u l=150000u
X14 D G S_uq1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=470000u l=150000u
X15 S_uq5 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=470000u l=150000u
.ends

.subckt pmos_m16_w1_420_sli_dli_da_p S S_uq0 S_uq1 S_uq3 S_uq2 S_uq4 S_uq5 S_uq6 S_uq7
+ w_n59_58# gnd D G
X0 D G S_uq6 w_n59_58# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.42e+06u l=150000u
X1 S_uq0 G D w_n59_58# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.42e+06u l=150000u
X2 D G S_uq3 w_n59_58# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.42e+06u l=150000u
X3 S_uq6 G D w_n59_58# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.42e+06u l=150000u
X4 D G S_uq2 w_n59_58# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.42e+06u l=150000u
X5 D G S w_n59_58# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.42e+06u l=150000u
X6 S_uq3 G D w_n59_58# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.42e+06u l=150000u
X7 S G D w_n59_58# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.42e+06u l=150000u
X8 S_uq2 G D w_n59_58# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.42e+06u l=150000u
X9 D G S_uq5 w_n59_58# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.42e+06u l=150000u
X10 D G S_uq4 w_n59_58# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.42e+06u l=150000u
X11 D G S_uq1 w_n59_58# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.42e+06u l=150000u
X12 S_uq5 G D w_n59_58# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.42e+06u l=150000u
X13 S_uq4 G D w_n59_58# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.42e+06u l=150000u
X14 D G S_uq7 w_n59_58# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.42e+06u l=150000u
X15 S_uq1 G D w_n59_58# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.42e+06u l=150000u
.ends

.subckt pinv_8 Z gnd vdd A
Xnmos_m16_w0_470_sli_dli_da_p_0 gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd Z A nmos_m16_w0_470_sli_dli_da_p
Xpmos_m16_w1_420_sli_dli_da_p_0 vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd gnd Z A pmos_m16_w1_420_sli_dli_da_p
.ends

.subckt pdriver_0 A Z gnd vdd
Xpinv_7_0 pinv_8_0/A gnd vdd pinv_7_0/A pinv_7
Xpinv_5_0 pinv_6_0/A A gnd vdd pinv_5
Xpinv_8_0 Z gnd vdd pinv_8_0/A pinv_8
Xpinv_6_0 vdd pinv_7_0/A gnd pinv_6_0/A pinv_6
.ends

.subckt control_logic_multiport p_en_bar clk web vdd csb wl_en w_en
Xdff_buf_array_0 vdd dff_buf_array_0/dout_0 dff_buf_array_0/dout_1 csb pand2_0/A pand2_2/B
+ web dff_buf_array
Xpinv_3_0 vdd pand2_2/A vdd pand2_2/vdd pinv_3
Xpdriver_1_0 pnand2_1_0/vdd wl_en vdd pand2_2/Z pdriver_1
Xpand2_0 pand2_1/vdd vdd w_en pand2_0/A pand2_2/Z pand2
Xpand2_1 pand2_1/vdd vdd pand2_1/Z vdd pand2_2/B pand2
Xpnand2_1_0 pnand2_1_0/Z vdd pnand2_1_0/vdd pand2_1/Z pnand2_1
Xpdriver_2_0 p_en_bar vdd pnand2_1_0/vdd pnand2_1_0/Z pdriver_2
Xpand2_2 pand2_2/vdd vdd pand2_2/Z pand2_2/A pand2_2/B pand2
Xpdriver_0_0 clk vdd vdd pand2_2/vdd pdriver_0
.ends

.subckt data_dff vdd clk gnd din_0 din_1 din_2 din_3
Xdff_0 clk vdd gnd din_3 dout_3 dff
Xdff_1 clk vdd gnd din_2 dout_2 dff
Xdff_2 clk vdd gnd din_1 dout_1 dff
Xdff_3 clk vdd gnd din_0 dout_0 dff
.ends

.subckt row_addr_dff vdd_uq0 vdd_uq1 vdd_uq2 clk dout_0 dout_1 dout_3 dout_2 gnd dout_4
+ dout_5 vdd din_0 din_1 din_2 din_3 din_4 din_5
Xdff_0 clk vdd_uq2 gnd din_7 dout_7 dff
Xdff_1 clk vdd_uq2 gnd din_6 dout_6 dff
Xdff_2 clk vdd_uq1 gnd din_5 dout_5 dff
Xdff_3 clk vdd_uq1 gnd din_4 dout_4 dff
Xdff_4 clk vdd gnd din_3 dout_3 dff
Xdff_5 clk vdd gnd din_2 dout_2 dff
Xdff_6 clk vdd_uq0 gnd din_1 dout_1 dff
Xdff_7 clk vdd_uq0 gnd din_0 dout_0 dff
.ends

.subckt sense_amp_multiport vdd gnd rbl dout
X0 dout rbl gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 dout rbl vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.7e+06u l=150000u
.ends

.subckt sense_amp_array vdd_uq2 vdd_uq4 vdd_uq6 gnd data_0 data_1 data_2 data_3 vdd
Xsense_amp_multiport_0 vdd gnd rbl_7 data_7 sense_amp_multiport
Xsense_amp_multiport_1 vdd gnd rbl_6 data_6 sense_amp_multiport
Xsense_amp_multiport_2 vdd_uq2 gnd rbl_5 data_5 sense_amp_multiport
Xsense_amp_multiport_3 vdd_uq2 gnd rbl_4 data_4 sense_amp_multiport
Xsense_amp_multiport_4 vdd_uq4 gnd rbl_3 data_3 sense_amp_multiport
Xsense_amp_multiport_5 vdd_uq4 gnd rbl_2 data_2 sense_amp_multiport
Xsense_amp_multiport_6 vdd_uq6 gnd rbl_1 data_1 sense_amp_multiport
Xsense_amp_multiport_7 vdd_uq6 gnd rbl_0 data_0 sense_amp_multiport
.ends

.subckt write_driver_multiport din vdd gnd en wbl
X0 net2 net1 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.35e+06u l=150000u
X1 net1 din gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 wbl en a_478_138# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 gnd en enb gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_478_138# net1 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 net1 din vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.35e+06u l=150000u
X6 wbl enb net2 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.35e+06u l=150000u
X7 vdd en enb vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.35e+06u l=150000u
.ends

.subckt write_driver_array vdd_uq0 vdd_uq1 vdd_uq2 en wbl0_0 gnd din_2 vdd din_0 din_1
+ din_3
Xwrite_driver_multiport_0 din_3 vdd_uq0 gnd en wbl0_3 write_driver_multiport
Xwrite_driver_multiport_1 din_2 vdd gnd en wbl0_2 write_driver_multiport
Xwrite_driver_multiport_2 din_1 vdd_uq1 gnd en wbl0_1 write_driver_multiport
Xwrite_driver_multiport_3 din_0 vdd_uq2 gnd en wbl0_0 write_driver_multiport
.ends

.subckt precharge_multiport_0 en_bar rbl1 gnd rbl0 vdd
Xpmos_m1_w1_260_sli_dli_0 vdd vdd gnd rbl1 en_bar pmos_m1_w1_260_sli_dli
Xpmos_m1_w1_260_sli_dli_1 vdd rbl0 gnd vdd en_bar pmos_m1_w1_260_sli_dli
Xpmos_m1_w1_260_sli_dli_2 vdd rbl0 gnd rbl1 en_bar pmos_m1_w1_260_sli_dli
.ends

.subckt precharge_array_multiport rbl0_0 rbl0_1 rbl0_2 rbl0_3 vdd en_bar rbl1_4 rbl1_0
+ rbl1_1 rbl1_2 rbl1_3 gnd
Xprecharge_multiport_0_1 en_bar rbl1_3 gnd rbl0_3 vdd precharge_multiport_0
Xprecharge_multiport_0_2 en_bar rbl1_2 gnd rbl0_2 vdd precharge_multiport_0
Xprecharge_multiport_0_3 en_bar rbl1_1 gnd rbl0_1 vdd precharge_multiport_0
Xprecharge_multiport_0_4 en_bar rbl1_0 gnd rbl0_0 vdd precharge_multiport_0
Xprecharge_multiport_0_0 en_bar rbl1_4 gnd rbl0_4 vdd precharge_multiport_0
.ends

.subckt port_data p_en_bar vdd vdd_uq5 vdd_uq7 dout1_0 vdd_uq9 dout1_1 dout1_2 dout1_3
+ w_en precharge_array_multiport_0/rbl1_4 gnd vdd_uq11 vdd_uq12 vdd_uq13 vdd_uq14
+ vdd_uq15 din0_0 din0_1 din0_2 din0_3
Xsense_amp_array_0 vdd_uq7 vdd_uq9 vdd_uq11 gnd dout1_0 dout1_1 dout1_2 dout1_3 vdd_uq5
+ sense_amp_array
Xwrite_driver_array_0 vdd_uq12 vdd_uq14 vdd_uq15 w_en wbl0_0 gnd din0_2 vdd_uq13 din0_0
+ din0_1 din0_3 write_driver_array
Xprecharge_array_multiport_0 rbl0_0 rbl0_1 rbl0_2 rbl0_3 vdd p_en_bar precharge_array_multiport_0/rbl1_4
+ rbl1_0 rbl1_1 rbl1_2 rbl1_3 gnd precharge_array_multiport
.ends

.subckt pinv Z A vdd gnd
Xnmos_m1_w0_420_sli_dli_da_p_0 gnd gnd Z A nmos_m1_w0_420_sli_dli_da_p
Xpmos_m1_w1_260_sli_dli_da_p_0 vdd vdd gnd Z A pmos_m1_w1_260_sli_dli_da_p
.ends

.subckt pnand2 Z gnd vdd A B
Xpmos_m1_w1_260_sli_dli_0 vdd Z gnd vdd B pmos_m1_w1_260_sli_dli
Xpmos_m1_w1_260_sli_dli_1 vdd vdd gnd Z A pmos_m1_w1_260_sli_dli
Xnmos_m1_w0_840_sli_dactive_0 gnd gnd A nmos_m1_w0_840_sactive_dli_0/a_0_0# nmos_m1_w0_840_sli_dactive
Xnmos_m1_w0_840_sactive_dli_0 nmos_m1_w0_840_sactive_dli_0/a_0_0# gnd Z B nmos_m1_w0_840_sactive_dli
.ends

.subckt and2_dec Z gnd vdd A B
Xpinv_0 Z pinv_0/A vdd gnd pinv
Xpnand2_0 pinv_0/A gnd vdd A B pnand2
.ends

.subckt hierarchical_predecode2x4 in_1 vdd_uq0 gnd out_0 out_1 out_2 out_3 in_0 vdd
Xand2_dec_0 out_3 gnd vdd in_0 in_1 and2_dec
Xand2_dec_1 out_2 gnd vdd pinv_1/Z in_1 and2_dec
Xpinv_0 pinv_0/Z in_1 vdd_uq0 gnd pinv
Xand2_dec_2 out_1 gnd vdd_uq0 in_0 pinv_0/Z and2_dec
Xpinv_1 pinv_1/Z in_0 vdd_uq0 gnd pinv
Xand2_dec_3 out_0 gnd vdd_uq0 pinv_1/Z pinv_0/Z and2_dec
.ends

.subckt dec_cell3_2r1w A0 B0 C0 A1 B1 C1 A2 B2 C2 OUT2 vdd gnd OUT0 OUT1
X0 vdd A2 net9 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_124_132# A0 net3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 net6 A1 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 OUT2 net9 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.35e+06u l=150000u
X4 OUT2 net9 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 vdd C0 net3 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 net6 C1 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 vdd C2 net9 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 OUT0 net6 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.35e+06u l=150000u
X9 a_220_132# B0 a_124_132# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_412_132# A1 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 gnd net3 OUT1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 OUT0 net6 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 gnd C0 a_220_132# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_508_132# B1 a_412_132# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 net6 C1 a_508_132# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 vdd B1 net6 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 vdd A0 net3 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 net9 B2 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 vdd net3 OUT1 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.35e+06u l=150000u
X20 a_808_132# A2 net9 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 a_904_132# B2 a_808_132# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 gnd C2 a_904_132# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 net3 B0 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt hierarchical_decoder addr_0 decode0_6 decode2_9 decode1_10 gnd addr_1 vdd_uq4
+ decode0_7 decode1_11 vdd addr_2 vdd_uq2 decode0_8 decode1_12 addr_3 decode0_9 decode1_13
+ addr_4 decode1_14 addr_5 decode1_15 vdd_uq6 vdd_uq8 vdd_uq9 decode1_0 decode1_1
+ decode2_10 decode1_2 decode1_3 decode2_11 decode2_12 decode1_4 decode1_5 decode2_13
+ decode2_14 decode1_6 decode2_15 decode1_7 decode1_8 decode1_9 decode0_10 decode0_11
+ vdd_uq11 decode0_12 vdd_uq12 decode2_0 decode0_13 vdd_uq13 decode2_1 decode0_14
+ vdd_uq14 decode0_15 decode2_2 vdd_uq15 decode0_0 decode2_3 vdd_uq16 decode2_4 decode0_1
+ vdd_uq17 decode0_2 decode2_5 vdd_uq18 decode2_6 decode0_3 decode0_4 decode2_7 decode2_8
+ decode0_5
Xhierarchical_predecode2x4_0 addr_5 vdd_uq8 gnd predecode_8 predecode_9 predecode_10
+ predecode_11 addr_4 vdd_uq9 hierarchical_predecode2x4
Xhierarchical_predecode2x4_1 addr_3 vdd_uq4 gnd predecode_4 predecode_5 predecode_6
+ predecode_7 addr_2 vdd_uq6 hierarchical_predecode2x4
Xhierarchical_predecode2x4_2 addr_1 vdd gnd predecode_0 predecode_1 predecode_2 predecode_3
+ addr_0 vdd_uq2 hierarchical_predecode2x4
Xdec_cell3_2r1w_0 predecode_0 predecode_7 predecode_10 predecode_1 predecode_7 predecode_10
+ predecode_2 predecode_7 predecode_10 decode2_15 vdd_uq18 gnd decode0_15 decode1_15
+ dec_cell3_2r1w
Xdec_cell3_2r1w_1 predecode_1 predecode_6 predecode_10 predecode_2 predecode_6 predecode_10
+ predecode_3 predecode_6 predecode_10 decode2_14 vdd_uq18 gnd decode0_14 decode1_14
+ dec_cell3_2r1w
Xdec_cell3_2r1w_2 predecode_2 predecode_5 predecode_10 predecode_3 predecode_5 predecode_10
+ predecode_0 predecode_6 predecode_10 decode2_13 vdd_uq17 gnd decode0_13 decode1_13
+ dec_cell3_2r1w
Xdec_cell3_2r1w_10 predecode_2 predecode_7 predecode_8 predecode_3 predecode_7 predecode_8
+ predecode_0 predecode_4 predecode_9 decode2_5 vdd_uq13 gnd decode0_5 decode1_5 dec_cell3_2r1w
Xdec_cell3_2r1w_3 predecode_3 predecode_4 predecode_10 predecode_0 predecode_5 predecode_10
+ predecode_1 predecode_5 predecode_10 decode2_12 vdd_uq17 gnd decode0_12 decode1_12
+ dec_cell3_2r1w
Xdec_cell3_2r1w_11 predecode_3 predecode_6 predecode_8 predecode_0 predecode_7 predecode_8
+ predecode_1 predecode_7 predecode_8 decode2_4 vdd_uq13 gnd decode0_4 decode1_4 dec_cell3_2r1w
Xdec_cell3_2r1w_4 predecode_0 predecode_4 predecode_10 predecode_1 predecode_4 predecode_10
+ predecode_2 predecode_4 predecode_10 decode2_11 vdd_uq16 gnd decode0_11 decode1_11
+ dec_cell3_2r1w
Xdec_cell3_2r1w_12 predecode_0 predecode_6 predecode_8 predecode_1 predecode_6 predecode_8
+ predecode_2 predecode_6 predecode_8 decode2_3 vdd_uq12 gnd decode0_3 decode1_3 dec_cell3_2r1w
Xdec_cell3_2r1w_13 predecode_1 predecode_5 predecode_8 predecode_2 predecode_5 predecode_8
+ predecode_3 predecode_5 predecode_8 decode2_2 vdd_uq12 gnd decode0_2 decode1_2 dec_cell3_2r1w
Xdec_cell3_2r1w_5 predecode_1 predecode_7 predecode_9 predecode_2 predecode_7 predecode_9
+ predecode_3 predecode_7 predecode_9 decode2_10 vdd_uq16 gnd decode0_10 decode1_10
+ dec_cell3_2r1w
Xdec_cell3_2r1w_6 predecode_2 predecode_6 predecode_9 predecode_3 predecode_6 predecode_9
+ predecode_0 predecode_7 predecode_9 decode2_9 vdd_uq15 gnd decode0_9 decode1_9 dec_cell3_2r1w
Xdec_cell3_2r1w_14 predecode_2 predecode_4 predecode_8 predecode_3 predecode_4 predecode_8
+ predecode_0 predecode_5 predecode_8 decode2_1 vdd_uq11 gnd decode0_1 decode1_1 dec_cell3_2r1w
Xdec_cell3_2r1w_15 dec_cell3_2r1w_15/A0 dec_cell3_2r1w_15/B0 dec_cell3_2r1w_15/C0
+ predecode_0 predecode_4 predecode_8 predecode_1 predecode_4 predecode_8 decode2_0
+ vdd_uq11 gnd decode0_0 decode1_0 dec_cell3_2r1w
Xdec_cell3_2r1w_7 predecode_3 predecode_5 predecode_9 predecode_0 predecode_6 predecode_9
+ predecode_1 predecode_6 predecode_9 decode2_8 vdd_uq15 gnd decode0_8 decode1_8 dec_cell3_2r1w
Xdec_cell3_2r1w_8 predecode_0 predecode_5 predecode_9 predecode_1 predecode_5 predecode_9
+ predecode_2 predecode_5 predecode_9 decode2_7 vdd_uq14 gnd decode0_7 decode1_7 dec_cell3_2r1w
Xdec_cell3_2r1w_9 predecode_1 predecode_4 predecode_9 predecode_2 predecode_4 predecode_9
+ predecode_3 predecode_4 predecode_9 decode2_6 vdd_uq14 gnd decode0_6 decode1_6 dec_cell3_2r1w
.ends

.subckt wordline_driver_cell A0 vdd gnd wl_en A1 A2 rwl0 wwl0 rwl1
X0 gnd wl_en a_124_308# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X1 net4 wl_en a_316_308# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X2 a_316_308# A1 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X3 vdd wl_en net4 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 vdd net4 rwl0 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.35e+06u l=150000u
X5 a_616_308# A2 net6 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X6 gnd wl_en a_616_308# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X7 wwl0 net6 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 net4 A1 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 vdd wl_en net6 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_124_308# A0 net2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X11 net6 A2 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 wwl0 net6 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.35e+06u l=150000u
X13 gnd net4 rwl0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 net2 A0 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 rwl1 net2 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 vdd wl_en net2 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 rwl1 net2 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.35e+06u l=150000u
.ends

.subckt wordline_driver_array wl_en wwl0_0 rwl1_0 rwl1_11 rwl1_1 wwl0_1 rwl1_12 vdd_uq0
+ wwl0_2 rwl1_2 vdd_uq1 rwl1_13 rwl1_3 wwl0_3 vdd_uq2 in2_10 rwl1_14 in2_11 wwl0_4
+ rwl1_4 vdd_uq3 rwl1_15 rwl1_5 wwl0_5 in2_12 vdd_uq4 in1_0 in2_13 vdd_uq5 wwl0_6
+ rwl1_6 in1_1 rwl1_7 vdd_uq6 in2_14 wwl0_7 in1_2 in2_15 wwl0_8 rwl1_8 in1_3 rwl1_9
+ wwl0_9 in1_4 in1_5 in1_6 in1_7 in1_8 in1_9 in0_10 in0_11 in0_12 wwl0_10 gnd in0_13
+ wwl0_11 in0_14 wwl0_12 in0_15 rwl0_0 wwl0_13 wwl0_14 rwl0_1 rwl0_2 wwl0_15 in2_0
+ rwl0_3 in2_1 rwl0_10 rwl0_4 in2_2 rwl0_11 rwl0_5 in0_0 in2_3 rwl0_12 in2_4 rwl0_6
+ in0_1 rwl0_13 rwl0_7 in2_5 in1_10 rwl0_14 in0_2 vdd in2_6 rwl0_8 in1_11 in0_3 rwl0_15
+ rwl0_9 in1_12 in2_7 in0_4 in1_13 in0_5 in2_8 in1_14 in2_9 in0_6 in1_15 in0_7 in0_8
+ in0_9 rwl1_10
Xwordline_driver_cell_0 in0_15 vdd_uq6 gnd wl_en in1_15 in2_15 rwl0_15 wwl0_15 rwl1_15
+ wordline_driver_cell
Xwordline_driver_cell_1 in0_14 vdd_uq6 gnd wl_en in1_14 in2_14 rwl0_14 wwl0_14 rwl1_14
+ wordline_driver_cell
Xwordline_driver_cell_2 in0_13 vdd_uq5 gnd wl_en in1_13 in2_13 rwl0_13 wwl0_13 rwl1_13
+ wordline_driver_cell
Xwordline_driver_cell_3 in0_12 vdd_uq5 gnd wl_en in1_12 in2_12 rwl0_12 wwl0_12 rwl1_12
+ wordline_driver_cell
Xwordline_driver_cell_4 in0_11 vdd_uq4 gnd wl_en in1_11 in2_11 rwl0_11 wwl0_11 rwl1_11
+ wordline_driver_cell
Xwordline_driver_cell_5 in0_10 vdd_uq4 gnd wl_en in1_10 in2_10 rwl0_10 wwl0_10 rwl1_10
+ wordline_driver_cell
Xwordline_driver_cell_6 in0_9 vdd_uq3 gnd wl_en in1_9 in2_9 rwl0_9 wwl0_9 rwl1_9 wordline_driver_cell
Xwordline_driver_cell_7 in0_8 vdd_uq3 gnd wl_en in1_8 in2_8 rwl0_8 wwl0_8 rwl1_8 wordline_driver_cell
Xwordline_driver_cell_10 in0_5 vdd_uq1 gnd wl_en in1_5 in2_5 rwl0_5 wwl0_5 rwl1_5
+ wordline_driver_cell
Xwordline_driver_cell_8 in0_7 vdd_uq2 gnd wl_en in1_7 in2_7 rwl0_7 wwl0_7 rwl1_7 wordline_driver_cell
Xwordline_driver_cell_11 in0_4 vdd_uq1 gnd wl_en in1_4 in2_4 rwl0_4 wwl0_4 rwl1_4
+ wordline_driver_cell
Xwordline_driver_cell_12 in0_3 vdd gnd wl_en in1_3 in2_3 rwl0_3 wwl0_3 rwl1_3 wordline_driver_cell
Xwordline_driver_cell_9 in0_6 vdd_uq2 gnd wl_en in1_6 in2_6 rwl0_6 wwl0_6 rwl1_6 wordline_driver_cell
Xwordline_driver_cell_13 in0_2 vdd gnd wl_en in1_2 in2_2 rwl0_2 wwl0_2 rwl1_2 wordline_driver_cell
Xwordline_driver_cell_14 in0_1 vdd_uq0 gnd wl_en in1_1 in2_1 rwl0_1 wwl0_1 rwl1_1
+ wordline_driver_cell
Xwordline_driver_cell_15 in0_0 vdd_uq0 gnd wl_en in1_0 in2_0 rwl0_0 wwl0_0 rwl1_0
+ wordline_driver_cell
.ends

.subckt port_address addr2 vdd_uq26 wwl0_0 rwl1_0 gnd rwl1_11 addr3 rwl1_1 wwl0_1
+ rwl1_12 vdd_uq0 addr4 vdd_uq9 vdd_uq2 wwl0_2 rwl1_2 rwl1_13 addr5 rwl1_3 wwl0_3
+ rwl1_14 rwl1_4 wwl0_4 vdd_uq3 rwl1_15 vdd_uq19 wwl0_5 rwl1_5 vdd_uq4 rwl1_6 wwl0_6
+ vdd_uq6 vdd rwl1_7 wwl0_7 vdd_uq22 rwl1_8 wwl0_8 vdd_uq7 vdd_uq8 wwl0_9 rwl1_9 vdd_uq10
+ vdd_uq14 vdd_uq18 vdd_uq20 vdd_uq24 wl_en vdd_uq12 wwl0_10 wwl0_11 wwl0_12 rwl0_0
+ wwl0_13 wwl0_14 rwl0_1 rwl0_2 wwl0_15 rwl0_3 rwl0_10 rwl0_4 rwl0_11 rwl0_5 rwl0_12
+ rwl0_6 rwl0_13 vdd_uq23 vdd_uq16 rwl0_7 rwl0_14 vdd_uq13 rwl0_8 rwl0_15 rwl0_9 addr0
+ addr1 vdd_uq17 rwl1_10
Xhierarchical_decoder_0 addr0 wordline_driver_array_0/in0_6 wordline_driver_array_0/in2_9
+ wordline_driver_array_0/in1_10 gnd addr1 vdd_uq12 wordline_driver_array_0/in0_7
+ wordline_driver_array_0/in1_11 vdd_uq2 addr2 vdd_uq6 wordline_driver_array_0/in0_8
+ wordline_driver_array_0/in1_12 addr3 wordline_driver_array_0/in0_9 wordline_driver_array_0/in1_13
+ addr4 wordline_driver_array_0/in1_14 addr5 wordline_driver_array_0/in1_15 vdd_uq16
+ vdd_uq22 vdd_uq26 wordline_driver_array_0/in1_0 wordline_driver_array_0/in1_1 wordline_driver_array_0/in2_10
+ wordline_driver_array_0/in1_2 wordline_driver_array_0/in1_3 wordline_driver_array_0/in2_11
+ wordline_driver_array_0/in2_12 wordline_driver_array_0/in1_4 wordline_driver_array_0/in1_5
+ wordline_driver_array_0/in2_13 wordline_driver_array_0/in2_14 wordline_driver_array_0/in1_6
+ wordline_driver_array_0/in2_15 wordline_driver_array_0/in1_7 wordline_driver_array_0/in1_8
+ wordline_driver_array_0/in1_9 wordline_driver_array_0/in0_10 wordline_driver_array_0/in0_11
+ vdd wordline_driver_array_0/in0_12 vdd_uq4 wordline_driver_array_0/in2_0 wordline_driver_array_0/in0_13
+ vdd_uq8 wordline_driver_array_0/in2_1 wordline_driver_array_0/in0_14 vdd_uq10 wordline_driver_array_0/in0_15
+ wordline_driver_array_0/in2_2 vdd_uq14 wordline_driver_array_0/in0_0 wordline_driver_array_0/in2_3
+ vdd_uq18 wordline_driver_array_0/in2_4 wordline_driver_array_0/in0_1 vdd_uq20 wordline_driver_array_0/in0_2
+ wordline_driver_array_0/in2_5 vdd_uq24 wordline_driver_array_0/in2_6 wordline_driver_array_0/in0_3
+ wordline_driver_array_0/in0_4 wordline_driver_array_0/in2_7 wordline_driver_array_0/in2_8
+ wordline_driver_array_0/in0_5 hierarchical_decoder
Xwordline_driver_array_0 wl_en wwl0_0 rwl1_0 rwl1_11 rwl1_1 wwl0_1 rwl1_12 vdd_uq0
+ wwl0_2 rwl1_2 vdd_uq7 rwl1_13 rwl1_3 wwl0_3 vdd_uq9 wordline_driver_array_0/in2_10
+ rwl1_14 wordline_driver_array_0/in2_11 wwl0_4 rwl1_4 vdd_uq13 rwl1_15 rwl1_5 wwl0_5
+ wordline_driver_array_0/in2_12 vdd_uq17 wordline_driver_array_0/in1_0 wordline_driver_array_0/in2_13
+ vdd_uq19 wwl0_6 rwl1_6 wordline_driver_array_0/in1_1 rwl1_7 vdd_uq23 wordline_driver_array_0/in2_14
+ wwl0_7 wordline_driver_array_0/in1_2 wordline_driver_array_0/in2_15 wwl0_8 rwl1_8
+ wordline_driver_array_0/in1_3 rwl1_9 wwl0_9 wordline_driver_array_0/in1_4 wordline_driver_array_0/in1_5
+ wordline_driver_array_0/in1_6 wordline_driver_array_0/in1_7 wordline_driver_array_0/in1_8
+ wordline_driver_array_0/in1_9 wordline_driver_array_0/in0_10 wordline_driver_array_0/in0_11
+ wordline_driver_array_0/in0_12 wwl0_10 gnd wordline_driver_array_0/in0_13 wwl0_11
+ wordline_driver_array_0/in0_14 wwl0_12 wordline_driver_array_0/in0_15 rwl0_0 wwl0_13
+ wwl0_14 rwl0_1 rwl0_2 wwl0_15 wordline_driver_array_0/in2_0 rwl0_3 wordline_driver_array_0/in2_1
+ rwl0_10 rwl0_4 wordline_driver_array_0/in2_2 rwl0_11 rwl0_5 wordline_driver_array_0/in0_0
+ wordline_driver_array_0/in2_3 rwl0_12 wordline_driver_array_0/in2_4 rwl0_6 wordline_driver_array_0/in0_1
+ rwl0_13 rwl0_7 wordline_driver_array_0/in2_5 wordline_driver_array_0/in1_10 rwl0_14
+ wordline_driver_array_0/in0_2 vdd_uq3 wordline_driver_array_0/in2_6 rwl0_8 wordline_driver_array_0/in1_11
+ wordline_driver_array_0/in0_3 rwl0_15 rwl0_9 wordline_driver_array_0/in1_12 wordline_driver_array_0/in2_7
+ wordline_driver_array_0/in0_4 wordline_driver_array_0/in1_13 wordline_driver_array_0/in0_5
+ wordline_driver_array_0/in2_8 wordline_driver_array_0/in1_14 wordline_driver_array_0/in2_9
+ wordline_driver_array_0/in0_6 wordline_driver_array_0/in1_15 wordline_driver_array_0/in0_7
+ wordline_driver_array_0/in0_8 wordline_driver_array_0/in0_9 rwl1_10 wordline_driver_array
.ends

.subckt cell_2r1w vdd gnd rbl0 rbl1 wbl0 wwl0 rwl1 rwl0
X0 q qbar vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X1 net2 q gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X2 gnd qbar q gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 wbl0 wwl0 q gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X4 net1 wwl0 qbar gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X5 rbl1 rwl1 net3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X6 vdd q qbar vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X7 rbl0 rwl0 net2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X8 gnd q net3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X9 net1 wbl0 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X10 qbar q gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 net1 wbl0 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt bitcell_array write_bl_0_3 read_bl_0_3 read_bl_0_1 read_bl_0_0 rwl_0_3 write_bl_0_1
+ rwl_1_14 read_bl_1_1 read_bl_1_3 read_bl_1_0 wwl_0_0 rwl_0_4 rwl_0_5 rwl_0_1 write_bl_0_0
+ rwl_0_6 wwl_0_10 rwl_1_1 read_bl_0_2 rwl_0_7 rwl_0_11 write_bl_0_2 wwl_0_11 rwl_0_14
+ wwl_0_15 rwl_1_11 rwl_0_8 wwl_0_12 rwl_0_9 wwl_0_13 rwl_0_10 wwl_0_14 rwl_1_8 rwl_0_12
+ read_bl_1_2 wwl_0_4 wwl_0_9 rwl_0_13 rwl_1_5 rwl_1_3 rwl_0_15 rwl_1_15 rwl_0_0 wwl_0_1
+ wwl_0_6 rwl_1_0 rwl_0_2 rwl_1_2 rwl_1_12 rwl_1_4 rwl_1_9 rwl_1_6 rwl_1_10 wwl_0_5
+ rwl_1_7 rwl_1_13 wwl_0_2 wwl_0_7 gnd wwl_0_3 wwl_0_8
Xcell_2r1w_60 vdd gnd read_bl_0_0 read_bl_1_0 write_bl_0_0 wwl_0_3 rwl_1_3 rwl_0_3
+ cell_2r1w
Xcell_2r1w_50 vdd_uq5 gnd read_bl_0_0 read_bl_1_0 write_bl_0_0 wwl_0_13 rwl_1_13 rwl_0_13
+ cell_2r1w
Xcell_2r1w_61 vdd gnd read_bl_0_0 read_bl_1_0 write_bl_0_0 wwl_0_2 rwl_1_2 rwl_0_2
+ cell_2r1w
Xcell_2r1w_51 vdd_uq5 gnd read_bl_0_0 read_bl_1_0 write_bl_0_0 wwl_0_12 rwl_1_12 rwl_0_12
+ cell_2r1w
Xcell_2r1w_52 vdd_uq4 gnd read_bl_0_0 read_bl_1_0 write_bl_0_0 wwl_0_11 rwl_1_11 rwl_0_11
+ cell_2r1w
Xcell_2r1w_40 vdd_uq2 gnd read_bl_0_1 read_bl_1_1 write_bl_0_1 wwl_0_7 rwl_1_7 rwl_0_7
+ cell_2r1w
Xcell_2r1w_41 vdd_uq2 gnd read_bl_0_1 read_bl_1_1 write_bl_0_1 wwl_0_6 rwl_1_6 rwl_0_6
+ cell_2r1w
Xcell_2r1w_30 vdd_uq0 gnd read_bl_0_2 read_bl_1_2 write_bl_0_2 wwl_0_1 rwl_1_1 rwl_0_1
+ cell_2r1w
Xcell_2r1w_62 vdd_uq0 gnd read_bl_0_0 read_bl_1_0 write_bl_0_0 wwl_0_1 rwl_1_1 rwl_0_1
+ cell_2r1w
Xcell_2r1w_63 vdd_uq0 gnd read_bl_0_0 read_bl_1_0 write_bl_0_0 wwl_0_0 rwl_1_0 rwl_0_0
+ cell_2r1w
Xcell_2r1w_20 vdd_uq4 gnd read_bl_0_2 read_bl_1_2 write_bl_0_2 wwl_0_11 rwl_1_11 rwl_0_11
+ cell_2r1w
Xcell_2r1w_53 vdd_uq4 gnd read_bl_0_0 read_bl_1_0 write_bl_0_0 wwl_0_10 rwl_1_10 rwl_0_10
+ cell_2r1w
Xcell_2r1w_42 vdd_uq1 gnd read_bl_0_1 read_bl_1_1 write_bl_0_1 wwl_0_5 rwl_1_5 rwl_0_5
+ cell_2r1w
Xcell_2r1w_31 vdd_uq0 gnd read_bl_0_2 read_bl_1_2 write_bl_0_2 wwl_0_0 rwl_1_0 rwl_0_0
+ cell_2r1w
Xcell_2r1w_0 vdd_uq6 gnd read_bl_0_3 read_bl_1_3 write_bl_0_3 wwl_0_15 rwl_1_15 rwl_0_15
+ cell_2r1w
Xcell_2r1w_32 vdd_uq6 gnd read_bl_0_1 read_bl_1_1 write_bl_0_1 wwl_0_15 rwl_1_15 rwl_0_15
+ cell_2r1w
Xcell_2r1w_21 vdd_uq4 gnd read_bl_0_2 read_bl_1_2 write_bl_0_2 wwl_0_10 rwl_1_10 rwl_0_10
+ cell_2r1w
Xcell_2r1w_54 vdd_uq3 gnd read_bl_0_0 read_bl_1_0 write_bl_0_0 wwl_0_9 rwl_1_9 rwl_0_9
+ cell_2r1w
Xcell_2r1w_10 vdd_uq1 gnd read_bl_0_3 read_bl_1_3 write_bl_0_3 wwl_0_5 rwl_1_5 rwl_0_5
+ cell_2r1w
Xcell_2r1w_43 vdd_uq1 gnd read_bl_0_1 read_bl_1_1 write_bl_0_1 wwl_0_4 rwl_1_4 rwl_0_4
+ cell_2r1w
Xcell_2r1w_1 vdd_uq6 gnd read_bl_0_3 read_bl_1_3 write_bl_0_3 wwl_0_14 rwl_1_14 rwl_0_14
+ cell_2r1w
Xcell_2r1w_33 vdd_uq6 gnd read_bl_0_1 read_bl_1_1 write_bl_0_1 wwl_0_14 rwl_1_14 rwl_0_14
+ cell_2r1w
Xcell_2r1w_22 vdd_uq3 gnd read_bl_0_2 read_bl_1_2 write_bl_0_2 wwl_0_9 rwl_1_9 rwl_0_9
+ cell_2r1w
Xcell_2r1w_55 vdd_uq3 gnd read_bl_0_0 read_bl_1_0 write_bl_0_0 wwl_0_8 rwl_1_8 rwl_0_8
+ cell_2r1w
Xcell_2r1w_11 vdd_uq1 gnd read_bl_0_3 read_bl_1_3 write_bl_0_3 wwl_0_4 rwl_1_4 rwl_0_4
+ cell_2r1w
Xcell_2r1w_44 vdd gnd read_bl_0_1 read_bl_1_1 write_bl_0_1 wwl_0_3 rwl_1_3 rwl_0_3
+ cell_2r1w
Xcell_2r1w_2 vdd_uq5 gnd read_bl_0_3 read_bl_1_3 write_bl_0_3 wwl_0_13 rwl_1_13 rwl_0_13
+ cell_2r1w
Xcell_2r1w_34 vdd_uq5 gnd read_bl_0_1 read_bl_1_1 write_bl_0_1 wwl_0_13 rwl_1_13 rwl_0_13
+ cell_2r1w
Xcell_2r1w_23 vdd_uq3 gnd read_bl_0_2 read_bl_1_2 write_bl_0_2 wwl_0_8 rwl_1_8 rwl_0_8
+ cell_2r1w
Xcell_2r1w_56 vdd_uq2 gnd read_bl_0_0 read_bl_1_0 write_bl_0_0 wwl_0_7 rwl_1_7 rwl_0_7
+ cell_2r1w
Xcell_2r1w_12 vdd gnd read_bl_0_3 read_bl_1_3 write_bl_0_3 wwl_0_3 rwl_1_3 rwl_0_3
+ cell_2r1w
Xcell_2r1w_45 vdd gnd read_bl_0_1 read_bl_1_1 write_bl_0_1 wwl_0_2 rwl_1_2 rwl_0_2
+ cell_2r1w
Xcell_2r1w_3 vdd_uq5 gnd read_bl_0_3 read_bl_1_3 write_bl_0_3 wwl_0_12 rwl_1_12 rwl_0_12
+ cell_2r1w
Xcell_2r1w_35 vdd_uq5 gnd read_bl_0_1 read_bl_1_1 write_bl_0_1 wwl_0_12 rwl_1_12 rwl_0_12
+ cell_2r1w
Xcell_2r1w_24 vdd_uq2 gnd read_bl_0_2 read_bl_1_2 write_bl_0_2 wwl_0_7 rwl_1_7 rwl_0_7
+ cell_2r1w
Xcell_2r1w_57 vdd_uq2 gnd read_bl_0_0 read_bl_1_0 write_bl_0_0 wwl_0_6 rwl_1_6 rwl_0_6
+ cell_2r1w
Xcell_2r1w_13 vdd gnd read_bl_0_3 read_bl_1_3 write_bl_0_3 wwl_0_2 rwl_1_2 rwl_0_2
+ cell_2r1w
Xcell_2r1w_46 vdd_uq0 gnd read_bl_0_1 read_bl_1_1 write_bl_0_1 wwl_0_1 rwl_1_1 rwl_0_1
+ cell_2r1w
Xcell_2r1w_4 vdd_uq4 gnd read_bl_0_3 read_bl_1_3 write_bl_0_3 wwl_0_11 rwl_1_11 rwl_0_11
+ cell_2r1w
Xcell_2r1w_36 vdd_uq4 gnd read_bl_0_1 read_bl_1_1 write_bl_0_1 wwl_0_11 rwl_1_11 rwl_0_11
+ cell_2r1w
Xcell_2r1w_25 vdd_uq2 gnd read_bl_0_2 read_bl_1_2 write_bl_0_2 wwl_0_6 rwl_1_6 rwl_0_6
+ cell_2r1w
Xcell_2r1w_58 vdd_uq1 gnd read_bl_0_0 read_bl_1_0 write_bl_0_0 wwl_0_5 rwl_1_5 rwl_0_5
+ cell_2r1w
Xcell_2r1w_14 vdd_uq0 gnd read_bl_0_3 read_bl_1_3 write_bl_0_3 wwl_0_1 rwl_1_1 rwl_0_1
+ cell_2r1w
Xcell_2r1w_47 vdd_uq0 gnd read_bl_0_1 read_bl_1_1 write_bl_0_1 wwl_0_0 rwl_1_0 rwl_0_0
+ cell_2r1w
Xcell_2r1w_48 vdd_uq6 gnd read_bl_0_0 read_bl_1_0 write_bl_0_0 wwl_0_15 rwl_1_15 rwl_0_15
+ cell_2r1w
Xcell_2r1w_5 vdd_uq4 gnd read_bl_0_3 read_bl_1_3 write_bl_0_3 wwl_0_10 rwl_1_10 rwl_0_10
+ cell_2r1w
Xcell_2r1w_37 vdd_uq4 gnd read_bl_0_1 read_bl_1_1 write_bl_0_1 wwl_0_10 rwl_1_10 rwl_0_10
+ cell_2r1w
Xcell_2r1w_26 vdd_uq1 gnd read_bl_0_2 read_bl_1_2 write_bl_0_2 wwl_0_5 rwl_1_5 rwl_0_5
+ cell_2r1w
Xcell_2r1w_59 vdd_uq1 gnd read_bl_0_0 read_bl_1_0 write_bl_0_0 wwl_0_4 rwl_1_4 rwl_0_4
+ cell_2r1w
Xcell_2r1w_15 vdd_uq0 gnd read_bl_0_3 read_bl_1_3 write_bl_0_3 wwl_0_0 rwl_1_0 rwl_0_0
+ cell_2r1w
Xcell_2r1w_16 vdd_uq6 gnd read_bl_0_2 read_bl_1_2 write_bl_0_2 wwl_0_15 rwl_1_15 rwl_0_15
+ cell_2r1w
Xcell_2r1w_17 vdd_uq6 gnd read_bl_0_2 read_bl_1_2 write_bl_0_2 wwl_0_14 rwl_1_14 rwl_0_14
+ cell_2r1w
Xcell_2r1w_49 vdd_uq6 gnd read_bl_0_0 read_bl_1_0 write_bl_0_0 wwl_0_14 rwl_1_14 rwl_0_14
+ cell_2r1w
Xcell_2r1w_6 vdd_uq3 gnd read_bl_0_3 read_bl_1_3 write_bl_0_3 wwl_0_9 rwl_1_9 rwl_0_9
+ cell_2r1w
Xcell_2r1w_38 vdd_uq3 gnd read_bl_0_1 read_bl_1_1 write_bl_0_1 wwl_0_9 rwl_1_9 rwl_0_9
+ cell_2r1w
Xcell_2r1w_39 vdd_uq3 gnd read_bl_0_1 read_bl_1_1 write_bl_0_1 wwl_0_8 rwl_1_8 rwl_0_8
+ cell_2r1w
Xcell_2r1w_27 vdd_uq1 gnd read_bl_0_2 read_bl_1_2 write_bl_0_2 wwl_0_4 rwl_1_4 rwl_0_4
+ cell_2r1w
Xcell_2r1w_28 vdd gnd read_bl_0_2 read_bl_1_2 write_bl_0_2 wwl_0_3 rwl_1_3 rwl_0_3
+ cell_2r1w
Xcell_2r1w_18 vdd_uq5 gnd read_bl_0_2 read_bl_1_2 write_bl_0_2 wwl_0_13 rwl_1_13 rwl_0_13
+ cell_2r1w
Xcell_2r1w_7 vdd_uq3 gnd read_bl_0_3 read_bl_1_3 write_bl_0_3 wwl_0_8 rwl_1_8 rwl_0_8
+ cell_2r1w
Xcell_2r1w_8 vdd_uq2 gnd read_bl_0_3 read_bl_1_3 write_bl_0_3 wwl_0_7 rwl_1_7 rwl_0_7
+ cell_2r1w
Xcell_2r1w_29 vdd gnd read_bl_0_2 read_bl_1_2 write_bl_0_2 wwl_0_2 rwl_1_2 rwl_0_2
+ cell_2r1w
Xcell_2r1w_19 vdd_uq5 gnd read_bl_0_2 read_bl_1_2 write_bl_0_2 wwl_0_12 rwl_1_12 rwl_0_12
+ cell_2r1w
Xcell_2r1w_9 vdd_uq2 gnd read_bl_0_3 read_bl_1_3 write_bl_0_3 wwl_0_6 rwl_1_6 rwl_0_6
+ cell_2r1w
.ends

.subckt replica_bitcell_array rwl_0_10 rwl_1_0 rwl_1_10 wwl_0_10 rwl_0_7 wwl_0_11
+ rwl_1_7 wwl_0_12 rwl_0_4 wwl_0_13 rwl_0_14 rwl_1_4 wwl_0_14 rwl_1_14 wwl_0_15 rwl_0_1
+ rwl_1_1 rwl_0_11 rwl_1_11 rwl_0_8 rwl_1_2 rwl_1_8 rwl_1_3 rwl_0_5 rwl_0_15 rwl_1_5
+ rwl_1_15 rwl_1_6 rwl_0_2 rwl_1_13 rwl_1_12 rwl_0_12 rwl_1_9 gnd rwl_0_9 wwl_0_0
+ wwl_0_1 rwl_0_6 wwl_0_2 wwl_0_3 wwl_0_4 wwl_0_5 rwl_0_3 wwl_0_7 wwl_0_6 rwl_0_0
+ rwl_0_13 wwl_0_8 wwl_0_9
Xbitcell_array_0 write_bl_0_3 read_bl_0_3 read_bl_0_1 read_bl_0_0 rwl_0_3 write_bl_0_1
+ rwl_1_14 read_bl_1_1 read_bl_1_3 read_bl_1_0 wwl_0_0 rwl_0_4 rwl_0_5 rwl_0_1 write_bl_0_0
+ rwl_0_6 wwl_0_10 rwl_1_1 read_bl_0_2 rwl_0_7 rwl_0_11 write_bl_0_2 wwl_0_11 rwl_0_14
+ wwl_0_15 rwl_1_11 rwl_0_8 wwl_0_12 rwl_0_9 wwl_0_13 rwl_0_10 wwl_0_14 rwl_1_8 rwl_0_12
+ read_bl_1_2 wwl_0_4 wwl_0_9 rwl_0_13 rwl_1_5 rwl_1_3 rwl_0_15 rwl_1_15 rwl_0_0 wwl_0_1
+ wwl_0_6 rwl_1_0 rwl_0_2 rwl_1_2 rwl_1_12 rwl_1_4 rwl_1_9 rwl_1_6 rwl_1_10 wwl_0_5
+ rwl_1_7 rwl_1_13 wwl_0_2 wwl_0_7 gnd wwl_0_3 wwl_0_8 bitcell_array
.ends

.subckt bank addr2 wl_en addr0 addr3 addr1 vdd addr4 gnd p_en_bar addr5 vdd_uq5 vdd_uq7
+ w_en vdd_uq29 dout1_0 vdd_uq9 vdd_uq23 dout1_1 dout1_2 dout1_3 vdd_uq39 vdd_uq33
+ vdd_uq40 vdd_uq30 vdd_uq41 vdd_uq20 vdd_uq31 vdd_uq43 vdd_uq11 vdd_uq21 vdd_uq12
+ vdd_uq34 vdd_uq13 vdd_uq24 vdd_uq35 vdd_uq14 vdd_uq25 vdd_uq36 vdd_uq15 vdd_uq26
+ vdd_uq37 vdd_uq16 vdd_uq27 vdd_uq17 vdd_uq19
Xport_data_0 p_en_bar vdd vdd_uq5 vdd_uq7 dout1_0 vdd_uq9 dout1_1 dout1_2 dout1_3
+ w_en p_en_bar gnd vdd_uq11 vdd_uq12 vdd_uq13 vdd_uq14 vdd_uq15 din0_0 din0_1 din0_2
+ din0_3 port_data
Xport_address_0 addr2 vdd_uq43 port_address_0/wwl0_0 port_address_0/rwl1_0 gnd port_address_0/rwl1_11
+ addr3 port_address_0/rwl1_1 port_address_0/wwl0_1 port_address_0/rwl1_12 vdd_uq16
+ addr4 vdd_uq26 vdd_uq19 port_address_0/wwl0_2 port_address_0/rwl1_2 port_address_0/rwl1_13
+ addr5 port_address_0/rwl1_3 port_address_0/wwl0_3 port_address_0/rwl1_14 port_address_0/rwl1_4
+ port_address_0/wwl0_4 vdd_uq20 port_address_0/rwl1_15 vdd_uq36 port_address_0/wwl0_5
+ port_address_0/rwl1_5 vdd_uq21 port_address_0/rwl1_6 port_address_0/wwl0_6 vdd_uq23
+ vdd_uq17 port_address_0/rwl1_7 port_address_0/wwl0_7 vdd_uq39 port_address_0/rwl1_8
+ port_address_0/wwl0_8 vdd_uq24 vdd_uq25 port_address_0/wwl0_9 port_address_0/rwl1_9
+ vdd_uq27 vdd_uq31 vdd_uq35 vdd_uq37 vdd_uq41 wl_en vdd_uq29 port_address_0/wwl0_10
+ port_address_0/wwl0_11 port_address_0/wwl0_12 port_address_0/rwl0_0 port_address_0/wwl0_13
+ port_address_0/wwl0_14 port_address_0/rwl0_1 port_address_0/rwl0_2 port_address_0/wwl0_15
+ port_address_0/rwl0_3 port_address_0/rwl0_10 port_address_0/rwl0_4 port_address_0/rwl0_11
+ port_address_0/rwl0_5 port_address_0/rwl0_12 port_address_0/rwl0_6 port_address_0/rwl0_13
+ vdd_uq40 vdd_uq33 port_address_0/rwl0_7 port_address_0/rwl0_14 vdd_uq30 port_address_0/rwl0_8
+ port_address_0/rwl0_15 port_address_0/rwl0_9 addr0 addr1 vdd_uq34 port_address_0/rwl1_10
+ port_address
Xreplica_bitcell_array_0 port_address_0/rwl0_10 port_address_0/rwl1_0 port_address_0/rwl1_10
+ port_address_0/wwl0_10 port_address_0/rwl0_7 port_address_0/wwl0_11 port_address_0/rwl1_7
+ port_address_0/wwl0_12 port_address_0/rwl0_4 port_address_0/wwl0_13 port_address_0/rwl0_14
+ port_address_0/rwl1_4 port_address_0/wwl0_14 port_address_0/rwl1_14 port_address_0/wwl0_15
+ port_address_0/rwl0_1 port_address_0/rwl1_1 port_address_0/rwl0_11 port_address_0/rwl1_11
+ port_address_0/rwl0_8 port_address_0/rwl1_2 port_address_0/rwl1_8 port_address_0/rwl1_3
+ port_address_0/rwl0_5 port_address_0/rwl0_15 port_address_0/rwl1_5 port_address_0/rwl1_15
+ port_address_0/rwl1_6 port_address_0/rwl0_2 port_address_0/rwl1_13 port_address_0/rwl1_12
+ port_address_0/rwl0_12 port_address_0/rwl1_9 gnd port_address_0/rwl0_9 port_address_0/wwl0_0
+ port_address_0/wwl0_1 port_address_0/rwl0_6 port_address_0/wwl0_2 port_address_0/wwl0_3
+ port_address_0/wwl0_4 port_address_0/wwl0_5 port_address_0/rwl0_3 port_address_0/wwl0_7
+ port_address_0/wwl0_6 port_address_0/rwl0_0 port_address_0/rwl0_13 port_address_0/wwl0_8
+ port_address_0/wwl0_9 replica_bitcell_array
.ends

.subckt sram_0rw2r1w_4_16_sky130A
Xcontrol_logic_multiport_0 vdd clk web vdd csb vdd vdd control_logic_multiport
Xdata_dff_0 vdd vdd vdd vdd vdd vdd vdd data_dff
Xrow_addr_dff_0 vdd vdd vdd vdd bank_0/addr0 bank_0/addr1 bank_0/addr3 bank_0/addr2
+ vdd bank_0/addr4 bank_0/addr5 vdd vdd addr1[1] addr1[2] addr1[3] addr1[4] addr1[5]
+ row_addr_dff
Xbank_0 bank_0/addr2 vdd bank_0/addr0 bank_0/addr3 bank_0/addr1 vdd bank_0/addr4 vdd
+ vdd bank_0/addr5 vdd vdd vdd vdd dout1[0] vdd vdd dout1[1] dout1[2] dout1[3] vdd
+ vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd
+ vdd vdd vdd vdd bank
.ends

