magic
tech sky130A
magscale 1 2
timestamp 1644969367
<< checkpaint >>
rect -1326 -1302 16788 7166
<< locali >>
rect 3995 4734 4214 4768
rect 4180 4550 4214 4734
rect 3977 2207 4162 2241
rect 3977 2154 4011 2207
rect 3844 2120 4011 2154
<< viali >>
rect 3712 5472 3746 5506
rect 6447 5479 6481 5513
rect 6915 4543 6949 4577
rect 3760 4463 3794 4497
rect 3760 3883 3794 3917
rect 5937 3804 5971 3838
rect 3860 3759 3894 3793
rect 3860 2911 3894 2945
rect 4747 2870 4781 2904
rect 3760 2787 3794 2821
rect 3712 2120 3746 2154
rect 5115 2124 5149 2158
rect 4228 2083 4262 2117
rect 3712 1198 3746 1232
rect 11933 1190 11967 1224
<< metal1 >>
rect 2958 5463 2964 5515
rect 3016 5503 3022 5515
rect 3700 5506 3758 5512
rect 3700 5503 3712 5506
rect 3016 5475 3712 5503
rect 3016 5463 3022 5475
rect 3700 5472 3712 5475
rect 3746 5472 3758 5506
rect 3700 5466 3758 5472
rect 6432 5470 6438 5522
rect 6490 5470 6496 5522
rect 6900 4534 6906 4586
rect 6958 4534 6964 4586
rect 3042 4454 3048 4506
rect 3100 4494 3106 4506
rect 3748 4497 3806 4503
rect 3748 4494 3760 4497
rect 3100 4466 3760 4494
rect 3100 4454 3106 4466
rect 3748 4463 3760 4466
rect 3794 4463 3806 4497
rect 3748 4457 3806 4463
rect 3126 3874 3132 3926
rect 3184 3914 3190 3926
rect 3748 3917 3806 3923
rect 3748 3914 3760 3917
rect 3184 3886 3760 3914
rect 3184 3874 3190 3886
rect 3748 3883 3760 3886
rect 3794 3883 3806 3917
rect 3748 3877 3806 3883
rect 2958 3750 2964 3802
rect 3016 3790 3022 3802
rect 3848 3793 3906 3799
rect 5922 3795 5928 3847
rect 5980 3795 5986 3847
rect 3848 3790 3860 3793
rect 3016 3762 3860 3790
rect 3016 3750 3022 3762
rect 3848 3759 3860 3762
rect 3894 3759 3906 3793
rect 3848 3753 3906 3759
rect -18 3246 -12 3298
rect 40 3286 46 3298
rect 3294 3286 3300 3298
rect 40 3258 3300 3286
rect 40 3246 46 3258
rect 3294 3246 3300 3258
rect 3352 3246 3358 3298
rect 3378 2902 3384 2954
rect 3436 2942 3442 2954
rect 3848 2945 3906 2951
rect 3848 2942 3860 2945
rect 3436 2914 3860 2942
rect 3436 2902 3442 2914
rect 3848 2911 3860 2914
rect 3894 2911 3906 2945
rect 3848 2905 3906 2911
rect 4732 2861 4738 2913
rect 4790 2861 4796 2913
rect 3294 2778 3300 2830
rect 3352 2818 3358 2830
rect 3748 2821 3806 2827
rect 3748 2818 3760 2821
rect 3352 2790 3760 2818
rect 3352 2778 3358 2790
rect 3748 2787 3760 2790
rect 3794 2787 3806 2821
rect 3748 2781 3806 2787
rect 3294 2111 3300 2163
rect 3352 2151 3358 2163
rect 3700 2154 3758 2160
rect 3700 2151 3712 2154
rect 3352 2123 3712 2151
rect 3352 2111 3358 2123
rect 3700 2120 3712 2123
rect 3746 2120 3758 2154
rect 3700 2114 3758 2120
rect 4213 2074 4219 2126
rect 4271 2074 4277 2126
rect 5100 2115 5106 2167
rect 5158 2115 5164 2167
rect 3697 1189 3703 1241
rect 3755 1189 3761 1241
rect 11918 1181 11924 1233
rect 11976 1181 11982 1233
<< via1 >>
rect 2964 5463 3016 5515
rect 6438 5513 6490 5522
rect 6438 5479 6447 5513
rect 6447 5479 6481 5513
rect 6481 5479 6490 5513
rect 6438 5470 6490 5479
rect 6906 4577 6958 4586
rect 6906 4543 6915 4577
rect 6915 4543 6949 4577
rect 6949 4543 6958 4577
rect 6906 4534 6958 4543
rect 3048 4454 3100 4506
rect 3132 3874 3184 3926
rect 2964 3750 3016 3802
rect 5928 3838 5980 3847
rect 5928 3804 5937 3838
rect 5937 3804 5971 3838
rect 5971 3804 5980 3838
rect 5928 3795 5980 3804
rect -12 3246 40 3298
rect 3300 3246 3352 3298
rect 3384 2902 3436 2954
rect 4738 2904 4790 2913
rect 4738 2870 4747 2904
rect 4747 2870 4781 2904
rect 4781 2870 4790 2904
rect 4738 2861 4790 2870
rect 3300 2778 3352 2830
rect 3300 2111 3352 2163
rect 4219 2117 4271 2126
rect 4219 2083 4228 2117
rect 4228 2083 4262 2117
rect 4262 2083 4271 2117
rect 4219 2074 4271 2083
rect 5106 2158 5158 2167
rect 5106 2124 5115 2158
rect 5115 2124 5149 2158
rect 5149 2124 5158 2158
rect 5106 2115 5158 2124
rect 3703 1232 3755 1241
rect 3703 1198 3712 1232
rect 3712 1198 3746 1232
rect 3746 1198 3755 1232
rect 3703 1189 3755 1198
rect 11924 1224 11976 1233
rect 11924 1190 11933 1224
rect 11933 1190 11967 1224
rect 11967 1190 11976 1224
rect 11924 1181 11976 1190
<< metal2 >>
rect 2976 5521 3004 5906
rect 2964 5515 3016 5521
rect 2964 5457 3016 5463
rect 2976 3808 3004 5457
rect 3060 4512 3088 5906
rect 3048 4506 3100 4512
rect 3048 4448 3100 4454
rect 2964 3802 3016 3808
rect 2964 3744 3016 3750
rect -12 3298 40 3304
rect -12 3240 40 3246
rect 0 1676 28 3240
rect 2976 1843 3004 3744
rect 3060 2924 3088 4448
rect 3144 3932 3172 5906
rect 3132 3926 3184 3932
rect 3132 3868 3184 3874
rect 3046 2915 3102 2924
rect 3046 2850 3102 2859
rect 2962 1834 3018 1843
rect 2962 1769 3018 1778
rect 2666 1531 2722 1540
rect 2666 1466 2722 1475
rect 180 1416 234 1444
rect 2158 1123 2214 1132
rect 2158 1058 2214 1067
rect 2158 609 2214 618
rect 2158 544 2214 553
rect 180 232 234 260
rect 2666 201 2722 210
rect 2666 136 2722 145
rect 2976 0 3004 1769
rect 3060 0 3088 2850
rect 3144 618 3172 3868
rect 3130 609 3186 618
rect 3130 544 3186 553
rect 3144 0 3172 544
rect 3228 210 3256 5906
rect 3312 3304 3340 5906
rect 3300 3298 3352 3304
rect 3300 3240 3352 3246
rect 3312 2836 3340 3240
rect 3396 2960 3424 5906
rect 3384 2954 3436 2960
rect 3384 2896 3436 2902
rect 3300 2830 3352 2836
rect 3300 2772 3352 2778
rect 3312 2169 3340 2772
rect 3300 2163 3352 2169
rect 3396 2137 3424 2896
rect 3300 2105 3352 2111
rect 3382 2128 3438 2137
rect 3312 909 3340 2105
rect 3382 2063 3438 2072
rect 3396 1132 3424 2063
rect 3480 1540 3508 5906
rect 6438 5522 6490 5528
rect 6490 5482 15528 5510
rect 6438 5464 6490 5470
rect 6906 4586 6958 4592
rect 6958 4546 15528 4574
rect 6906 4528 6958 4534
rect 5928 3847 5980 3853
rect 5980 3807 15528 3835
rect 5928 3789 5980 3795
rect 4736 2915 4792 2924
rect 4736 2850 4792 2859
rect 5106 2167 5158 2173
rect 4217 2128 4273 2137
rect 5106 2109 5158 2115
rect 4217 2063 4273 2072
rect 5118 1843 5146 2109
rect 5104 1834 5160 1843
rect 5104 1769 5160 1778
rect 3466 1531 3522 1540
rect 3466 1466 3522 1475
rect 3382 1123 3438 1132
rect 3382 1058 3438 1067
rect 3298 900 3354 909
rect 3298 835 3354 844
rect 3214 201 3270 210
rect 3214 136 3270 145
rect 3228 0 3256 136
rect 3312 0 3340 835
rect 3396 0 3424 1058
rect 3480 0 3508 1466
rect 3703 1241 3755 1247
rect 3703 1183 3755 1189
rect 11924 1233 11976 1239
rect 11976 1193 15528 1221
rect 11924 1175 11976 1181
rect 11936 909 11964 1175
rect 11922 900 11978 909
rect 11922 835 11978 844
<< via2 >>
rect 3046 2859 3102 2915
rect 2962 1778 3018 1834
rect 2666 1475 2722 1531
rect 2158 1067 2214 1123
rect 2158 553 2214 609
rect 2666 145 2722 201
rect 3130 553 3186 609
rect 3382 2072 3438 2128
rect 4736 2913 4792 2915
rect 4736 2861 4738 2913
rect 4738 2861 4790 2913
rect 4790 2861 4792 2913
rect 4736 2859 4792 2861
rect 4217 2126 4273 2128
rect 4217 2074 4219 2126
rect 4219 2074 4271 2126
rect 4271 2074 4273 2126
rect 4217 2072 4273 2074
rect 5104 1778 5160 1834
rect 3466 1475 3522 1531
rect 3382 1067 3438 1123
rect 3298 844 3354 900
rect 3214 145 3270 201
rect 11922 844 11978 900
<< metal3 >>
rect 3008 2917 3140 2920
rect 4698 2917 4830 2920
rect 3008 2915 4830 2917
rect 3008 2859 3046 2915
rect 3102 2859 4736 2915
rect 4792 2859 4830 2915
rect 3008 2857 4830 2859
rect 3008 2854 3140 2857
rect 4698 2854 4830 2857
rect 3344 2130 3476 2133
rect 4179 2130 4311 2133
rect 3344 2128 4311 2130
rect 3344 2072 3382 2128
rect 3438 2072 4217 2128
rect 4273 2072 4311 2128
rect 3344 2070 4311 2072
rect 3344 2067 3476 2070
rect 4179 2067 4311 2070
rect 2924 1836 3056 1839
rect 5066 1836 5198 1839
rect 2924 1834 5198 1836
rect 2924 1778 2962 1834
rect 3018 1778 5104 1834
rect 5160 1778 5198 1834
rect 2924 1776 5198 1778
rect 2924 1773 3056 1776
rect 5066 1773 5198 1776
rect -66 1639 66 1713
rect 2628 1533 2760 1536
rect 3428 1533 3560 1536
rect 2628 1531 3560 1533
rect 2628 1475 2666 1531
rect 2722 1475 3466 1531
rect 3522 1475 3560 1531
rect 2628 1473 3560 1475
rect 2628 1470 2760 1473
rect 3428 1470 3560 1473
rect 2120 1125 2252 1128
rect 3344 1125 3476 1128
rect 2120 1123 3476 1125
rect 2120 1067 2158 1123
rect 2214 1067 3382 1123
rect 3438 1067 3476 1123
rect 2120 1065 3476 1067
rect 2120 1062 2252 1065
rect 3344 1062 3476 1065
rect 3260 902 3392 905
rect 11884 902 12016 905
rect 3260 900 12016 902
rect -66 801 66 875
rect 3260 844 3298 900
rect 3354 844 11922 900
rect 11978 844 12016 900
rect 3260 842 12016 844
rect 3260 839 3392 842
rect 11884 839 12016 842
rect 2120 611 2252 614
rect 3092 611 3224 614
rect 2120 609 3224 611
rect 2120 553 2158 609
rect 2214 553 3130 609
rect 3186 553 3224 609
rect 2120 551 3224 553
rect 2120 548 2252 551
rect 3092 548 3224 551
rect 2628 203 2760 206
rect 3176 203 3308 206
rect 2628 201 3308 203
rect 2628 145 2666 201
rect 2722 145 3214 201
rect 3270 145 3308 201
rect 2628 143 3308 145
rect 2628 140 2760 143
rect 3176 140 3308 143
rect -66 -37 66 37
use contact_17  contact_17_0
timestamp 1644969367
transform 1 0 4732 0 1 2855
box 0 0 1 1
use contact_13  contact_13_0
timestamp 1644969367
transform 1 0 4735 0 1 2864
box 0 0 1 1
use contact_18  contact_18_0
timestamp 1644969367
transform 1 0 4698 0 1 2850
box 0 0 1 1
use contact_17  contact_17_1
timestamp 1644969367
transform 1 0 4732 0 1 2855
box 0 0 1 1
use contact_13  contact_13_1
timestamp 1644969367
transform 1 0 4735 0 1 2864
box 0 0 1 1
use contact_30  contact_30_0
timestamp 1644969367
transform 1 0 3008 0 1 2850
box 0 0 1 1
use contact_13  contact_13_2
timestamp 1644969367
transform 1 0 3848 0 1 2905
box 0 0 1 1
use contact_17  contact_17_2
timestamp 1644969367
transform 1 0 3378 0 1 2896
box 0 0 1 1
use contact_13  contact_13_3
timestamp 1644969367
transform 1 0 3748 0 1 2781
box 0 0 1 1
use contact_17  contact_17_3
timestamp 1644969367
transform 1 0 3294 0 1 2772
box 0 0 1 1
use contact_17  contact_17_4
timestamp 1644969367
transform 1 0 5100 0 1 2109
box 0 0 1 1
use contact_13  contact_13_4
timestamp 1644969367
transform 1 0 5103 0 1 2118
box 0 0 1 1
use contact_30  contact_30_1
timestamp 1644969367
transform 1 0 2924 0 1 1769
box 0 0 1 1
use contact_30  contact_30_2
timestamp 1644969367
transform 1 0 5066 0 1 1769
box 0 0 1 1
use contact_18  contact_18_1
timestamp 1644969367
transform 1 0 4179 0 1 2063
box 0 0 1 1
use contact_17  contact_17_5
timestamp 1644969367
transform 1 0 4213 0 1 2068
box 0 0 1 1
use contact_13  contact_13_5
timestamp 1644969367
transform 1 0 4216 0 1 2077
box 0 0 1 1
use contact_18  contact_18_2
timestamp 1644969367
transform 1 0 4179 0 1 2063
box 0 0 1 1
use contact_17  contact_17_6
timestamp 1644969367
transform 1 0 4213 0 1 2068
box 0 0 1 1
use contact_13  contact_13_6
timestamp 1644969367
transform 1 0 4216 0 1 2077
box 0 0 1 1
use contact_30  contact_30_3
timestamp 1644969367
transform 1 0 3344 0 1 2063
box 0 0 1 1
use contact_13  contact_13_7
timestamp 1644969367
transform 1 0 3700 0 1 2114
box 0 0 1 1
use contact_17  contact_17_7
timestamp 1644969367
transform 1 0 3294 0 1 2105
box 0 0 1 1
use contact_17  contact_17_8
timestamp 1644969367
transform 1 0 11918 0 1 1175
box 0 0 1 1
use contact_13  contact_13_8
timestamp 1644969367
transform 1 0 11921 0 1 1184
box 0 0 1 1
use contact_17  contact_17_9
timestamp 1644969367
transform 1 0 11918 0 1 1175
box 0 0 1 1
use contact_13  contact_13_9
timestamp 1644969367
transform 1 0 11921 0 1 1184
box 0 0 1 1
use contact_30  contact_30_4
timestamp 1644969367
transform 1 0 3260 0 1 835
box 0 0 1 1
use contact_30  contact_30_5
timestamp 1644969367
transform 1 0 11884 0 1 835
box 0 0 1 1
use contact_17  contact_17_10
timestamp 1644969367
transform 1 0 3697 0 1 1183
box 0 0 1 1
use contact_13  contact_13_10
timestamp 1644969367
transform 1 0 3700 0 1 1192
box 0 0 1 1
use contact_17  contact_17_11
timestamp 1644969367
transform 1 0 6900 0 1 4528
box 0 0 1 1
use contact_13  contact_13_11
timestamp 1644969367
transform 1 0 6903 0 1 4537
box 0 0 1 1
use contact_13  contact_13_12
timestamp 1644969367
transform 1 0 3748 0 1 4457
box 0 0 1 1
use contact_17  contact_17_12
timestamp 1644969367
transform 1 0 3042 0 1 4448
box 0 0 1 1
use contact_17  contact_17_13
timestamp 1644969367
transform 1 0 5922 0 1 3789
box 0 0 1 1
use contact_13  contact_13_13
timestamp 1644969367
transform 1 0 5925 0 1 3798
box 0 0 1 1
use contact_13  contact_13_14
timestamp 1644969367
transform 1 0 3848 0 1 3753
box 0 0 1 1
use contact_17  contact_17_14
timestamp 1644969367
transform 1 0 2958 0 1 3744
box 0 0 1 1
use contact_13  contact_13_15
timestamp 1644969367
transform 1 0 3748 0 1 3877
box 0 0 1 1
use contact_17  contact_17_15
timestamp 1644969367
transform 1 0 3126 0 1 3868
box 0 0 1 1
use contact_17  contact_17_16
timestamp 1644969367
transform 1 0 6432 0 1 5464
box 0 0 1 1
use contact_13  contact_13_16
timestamp 1644969367
transform 1 0 6435 0 1 5473
box 0 0 1 1
use contact_13  contact_13_17
timestamp 1644969367
transform 1 0 3700 0 1 5466
box 0 0 1 1
use contact_17  contact_17_17
timestamp 1644969367
transform 1 0 2958 0 1 5457
box 0 0 1 1
use contact_17  contact_17_18
timestamp 1644969367
transform 1 0 3294 0 1 3240
box 0 0 1 1
use contact_17  contact_17_19
timestamp 1644969367
transform 1 0 -18 0 1 3240
box 0 0 1 1
use contact_18  contact_18_3
timestamp 1644969367
transform 1 0 2628 0 1 1466
box 0 0 1 1
use contact_30  contact_30_6
timestamp 1644969367
transform 1 0 3428 0 1 1466
box 0 0 1 1
use contact_18  contact_18_4
timestamp 1644969367
transform 1 0 2120 0 1 1058
box 0 0 1 1
use contact_30  contact_30_7
timestamp 1644969367
transform 1 0 3344 0 1 1058
box 0 0 1 1
use contact_18  contact_18_5
timestamp 1644969367
transform 1 0 2628 0 1 136
box 0 0 1 1
use contact_30  contact_30_8
timestamp 1644969367
transform 1 0 3176 0 1 136
box 0 0 1 1
use contact_18  contact_18_6
timestamp 1644969367
transform 1 0 2120 0 1 544
box 0 0 1 1
use contact_30  contact_30_9
timestamp 1644969367
transform 1 0 3092 0 1 544
box 0 0 1 1
use pdriver_1  pdriver_1_0
timestamp 1644969367
transform 1 0 4116 0 1 4190
box -36 -17 3992 895
use pnand2_1  pnand2_1_0
timestamp 1644969367
transform 1 0 3648 0 1 4190
box -36 -17 504 895
use pand2_0  pand2_0_0
timestamp 1644969367
transform 1 0 3648 0 -1 4190
box -36 -17 4346 895
use pdriver_1  pdriver_1_1
timestamp 1644969367
transform 1 0 3648 0 -1 5866
box -36 -17 3992 895
use pand2  pand2_0
timestamp 1644969367
transform 1 0 3648 0 1 2514
box -36 -17 1862 895
use pand2  pand2_1
timestamp 1644969367
transform 1 0 4016 0 -1 2514
box -36 -17 1862 895
use pinv_0  pinv_0_0
timestamp 1644969367
transform 1 0 3648 0 -1 2514
box -36 -17 404 895
use pdriver_0  pdriver_0_0
timestamp 1644969367
transform 1 0 3648 0 1 838
box -36 -17 11748 895
use dff_buf_array  dff_buf_array_0
timestamp 1644969367
transform 1 0 0 0 1 0
box -66 -42 3012 1718
<< labels >>
rlabel metal2 s 180 1416 234 1444 4 csb
rlabel metal2 s 180 232 234 260 4 web
rlabel metal2 s 6464 5482 15528 5510 4 wl_en
rlabel metal2 s 5954 3807 15528 3835 4 w_en
rlabel metal2 s 6932 4546 15528 4574 4 p_en_bar
rlabel metal2 s 3715 1201 3743 1229 4 clk
rlabel metal2 s 11950 1193 15528 1221 4 clk_buf
rlabel metal3 s -66 -37 66 37 4 gnd
rlabel metal3 s -66 1639 66 1713 4 gnd
rlabel metal3 s -66 801 66 875 4 vdd
<< properties >>
string FIXED_BBOX 0 0 15528 160
string GDS_FILE sram_0rw2r1w_32_128_sky130A.gds
string GDS_END 3276626
string GDS_START 3267916
<< end >>
