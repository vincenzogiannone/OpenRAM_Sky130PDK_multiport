magic
tech sky130A
magscale 1 2
timestamp 1644951705
<< checkpaint >>
rect -1260 -1260 59706 57160
<< viali >>
rect 5910 5094 5944 5128
rect 5910 4172 5944 4206
rect 5910 3418 5944 3452
rect 5910 2496 5944 2530
<< metal1 >>
rect 7735 55144 7876 55172
rect 7735 55100 7763 55144
rect 7586 55072 7763 55100
rect 7735 55018 7876 55046
rect 7735 54974 7763 55018
rect 7586 54946 7763 54974
rect 7735 54792 7876 54820
rect 7735 54748 7763 54792
rect 7586 54720 7763 54748
rect 7735 53732 7876 53760
rect 7735 53708 7763 53732
rect 7586 53680 7763 53708
rect 7735 53506 7876 53534
rect 7735 53482 7763 53506
rect 7586 53454 7763 53482
rect 7735 53380 7876 53408
rect 7735 53356 7763 53380
rect 7586 53328 7763 53356
rect 7735 52064 7876 52092
rect 7735 52024 7763 52064
rect 7586 51996 7763 52024
rect 7735 51938 7876 51966
rect 7735 51898 7763 51938
rect 7586 51870 7763 51898
rect 7735 51712 7876 51740
rect 7735 51672 7763 51712
rect 7586 51644 7763 51672
rect 7735 50652 7876 50680
rect 7735 50632 7763 50652
rect 7586 50604 7763 50632
rect 7735 50426 7876 50454
rect 7735 50406 7763 50426
rect 7586 50378 7763 50406
rect 7735 50300 7876 50328
rect 7735 50280 7763 50300
rect 7586 50252 7763 50280
rect 7735 48984 7876 49012
rect 7735 48948 7763 48984
rect 7586 48920 7763 48948
rect 7735 48858 7876 48886
rect 7735 48822 7763 48858
rect 7586 48794 7763 48822
rect 7735 48632 7876 48660
rect 7735 48596 7763 48632
rect 7586 48568 7763 48596
rect 7735 47572 7876 47600
rect 7735 47556 7763 47572
rect 7586 47528 7763 47556
rect 7735 47346 7876 47374
rect 7735 47330 7763 47346
rect 7586 47302 7763 47330
rect 7735 47220 7876 47248
rect 7735 47204 7763 47220
rect 7586 47176 7763 47204
rect 7735 45904 7876 45932
rect 7735 45872 7763 45904
rect 7586 45844 7763 45872
rect 7735 45778 7876 45806
rect 7735 45746 7763 45778
rect 7586 45718 7763 45746
rect 7735 45552 7876 45580
rect 7735 45520 7763 45552
rect 7586 45492 7763 45520
rect 7735 44492 7876 44520
rect 7735 44480 7763 44492
rect 7586 44452 7763 44480
rect 7735 44266 7876 44294
rect 7735 44254 7763 44266
rect 7586 44226 7763 44254
rect 7735 44140 7876 44168
rect 7735 44128 7763 44140
rect 7586 44100 7763 44128
rect 7735 42824 7876 42852
rect 7735 42796 7763 42824
rect 7586 42768 7763 42796
rect 7735 42698 7876 42726
rect 7735 42670 7763 42698
rect 7586 42642 7763 42670
rect 7735 42472 7876 42500
rect 7735 42444 7763 42472
rect 7586 42416 7763 42444
rect 7735 41412 7876 41440
rect 7735 41404 7763 41412
rect 7586 41376 7763 41404
rect 7735 41186 7876 41214
rect 7735 41178 7763 41186
rect 7586 41150 7763 41178
rect 7735 41060 7876 41088
rect 7735 41052 7763 41060
rect 7586 41024 7763 41052
rect 7735 39744 7876 39772
rect 7735 39720 7763 39744
rect 7586 39692 7763 39720
rect 7735 39618 7876 39646
rect 7735 39594 7763 39618
rect 7586 39566 7763 39594
rect 7735 39392 7876 39420
rect 7735 39368 7763 39392
rect 7586 39340 7763 39368
rect 7735 38332 7876 38360
rect 7735 38328 7763 38332
rect 7586 38300 7763 38328
rect 7735 38106 7876 38134
rect 7735 38102 7763 38106
rect 7586 38074 7763 38102
rect 7735 37980 7876 38008
rect 7735 37976 7763 37980
rect 7586 37948 7763 37976
rect 7735 36664 7876 36692
rect 7735 36644 7763 36664
rect 7586 36616 7763 36644
rect 7735 36538 7876 36566
rect 7735 36518 7763 36538
rect 7586 36490 7763 36518
rect 7735 36312 7876 36340
rect 7735 36292 7763 36312
rect 7586 36264 7763 36292
rect 7735 35252 7876 35280
rect 7586 35224 7763 35252
rect 7735 35026 7876 35054
rect 7586 34998 7763 35026
rect 7735 34900 7876 34928
rect 7586 34872 7763 34900
rect 7735 33584 7876 33612
rect 7735 33568 7763 33584
rect 7586 33540 7763 33568
rect 7735 33458 7876 33486
rect 7735 33442 7763 33458
rect 7586 33414 7763 33442
rect 7735 33232 7876 33260
rect 7735 33216 7763 33232
rect 7586 33188 7763 33216
rect 7735 32176 7876 32200
rect 7586 32172 7876 32176
rect 7586 32148 7763 32172
rect 7735 31950 7876 31974
rect 7586 31946 7876 31950
rect 7586 31922 7763 31946
rect 7735 31824 7876 31848
rect 7586 31820 7876 31824
rect 7586 31796 7763 31820
rect 7735 30504 7876 30532
rect 7735 30492 7763 30504
rect 7586 30464 7763 30492
rect 7735 30378 7876 30406
rect 7735 30366 7763 30378
rect 7586 30338 7763 30366
rect 7735 30152 7876 30180
rect 7735 30140 7763 30152
rect 7586 30112 7763 30140
rect 7735 29100 7876 29120
rect 7586 29092 7876 29100
rect 7586 29072 7763 29092
rect 7735 28874 7876 28894
rect 7586 28866 7876 28874
rect 7586 28846 7763 28866
rect 7735 28748 7876 28768
rect 7586 28740 7876 28748
rect 7586 28720 7763 28740
rect 7735 27424 7876 27452
rect 7735 27416 7763 27424
rect 7586 27388 7763 27416
rect 7735 27298 7876 27326
rect 7735 27290 7763 27298
rect 7586 27262 7763 27290
rect 7735 27072 7876 27100
rect 7735 27064 7763 27072
rect 7586 27036 7763 27064
rect 7735 26024 7876 26040
rect 7586 26012 7876 26024
rect 7586 25996 7763 26012
rect 7735 25798 7876 25814
rect 7586 25786 7876 25798
rect 7586 25770 7763 25786
rect 7735 25672 7876 25688
rect 7586 25660 7876 25672
rect 7586 25644 7763 25660
rect 7735 24344 7876 24372
rect 7735 24340 7763 24344
rect 7586 24312 7763 24340
rect 7735 24218 7876 24246
rect 7735 24214 7763 24218
rect 7586 24186 7763 24214
rect 7735 23992 7876 24020
rect 7735 23988 7763 23992
rect 7586 23960 7763 23988
rect 7735 22948 7876 22960
rect 7586 22932 7876 22948
rect 7586 22920 7763 22932
rect 7735 22722 7876 22734
rect 7586 22706 7876 22722
rect 7586 22694 7763 22706
rect 7735 22596 7876 22608
rect 7586 22580 7876 22596
rect 7586 22568 7763 22580
rect 7735 21264 7876 21292
rect 7586 21236 7763 21264
rect 7735 21138 7876 21166
rect 7586 21110 7763 21138
rect 7735 20912 7876 20940
rect 7586 20884 7763 20912
rect 7735 19872 7876 19880
rect 7586 19852 7876 19872
rect 7586 19844 7763 19852
rect 7735 19646 7876 19654
rect 7586 19626 7876 19646
rect 7586 19618 7763 19626
rect 7735 19520 7876 19528
rect 7586 19500 7876 19520
rect 7586 19492 7763 19500
rect 7735 18188 7876 18212
rect 7586 18184 7876 18188
rect 7586 18160 7763 18184
rect 7735 18062 7876 18086
rect 7586 18058 7876 18062
rect 7586 18034 7763 18058
rect 7735 17836 7876 17860
rect 7586 17832 7876 17836
rect 7586 17808 7763 17832
rect 7735 16796 7876 16800
rect 7586 16772 7876 16796
rect 7586 16768 7763 16772
rect 7735 16570 7876 16574
rect 7586 16546 7876 16570
rect 7586 16542 7763 16546
rect 7735 16444 7876 16448
rect 7586 16420 7876 16444
rect 7586 16416 7763 16420
rect 7735 15112 7876 15132
rect 7586 15104 7876 15112
rect 7586 15084 7763 15104
rect 7735 14986 7876 15006
rect 7586 14978 7876 14986
rect 7586 14958 7763 14978
rect 7735 14760 7876 14780
rect 7586 14752 7876 14760
rect 7586 14732 7763 14752
rect 7586 13692 7876 13720
rect 7586 13466 7876 13494
rect 7586 13340 7876 13368
rect 7735 12036 7876 12052
rect 7586 12024 7876 12036
rect 7586 12008 7763 12024
rect 7735 11910 7876 11926
rect 7586 11898 7876 11910
rect 7586 11882 7763 11898
rect 7735 11684 7876 11700
rect 7586 11672 7876 11684
rect 7586 11656 7763 11672
rect 7586 10640 7763 10644
rect 7586 10616 7876 10640
rect 7735 10612 7876 10616
rect 7586 10414 7763 10418
rect 7586 10390 7876 10414
rect 7735 10386 7876 10390
rect 7586 10288 7763 10292
rect 7586 10264 7876 10288
rect 7735 10260 7876 10264
rect 7735 8960 7876 8972
rect 7586 8944 7876 8960
rect 7586 8932 7763 8944
rect 7735 8834 7876 8846
rect 7586 8818 7876 8834
rect 7586 8806 7763 8818
rect 7735 8608 7876 8620
rect 7586 8592 7876 8608
rect 7586 8580 7763 8592
rect 7586 7560 7763 7568
rect 7586 7540 7876 7560
rect 7735 7532 7876 7540
rect 7586 7334 7763 7342
rect 7586 7314 7876 7334
rect 7735 7306 7876 7314
rect 7586 7208 7763 7216
rect 7586 7188 7876 7208
rect 7735 7180 7876 7188
rect 7486 5972 7492 6024
rect 7544 6012 7550 6024
rect 7544 5984 31760 6012
rect 7544 5972 7550 5984
rect 3494 5085 3500 5137
rect 3552 5125 3558 5137
rect 5898 5128 5956 5134
rect 5898 5125 5910 5128
rect 3552 5097 5910 5125
rect 3552 5085 3558 5097
rect 5898 5094 5910 5097
rect 5944 5094 5956 5128
rect 5898 5088 5956 5094
rect 3586 4163 3592 4215
rect 3644 4203 3650 4215
rect 5898 4206 5956 4212
rect 5898 4203 5910 4206
rect 3644 4175 5910 4203
rect 3644 4163 3650 4175
rect 5898 4172 5910 4175
rect 5944 4172 5956 4206
rect 5898 4166 5956 4172
rect 3310 3582 3316 3634
rect 3368 3622 3374 3634
rect 3368 3594 7890 3622
rect 3368 3582 3374 3594
rect 3420 3514 7890 3542
rect 3420 3449 3448 3514
rect 3586 3449 3592 3474
rect 3420 3422 3592 3449
rect 3644 3462 3650 3474
rect 3644 3452 7890 3462
rect 3644 3422 5910 3452
rect 3420 3421 5910 3422
rect 5898 3418 5910 3421
rect 5944 3434 7890 3452
rect 5944 3418 5956 3434
rect 5898 3412 5956 3418
rect 3494 3342 3500 3394
rect 3552 3382 3558 3394
rect 3552 3354 7890 3382
rect 3552 3342 3558 3354
rect 3310 2487 3316 2539
rect 3368 2527 3374 2539
rect 5898 2530 5956 2536
rect 5898 2527 5910 2530
rect 3368 2499 5910 2527
rect 3368 2487 3374 2499
rect 5898 2496 5910 2499
rect 5944 2496 5956 2530
rect 5898 2490 5956 2496
rect 57960 1531 57966 1543
rect 33161 1503 57966 1531
rect 57960 1491 57966 1503
rect 58018 1491 58024 1543
<< via1 >>
rect 7492 5972 7544 6024
rect 3500 5085 3552 5137
rect 3592 4163 3644 4215
rect 3316 3582 3368 3634
rect 3592 3422 3644 3474
rect 3500 3342 3552 3394
rect 3316 2487 3368 2539
rect 57966 1491 58018 1543
<< metal2 >>
rect 6382 55738 6410 55766
rect 18 6536 46 37328
rect 102 6536 130 37328
rect 186 6536 214 37328
rect 270 6536 298 37328
rect 354 6536 382 37328
rect 438 6536 466 37328
rect 522 6536 550 37328
rect 7504 6030 7532 6116
rect 8461 6068 8515 6096
rect 11573 6068 11627 6096
rect 14685 6068 14739 6096
rect 17797 6068 17851 6096
rect 20909 6068 20963 6096
rect 24021 6068 24075 6096
rect 27133 6068 27187 6096
rect 30245 6068 30299 6096
rect 33357 6068 33411 6096
rect 36469 6068 36523 6096
rect 39581 6068 39635 6096
rect 42693 6068 42747 6096
rect 45805 6068 45859 6096
rect 48917 6068 48971 6096
rect 52029 6068 52083 6096
rect 55141 6068 55195 6096
rect 7492 6024 7544 6030
rect 7492 5966 7544 5972
rect 3500 5137 3552 5143
rect 3500 5079 3552 5085
rect 3316 3634 3368 3640
rect 3316 3576 3368 3582
rect 3328 2545 3356 3576
rect 3512 3400 3540 5079
rect 3592 4215 3644 4221
rect 3592 4157 3644 4163
rect 3604 3480 3632 4157
rect 3592 3474 3644 3480
rect 3592 3416 3644 3422
rect 3998 3403 4050 3467
rect 3500 3394 3552 3400
rect 3500 3336 3552 3342
rect 3316 2539 3368 2545
rect 3316 2481 3368 2487
rect 3874 2481 3926 2545
rect 7504 0 7532 5966
rect 8195 4924 8223 5164
rect 8467 4924 8495 5164
rect 11307 4924 11335 5164
rect 11579 4924 11607 5164
rect 14419 4924 14447 5164
rect 14691 4924 14719 5164
rect 17531 4924 17559 5164
rect 17803 4924 17831 5164
rect 20643 4924 20671 5164
rect 20915 4924 20943 5164
rect 23755 4924 23783 5164
rect 24027 4924 24055 5164
rect 26867 4924 26895 5164
rect 27139 4924 27167 5164
rect 29979 4924 30007 5164
rect 30251 4924 30279 5164
rect 57978 1549 58006 55900
rect 57966 1543 58018 1549
rect 57966 1485 58018 1491
rect 57978 0 58006 1485
<< metal3 >>
rect 5980 55715 6112 55789
rect 7520 55715 7652 55789
rect 5980 54177 6112 54251
rect 7520 54177 7652 54251
rect 5980 52639 6112 52713
rect 7520 52639 7652 52713
rect 5980 51101 6112 51175
rect 7520 51101 7652 51175
rect 5980 49563 6112 49637
rect 7520 49563 7652 49637
rect 5980 48025 6112 48099
rect 7520 48025 7652 48099
rect 5980 46487 6112 46561
rect 7520 46487 7652 46561
rect 5980 44949 6112 45023
rect 7520 44949 7652 45023
rect 5980 43411 6112 43485
rect 7520 43411 7652 43485
rect 5980 41873 6112 41947
rect 7520 41873 7652 41947
rect 5980 40335 6112 40409
rect 7520 40335 7652 40409
rect 5980 38797 6112 38871
rect 7520 38797 7652 38871
rect 960 37291 1092 37365
rect 2000 37291 2132 37365
rect 5980 37259 6112 37333
rect 7520 37259 7652 37333
rect 960 35751 1092 35825
rect 2000 35751 2132 35825
rect 5980 35721 6112 35795
rect 7520 35721 7652 35795
rect 960 34211 1092 34285
rect 2000 34211 2132 34285
rect 5980 34183 6112 34257
rect 7520 34183 7652 34257
rect 960 32671 1092 32745
rect 2000 32671 2132 32745
rect 5980 32645 6112 32719
rect 7520 32645 7652 32719
rect 960 31131 1092 31205
rect 2000 31131 2132 31205
rect 5980 31107 6112 31181
rect 7520 31107 7652 31181
rect 960 29591 1092 29665
rect 2000 29591 2132 29665
rect 5980 29569 6112 29643
rect 7520 29569 7652 29643
rect 960 28051 1092 28125
rect 2000 28051 2132 28125
rect 5980 28031 6112 28105
rect 7520 28031 7652 28105
rect 960 26511 1092 26585
rect 2000 26511 2132 26585
rect 5980 26493 6112 26567
rect 7520 26493 7652 26567
rect 960 24971 1092 25045
rect 2000 24971 2132 25045
rect 5980 24955 6112 25029
rect 7520 24955 7652 25029
rect 5980 23417 6112 23491
rect 7520 23417 7652 23491
rect 1308 21895 1440 21969
rect 2180 21895 2312 21969
rect 5980 21879 6112 21953
rect 7520 21879 7652 21953
rect 1308 20355 1440 20429
rect 2180 20355 2312 20429
rect 5980 20341 6112 20415
rect 7520 20341 7652 20415
rect 1308 18815 1440 18889
rect 2180 18815 2312 18889
rect 5980 18803 6112 18877
rect 7520 18803 7652 18877
rect 1308 17275 1440 17349
rect 2180 17275 2312 17349
rect 5980 17265 6112 17339
rect 7520 17265 7652 17339
rect 1308 15735 1440 15809
rect 2180 15735 2312 15809
rect 5980 15727 6112 15801
rect 7520 15727 7652 15801
rect 5980 14189 6112 14263
rect 7520 14189 7652 14263
rect 1308 12659 1440 12733
rect 2180 12659 2312 12733
rect 5980 12651 6112 12725
rect 7520 12651 7652 12725
rect 1308 11119 1440 11193
rect 2180 11119 2312 11193
rect 5980 11113 6112 11187
rect 7520 11113 7652 11187
rect 1308 9579 1440 9653
rect 2180 9579 2312 9653
rect 5980 9575 6112 9649
rect 7520 9575 7652 9649
rect 1308 8039 1440 8113
rect 2180 8039 2312 8113
rect 5980 8037 6112 8111
rect 7520 8037 7652 8111
rect 1308 6499 1440 6573
rect 2180 6499 2312 6573
rect 5980 6499 6112 6573
rect 7520 6499 7652 6573
rect 8581 6260 8647 6392
rect 11693 6260 11759 6392
rect 14805 6260 14871 6392
rect 17917 6260 17983 6392
rect 21029 6260 21095 6392
rect 24141 6260 24207 6392
rect 27253 6260 27319 6392
rect 30365 6260 30431 6392
rect 33477 6260 33543 6392
rect 36589 6260 36655 6392
rect 39701 6260 39767 6392
rect 42813 6260 42879 6392
rect 45925 6260 45991 6392
rect 49037 6260 49103 6392
rect 52149 6260 52215 6392
rect 55261 6260 55327 6392
rect 4132 5451 4264 5525
rect 5244 5451 5376 5525
rect 8581 5428 8647 5560
rect 11693 5428 11759 5560
rect 14805 5428 14871 5560
rect 17917 5428 17983 5560
rect 21029 5428 21095 5560
rect 24141 5428 24207 5560
rect 27253 5428 27319 5560
rect 30365 5428 30431 5560
rect 33477 5428 33543 5560
rect 36589 5428 36655 5560
rect 39701 5428 39767 5560
rect 42813 5428 42879 5560
rect 45925 5428 45991 5560
rect 49037 5428 49103 5560
rect 52149 5428 52215 5560
rect 55261 5428 55327 5560
rect 8063 5093 8195 5167
rect 8335 5093 8467 5167
rect 11175 5093 11307 5167
rect 11447 5093 11579 5167
rect 14287 5093 14419 5167
rect 14559 5093 14691 5167
rect 17399 5093 17531 5167
rect 17671 5093 17803 5167
rect 20511 5093 20643 5167
rect 20783 5093 20915 5167
rect 23623 5093 23755 5167
rect 23895 5093 24027 5167
rect 26735 5093 26867 5167
rect 27007 5093 27139 5167
rect 29847 5093 29979 5167
rect 30119 5093 30251 5167
rect 32959 5093 33091 5167
rect 33231 5093 33363 5167
rect 36071 5093 36203 5167
rect 36343 5093 36475 5167
rect 39183 5093 39315 5167
rect 39455 5093 39587 5167
rect 42295 5093 42427 5167
rect 42567 5093 42699 5167
rect 45407 5093 45539 5167
rect 45679 5093 45811 5167
rect 48519 5093 48651 5167
rect 48791 5093 48923 5167
rect 51631 5093 51763 5167
rect 51903 5093 52035 5167
rect 54743 5093 54875 5167
rect 55015 5093 55147 5167
rect 4132 4613 4264 4687
rect 5244 4613 5376 4687
rect 8063 4147 8195 4221
rect 8335 4147 8467 4221
rect 11175 4147 11307 4221
rect 11447 4147 11579 4221
rect 14287 4147 14419 4221
rect 14559 4147 14691 4221
rect 17399 4147 17531 4221
rect 17671 4147 17803 4221
rect 20511 4147 20643 4221
rect 20783 4147 20915 4221
rect 23623 4147 23755 4221
rect 23895 4147 24027 4221
rect 26735 4147 26867 4221
rect 27007 4147 27139 4221
rect 29847 4147 29979 4221
rect 30119 4147 30251 4221
rect 32959 4147 33091 4221
rect 33231 4147 33363 4221
rect 36071 4147 36203 4221
rect 36343 4147 36475 4221
rect 39183 4147 39315 4221
rect 39455 4147 39587 4221
rect 42295 4147 42427 4221
rect 42567 4147 42699 4221
rect 45407 4147 45539 4221
rect 45679 4147 45811 4221
rect 48519 4147 48651 4221
rect 48791 4147 48923 4221
rect 51631 4147 51763 4221
rect 51903 4147 52035 4221
rect 54743 4147 54875 4221
rect 55015 4147 55147 4221
rect 4132 3775 4264 3849
rect 5244 3775 5376 3849
rect 4132 2937 4264 3011
rect 5244 2937 5376 3011
rect 8588 2506 8720 2580
rect 9366 2506 9498 2580
rect 10144 2506 10276 2580
rect 10922 2506 11054 2580
rect 11700 2506 11832 2580
rect 12478 2506 12610 2580
rect 13256 2506 13388 2580
rect 14034 2506 14166 2580
rect 14812 2506 14944 2580
rect 15590 2506 15722 2580
rect 16368 2506 16500 2580
rect 17146 2506 17278 2580
rect 17924 2506 18056 2580
rect 18702 2506 18834 2580
rect 19480 2506 19612 2580
rect 20258 2506 20390 2580
rect 21036 2506 21168 2580
rect 21814 2506 21946 2580
rect 22592 2506 22724 2580
rect 23370 2506 23502 2580
rect 24148 2506 24280 2580
rect 24926 2506 25058 2580
rect 25704 2506 25836 2580
rect 26482 2506 26614 2580
rect 27260 2506 27392 2580
rect 28038 2506 28170 2580
rect 28816 2506 28948 2580
rect 29594 2506 29726 2580
rect 30372 2506 30504 2580
rect 31150 2506 31282 2580
rect 31928 2506 32060 2580
rect 32706 2506 32838 2580
rect 33484 2506 33616 2580
rect 34262 2506 34394 2580
rect 35040 2506 35172 2580
rect 35818 2506 35950 2580
rect 36596 2506 36728 2580
rect 37374 2506 37506 2580
rect 38152 2506 38284 2580
rect 38930 2506 39062 2580
rect 39708 2506 39840 2580
rect 40486 2506 40618 2580
rect 41264 2506 41396 2580
rect 42042 2506 42174 2580
rect 42820 2506 42952 2580
rect 43598 2506 43730 2580
rect 44376 2506 44508 2580
rect 45154 2506 45286 2580
rect 45932 2506 46064 2580
rect 46710 2506 46842 2580
rect 47488 2506 47620 2580
rect 48266 2506 48398 2580
rect 49044 2506 49176 2580
rect 49822 2506 49954 2580
rect 50600 2506 50732 2580
rect 51378 2506 51510 2580
rect 52156 2506 52288 2580
rect 52934 2506 53066 2580
rect 53712 2506 53844 2580
rect 54490 2506 54622 2580
rect 55268 2506 55400 2580
rect 56046 2506 56178 2580
rect 56824 2506 56956 2580
rect 57602 2506 57734 2580
rect 4132 2099 4264 2173
rect 5244 2099 5376 2173
rect 8036 548 8102 680
rect 8814 548 8880 680
rect 9592 548 9658 680
rect 10370 548 10436 680
rect 11148 548 11214 680
rect 11926 548 11992 680
rect 12704 548 12770 680
rect 13482 548 13548 680
rect 14260 548 14326 680
rect 15038 548 15104 680
rect 15816 548 15882 680
rect 16594 548 16660 680
rect 17372 548 17438 680
rect 18150 548 18216 680
rect 18928 548 18994 680
rect 19706 548 19772 680
rect 20484 548 20550 680
rect 21262 548 21328 680
rect 22040 548 22106 680
rect 22818 548 22884 680
rect 23596 548 23662 680
rect 24374 548 24440 680
rect 25152 548 25218 680
rect 25930 548 25996 680
rect 26708 548 26774 680
rect 27486 548 27552 680
rect 28264 548 28330 680
rect 29042 548 29108 680
rect 29820 548 29886 680
rect 30598 548 30664 680
rect 31376 548 31442 680
rect 32154 548 32220 680
rect 32932 548 32998 680
rect 33710 548 33776 680
rect 34488 548 34554 680
rect 35266 548 35332 680
rect 36044 548 36110 680
rect 36822 548 36888 680
rect 37600 548 37666 680
rect 38378 548 38444 680
rect 39156 548 39222 680
rect 39934 548 40000 680
rect 40712 548 40778 680
rect 41490 548 41556 680
rect 42268 548 42334 680
rect 43046 548 43112 680
rect 43824 548 43890 680
rect 44602 548 44668 680
rect 45380 548 45446 680
rect 46158 548 46224 680
rect 46936 548 47002 680
rect 47714 548 47780 680
rect 48492 548 48558 680
rect 49270 548 49336 680
rect 50048 548 50114 680
rect 50826 548 50892 680
rect 51604 548 51670 680
rect 52382 548 52448 680
rect 53160 548 53226 680
rect 53938 548 54004 680
rect 54716 548 54782 680
rect 55494 548 55560 680
rect 56272 548 56338 680
rect 57050 548 57116 680
rect 57828 548 57894 680
use contact_17  contact_17_0
timestamp 1644951705
transform 1 0 57960 0 1 1485
box 0 0 1 1
use contact_17  contact_17_1
timestamp 1644951705
transform 1 0 7486 0 1 5966
box 0 0 1 1
use contact_17  contact_17_2
timestamp 1644951705
transform 1 0 3586 0 1 3416
box 0 0 1 1
use contact_13  contact_13_0
timestamp 1644951705
transform 1 0 5898 0 1 4166
box 0 0 1 1
use contact_17  contact_17_3
timestamp 1644951705
transform 1 0 3586 0 1 4157
box 0 0 1 1
use contact_17  contact_17_4
timestamp 1644951705
transform 1 0 3494 0 1 3336
box 0 0 1 1
use contact_13  contact_13_1
timestamp 1644951705
transform 1 0 5898 0 1 5088
box 0 0 1 1
use contact_17  contact_17_5
timestamp 1644951705
transform 1 0 3494 0 1 5079
box 0 0 1 1
use contact_13  contact_13_2
timestamp 1644951705
transform 1 0 5898 0 1 3412
box 0 0 1 1
use contact_17  contact_17_6
timestamp 1644951705
transform 1 0 3310 0 1 3576
box 0 0 1 1
use contact_13  contact_13_3
timestamp 1644951705
transform 1 0 5898 0 1 2490
box 0 0 1 1
use contact_17  contact_17_7
timestamp 1644951705
transform 1 0 3310 0 1 2481
box 0 0 1 1
use hierarchical_predecode2x4_0  hierarchical_predecode2x4_0_0
timestamp 1644951705
transform 1 0 3762 0 1 2136
box 0 -37 2390 3389
use port_address  port_address_0
timestamp 1644951705
transform 1 0 0 0 1 6536
box 0 -42 7652 49258
use port_data  port_data_0
timestamp 1644951705
transform 1 0 7876 0 1 0
box 0 490 50570 6392
use replica_bitcell_array  replica_bitcell_array_0
timestamp 1644951705
transform 1 0 7876 0 1 6536
box 0 -42 49792 49322
<< labels >>
rlabel metal2 s 7504 0 7532 6116 4 w_en
rlabel metal2 s 6382 55738 6410 55766 4 wl_en
rlabel metal2 s 57978 0 58006 55900 4 p_en_bar
rlabel metal2 s 8460 6068 8514 6096 4 din0_0
rlabel metal2 s 11572 6068 11626 6096 4 din0_1
rlabel metal2 s 14684 6068 14738 6096 4 din0_2
rlabel metal2 s 17796 6068 17850 6096 4 din0_3
rlabel metal2 s 20908 6068 20962 6096 4 din0_4
rlabel metal2 s 24020 6068 24074 6096 4 din0_5
rlabel metal2 s 27132 6068 27186 6096 4 din0_6
rlabel metal2 s 30244 6068 30298 6096 4 din0_7
rlabel metal2 s 33356 6068 33410 6096 4 din0_8
rlabel metal2 s 36468 6068 36522 6096 4 din0_9
rlabel metal2 s 39580 6068 39634 6096 4 din0_10
rlabel metal2 s 42692 6068 42746 6096 4 din0_11
rlabel metal2 s 45804 6068 45858 6096 4 din0_12
rlabel metal2 s 48916 6068 48970 6096 4 din0_13
rlabel metal2 s 52028 6068 52082 6096 4 din0_14
rlabel metal2 s 55140 6068 55194 6096 4 din0_15
rlabel metal2 s 8194 4924 8222 5164 4 dout0_0
rlabel metal2 s 8209 5044 8209 5044 4 dout1_0
rlabel metal2 s 8466 4924 8494 5164 4 dout0_1
rlabel metal2 s 8481 5044 8481 5044 4 dout1_1
rlabel metal2 s 11306 4924 11334 5164 4 dout0_2
rlabel metal2 s 11321 5044 11321 5044 4 dout1_2
rlabel metal2 s 11578 4924 11606 5164 4 dout0_3
rlabel metal2 s 11593 5044 11593 5044 4 dout1_3
rlabel metal2 s 14418 4924 14446 5164 4 dout0_4
rlabel metal2 s 14433 5044 14433 5044 4 dout1_4
rlabel metal2 s 14690 4924 14718 5164 4 dout0_5
rlabel metal2 s 14705 5044 14705 5044 4 dout1_5
rlabel metal2 s 17530 4924 17558 5164 4 dout0_6
rlabel metal2 s 17545 5044 17545 5044 4 dout1_6
rlabel metal2 s 17802 4924 17830 5164 4 dout0_7
rlabel metal2 s 17817 5044 17817 5044 4 dout1_7
rlabel metal2 s 20642 4924 20670 5164 4 dout0_8
rlabel metal2 s 20657 5044 20657 5044 4 dout1_8
rlabel metal2 s 20914 4924 20942 5164 4 dout0_9
rlabel metal2 s 20929 5044 20929 5044 4 dout1_9
rlabel metal2 s 23754 4924 23782 5164 4 dout0_10
rlabel metal2 s 23769 5044 23769 5044 4 dout1_10
rlabel metal2 s 24026 4924 24054 5164 4 dout0_11
rlabel metal2 s 24041 5044 24041 5044 4 dout1_11
rlabel metal2 s 26866 4924 26894 5164 4 dout0_12
rlabel metal2 s 26881 5044 26881 5044 4 dout1_12
rlabel metal2 s 27138 4924 27166 5164 4 dout0_13
rlabel metal2 s 27153 5044 27153 5044 4 dout1_13
rlabel metal2 s 29978 4924 30006 5164 4 dout0_14
rlabel metal2 s 29993 5044 29993 5044 4 dout1_14
rlabel metal2 s 30250 4924 30278 5164 4 dout0_15
rlabel metal2 s 30265 5044 30265 5044 4 dout1_15
rlabel metal2 s 18 6536 46 37328 4 addr2
rlabel metal2 s 102 6536 130 37328 4 addr3
rlabel metal2 s 186 6536 214 37328 4 addr4
rlabel metal2 s 270 6536 298 37328 4 addr5
rlabel metal2 s 354 6536 382 37328 4 addr6
rlabel metal2 s 438 6536 466 37328 4 addr7
rlabel metal2 s 522 6536 550 37328 4 addr8
rlabel metal2 s 3874 2480 3926 2544 4 addr0
rlabel metal2 s 3998 3402 4050 3466 4 addr1
rlabel metal3 s 56272 548 56338 680 4 vdd
rlabel metal3 s 29820 548 29886 680 4 vdd
rlabel metal3 s 5980 51100 6112 51174 4 vdd
rlabel metal3 s 51604 548 51670 680 4 vdd
rlabel metal3 s 54742 4146 54874 4220 4 vdd
rlabel metal3 s 15816 548 15882 680 4 vdd
rlabel metal3 s 4132 2936 4264 3010 4 vdd
rlabel metal3 s 11926 548 11992 680 4 vdd
rlabel metal3 s 7520 51100 7652 51174 4 vdd
rlabel metal3 s 36822 548 36888 680 4 vdd
rlabel metal3 s 5980 14188 6112 14262 4 vdd
rlabel metal3 s 33476 5428 33542 5560 4 vdd
rlabel metal3 s 43824 548 43890 680 4 vdd
rlabel metal3 s 26708 548 26774 680 4 vdd
rlabel metal3 s 14804 5428 14870 5560 4 vdd
rlabel metal3 s 40712 548 40778 680 4 vdd
rlabel metal3 s 39934 548 40000 680 4 vdd
rlabel metal3 s 52382 548 52448 680 4 vdd
rlabel metal3 s 5980 17264 6112 17338 4 vdd
rlabel metal3 s 25152 548 25218 680 4 vdd
rlabel metal3 s 5980 48024 6112 48098 4 vdd
rlabel metal3 s 35266 548 35332 680 4 vdd
rlabel metal3 s 960 26510 1092 26584 4 vdd
rlabel metal3 s 7520 32644 7652 32718 4 vdd
rlabel metal3 s 2000 26510 2132 26584 4 vdd
rlabel metal3 s 2180 17274 2312 17348 4 vdd
rlabel metal3 s 17398 4146 17530 4220 4 vdd
rlabel metal3 s 24374 548 24440 680 4 vdd
rlabel metal3 s 5980 23416 6112 23490 4 vdd
rlabel metal3 s 5244 4612 5376 4686 4 vdd
rlabel metal3 s 24140 5428 24206 5560 4 vdd
rlabel metal3 s 33710 548 33776 680 4 vdd
rlabel metal3 s 30598 548 30664 680 4 vdd
rlabel metal3 s 960 29590 1092 29664 4 vdd
rlabel metal3 s 7520 29568 7652 29642 4 vdd
rlabel metal3 s 11148 548 11214 680 4 vdd
rlabel metal3 s 45380 548 45446 680 4 vdd
rlabel metal3 s 22040 548 22106 680 4 vdd
rlabel metal3 s 47714 548 47780 680 4 vdd
rlabel metal3 s 55014 4146 55146 4220 4 vdd
rlabel metal3 s 5980 35720 6112 35794 4 vdd
rlabel metal3 s 43046 548 43112 680 4 vdd
rlabel metal3 s 37600 548 37666 680 4 vdd
rlabel metal3 s 32154 548 32220 680 4 vdd
rlabel metal3 s 44602 548 44668 680 4 vdd
rlabel metal3 s 32932 548 32998 680 4 vdd
rlabel metal3 s 5980 54176 6112 54250 4 vdd
rlabel metal3 s 5980 8036 6112 8110 4 vdd
rlabel metal3 s 23596 548 23662 680 4 vdd
rlabel metal3 s 9592 548 9658 680 4 vdd
rlabel metal3 s 2180 20354 2312 20428 4 vdd
rlabel metal3 s 54716 548 54782 680 4 vdd
rlabel metal3 s 19706 548 19772 680 4 vdd
rlabel metal3 s 45678 4146 45810 4220 4 vdd
rlabel metal3 s 27252 5428 27318 5560 4 vdd
rlabel metal3 s 32958 4146 33090 4220 4 vdd
rlabel metal3 s 42268 548 42334 680 4 vdd
rlabel metal3 s 7520 44948 7652 45022 4 vdd
rlabel metal3 s 36342 4146 36474 4220 4 vdd
rlabel metal3 s 33230 4146 33362 4220 4 vdd
rlabel metal3 s 55494 548 55560 680 4 vdd
rlabel metal3 s 7520 8036 7652 8110 4 vdd
rlabel metal3 s 51630 4146 51762 4220 4 vdd
rlabel metal3 s 48518 4146 48650 4220 4 vdd
rlabel metal3 s 27006 4146 27138 4220 4 vdd
rlabel metal3 s 39700 5428 39766 5560 4 vdd
rlabel metal3 s 7520 41872 7652 41946 4 vdd
rlabel metal3 s 20510 4146 20642 4220 4 vdd
rlabel metal3 s 18150 548 18216 680 4 vdd
rlabel metal3 s 20484 548 20550 680 4 vdd
rlabel metal3 s 36044 548 36110 680 4 vdd
rlabel metal3 s 49270 548 49336 680 4 vdd
rlabel metal3 s 2000 29590 2132 29664 4 vdd
rlabel metal3 s 53938 548 54004 680 4 vdd
rlabel metal3 s 7520 54176 7652 54250 4 vdd
rlabel metal3 s 34488 548 34554 680 4 vdd
rlabel metal3 s 7520 20340 7652 20414 4 vdd
rlabel metal3 s 42294 4146 42426 4220 4 vdd
rlabel metal3 s 8334 4146 8466 4220 4 vdd
rlabel metal3 s 1308 20354 1440 20428 4 vdd
rlabel metal3 s 50048 548 50114 680 4 vdd
rlabel metal3 s 39454 4146 39586 4220 4 vdd
rlabel metal3 s 53160 548 53226 680 4 vdd
rlabel metal3 s 14558 4146 14690 4220 4 vdd
rlabel metal3 s 21262 548 21328 680 4 vdd
rlabel metal3 s 5980 41872 6112 41946 4 vdd
rlabel metal3 s 5244 2936 5376 3010 4 vdd
rlabel metal3 s 14260 548 14326 680 4 vdd
rlabel metal3 s 42812 5428 42878 5560 4 vdd
rlabel metal3 s 5980 44948 6112 45022 4 vdd
rlabel metal3 s 27486 548 27552 680 4 vdd
rlabel metal3 s 12704 548 12770 680 4 vdd
rlabel metal3 s 21028 5428 21094 5560 4 vdd
rlabel metal3 s 55260 5428 55326 5560 4 vdd
rlabel metal3 s 31376 548 31442 680 4 vdd
rlabel metal3 s 45406 4146 45538 4220 4 vdd
rlabel metal3 s 15038 548 15104 680 4 vdd
rlabel metal3 s 13482 548 13548 680 4 vdd
rlabel metal3 s 7520 38796 7652 38870 4 vdd
rlabel metal3 s 10370 548 10436 680 4 vdd
rlabel metal3 s 7520 35720 7652 35794 4 vdd
rlabel metal3 s 5980 38796 6112 38870 4 vdd
rlabel metal3 s 4132 4612 4264 4686 4 vdd
rlabel metal3 s 51902 4146 52034 4220 4 vdd
rlabel metal3 s 8580 5428 8646 5560 4 vdd
rlabel metal3 s 45924 5428 45990 5560 4 vdd
rlabel metal3 s 11174 4146 11306 4220 4 vdd
rlabel metal3 s 16594 548 16660 680 4 vdd
rlabel metal3 s 28264 548 28330 680 4 vdd
rlabel metal3 s 5980 26492 6112 26566 4 vdd
rlabel metal3 s 5980 20340 6112 20414 4 vdd
rlabel metal3 s 20782 4146 20914 4220 4 vdd
rlabel metal3 s 57050 548 57116 680 4 vdd
rlabel metal3 s 7520 11112 7652 11186 4 vdd
rlabel metal3 s 7520 17264 7652 17338 4 vdd
rlabel metal3 s 2000 32670 2132 32744 4 vdd
rlabel metal3 s 17670 4146 17802 4220 4 vdd
rlabel metal3 s 30118 4146 30250 4220 4 vdd
rlabel metal3 s 46936 548 47002 680 4 vdd
rlabel metal3 s 1308 17274 1440 17348 4 vdd
rlabel metal3 s 17372 548 17438 680 4 vdd
rlabel metal3 s 7520 23416 7652 23490 4 vdd
rlabel metal3 s 39156 548 39222 680 4 vdd
rlabel metal3 s 11446 4146 11578 4220 4 vdd
rlabel metal3 s 29846 4146 29978 4220 4 vdd
rlabel metal3 s 23622 4146 23754 4220 4 vdd
rlabel metal3 s 960 35750 1092 35824 4 vdd
rlabel metal3 s 41490 548 41556 680 4 vdd
rlabel metal3 s 5980 11112 6112 11186 4 vdd
rlabel metal3 s 17916 5428 17982 5560 4 vdd
rlabel metal3 s 29042 548 29108 680 4 vdd
rlabel metal3 s 7520 26492 7652 26566 4 vdd
rlabel metal3 s 1308 8038 1440 8112 4 vdd
rlabel metal3 s 23894 4146 24026 4220 4 vdd
rlabel metal3 s 960 32670 1092 32744 4 vdd
rlabel metal3 s 50826 548 50892 680 4 vdd
rlabel metal3 s 30364 5428 30430 5560 4 vdd
rlabel metal3 s 2180 11118 2312 11192 4 vdd
rlabel metal3 s 57828 548 57894 680 4 vdd
rlabel metal3 s 1308 11118 1440 11192 4 vdd
rlabel metal3 s 14286 4146 14418 4220 4 vdd
rlabel metal3 s 48492 548 48558 680 4 vdd
rlabel metal3 s 5980 29568 6112 29642 4 vdd
rlabel metal3 s 39182 4146 39314 4220 4 vdd
rlabel metal3 s 46158 548 46224 680 4 vdd
rlabel metal3 s 52148 5428 52214 5560 4 vdd
rlabel metal3 s 2000 35750 2132 35824 4 vdd
rlabel metal3 s 25930 548 25996 680 4 vdd
rlabel metal3 s 18928 548 18994 680 4 vdd
rlabel metal3 s 22818 548 22884 680 4 vdd
rlabel metal3 s 8036 548 8102 680 4 vdd
rlabel metal3 s 49036 5428 49102 5560 4 vdd
rlabel metal3 s 8814 548 8880 680 4 vdd
rlabel metal3 s 7520 48024 7652 48098 4 vdd
rlabel metal3 s 11692 5428 11758 5560 4 vdd
rlabel metal3 s 7520 14188 7652 14262 4 vdd
rlabel metal3 s 36070 4146 36202 4220 4 vdd
rlabel metal3 s 8062 4146 8194 4220 4 vdd
rlabel metal3 s 42566 4146 42698 4220 4 vdd
rlabel metal3 s 26734 4146 26866 4220 4 vdd
rlabel metal3 s 5980 32644 6112 32718 4 vdd
rlabel metal3 s 48790 4146 48922 4220 4 vdd
rlabel metal3 s 36588 5428 36654 5560 4 vdd
rlabel metal3 s 38378 548 38444 680 4 vdd
rlabel metal3 s 2180 8038 2312 8112 4 vdd
rlabel metal3 s 14804 6260 14870 6392 4 gnd
rlabel metal3 s 39182 5092 39314 5166 4 gnd
rlabel metal3 s 7520 9574 7652 9648 4 gnd
rlabel metal3 s 5980 18802 6112 18876 4 gnd
rlabel metal3 s 7520 28030 7652 28104 4 gnd
rlabel metal3 s 8062 5092 8194 5166 4 gnd
rlabel metal3 s 5980 28030 6112 28104 4 gnd
rlabel metal3 s 45924 6260 45990 6392 4 gnd
rlabel metal3 s 42294 5092 42426 5166 4 gnd
rlabel metal3 s 2000 28050 2132 28124 4 gnd
rlabel metal3 s 51902 5092 52034 5166 4 gnd
rlabel metal3 s 10922 2506 11054 2580 4 gnd
rlabel metal3 s 29594 2506 29726 2580 4 gnd
rlabel metal3 s 35040 2506 35172 2580 4 gnd
rlabel metal3 s 5980 9574 6112 9648 4 gnd
rlabel metal3 s 30364 6260 30430 6392 4 gnd
rlabel metal3 s 11446 5092 11578 5166 4 gnd
rlabel metal3 s 42812 6260 42878 6392 4 gnd
rlabel metal3 s 5980 49562 6112 49636 4 gnd
rlabel metal3 s 11174 5092 11306 5166 4 gnd
rlabel metal3 s 54490 2506 54622 2580 4 gnd
rlabel metal3 s 5244 2098 5376 2172 4 gnd
rlabel metal3 s 36070 5092 36202 5166 4 gnd
rlabel metal3 s 2180 15734 2312 15808 4 gnd
rlabel metal3 s 5244 5450 5376 5524 4 gnd
rlabel metal3 s 7520 37258 7652 37332 4 gnd
rlabel metal3 s 57602 2506 57734 2580 4 gnd
rlabel metal3 s 21028 6260 21094 6392 4 gnd
rlabel metal3 s 2180 6498 2312 6572 4 gnd
rlabel metal3 s 8334 5092 8466 5166 4 gnd
rlabel metal3 s 56046 2506 56178 2580 4 gnd
rlabel metal3 s 14812 2506 14944 2580 4 gnd
rlabel metal3 s 32706 2506 32838 2580 4 gnd
rlabel metal3 s 52934 2506 53066 2580 4 gnd
rlabel metal3 s 2180 12658 2312 12732 4 gnd
rlabel metal3 s 2180 18814 2312 18888 4 gnd
rlabel metal3 s 9366 2506 9498 2580 4 gnd
rlabel metal3 s 17924 2506 18056 2580 4 gnd
rlabel metal3 s 38930 2506 39062 2580 4 gnd
rlabel metal3 s 26734 5092 26866 5166 4 gnd
rlabel metal3 s 45154 2506 45286 2580 4 gnd
rlabel metal3 s 20510 5092 20642 5166 4 gnd
rlabel metal3 s 30372 2506 30504 2580 4 gnd
rlabel metal3 s 5980 12650 6112 12724 4 gnd
rlabel metal3 s 49036 6260 49102 6392 4 gnd
rlabel metal3 s 27260 2506 27392 2580 4 gnd
rlabel metal3 s 30118 5092 30250 5166 4 gnd
rlabel metal3 s 23622 5092 23754 5166 4 gnd
rlabel metal3 s 2000 34210 2132 34284 4 gnd
rlabel metal3 s 55014 5092 55146 5166 4 gnd
rlabel metal3 s 12478 2506 12610 2580 4 gnd
rlabel metal3 s 21814 2506 21946 2580 4 gnd
rlabel metal3 s 14558 5092 14690 5166 4 gnd
rlabel metal3 s 5980 37258 6112 37332 4 gnd
rlabel metal3 s 1308 18814 1440 18888 4 gnd
rlabel metal3 s 5980 24954 6112 25028 4 gnd
rlabel metal3 s 7520 49562 7652 49636 4 gnd
rlabel metal3 s 1308 15734 1440 15808 4 gnd
rlabel metal3 s 31150 2506 31282 2580 4 gnd
rlabel metal3 s 29846 5092 29978 5166 4 gnd
rlabel metal3 s 37374 2506 37506 2580 4 gnd
rlabel metal3 s 51378 2506 51510 2580 4 gnd
rlabel metal3 s 11692 6260 11758 6392 4 gnd
rlabel metal3 s 39700 6260 39766 6392 4 gnd
rlabel metal3 s 23894 5092 24026 5166 4 gnd
rlabel metal3 s 1308 9578 1440 9652 4 gnd
rlabel metal3 s 960 28050 1092 28124 4 gnd
rlabel metal3 s 48266 2506 48398 2580 4 gnd
rlabel metal3 s 53712 2506 53844 2580 4 gnd
rlabel metal3 s 5980 55714 6112 55788 4 gnd
rlabel metal3 s 20258 2506 20390 2580 4 gnd
rlabel metal3 s 33476 6260 33542 6392 4 gnd
rlabel metal3 s 14034 2506 14166 2580 4 gnd
rlabel metal3 s 15590 2506 15722 2580 4 gnd
rlabel metal3 s 20782 5092 20914 5166 4 gnd
rlabel metal3 s 17916 6260 17982 6392 4 gnd
rlabel metal3 s 5244 3774 5376 3848 4 gnd
rlabel metal3 s 13256 2506 13388 2580 4 gnd
rlabel metal3 s 24140 6260 24206 6392 4 gnd
rlabel metal3 s 39708 2506 39840 2580 4 gnd
rlabel metal3 s 4132 3774 4264 3848 4 gnd
rlabel metal3 s 21036 2506 21168 2580 4 gnd
rlabel metal3 s 40486 2506 40618 2580 4 gnd
rlabel metal3 s 7520 34182 7652 34256 4 gnd
rlabel metal3 s 17670 5092 17802 5166 4 gnd
rlabel metal3 s 7520 40334 7652 40408 4 gnd
rlabel metal3 s 7520 18802 7652 18876 4 gnd
rlabel metal3 s 42566 5092 42698 5166 4 gnd
rlabel metal3 s 4132 5450 4264 5524 4 gnd
rlabel metal3 s 960 31130 1092 31204 4 gnd
rlabel metal3 s 7520 6498 7652 6572 4 gnd
rlabel metal3 s 33230 5092 33362 5166 4 gnd
rlabel metal3 s 54742 5092 54874 5166 4 gnd
rlabel metal3 s 42820 2506 42952 2580 4 gnd
rlabel metal3 s 47488 2506 47620 2580 4 gnd
rlabel metal3 s 38152 2506 38284 2580 4 gnd
rlabel metal3 s 14286 5092 14418 5166 4 gnd
rlabel metal3 s 7520 55714 7652 55788 4 gnd
rlabel metal3 s 52156 2506 52288 2580 4 gnd
rlabel metal3 s 52148 6260 52214 6392 4 gnd
rlabel metal3 s 34262 2506 34394 2580 4 gnd
rlabel metal3 s 48790 5092 48922 5166 4 gnd
rlabel metal3 s 27252 6260 27318 6392 4 gnd
rlabel metal3 s 45406 5092 45538 5166 4 gnd
rlabel metal3 s 1308 21894 1440 21968 4 gnd
rlabel metal3 s 55268 2506 55400 2580 4 gnd
rlabel metal3 s 36596 2506 36728 2580 4 gnd
rlabel metal3 s 7520 43410 7652 43484 4 gnd
rlabel metal3 s 17398 5092 17530 5166 4 gnd
rlabel metal3 s 45678 5092 45810 5166 4 gnd
rlabel metal3 s 44376 2506 44508 2580 4 gnd
rlabel metal3 s 36342 5092 36474 5166 4 gnd
rlabel metal3 s 22592 2506 22724 2580 4 gnd
rlabel metal3 s 32958 5092 33090 5166 4 gnd
rlabel metal3 s 36588 6260 36654 6392 4 gnd
rlabel metal3 s 5980 31106 6112 31180 4 gnd
rlabel metal3 s 8580 6260 8646 6392 4 gnd
rlabel metal3 s 7520 46486 7652 46560 4 gnd
rlabel metal3 s 50600 2506 50732 2580 4 gnd
rlabel metal3 s 43598 2506 43730 2580 4 gnd
rlabel metal3 s 5980 46486 6112 46560 4 gnd
rlabel metal3 s 26482 2506 26614 2580 4 gnd
rlabel metal3 s 960 34210 1092 34284 4 gnd
rlabel metal3 s 48518 5092 48650 5166 4 gnd
rlabel metal3 s 5980 43410 6112 43484 4 gnd
rlabel metal3 s 49044 2506 49176 2580 4 gnd
rlabel metal3 s 17146 2506 17278 2580 4 gnd
rlabel metal3 s 33484 2506 33616 2580 4 gnd
rlabel metal3 s 45932 2506 46064 2580 4 gnd
rlabel metal3 s 31928 2506 32060 2580 4 gnd
rlabel metal3 s 35818 2506 35950 2580 4 gnd
rlabel metal3 s 960 37290 1092 37364 4 gnd
rlabel metal3 s 2000 37290 2132 37364 4 gnd
rlabel metal3 s 55260 6260 55326 6392 4 gnd
rlabel metal3 s 28038 2506 28170 2580 4 gnd
rlabel metal3 s 46710 2506 46842 2580 4 gnd
rlabel metal3 s 960 24970 1092 25044 4 gnd
rlabel metal3 s 2180 9578 2312 9652 4 gnd
rlabel metal3 s 2000 24970 2132 25044 4 gnd
rlabel metal3 s 27006 5092 27138 5166 4 gnd
rlabel metal3 s 16368 2506 16500 2580 4 gnd
rlabel metal3 s 4132 2098 4264 2172 4 gnd
rlabel metal3 s 24148 2506 24280 2580 4 gnd
rlabel metal3 s 11700 2506 11832 2580 4 gnd
rlabel metal3 s 18702 2506 18834 2580 4 gnd
rlabel metal3 s 41264 2506 41396 2580 4 gnd
rlabel metal3 s 2000 31130 2132 31204 4 gnd
rlabel metal3 s 24926 2506 25058 2580 4 gnd
rlabel metal3 s 28816 2506 28948 2580 4 gnd
rlabel metal3 s 25704 2506 25836 2580 4 gnd
rlabel metal3 s 7520 31106 7652 31180 4 gnd
rlabel metal3 s 7520 12650 7652 12724 4 gnd
rlabel metal3 s 7520 24954 7652 25028 4 gnd
rlabel metal3 s 7520 21878 7652 21952 4 gnd
rlabel metal3 s 5980 6498 6112 6572 4 gnd
rlabel metal3 s 1308 6498 1440 6572 4 gnd
rlabel metal3 s 5980 21878 6112 21952 4 gnd
rlabel metal3 s 7520 52638 7652 52712 4 gnd
rlabel metal3 s 56824 2506 56956 2580 4 gnd
rlabel metal3 s 39454 5092 39586 5166 4 gnd
rlabel metal3 s 42042 2506 42174 2580 4 gnd
rlabel metal3 s 10144 2506 10276 2580 4 gnd
rlabel metal3 s 49822 2506 49954 2580 4 gnd
rlabel metal3 s 7520 15726 7652 15800 4 gnd
rlabel metal3 s 23370 2506 23502 2580 4 gnd
rlabel metal3 s 5980 15726 6112 15800 4 gnd
rlabel metal3 s 51630 5092 51762 5166 4 gnd
rlabel metal3 s 8588 2506 8720 2580 4 gnd
rlabel metal3 s 2180 21894 2312 21968 4 gnd
rlabel metal3 s 5980 40334 6112 40408 4 gnd
rlabel metal3 s 1308 12658 1440 12732 4 gnd
rlabel metal3 s 5980 52638 6112 52712 4 gnd
rlabel metal3 s 5980 34182 6112 34256 4 gnd
rlabel metal3 s 19480 2506 19612 2580 4 gnd
<< properties >>
string FIXED_BBOX 0 0 58530 55900
string GDS_FILE sram_0rw2r1w_16_128_sky130A.gds
string GDS_END 308464
string GDS_START 201826
<< end >>
