magic
tech sky130A
magscale 1 2
timestamp 1643593061
<< checkpaint >>
rect -1260 -1268 2038 2312
<< nwell >>
rect 0 0 778 1038
<< nsubdiff >>
rect 168 945 218 969
rect 168 911 176 945
rect 210 911 218 945
rect 168 887 218 911
<< nsubdiffcont >>
rect 176 911 210 945
<< poly >>
rect 128 502 258 532
rect 128 416 158 502
rect 128 58 158 112
rect 125 42 191 58
rect 125 8 141 42
rect 175 8 191 42
rect 125 -8 191 8
<< polycont >>
rect 141 8 175 42
<< locali >>
rect 176 945 210 961
rect 176 895 210 911
rect 125 42 191 58
rect 125 8 141 42
rect 175 8 191 42
rect 125 -8 191 8
<< viali >>
rect 176 911 210 945
rect 76 667 110 701
rect 176 667 210 701
rect 276 667 310 701
rect 76 247 110 281
rect 176 247 210 281
rect 141 8 175 42
<< metal1 >>
rect 0 1024 778 1052
rect 179 960 207 1024
rect 167 954 219 960
rect 161 902 167 954
rect 219 902 225 954
rect 167 896 219 902
rect 67 710 119 716
rect 179 713 207 896
rect 67 652 119 658
rect 170 701 216 713
rect 170 667 176 701
rect 210 667 216 701
rect 170 655 216 667
rect 267 710 319 716
rect 267 652 319 658
rect 67 290 119 296
rect 67 232 119 238
rect 167 290 219 296
rect 167 232 219 238
rect 129 42 187 48
rect 129 39 141 42
rect 0 11 141 39
rect 129 8 141 11
rect 175 39 187 42
rect 175 11 778 39
rect 175 8 187 11
rect 129 2 187 8
<< via1 >>
rect 167 945 219 954
rect 167 911 176 945
rect 176 911 210 945
rect 210 911 219 945
rect 167 902 219 911
rect 67 701 119 710
rect 67 667 76 701
rect 76 667 110 701
rect 110 667 119 701
rect 67 658 119 667
rect 267 701 319 710
rect 267 667 276 701
rect 276 667 310 701
rect 310 667 319 701
rect 267 658 319 667
rect 67 281 119 290
rect 67 247 76 281
rect 76 247 110 281
rect 110 247 119 281
rect 67 238 119 247
rect 167 281 219 290
rect 167 247 176 281
rect 176 247 210 281
rect 210 247 219 281
rect 167 238 219 247
<< metal2 >>
rect 70 710 98 1038
rect 532 717 560 1038
rect 293 710 560 717
rect 319 658 560 710
rect 70 290 98 658
rect 293 651 560 658
rect 532 297 560 651
rect 193 290 560 297
rect 219 238 560 290
rect 70 0 98 238
rect 193 231 560 238
rect 532 0 560 231
<< via2 >>
rect 165 954 221 956
rect 165 902 167 954
rect 167 902 219 954
rect 219 902 221 954
rect 165 900 221 902
<< metal3 >>
rect 163 956 223 958
rect 163 900 165 956
rect 221 900 223 956
rect 163 898 223 900
use contact_22  contact_22_0
timestamp 1643593061
transform 1 0 267 0 1 652
box 0 0 1 1
use contact_24  contact_24_0
timestamp 1643593061
transform 1 0 270 0 1 655
box 0 0 1 1
use contact_22  contact_22_1
timestamp 1643593061
transform 1 0 67 0 1 652
box 0 0 1 1
use contact_24  contact_24_1
timestamp 1643593061
transform 1 0 70 0 1 655
box 0 0 1 1
use contact_22  contact_22_2
timestamp 1643593061
transform 1 0 167 0 1 232
box 0 0 1 1
use contact_24  contact_24_2
timestamp 1643593061
transform 1 0 170 0 1 235
box 0 0 1 1
use contact_22  contact_22_3
timestamp 1643593061
transform 1 0 67 0 1 232
box 0 0 1 1
use contact_24  contact_24_3
timestamp 1643593061
transform 1 0 70 0 1 235
box 0 0 1 1
use contact_24  contact_24_4
timestamp 1643593061
transform 1 0 170 0 1 655
box 0 0 1 1
use contact_23  contact_23_0
timestamp 1643593061
transform 1 0 163 0 1 898
box 0 0 1 1
use contact_22  contact_22_4
timestamp 1643593061
transform 1 0 167 0 1 896
box 0 0 1 1
use contact_17  contact_17_0
timestamp 1643593061
transform 1 0 161 0 1 902
box 0 0 1 1
use contact_13  contact_13_0
timestamp 1643593061
transform 1 0 164 0 1 905
box 0 0 1 1
use contact_21  contact_21_0
timestamp 1643593061
transform 1 0 168 0 1 887
box 0 0 1 1
use contact_13  contact_13_1
timestamp 1643593061
transform 1 0 129 0 1 2
box 0 0 1 1
use contact_12  contact_12_0
timestamp 1643593061
transform 1 0 125 0 1 -8
box 0 0 1 1
use pmos_m1_w1_260_sli_dli  pmos_m1_w1_260_sli_dli_0
timestamp 1643593061
transform 1 0 168 0 1 558
box -59 -54 209 306
use pmos_m1_w1_260_sli_dli  pmos_m1_w1_260_sli_dli_1
timestamp 1643593061
transform 1 0 68 0 1 558
box -59 -54 209 306
use pmos_m1_w1_260_sli_dli  pmos_m1_w1_260_sli_dli_2
timestamp 1643593061
transform 1 0 68 0 1 138
box -59 -54 209 306
<< labels >>
rlabel metal1 s 0 10 778 38 4 en_bar
rlabel metal3 s 162 898 222 958 4 vdd
rlabel metal2 s 70 0 98 1038 4 rbl0
rlabel metal2 s 532 0 560 1038 4 rbl1
<< properties >>
string FIXED_BBOX 115 -18 201 0
string GDS_FILE sram_0rw2r1w_2_16_sky130A.gds
string GDS_END 247520
string GDS_START 244566
<< end >>
