magic
tech sky130A
magscale 1 2
timestamp 1643678851
<< checkpaint >>
rect -1260 -1302 2464 2876
<< nwell >>
rect 0 976 1204 1616
<< pwell >>
rect 184 -42 256 42
rect 438 -42 510 42
rect 694 -42 766 42
rect 948 -42 1020 42
<< nmos >>
rect 94 308 124 418
rect 190 308 220 418
rect 286 308 316 418
rect 382 308 412 418
rect 586 308 616 418
rect 682 308 712 418
rect 784 308 814 392
rect 984 308 1014 392
rect 1080 308 1110 392
<< pmos >>
rect 94 1012 124 1096
rect 190 1012 220 1096
rect 286 1012 316 1096
rect 382 1012 412 1096
rect 586 1012 616 1096
rect 682 1012 712 1096
rect 784 1012 814 1282
rect 984 1012 1014 1282
rect 1080 1012 1110 1282
<< ndiff >>
rect 36 382 94 418
rect 36 348 44 382
rect 78 348 94 382
rect 36 308 94 348
rect 124 308 190 418
rect 220 382 286 418
rect 220 348 236 382
rect 270 348 286 382
rect 220 308 286 348
rect 316 308 382 418
rect 412 382 470 418
rect 412 348 428 382
rect 462 348 470 382
rect 412 308 470 348
rect 528 382 586 418
rect 528 348 536 382
rect 570 348 586 382
rect 528 308 586 348
rect 616 308 682 418
rect 712 392 768 418
rect 712 382 784 392
rect 712 348 728 382
rect 762 348 784 382
rect 712 308 784 348
rect 814 368 872 392
rect 814 334 830 368
rect 864 334 872 368
rect 814 308 872 334
rect 926 368 984 392
rect 926 334 934 368
rect 968 334 984 368
rect 926 308 984 334
rect 1014 368 1080 392
rect 1014 334 1030 368
rect 1064 334 1080 368
rect 1014 308 1080 334
rect 1110 368 1168 392
rect 1110 334 1126 368
rect 1160 334 1168 368
rect 1110 308 1168 334
<< pdiff >>
rect 728 1250 784 1282
rect 728 1216 736 1250
rect 770 1216 784 1250
rect 728 1166 784 1216
rect 728 1132 736 1166
rect 770 1132 784 1166
rect 728 1096 784 1132
rect 36 1070 94 1096
rect 36 1036 44 1070
rect 78 1036 94 1070
rect 36 1012 94 1036
rect 124 1070 190 1096
rect 124 1036 140 1070
rect 174 1036 190 1070
rect 124 1012 190 1036
rect 220 1070 286 1096
rect 220 1036 236 1070
rect 270 1036 286 1070
rect 220 1012 286 1036
rect 316 1070 382 1096
rect 316 1036 332 1070
rect 366 1036 382 1070
rect 316 1012 382 1036
rect 412 1070 470 1096
rect 412 1036 428 1070
rect 462 1036 470 1070
rect 412 1012 470 1036
rect 528 1070 586 1096
rect 528 1036 536 1070
rect 570 1036 586 1070
rect 528 1012 586 1036
rect 616 1068 682 1096
rect 616 1034 632 1068
rect 666 1034 682 1068
rect 616 1012 682 1034
rect 712 1068 784 1096
rect 712 1034 732 1068
rect 766 1034 784 1068
rect 712 1012 784 1034
rect 814 1250 872 1282
rect 814 1216 830 1250
rect 864 1216 872 1250
rect 814 1166 872 1216
rect 814 1132 830 1166
rect 864 1132 872 1166
rect 814 1080 872 1132
rect 814 1046 830 1080
rect 864 1046 872 1080
rect 814 1012 872 1046
rect 926 1250 984 1282
rect 926 1216 934 1250
rect 968 1216 984 1250
rect 926 1166 984 1216
rect 926 1132 934 1166
rect 968 1132 984 1166
rect 926 1080 984 1132
rect 926 1046 934 1080
rect 968 1046 984 1080
rect 926 1012 984 1046
rect 1014 1250 1080 1282
rect 1014 1216 1030 1250
rect 1064 1216 1080 1250
rect 1014 1166 1080 1216
rect 1014 1132 1030 1166
rect 1064 1132 1080 1166
rect 1014 1080 1080 1132
rect 1014 1046 1030 1080
rect 1064 1046 1080 1080
rect 1014 1012 1080 1046
rect 1110 1250 1168 1282
rect 1110 1216 1126 1250
rect 1160 1216 1168 1250
rect 1110 1166 1168 1216
rect 1110 1132 1126 1166
rect 1160 1132 1168 1166
rect 1110 1080 1168 1132
rect 1110 1046 1126 1080
rect 1160 1046 1168 1080
rect 1110 1012 1168 1046
<< ndiffc >>
rect 44 348 78 382
rect 236 348 270 382
rect 428 348 462 382
rect 536 348 570 382
rect 728 348 762 382
rect 830 334 864 368
rect 934 334 968 368
rect 1030 334 1064 368
rect 1126 334 1160 368
<< pdiffc >>
rect 736 1216 770 1250
rect 736 1132 770 1166
rect 44 1036 78 1070
rect 140 1036 174 1070
rect 236 1036 270 1070
rect 332 1036 366 1070
rect 428 1036 462 1070
rect 536 1036 570 1070
rect 632 1034 666 1068
rect 732 1034 766 1068
rect 830 1216 864 1250
rect 830 1132 864 1166
rect 830 1046 864 1080
rect 934 1216 968 1250
rect 934 1132 968 1166
rect 934 1046 968 1080
rect 1030 1216 1064 1250
rect 1030 1132 1064 1166
rect 1030 1046 1064 1080
rect 1126 1216 1160 1250
rect 1126 1132 1160 1166
rect 1126 1046 1160 1080
<< psubdiff >>
rect 184 17 256 42
rect 184 -17 203 17
rect 237 -17 256 17
rect 184 -42 256 -17
rect 438 17 510 42
rect 438 -17 457 17
rect 491 -17 510 17
rect 438 -42 510 -17
rect 694 17 766 42
rect 694 -17 713 17
rect 747 -17 766 17
rect 694 -42 766 -17
rect 948 17 1020 42
rect 948 -17 966 17
rect 1000 -17 1020 17
rect 948 -42 1020 -17
<< nsubdiff >>
rect 184 1555 256 1580
rect 184 1521 203 1555
rect 237 1521 256 1555
rect 184 1496 256 1521
rect 438 1555 510 1580
rect 438 1521 457 1555
rect 491 1521 510 1555
rect 438 1496 510 1521
rect 694 1555 766 1580
rect 694 1521 713 1555
rect 747 1521 766 1555
rect 694 1496 766 1521
rect 948 1555 1020 1580
rect 948 1521 967 1555
rect 1001 1521 1020 1555
rect 948 1496 1020 1521
<< psubdiffcont >>
rect 203 -17 237 17
rect 457 -17 491 17
rect 713 -17 747 17
rect 966 -17 1000 17
<< nsubdiffcont >>
rect 203 1521 237 1555
rect 457 1521 491 1555
rect 713 1521 747 1555
rect 967 1521 1001 1555
<< poly >>
rect 784 1282 814 1308
rect 984 1282 1014 1308
rect 1080 1282 1110 1308
rect 94 1096 124 1122
rect 190 1096 220 1122
rect 286 1096 316 1122
rect 382 1096 412 1122
rect 586 1096 616 1122
rect 682 1096 712 1122
rect 94 914 124 1012
rect 70 898 124 914
rect 70 864 80 898
rect 114 864 124 898
rect 70 848 124 864
rect 190 858 220 1012
rect 94 418 124 848
rect 166 842 220 858
rect 166 808 176 842
rect 210 808 220 842
rect 166 792 220 808
rect 286 802 316 1012
rect 190 418 220 792
rect 262 786 316 802
rect 262 752 272 786
rect 306 752 316 786
rect 262 736 316 752
rect 382 746 412 1012
rect 286 418 316 736
rect 358 730 412 746
rect 358 696 368 730
rect 402 696 412 730
rect 358 680 412 696
rect 382 418 412 680
rect 586 638 616 1012
rect 562 622 616 638
rect 562 588 572 622
rect 606 588 616 622
rect 562 572 616 588
rect 682 582 712 1012
rect 784 700 814 1012
rect 760 684 814 700
rect 760 650 770 684
rect 804 650 814 684
rect 760 634 814 650
rect 586 418 616 572
rect 658 566 712 582
rect 658 532 668 566
rect 702 532 712 566
rect 658 516 712 532
rect 682 418 712 516
rect 784 392 814 634
rect 984 786 1014 1012
rect 1080 914 1110 1012
rect 1056 898 1110 914
rect 1056 864 1066 898
rect 1100 864 1110 898
rect 1056 848 1110 864
rect 984 770 1038 786
rect 984 736 994 770
rect 1028 736 1038 770
rect 984 720 1038 736
rect 984 392 1014 720
rect 1080 392 1110 848
rect 94 282 124 308
rect 190 282 220 308
rect 286 282 316 308
rect 382 282 412 308
rect 586 282 616 308
rect 682 282 712 308
rect 784 282 814 308
rect 984 282 1014 308
rect 1080 282 1110 308
<< polycont >>
rect 80 864 114 898
rect 176 808 210 842
rect 272 752 306 786
rect 368 696 402 730
rect 572 588 606 622
rect 770 650 804 684
rect 668 532 702 566
rect 1066 864 1100 898
rect 994 736 1028 770
<< locali >>
rect 44 1555 1160 1572
rect 44 1521 203 1555
rect 237 1521 457 1555
rect 491 1521 713 1555
rect 747 1521 967 1555
rect 1001 1521 1160 1555
rect 44 1504 1160 1521
rect 44 1096 78 1504
rect 236 1096 270 1504
rect 428 1096 462 1504
rect 536 1096 570 1504
rect 736 1282 770 1504
rect 1030 1282 1064 1504
rect 728 1250 774 1282
rect 728 1216 736 1250
rect 770 1216 774 1250
rect 728 1166 774 1216
rect 728 1132 736 1166
rect 770 1132 774 1166
rect 728 1096 774 1132
rect 36 1070 84 1096
rect 36 1036 44 1070
rect 78 1036 84 1070
rect 36 1012 84 1036
rect 134 1070 180 1096
rect 134 1036 140 1070
rect 174 1036 180 1070
rect 134 1012 180 1036
rect 230 1070 276 1096
rect 230 1036 236 1070
rect 270 1036 276 1070
rect 230 1012 276 1036
rect 326 1070 372 1096
rect 326 1036 332 1070
rect 366 1036 372 1070
rect 326 1012 372 1036
rect 422 1070 470 1096
rect 422 1036 428 1070
rect 462 1036 470 1070
rect 422 1012 470 1036
rect 528 1070 576 1096
rect 528 1036 536 1070
rect 570 1036 576 1070
rect 528 1012 576 1036
rect 626 1068 672 1096
rect 626 1034 632 1068
rect 666 1034 672 1068
rect 626 1012 672 1034
rect 722 1068 774 1096
rect 722 1034 732 1068
rect 766 1034 774 1068
rect 722 1012 774 1034
rect 824 1250 872 1282
rect 824 1216 830 1250
rect 864 1216 872 1250
rect 824 1166 872 1216
rect 824 1132 830 1166
rect 864 1132 872 1166
rect 824 1080 872 1132
rect 824 1046 830 1080
rect 864 1046 872 1080
rect 824 1012 872 1046
rect 338 978 372 1012
rect 338 944 538 978
rect 80 898 114 914
rect 80 848 114 864
rect 176 842 210 858
rect 464 808 470 842
rect 176 792 210 808
rect 272 786 306 802
rect 272 736 306 752
rect 368 730 402 746
rect 368 680 402 696
rect 436 646 470 808
rect 50 612 470 646
rect 504 806 538 944
rect 50 418 84 612
rect 504 578 538 772
rect 632 752 666 1012
rect 632 718 804 752
rect 760 684 804 718
rect 760 666 770 684
rect 436 544 538 578
rect 572 622 606 638
rect 770 634 804 650
rect 572 572 606 588
rect 838 596 872 1012
rect 668 566 702 582
rect 436 418 470 544
rect 668 516 702 532
rect 36 382 84 418
rect 36 348 44 382
rect 78 348 84 382
rect 36 308 84 348
rect 230 382 276 418
rect 230 348 236 382
rect 270 348 276 382
rect 230 308 276 348
rect 422 382 470 418
rect 422 348 428 382
rect 462 348 470 382
rect 422 308 470 348
rect 528 382 576 418
rect 528 348 536 382
rect 570 348 576 382
rect 528 308 576 348
rect 722 382 768 418
rect 838 392 872 562
rect 722 348 728 382
rect 762 348 768 382
rect 722 308 768 348
rect 824 368 872 392
rect 824 334 830 368
rect 864 334 872 368
rect 824 308 872 334
rect 926 1250 974 1282
rect 926 1216 934 1250
rect 968 1216 974 1250
rect 926 1166 974 1216
rect 926 1132 934 1166
rect 968 1132 974 1166
rect 926 1080 974 1132
rect 926 1046 934 1080
rect 968 1046 974 1080
rect 926 1012 974 1046
rect 1024 1250 1070 1282
rect 1024 1216 1030 1250
rect 1064 1216 1070 1250
rect 1024 1166 1070 1216
rect 1024 1132 1030 1166
rect 1064 1132 1070 1166
rect 1024 1080 1070 1132
rect 1024 1046 1030 1080
rect 1064 1046 1070 1080
rect 1024 1012 1070 1046
rect 1120 1250 1168 1282
rect 1120 1216 1126 1250
rect 1160 1216 1168 1250
rect 1120 1166 1168 1216
rect 1120 1132 1126 1166
rect 1160 1132 1168 1166
rect 1120 1080 1168 1132
rect 1120 1046 1126 1080
rect 1160 1046 1168 1080
rect 1120 1026 1168 1046
rect 1120 1012 1134 1026
rect 926 684 960 1012
rect 1066 898 1100 914
rect 1066 848 1100 864
rect 994 770 1028 786
rect 994 720 1028 736
rect 926 392 960 650
rect 1134 392 1168 992
rect 926 368 974 392
rect 926 334 934 368
rect 968 334 974 368
rect 926 308 974 334
rect 1024 368 1070 392
rect 1024 334 1030 368
rect 1064 334 1070 368
rect 1024 308 1070 334
rect 1120 368 1168 392
rect 1120 334 1126 368
rect 1160 334 1168 368
rect 1120 308 1168 334
rect 236 34 270 308
rect 728 34 762 308
rect 1030 34 1064 308
rect 138 17 1064 34
rect 138 -17 203 17
rect 237 -17 457 17
rect 491 -17 713 17
rect 747 -17 966 17
rect 1000 -17 1064 17
rect 138 -34 1064 -17
<< viali >>
rect 203 1521 237 1555
rect 457 1521 491 1555
rect 713 1521 747 1555
rect 967 1521 1001 1555
rect 140 1036 174 1070
rect 80 864 114 898
rect 176 808 210 842
rect 430 808 464 842
rect 272 752 306 786
rect 368 696 402 730
rect 504 772 538 806
rect 770 650 804 684
rect 572 588 606 622
rect 668 532 702 566
rect 838 562 872 596
rect 536 348 570 382
rect 1134 992 1168 1026
rect 1066 864 1100 898
rect 994 736 1028 770
rect 926 650 960 684
rect 203 -17 237 17
rect 457 -17 491 17
rect 713 -17 747 17
rect 966 -17 1000 17
<< metal1 >>
rect 0 1555 1204 1568
rect 0 1521 203 1555
rect 237 1521 457 1555
rect 491 1521 713 1555
rect 747 1521 967 1555
rect 1001 1521 1204 1555
rect 0 1508 1204 1521
rect 134 1070 180 1082
rect 134 1036 140 1070
rect 174 1052 180 1070
rect 174 1036 476 1052
rect 134 1024 476 1036
rect 448 950 476 1024
rect 1128 1032 1174 1038
rect 1128 1026 1204 1032
rect 1128 992 1134 1026
rect 1168 1004 1204 1026
rect 1168 992 1174 1004
rect 1128 980 1174 992
rect 442 922 1106 950
rect 72 898 126 912
rect 72 876 80 898
rect 56 864 80 876
rect 114 864 126 898
rect 56 848 126 864
rect 168 848 222 856
rect 442 854 470 922
rect 220 796 222 848
rect 424 842 470 854
rect 1058 898 1106 922
rect 1058 864 1066 898
rect 1100 864 1106 898
rect 1058 850 1106 864
rect 424 808 430 842
rect 464 808 470 842
rect 168 794 222 796
rect 168 790 220 794
rect 264 786 318 800
rect 424 796 470 808
rect 498 806 544 818
rect 264 766 272 786
rect 262 752 272 766
rect 306 752 318 786
rect 498 772 504 806
rect 538 788 544 806
rect 538 772 1034 788
rect 498 770 1034 772
rect 498 760 994 770
rect 262 730 318 752
rect 234 702 318 730
rect 360 738 414 744
rect 412 686 414 738
rect 988 736 994 760
rect 1028 736 1034 770
rect 988 724 1034 736
rect 1080 778 1204 806
rect 360 682 414 686
rect 742 684 812 698
rect 360 680 412 682
rect 742 650 770 684
rect 804 650 812 684
rect 742 638 812 650
rect 920 686 966 696
rect 1080 686 1108 778
rect 920 684 1108 686
rect 920 650 926 684
rect 960 658 1108 684
rect 960 650 966 658
rect 920 638 966 650
rect 1136 652 1204 680
rect 564 622 618 636
rect 564 610 572 622
rect 536 588 572 610
rect 606 588 618 622
rect 536 582 618 588
rect 564 574 618 582
rect 660 574 714 580
rect 712 522 714 574
rect 660 518 714 522
rect 660 516 712 518
rect 742 394 770 638
rect 1136 608 1164 652
rect 832 596 1164 608
rect 832 562 838 596
rect 872 580 1164 596
rect 872 562 878 580
rect 832 550 878 562
rect 530 382 770 394
rect 530 348 536 382
rect 570 366 770 382
rect 570 348 576 366
rect 530 336 576 348
rect 0 17 1204 30
rect 0 -17 203 17
rect 237 -17 457 17
rect 491 -17 713 17
rect 747 -17 966 17
rect 1000 -17 1204 17
rect 0 -30 1204 -17
<< via1 >>
rect 168 842 220 848
rect 168 808 176 842
rect 176 808 210 842
rect 210 808 220 842
rect 168 796 220 808
rect 360 730 412 738
rect 360 696 368 730
rect 368 696 402 730
rect 402 696 412 730
rect 360 686 412 696
rect 660 566 712 574
rect 660 532 668 566
rect 668 532 702 566
rect 702 532 712 566
rect 660 522 712 532
<< metal2 >>
rect 168 848 220 854
rect 168 790 220 796
rect 168 708 196 790
rect 360 738 412 744
rect 0 686 360 708
rect 0 680 412 686
rect 360 544 388 680
rect 660 574 712 580
rect 360 522 660 544
rect 360 516 712 522
<< labels >>
rlabel mvpsubdiff s 156 356 156 356 4 net1
rlabel mvpsubdiff s 348 354 348 354 4 net3
rlabel mvpsubdiff s 652 348 652 348 4 net5
rlabel metal1 s 756 562 756 562 4 net6
rlabel metal1 s 540 936 540 936 4 net2
rlabel metal1 s 560 774 560 774 4 net4
rlabel metal1 s 56 848 126 876 4 A0
port 1 nsew
rlabel metal1 s 0 1508 1204 1568 4 vdd
port 2 nsew
rlabel metal1 s 0 -30 1204 30 4 gnd
port 3 nsew
rlabel metal2 s 0 680 412 708 4 wl_en
port 4 nsew
rlabel metal1 s 234 702 318 730 4 A1
port 5 nsew
rlabel metal1 s 536 582 618 610 4 A2
port 6 nsew
rlabel metal1 s 1080 778 1204 806 4 rwl0
port 7 nsew
rlabel metal1 s 1136 652 1204 680 4 wwl0
port 8 nsew
rlabel metal1 s 1128 1004 1204 1032 4 rwl1
port 9 nsew
rlabel metal1 s 91 862 91 862 4 A0
rlabel metal1 s 276 716 276 716 4 A1
rlabel metal1 s 577 596 577 596 4 A2
rlabel metal2 s 206 694 206 694 4 wl_en
rlabel metal1 s 1142 792 1142 792 4 rwl0
rlabel metal1 s 1166 1018 1166 1018 4 rwl1
rlabel metal1 s 1170 666 1170 666 4 wwl0
rlabel metal1 s 602 1538 602 1538 4 vdd
rlabel metal1 s 602 0 602 0 4 gnd
<< properties >>
string FIXED_BBOX 0 -42 1204 1538
string GDS_FILE sram_0rw2r1w_16_128_sky130A.gds
string GDS_END 1983322
string GDS_START 1964078
<< end >>
