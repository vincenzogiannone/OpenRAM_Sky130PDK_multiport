magic
tech sky130A
magscale 1 2
timestamp 1644949024
<< checkpaint >>
rect -1296 -1277 2204 2155
<< nwell >>
rect -36 402 944 895
<< pwell >>
rect 798 51 848 133
<< psubdiff >>
rect 798 109 848 133
rect 798 75 806 109
rect 840 75 848 109
rect 798 51 848 75
<< nsubdiff >>
rect 798 763 848 787
rect 798 729 806 763
rect 840 729 848 763
rect 798 705 848 729
<< psubdiffcont >>
rect 806 75 840 109
<< nsubdiffcont >>
rect 806 729 840 763
<< poly >>
rect 114 410 144 479
rect 48 394 144 410
rect 48 360 64 394
rect 98 360 144 394
rect 48 344 144 360
rect 114 191 144 344
<< polycont >>
rect 64 360 98 394
<< locali >>
rect 0 821 908 855
rect 62 628 96 821
rect 274 628 308 821
rect 490 628 524 821
rect 702 628 736 821
rect 806 763 840 821
rect 806 713 840 729
rect 48 394 114 410
rect 48 360 64 394
rect 98 360 114 394
rect 48 344 114 360
rect 382 394 416 594
rect 382 360 433 394
rect 382 160 416 360
rect 806 109 840 125
rect 62 17 96 60
rect 274 17 308 60
rect 490 17 524 60
rect 702 17 736 60
rect 806 17 840 75
rect 0 -17 908 17
use contact_12  contact_12_0
timestamp 1644949024
transform 1 0 48 0 1 344
box 0 0 1 1
use contact_11  contact_11_0
timestamp 1644949024
transform 1 0 798 0 1 51
box 0 0 1 1
use contact_10  contact_10_0
timestamp 1644949024
transform 1 0 798 0 1 705
box 0 0 1 1
use nmos_m6_w0_420_sli_dli_da_p  nmos_m6_w0_420_sli_dli_da_p_0
timestamp 1644949024
transform 1 0 54 0 1 51
box 0 -26 690 143
use pmos_m6_w1_260_sli_dli_da_p  pmos_m6_w1_260_sli_dli_da_p_0
timestamp 1644949024
transform 1 0 54 0 1 535
box -59 -56 749 306
<< labels >>
rlabel locali s 81 377 81 377 4 A
rlabel locali s 416 377 416 377 4 Z
rlabel locali s 454 0 454 0 4 gnd
rlabel locali s 454 838 454 838 4 vdd
<< properties >>
string FIXED_BBOX 0 0 908 838
string GDS_FILE sram_0rw2r1w_4_16_sky130A.gds
string GDS_END 470228
string GDS_START 468352
<< end >>
