magic
tech sky130A
magscale 1 2
timestamp 1644969367
<< checkpaint >>
rect -1260 -1260 80700 114196
<< metal2 >>
rect 16837 18830 16893 18839
rect 16837 18765 16893 18774
rect 17917 18834 17973 18843
rect 17917 18769 17973 18778
rect 16837 17646 16893 17655
rect 16837 17581 16893 17590
rect 17917 17642 17973 17651
rect 17917 17577 17973 17586
rect 16837 17154 16893 17163
rect 16837 17089 16893 17098
rect 17917 17158 17973 17167
rect 17917 17093 17973 17102
rect 16837 15970 16893 15979
rect 16837 15905 16893 15914
rect 17917 15966 17973 15975
rect 17917 15901 17973 15910
rect 16837 15478 16893 15487
rect 16837 15413 16893 15422
rect 17917 15482 17973 15491
rect 17917 15417 17973 15426
rect 16837 14294 16893 14303
rect 16837 14229 16893 14238
rect 17917 14290 17973 14299
rect 17917 14225 17973 14234
rect 16837 13802 16893 13811
rect 16837 13737 16893 13746
rect 17917 13806 17973 13815
rect 17917 13741 17973 13750
rect 16546 12680 16602 12689
rect 16546 12615 16602 12624
rect 16837 12618 16893 12627
rect 18326 12623 18354 30652
rect 18410 13815 18438 30652
rect 18494 14299 18522 30652
rect 18578 15491 18606 30652
rect 18662 15975 18690 30652
rect 18746 17167 18774 30652
rect 18830 17651 18858 30652
rect 18914 18843 18942 30652
rect 18900 18834 18956 18843
rect 18900 18769 18956 18778
rect 18816 17642 18872 17651
rect 18816 17577 18872 17586
rect 18732 17158 18788 17167
rect 18732 17093 18788 17102
rect 18648 15966 18704 15975
rect 18648 15901 18704 15910
rect 18564 15482 18620 15491
rect 18564 15417 18620 15426
rect 18480 14290 18536 14299
rect 18480 14225 18536 14234
rect 18396 13806 18452 13815
rect 18396 13741 18452 13750
rect 2791 7644 2847 7653
rect 2791 7579 2847 7588
rect 6313 7429 6369 7438
rect 16560 7407 16588 12615
rect 16837 12553 16893 12562
rect 17917 12614 17973 12623
rect 17917 12549 17973 12558
rect 18312 12614 18368 12623
rect 18312 12549 18368 12558
rect 25110 11719 25138 110608
rect 18112 11710 18168 11719
rect 18112 11645 18168 11654
rect 25096 11710 25152 11719
rect 25096 11645 25152 11654
rect 18112 10774 18168 10783
rect 18112 10709 18168 10718
rect 26232 10044 26260 11770
rect 76692 10774 76748 10783
rect 26909 10712 26965 10721
rect 26909 10647 26965 10656
rect 27181 10712 27237 10721
rect 27181 10647 27237 10656
rect 28465 10712 28521 10721
rect 28465 10647 28521 10656
rect 28737 10712 28793 10721
rect 28737 10647 28793 10656
rect 30021 10712 30077 10721
rect 30021 10647 30077 10656
rect 30293 10712 30349 10721
rect 30293 10647 30349 10656
rect 31577 10712 31633 10721
rect 31577 10647 31633 10656
rect 31849 10712 31905 10721
rect 31849 10647 31905 10656
rect 33133 10712 33189 10721
rect 33133 10647 33189 10656
rect 33405 10712 33461 10721
rect 33405 10647 33461 10656
rect 34689 10712 34745 10721
rect 34689 10647 34745 10656
rect 34961 10712 35017 10721
rect 34961 10647 35017 10656
rect 36245 10712 36301 10721
rect 36245 10647 36301 10656
rect 36517 10712 36573 10721
rect 36517 10647 36573 10656
rect 37801 10712 37857 10721
rect 37801 10647 37857 10656
rect 38073 10712 38129 10721
rect 38073 10647 38129 10656
rect 39357 10712 39413 10721
rect 39357 10647 39413 10656
rect 39629 10712 39685 10721
rect 39629 10647 39685 10656
rect 40913 10712 40969 10721
rect 40913 10647 40969 10656
rect 41185 10712 41241 10721
rect 41185 10647 41241 10656
rect 42469 10712 42525 10721
rect 42469 10647 42525 10656
rect 42741 10712 42797 10721
rect 42741 10647 42797 10656
rect 44025 10712 44081 10721
rect 44025 10647 44081 10656
rect 44297 10712 44353 10721
rect 44297 10647 44353 10656
rect 45581 10712 45637 10721
rect 45581 10647 45637 10656
rect 45853 10712 45909 10721
rect 45853 10647 45909 10656
rect 47137 10712 47193 10721
rect 47137 10647 47193 10656
rect 47409 10712 47465 10721
rect 47409 10647 47465 10656
rect 48693 10712 48749 10721
rect 48693 10647 48749 10656
rect 48965 10712 49021 10721
rect 48965 10647 49021 10656
rect 50249 10712 50305 10721
rect 50249 10647 50305 10656
rect 50521 10712 50577 10721
rect 76692 10709 76748 10718
rect 50521 10647 50577 10656
rect 18112 10035 18168 10044
rect 18112 9970 18168 9979
rect 26218 10035 26274 10044
rect 26218 9970 26274 9979
rect 14562 7393 16588 7407
rect 14562 7379 16640 7393
rect 6313 7364 6369 7373
rect 2791 6460 2847 6469
rect 2791 6395 2847 6404
rect 16508 3102 16640 7379
rect 76706 5786 76734 10709
rect 16508 3074 16546 3102
rect 16602 3074 16640 3102
rect 16546 3037 16602 3046
rect 19801 3040 19857 3049
rect 19801 2975 19857 2984
rect 21283 3040 21339 3049
rect 21283 2975 21339 2984
rect 22765 3040 22821 3049
rect 22765 2975 22821 2984
rect 24247 3040 24303 3049
rect 24247 2975 24303 2984
rect 25729 3040 25785 3049
rect 25729 2975 25785 2984
rect 27211 3040 27267 3049
rect 27211 2975 27267 2984
rect 28693 3040 28749 3049
rect 28693 2975 28749 2984
rect 30175 3040 30231 3049
rect 30175 2975 30231 2984
rect 31657 3040 31713 3049
rect 31657 2975 31713 2984
rect 33139 3040 33195 3049
rect 33139 2975 33195 2984
rect 34621 3040 34677 3049
rect 34621 2975 34677 2984
rect 36103 3040 36159 3049
rect 36103 2975 36159 2984
rect 37585 3040 37641 3049
rect 37585 2975 37641 2984
rect 39067 3040 39123 3049
rect 39067 2975 39123 2984
rect 40549 3040 40605 3049
rect 40549 2975 40605 2984
rect 42031 3040 42087 3049
rect 42031 2975 42087 2984
rect 43513 3040 43569 3049
rect 43513 2975 43569 2984
rect 44995 3040 45051 3049
rect 44995 2975 45051 2984
rect 46477 3040 46533 3049
rect 46477 2975 46533 2984
rect 47959 3040 48015 3049
rect 47959 2975 48015 2984
rect 49441 3040 49497 3049
rect 49441 2975 49497 2984
rect 50923 3040 50979 3049
rect 50923 2975 50979 2984
rect 52405 3040 52461 3049
rect 52405 2975 52461 2984
rect 53887 3040 53943 3049
rect 53887 2975 53943 2984
rect 55369 3040 55425 3049
rect 55369 2975 55425 2984
rect 56851 3040 56907 3049
rect 56851 2975 56907 2984
rect 58333 3040 58389 3049
rect 58333 2975 58389 2984
rect 59815 3040 59871 3049
rect 59815 2975 59871 2984
rect 61297 3040 61353 3049
rect 61297 2975 61353 2984
rect 62779 3040 62835 3049
rect 62779 2975 62835 2984
rect 64261 3040 64317 3049
rect 64261 2975 64317 2984
rect 65743 3040 65799 3049
rect 65743 2975 65799 2984
rect 67225 3040 67281 3049
rect 67225 2975 67281 2984
<< via2 >>
rect 16837 18774 16893 18830
rect 17917 18778 17973 18834
rect 16837 17590 16893 17646
rect 17917 17586 17973 17642
rect 16837 17098 16893 17154
rect 17917 17102 17973 17158
rect 16837 15914 16893 15970
rect 17917 15910 17973 15966
rect 16837 15422 16893 15478
rect 17917 15426 17973 15482
rect 16837 14238 16893 14294
rect 17917 14234 17973 14290
rect 16837 13746 16893 13802
rect 17917 13750 17973 13806
rect 16546 12624 16602 12680
rect 18900 18778 18956 18834
rect 18816 17586 18872 17642
rect 18732 17102 18788 17158
rect 18648 15910 18704 15966
rect 18564 15426 18620 15482
rect 18480 14234 18536 14290
rect 18396 13750 18452 13806
rect 2791 7588 2847 7644
rect 6313 7373 6369 7429
rect 16837 12562 16893 12618
rect 17917 12558 17973 12614
rect 18312 12558 18368 12614
rect 18112 11654 18168 11710
rect 25096 11654 25152 11710
rect 18112 10718 18168 10774
rect 26909 10656 26965 10712
rect 27181 10656 27237 10712
rect 28465 10656 28521 10712
rect 28737 10656 28793 10712
rect 30021 10656 30077 10712
rect 30293 10656 30349 10712
rect 31577 10656 31633 10712
rect 31849 10656 31905 10712
rect 33133 10656 33189 10712
rect 33405 10656 33461 10712
rect 34689 10656 34745 10712
rect 34961 10656 35017 10712
rect 36245 10656 36301 10712
rect 36517 10656 36573 10712
rect 37801 10656 37857 10712
rect 38073 10656 38129 10712
rect 39357 10656 39413 10712
rect 39629 10656 39685 10712
rect 40913 10656 40969 10712
rect 41185 10656 41241 10712
rect 42469 10656 42525 10712
rect 42741 10656 42797 10712
rect 44025 10656 44081 10712
rect 44297 10656 44353 10712
rect 45581 10656 45637 10712
rect 45853 10656 45909 10712
rect 47137 10656 47193 10712
rect 47409 10656 47465 10712
rect 48693 10656 48749 10712
rect 48965 10656 49021 10712
rect 50249 10656 50305 10712
rect 50521 10656 50577 10712
rect 76692 10718 76748 10774
rect 18112 9979 18168 10035
rect 26218 9979 26274 10035
rect 2791 6404 2847 6460
rect 16546 3046 16602 3102
rect 19801 2984 19857 3040
rect 21283 2984 21339 3040
rect 22765 2984 22821 3040
rect 24247 2984 24303 3040
rect 25729 2984 25785 3040
rect 27211 2984 27267 3040
rect 28693 2984 28749 3040
rect 30175 2984 30231 3040
rect 31657 2984 31713 3040
rect 33139 2984 33195 3040
rect 34621 2984 34677 3040
rect 36103 2984 36159 3040
rect 37585 2984 37641 3040
rect 39067 2984 39123 3040
rect 40549 2984 40605 3040
rect 42031 2984 42087 3040
rect 43513 2984 43569 3040
rect 44995 2984 45051 3040
rect 46477 2984 46533 3040
rect 47959 2984 48015 3040
rect 49441 2984 49497 3040
rect 50923 2984 50979 3040
rect 52405 2984 52461 3040
rect 53887 2984 53943 3040
rect 55369 2984 55425 3040
rect 56851 2984 56907 3040
rect 58333 2984 58389 3040
rect 59815 2984 59871 3040
rect 61297 2984 61353 3040
rect 62779 2984 62835 3040
rect 64261 2984 64317 3040
rect 65743 2984 65799 3040
rect 67225 2984 67281 3040
<< metal3 >>
rect 424 112892 79440 112936
rect 424 112828 468 112892
rect 532 112828 680 112892
rect 744 112828 892 112892
rect 956 112828 78908 112892
rect 78972 112828 79120 112892
rect 79184 112828 79332 112892
rect 79396 112828 79440 112892
rect 424 112680 79440 112828
rect 424 112616 468 112680
rect 532 112616 680 112680
rect 744 112616 892 112680
rect 956 112616 78908 112680
rect 78972 112616 79120 112680
rect 79184 112616 79332 112680
rect 79396 112616 79440 112680
rect 424 112468 79440 112616
rect 424 112404 468 112468
rect 532 112404 680 112468
rect 744 112404 892 112468
rect 956 112404 26332 112468
rect 26396 112404 78908 112468
rect 78972 112404 79120 112468
rect 79184 112404 79332 112468
rect 79396 112404 79440 112468
rect 424 112360 79440 112404
rect 1484 111832 78380 111876
rect 1484 111768 1528 111832
rect 1592 111768 1740 111832
rect 1804 111768 1952 111832
rect 2016 111768 77848 111832
rect 77912 111768 78060 111832
rect 78124 111768 78272 111832
rect 78336 111768 78380 111832
rect 1484 111620 78380 111768
rect 1484 111556 1528 111620
rect 1592 111556 1740 111620
rect 1804 111556 1952 111620
rect 2016 111556 77848 111620
rect 77912 111556 78060 111620
rect 78124 111556 78272 111620
rect 78336 111556 78380 111620
rect 1484 111408 78380 111556
rect 1484 111344 1528 111408
rect 1592 111344 1740 111408
rect 1804 111344 1952 111408
rect 2016 111344 24636 111408
rect 24700 111344 77848 111408
rect 77912 111344 78060 111408
rect 78124 111344 78272 111408
rect 78336 111344 78380 111408
rect 1484 111300 78380 111344
rect 24592 110604 24956 110816
rect 26076 110772 26440 110816
rect 26076 110708 26332 110772
rect 26396 110708 26440 110772
rect 26076 110604 26440 110708
rect 24592 110560 26440 110604
rect 24592 110496 24848 110560
rect 24912 110496 26440 110560
rect 24592 110452 26440 110496
rect 24592 109076 26440 109120
rect 24592 109012 24636 109076
rect 24700 109012 26332 109076
rect 26396 109012 26440 109076
rect 24592 108968 26440 109012
rect 24592 107592 26576 107636
rect 24592 107528 24848 107592
rect 24912 107528 26544 107592
rect 26608 107528 26652 107592
rect 24592 107484 26576 107528
rect 24592 106108 26440 106152
rect 24592 106044 26332 106108
rect 26396 106044 26440 106108
rect 24592 106000 26440 106044
rect 24592 105788 24956 106000
rect 26076 105896 26440 106000
rect 26076 105832 26120 105896
rect 26184 105832 26440 105896
rect 26076 105788 26440 105832
rect 24592 104624 26652 104668
rect 24592 104560 26544 104624
rect 26608 104560 26652 104624
rect 24592 104516 26652 104560
rect 24592 104412 24956 104516
rect 24592 104348 24848 104412
rect 24912 104348 24956 104412
rect 24592 104304 24956 104348
rect 26076 104304 26440 104516
rect 24592 102928 26440 102972
rect 24592 102864 24636 102928
rect 24700 102864 26120 102928
rect 26184 102864 26440 102928
rect 24592 102820 26440 102864
rect 24592 101444 26440 101488
rect 24592 101380 24848 101444
rect 24912 101380 26120 101444
rect 26184 101380 26440 101444
rect 24592 101336 26440 101380
rect 24592 99960 24956 100004
rect 24592 99896 24636 99960
rect 24700 99896 24956 99960
rect 24592 99792 24956 99896
rect 26076 99792 26440 100004
rect 24592 99748 26440 99792
rect 24592 99684 24636 99748
rect 24700 99684 26440 99748
rect 24592 99640 26440 99684
rect 24592 98308 24956 98520
rect 26076 98476 26440 98520
rect 26076 98412 26120 98476
rect 26184 98412 26440 98476
rect 26076 98308 26440 98412
rect 24380 98264 26440 98308
rect 24380 98200 24424 98264
rect 24488 98200 26440 98264
rect 24380 98156 26440 98200
rect 24592 96780 26440 96824
rect 24592 96716 24636 96780
rect 24700 96716 24848 96780
rect 24912 96716 26440 96780
rect 24592 96672 26440 96716
rect 24456 95296 26440 95340
rect 24380 95232 24424 95296
rect 24488 95232 26332 95296
rect 26396 95232 26440 95296
rect 24456 95188 26440 95232
rect 24592 93812 24956 93856
rect 24592 93748 24848 93812
rect 24912 93748 24956 93812
rect 24592 93644 24956 93748
rect 26076 93644 26440 93856
rect 24592 93600 26440 93644
rect 24592 93536 26120 93600
rect 26184 93536 26440 93600
rect 24592 93492 26440 93536
rect 24592 92328 26440 92372
rect 24592 92264 26332 92328
rect 26396 92264 26440 92328
rect 24592 92220 26440 92264
rect 24592 92008 24956 92220
rect 26076 92008 26440 92220
rect 24592 90632 26440 90676
rect 24592 90568 24636 90632
rect 24700 90568 26120 90632
rect 26184 90568 26440 90632
rect 24592 90524 26440 90568
rect 24592 89040 26440 89192
rect 24592 88828 24956 89040
rect 26076 88936 26440 89040
rect 26076 88872 26332 88936
rect 26396 88872 26440 88936
rect 26076 88828 26440 88872
rect 24592 87664 24956 87708
rect 24592 87600 24636 87664
rect 24700 87600 24956 87664
rect 24592 87496 24956 87600
rect 26076 87496 26440 87708
rect 24592 87452 26440 87496
rect 24592 87388 26120 87452
rect 26184 87388 26440 87452
rect 24592 87344 26440 87388
rect 24592 86012 24956 86224
rect 26076 86180 26440 86224
rect 26076 86116 26332 86180
rect 26396 86116 26440 86180
rect 26076 86012 26440 86116
rect 24592 85968 26440 86012
rect 24592 85904 24848 85968
rect 24912 85904 26440 85968
rect 24592 85860 26440 85904
rect 24592 84484 26440 84528
rect 24592 84420 26120 84484
rect 26184 84420 26332 84484
rect 26396 84420 26440 84484
rect 24592 84376 26440 84420
rect 24592 83000 26440 83044
rect 24592 82936 24848 83000
rect 24912 82936 26440 83000
rect 24592 82892 26440 82936
rect 24592 82680 24956 82892
rect 26076 82788 26440 82892
rect 26076 82724 26120 82788
rect 26184 82724 26440 82788
rect 26076 82680 26440 82724
rect 24592 81348 24956 81560
rect 26076 81516 26440 81560
rect 26076 81452 26332 81516
rect 26396 81452 26440 81516
rect 26076 81348 26440 81452
rect 24592 81304 26440 81348
rect 24592 81240 26332 81304
rect 26396 81240 26440 81304
rect 24592 81196 26440 81240
rect 24592 79864 24956 80076
rect 26076 80032 26440 80076
rect 26076 79968 26120 80032
rect 26184 79968 26440 80032
rect 26076 79864 26440 79968
rect 24592 79820 26576 79864
rect 24592 79756 26544 79820
rect 26608 79756 26652 79820
rect 24592 79712 26576 79756
rect 24592 78336 26440 78380
rect 24592 78272 26120 78336
rect 26184 78272 26332 78336
rect 26396 78272 26440 78336
rect 24592 78228 26440 78272
rect 24592 76852 26652 76896
rect 24592 76788 26544 76852
rect 26608 76788 26652 76852
rect 24592 76744 26652 76788
rect 24592 76640 24956 76744
rect 24592 76576 24848 76640
rect 24912 76576 24956 76640
rect 24592 76532 24956 76576
rect 26076 76532 26440 76744
rect 24592 75200 24956 75412
rect 26076 75368 26440 75412
rect 26076 75304 26120 75368
rect 26184 75304 26440 75368
rect 26076 75200 26440 75304
rect 24592 75156 26440 75200
rect 24592 75092 24636 75156
rect 24700 75092 26440 75156
rect 24592 75048 26440 75092
rect 24592 73884 26440 73928
rect 24592 73820 24848 73884
rect 24912 73820 26440 73884
rect 24592 73776 26440 73820
rect 24592 73672 24956 73776
rect 24592 73608 24848 73672
rect 24912 73608 24956 73672
rect 24592 73564 24956 73608
rect 26076 73564 26440 73776
rect 24592 72188 26440 72232
rect 24592 72124 24636 72188
rect 24700 72124 26120 72188
rect 26184 72124 26440 72188
rect 24592 72080 26440 72124
rect 24592 70704 24956 70748
rect 24592 70640 24848 70704
rect 24912 70640 24956 70704
rect 24592 70536 24956 70640
rect 26076 70536 26440 70748
rect 24592 70492 26440 70536
rect 24592 70428 26332 70492
rect 26396 70428 26440 70492
rect 24592 70384 26440 70428
rect 24592 69052 24956 69264
rect 26076 69220 26440 69264
rect 26076 69156 26120 69220
rect 26184 69156 26440 69220
rect 26076 69052 26440 69156
rect 24592 69008 26440 69052
rect 24592 68944 26120 69008
rect 26184 68944 26440 69008
rect 24592 68900 26440 68944
rect 24592 67568 24956 67780
rect 26076 67736 26440 67780
rect 26076 67672 26332 67736
rect 26396 67672 26440 67736
rect 26076 67568 26440 67672
rect 24592 67524 26652 67568
rect 24592 67460 26544 67524
rect 26608 67460 26652 67524
rect 24592 67416 26652 67460
rect 24592 66040 26440 66084
rect 24592 65976 26120 66040
rect 26184 65976 26332 66040
rect 26396 65976 26440 66040
rect 24592 65932 26440 65976
rect 24592 64556 26576 64600
rect 24592 64492 26544 64556
rect 26608 64492 26652 64556
rect 24592 64448 26576 64492
rect 24592 64236 24956 64448
rect 26076 64344 26440 64448
rect 26076 64280 26120 64344
rect 26184 64280 26440 64344
rect 26076 64236 26440 64280
rect 24592 63072 26440 63116
rect 24592 63008 26332 63072
rect 26396 63008 26440 63072
rect 24592 62964 26440 63008
rect 24592 62752 24956 62964
rect 26076 62860 26440 62964
rect 26076 62796 26332 62860
rect 26396 62796 26440 62860
rect 26076 62752 26440 62796
rect 24592 61420 24956 61632
rect 26076 61588 26440 61632
rect 26076 61524 26120 61588
rect 26184 61524 26440 61588
rect 26076 61420 26440 61524
rect 24592 61376 26440 61420
rect 24592 61312 24848 61376
rect 24912 61312 26440 61376
rect 24592 61268 26440 61312
rect 24592 59892 26440 59936
rect 24592 59828 26120 59892
rect 26184 59828 26332 59892
rect 26396 59828 26440 59892
rect 24592 59784 26440 59828
rect 24592 58408 26440 58452
rect 24592 58344 24848 58408
rect 24912 58344 26440 58408
rect 24592 58300 26440 58344
rect 24592 58196 24956 58300
rect 24592 58132 24848 58196
rect 24912 58132 24956 58196
rect 24592 58088 24956 58132
rect 26076 58088 26440 58300
rect 24592 56756 24956 56968
rect 26076 56924 26440 56968
rect 26076 56860 26120 56924
rect 26184 56860 26440 56924
rect 26076 56756 26440 56860
rect 24592 56712 26440 56756
rect 24592 56648 26120 56712
rect 26184 56648 26440 56712
rect 24592 56604 26440 56648
rect 24592 55440 26440 55484
rect 24592 55376 24848 55440
rect 24912 55376 26440 55440
rect 24592 55332 26440 55376
rect 24592 55228 24956 55332
rect 24592 55164 24636 55228
rect 24700 55164 24956 55228
rect 24592 55120 24956 55164
rect 26076 55120 26440 55332
rect 24592 53744 26440 53788
rect 24592 53680 26120 53744
rect 26184 53680 26332 53744
rect 26396 53680 26440 53744
rect 24592 53636 26440 53680
rect 24592 52260 24956 52304
rect 24592 52196 24636 52260
rect 24700 52196 24956 52260
rect 24592 52092 24956 52196
rect 26076 52092 26440 52304
rect 24592 52048 26652 52092
rect 24592 51984 26544 52048
rect 26608 51984 26652 52048
rect 24592 51940 26652 51984
rect 24592 50776 26440 50820
rect 24592 50712 26332 50776
rect 26396 50712 26440 50776
rect 24592 50668 26440 50712
rect 24592 50456 24956 50668
rect 26076 50564 26440 50668
rect 26076 50500 26120 50564
rect 26184 50500 26440 50564
rect 26076 50456 26440 50500
rect 19292 49184 20716 49336
rect 19292 48972 19656 49184
rect 20352 49124 20716 49184
rect 20216 49080 20716 49124
rect 20140 49016 20184 49080
rect 20248 49016 20716 49080
rect 20216 48972 20716 49016
rect 24592 49124 24956 49336
rect 26076 49292 26576 49336
rect 26076 49228 26544 49292
rect 26608 49228 26652 49292
rect 26076 49184 26576 49228
rect 26076 49124 26440 49184
rect 24592 49080 26440 49124
rect 24592 49016 24848 49080
rect 24912 49016 26440 49080
rect 24592 48972 26440 49016
rect 19292 47596 21140 47640
rect 19292 47532 19336 47596
rect 19400 47532 21140 47596
rect 19292 47488 21140 47532
rect 20988 47428 21140 47488
rect 24592 47596 26440 47640
rect 24592 47532 24636 47596
rect 24700 47532 26120 47596
rect 26184 47532 26440 47596
rect 24592 47488 26440 47532
rect 24592 47428 24744 47488
rect 20988 47276 24744 47428
rect 19504 46216 20504 46368
rect 19504 46156 19656 46216
rect 20352 46156 20504 46216
rect 19292 46112 20292 46156
rect 19292 46048 20184 46112
rect 20248 46048 20292 46112
rect 19292 46004 20292 46048
rect 20352 46004 20716 46156
rect 24592 46112 24956 46156
rect 24592 46048 24848 46112
rect 24912 46048 24956 46112
rect 19504 45944 19656 46004
rect 24592 45944 24956 46048
rect 26076 45944 26440 46156
rect 19504 45900 20504 45944
rect 19504 45836 20396 45900
rect 20460 45836 20504 45900
rect 19504 45792 20504 45836
rect 24592 45900 26440 45944
rect 24592 45836 24848 45900
rect 24912 45836 26440 45900
rect 24592 45792 26440 45836
rect 19292 44628 19656 44672
rect 19292 44564 19336 44628
rect 19400 44564 19656 44628
rect 19292 44460 19656 44564
rect 20352 44460 20716 44672
rect 19292 44416 20716 44460
rect 19292 44352 20608 44416
rect 20672 44352 20716 44416
rect 19292 44308 20716 44352
rect 24592 44628 26440 44672
rect 24592 44564 24636 44628
rect 24700 44564 26440 44628
rect 24592 44520 26440 44564
rect 24592 44308 24956 44520
rect 26076 44416 26440 44520
rect 26076 44352 26120 44416
rect 26184 44352 26440 44416
rect 26076 44308 26440 44352
rect 19292 42976 19656 43188
rect 20352 43144 20716 43188
rect 20352 43080 20396 43144
rect 20460 43080 20716 43144
rect 20352 42976 20716 43080
rect 19292 42932 20716 42976
rect 19292 42868 20396 42932
rect 20460 42868 20716 42932
rect 19292 42824 20716 42868
rect 24592 42932 26440 42976
rect 24592 42868 24848 42932
rect 24912 42868 26440 42932
rect 24592 42824 26440 42868
rect 24804 42720 24956 42824
rect 24804 42656 24848 42720
rect 24912 42656 24956 42720
rect 19292 41448 20716 41492
rect 19292 41384 19336 41448
rect 19400 41384 20608 41448
rect 20672 41384 20716 41448
rect 19292 41340 20716 41384
rect 24592 41448 26440 41492
rect 24592 41384 24636 41448
rect 24700 41384 26120 41448
rect 26184 41384 26440 41448
rect 24592 41340 26440 41384
rect 19504 40176 20504 40220
rect 19504 40112 20396 40176
rect 20460 40112 20504 40176
rect 19504 40068 20504 40112
rect 19504 40008 19656 40068
rect 19292 39856 20716 40008
rect 19292 39644 19656 39856
rect 20352 39752 20716 39856
rect 20352 39688 20608 39752
rect 20672 39688 20716 39752
rect 20352 39644 20716 39688
rect 24592 39964 26440 40008
rect 24592 39900 24848 39964
rect 24912 39900 26440 39964
rect 24592 39856 26440 39900
rect 24592 39644 24956 39856
rect 26076 39752 26440 39856
rect 26076 39688 26332 39752
rect 26396 39688 26440 39752
rect 26076 39644 26440 39688
rect 19292 38480 20716 38524
rect 19292 38416 19336 38480
rect 19400 38416 20716 38480
rect 19292 38372 20716 38416
rect 19292 38160 19656 38372
rect 20352 38160 20716 38372
rect 24592 38480 24956 38524
rect 24592 38416 24636 38480
rect 24700 38416 24956 38480
rect 24592 38312 24956 38416
rect 26076 38312 26440 38524
rect 24592 38268 26440 38312
rect 24592 38204 24848 38268
rect 24912 38204 26440 38268
rect 24592 38160 26440 38204
rect 19292 36996 20716 37040
rect 19292 36932 20608 36996
rect 20672 36932 20716 36996
rect 19292 36888 20716 36932
rect 19292 36676 19656 36888
rect 20352 36784 20716 36888
rect 20352 36720 20396 36784
rect 20460 36720 20716 36784
rect 20352 36676 20716 36720
rect 24592 36784 26440 36828
rect 24592 36720 26120 36784
rect 26184 36720 26332 36784
rect 26396 36720 26440 36784
rect 24592 36676 26440 36720
rect 24592 35300 26440 35344
rect 24592 35236 24848 35300
rect 24912 35236 26440 35300
rect 24592 35192 26440 35236
rect 19292 33816 20716 33860
rect 19292 33752 20396 33816
rect 20460 33752 20716 33816
rect 19292 33708 20716 33752
rect 19292 33648 19656 33708
rect 19292 33604 20292 33648
rect 19292 33540 20184 33604
rect 20248 33540 20292 33604
rect 19292 33496 20292 33540
rect 20352 33496 20716 33708
rect 24592 33648 24956 33860
rect 26076 33816 26440 33860
rect 26076 33752 26120 33816
rect 26184 33752 26440 33816
rect 26076 33648 26440 33752
rect 24592 33604 26440 33648
rect 24592 33540 26332 33604
rect 26396 33540 26440 33604
rect 24592 33496 26440 33540
rect 19292 32164 19656 32376
rect 20352 32164 20716 32376
rect 19292 32120 20716 32164
rect 19292 32056 20396 32120
rect 20460 32056 20716 32120
rect 19292 32012 20716 32056
rect 24592 32164 24956 32376
rect 26076 32164 26440 32376
rect 24592 32120 26440 32164
rect 24592 32056 24636 32120
rect 24700 32056 26440 32120
rect 24592 32012 26440 32056
rect 19292 30680 19656 30892
rect 20216 30848 20716 30892
rect 20140 30784 20184 30848
rect 20248 30784 20716 30848
rect 20216 30740 20716 30784
rect 20352 30680 20716 30740
rect 19292 30636 20928 30680
rect 19292 30572 20820 30636
rect 20884 30572 20928 30636
rect 19292 30528 20928 30572
rect 24592 30636 26440 30680
rect 24592 30572 26120 30636
rect 26184 30572 26332 30636
rect 26396 30572 26440 30636
rect 24592 30528 26440 30572
rect 19292 29152 20716 29196
rect 19292 29088 20396 29152
rect 20460 29088 20608 29152
rect 20672 29088 20716 29152
rect 19292 29044 20716 29088
rect 24592 29152 26440 29196
rect 24592 29088 24636 29152
rect 24700 29088 24848 29152
rect 24912 29088 26440 29152
rect 24592 29044 26440 29088
rect 19292 27500 19656 27712
rect 20352 27668 20852 27712
rect 20352 27604 20820 27668
rect 20884 27604 20928 27668
rect 20352 27560 20852 27604
rect 20352 27500 20716 27560
rect 19292 27456 20716 27500
rect 19292 27392 20396 27456
rect 20460 27392 20716 27456
rect 19292 27348 20716 27392
rect 24592 27500 24956 27712
rect 26076 27668 26440 27712
rect 26076 27604 26120 27668
rect 26184 27604 26440 27668
rect 26076 27500 26440 27604
rect 24592 27456 26440 27500
rect 24592 27392 24636 27456
rect 24700 27392 26440 27456
rect 24592 27348 26440 27392
rect 19292 26184 20716 26228
rect 19292 26120 20608 26184
rect 20672 26120 20716 26184
rect 19292 26076 20716 26120
rect 19292 25864 19656 26076
rect 20352 26016 20716 26076
rect 20216 25972 20716 26016
rect 20140 25908 20184 25972
rect 20248 25908 20716 25972
rect 20216 25864 20716 25908
rect 24592 26184 26440 26228
rect 24592 26120 24848 26184
rect 24912 26120 26440 26184
rect 24592 26076 26440 26120
rect 24592 25864 24956 26076
rect 26076 25972 26440 26076
rect 26076 25908 26120 25972
rect 26184 25908 26440 25972
rect 26076 25864 26440 25908
rect 19504 24592 20504 24744
rect 19504 24532 19656 24592
rect 20352 24532 20504 24592
rect 19292 24488 20080 24532
rect 19292 24424 19972 24488
rect 20036 24424 20080 24488
rect 19292 24380 20080 24424
rect 20352 24488 20716 24532
rect 20352 24424 20396 24488
rect 20460 24424 20716 24488
rect 20352 24380 20716 24424
rect 24592 24488 26576 24532
rect 24592 24424 24636 24488
rect 24700 24424 26544 24488
rect 26608 24424 26652 24488
rect 24592 24380 26576 24424
rect 19504 23108 20504 23260
rect 19504 23048 19656 23108
rect 20352 23048 20504 23108
rect 19292 23004 20292 23048
rect 19292 22940 19336 23004
rect 19400 22940 20184 23004
rect 20248 22940 20292 23004
rect 19292 22896 20292 22940
rect 20352 22896 21140 23048
rect 20988 22836 21140 22896
rect 24592 23004 26440 23048
rect 24592 22940 26120 23004
rect 26184 22940 26332 23004
rect 26396 22940 26440 23004
rect 24592 22896 26440 22940
rect 24592 22836 24744 22896
rect 20988 22684 24744 22836
rect 19292 21412 20716 21564
rect 19292 21200 19656 21412
rect 20352 21352 20716 21412
rect 20004 21308 20716 21352
rect 19928 21244 19972 21308
rect 20036 21244 20716 21308
rect 20004 21200 20716 21244
rect 24592 21520 26652 21564
rect 24592 21456 26544 21520
rect 26608 21456 26652 21520
rect 24592 21412 26652 21456
rect 24592 21308 24956 21412
rect 24592 21244 24848 21308
rect 24912 21244 24956 21308
rect 24592 21200 24956 21244
rect 26076 21200 26440 21412
rect 19292 20928 19444 21200
rect 17172 20776 19444 20928
rect 17172 20672 17536 20776
rect 17172 20608 17216 20672
rect 17280 20608 17536 20672
rect 17172 20564 17536 20608
rect 17172 20036 19444 20080
rect 17172 19972 19336 20036
rect 19400 19972 19444 20036
rect 17172 19928 19444 19972
rect 24592 20036 26440 20080
rect 24592 19972 26332 20036
rect 26396 19972 26440 20036
rect 24592 19928 26440 19972
rect 17172 19824 17536 19928
rect 17172 19760 17428 19824
rect 17492 19760 17536 19824
rect 17172 19716 17536 19760
rect 24592 19824 24956 19928
rect 24592 19760 24636 19824
rect 24700 19760 24956 19824
rect 24592 19716 24956 19760
rect 26076 19716 26440 19928
rect 17172 19188 17536 19232
rect 17172 19124 17216 19188
rect 17280 19124 17536 19188
rect 17172 19080 17536 19124
rect 17333 19020 17536 19080
rect 16748 18830 17112 19020
rect 17333 19011 17672 19020
rect 17384 18976 17672 19011
rect 17384 18912 17640 18976
rect 17704 18912 17748 18976
rect 17384 18868 17672 18912
rect 16748 18808 16837 18830
rect 0 18774 16837 18808
rect 16893 18774 17112 18830
rect 0 18656 17112 18774
rect 17879 18836 18011 18839
rect 18862 18836 18994 18839
rect 17879 18834 18994 18836
rect 17879 18778 17917 18834
rect 17973 18778 18900 18834
rect 18956 18778 18994 18834
rect 17879 18776 18994 18778
rect 17879 18773 18011 18776
rect 18862 18773 18994 18776
rect 24804 18552 24956 18596
rect 24804 18488 24848 18552
rect 24912 18488 24956 18552
rect 24804 18384 24956 18488
rect 17172 18340 17536 18384
rect 17172 18276 17428 18340
rect 17492 18276 17536 18340
rect 17172 18128 17536 18276
rect 19504 18340 20716 18384
rect 19504 18276 19548 18340
rect 19612 18276 20716 18340
rect 19504 18232 20716 18276
rect 24592 18340 26440 18384
rect 24592 18276 24848 18340
rect 24912 18276 26440 18340
rect 24592 18232 26440 18276
rect 17172 18064 17216 18128
rect 17280 18064 17536 18128
rect 17172 18020 17536 18064
rect 17460 17916 19656 17960
rect 17384 17852 17428 17916
rect 17492 17852 19548 17916
rect 19612 17852 19656 17916
rect 17460 17808 19656 17852
rect 0 17646 17112 17748
rect 0 17596 16837 17646
rect 16748 17590 16837 17596
rect 16893 17590 17112 17646
rect 16748 17384 17112 17590
rect 17879 17644 18011 17647
rect 18778 17644 18910 17647
rect 17879 17642 18910 17644
rect 17879 17586 17917 17642
rect 17973 17586 18816 17642
rect 18872 17586 18910 17642
rect 17879 17584 18910 17586
rect 17879 17581 18011 17584
rect 18778 17581 18910 17584
rect 17384 17492 17748 17536
rect 17384 17428 17428 17492
rect 17492 17428 17640 17492
rect 17704 17428 17748 17492
rect 17384 17409 17748 17428
rect 17333 17384 17748 17409
rect 17333 17335 17536 17384
rect 16748 17154 17112 17324
rect 17384 17280 17536 17335
rect 17384 17216 17428 17280
rect 17492 17216 17536 17280
rect 17384 17172 17536 17216
rect 16748 17112 16837 17154
rect 0 17098 16837 17112
rect 16893 17098 17112 17154
rect 0 16960 17112 17098
rect 17879 17160 18011 17163
rect 18694 17160 18826 17163
rect 17879 17158 18826 17160
rect 17879 17102 17917 17158
rect 17973 17102 18732 17158
rect 18788 17102 18826 17158
rect 17879 17100 18826 17102
rect 17879 17097 18011 17100
rect 18694 17097 18826 17100
rect 19504 16748 20716 16900
rect 24592 16856 26440 16900
rect 24592 16792 24636 16856
rect 24700 16792 26120 16856
rect 26184 16792 26440 16856
rect 24592 16748 26440 16792
rect 19504 16688 19656 16748
rect 17172 16644 19656 16688
rect 17172 16580 17216 16644
rect 17280 16580 19656 16644
rect 17172 16536 19656 16580
rect 17172 16476 17536 16536
rect 16960 16432 17536 16476
rect 16960 16368 17004 16432
rect 17068 16368 17536 16432
rect 16960 16324 17536 16368
rect 16324 16008 17112 16052
rect 16324 15944 16368 16008
rect 16432 15970 17112 16008
rect 16432 15944 16837 15970
rect 16324 15914 16837 15944
rect 16893 15914 17112 15970
rect 16324 15900 17112 15914
rect 17384 16008 17748 16052
rect 17384 15944 17640 16008
rect 17704 15944 17748 16008
rect 17384 15900 17748 15944
rect 17879 15968 18011 15971
rect 18610 15968 18742 15971
rect 17879 15966 18742 15968
rect 17879 15910 17917 15966
rect 17973 15910 18648 15966
rect 18704 15910 18742 15966
rect 17879 15908 18742 15910
rect 17879 15905 18011 15908
rect 18610 15905 18742 15908
rect 17384 15840 17536 15900
rect 17384 15796 17960 15840
rect 17384 15733 17428 15796
rect 17333 15732 17428 15733
rect 17492 15732 17852 15796
rect 17916 15732 17960 15796
rect 17333 15688 17960 15732
rect 17333 15659 17465 15688
rect 16748 15478 17112 15628
rect 16748 15422 16837 15478
rect 16893 15422 17112 15478
rect 16748 15416 17112 15422
rect 17879 15484 18011 15487
rect 18526 15484 18658 15487
rect 17879 15482 18658 15484
rect 17879 15426 17917 15482
rect 17973 15426 18564 15482
rect 18620 15426 18658 15482
rect 17879 15424 18658 15426
rect 17879 15421 18011 15424
rect 18526 15421 18658 15424
rect 16748 15372 17324 15416
rect 16748 15308 17216 15372
rect 17280 15308 17324 15372
rect 16748 15264 17324 15308
rect 19504 15264 20716 15416
rect 19504 15204 19868 15264
rect 17672 15160 19868 15204
rect 17596 15096 17640 15160
rect 17704 15096 19868 15160
rect 17672 15052 19868 15096
rect 20564 15052 20716 15264
rect 24592 15372 24956 15416
rect 24592 15308 24848 15372
rect 24912 15308 24956 15372
rect 24592 15204 24956 15308
rect 26076 15204 26440 15416
rect 24592 15160 26440 15204
rect 24592 15096 26332 15160
rect 26396 15096 26440 15160
rect 24592 15052 26440 15096
rect 17036 14948 17536 14992
rect 16960 14884 17004 14948
rect 17068 14884 17536 14948
rect 17036 14840 17536 14884
rect 17172 14780 17536 14840
rect 17172 14736 17748 14780
rect 17172 14672 17640 14736
rect 17704 14672 17748 14736
rect 17172 14628 17748 14672
rect 17384 14524 18096 14568
rect 17384 14460 18064 14524
rect 18128 14460 18172 14524
rect 17384 14416 18096 14460
rect 16536 14312 17112 14356
rect 16536 14248 16580 14312
rect 16644 14294 17112 14312
rect 16644 14248 16837 14294
rect 16536 14238 16837 14248
rect 16893 14238 17112 14294
rect 16536 14204 17112 14238
rect 17384 14144 17536 14416
rect 17879 14292 18011 14295
rect 18442 14292 18574 14295
rect 17879 14290 18574 14292
rect 17879 14234 17917 14290
rect 17973 14234 18480 14290
rect 18536 14234 18574 14290
rect 17879 14232 18574 14234
rect 17879 14229 18011 14232
rect 18442 14229 18574 14232
rect 17384 14100 17884 14144
rect 17384 14057 17852 14100
rect 17333 14036 17852 14057
rect 17916 14036 17960 14100
rect 17333 13992 17884 14036
rect 17333 13983 17536 13992
rect 16748 13802 17112 13932
rect 16748 13746 16837 13802
rect 16893 13746 17112 13802
rect 17384 13780 17536 13983
rect 17879 13808 18011 13811
rect 18358 13808 18490 13811
rect 17879 13806 18490 13808
rect 16748 13676 17112 13746
rect 17879 13750 17917 13806
rect 17973 13750 18396 13806
rect 18452 13750 18490 13806
rect 17879 13748 18490 13750
rect 17879 13745 18011 13748
rect 18358 13745 18490 13748
rect 16748 13612 17004 13676
rect 17068 13612 17112 13676
rect 16748 13568 17112 13612
rect 19504 13720 19868 13932
rect 20564 13720 20716 13932
rect 19504 13568 20716 13720
rect 24592 13720 24956 13932
rect 26076 13888 26440 13932
rect 26076 13824 26120 13888
rect 26184 13824 26440 13888
rect 26076 13720 26440 13824
rect 24592 13676 27288 13720
rect 24592 13612 27180 13676
rect 27244 13612 27288 13676
rect 24592 13568 27288 13612
rect 19504 13508 19656 13568
rect 17384 13356 19656 13508
rect 17384 13296 17536 13356
rect 17172 13252 17672 13296
rect 17172 13188 17640 13252
rect 17704 13188 17748 13252
rect 17172 13144 17672 13188
rect 16574 12685 16658 12689
rect 16508 12680 16658 12685
rect 16508 12624 16546 12680
rect 16602 12624 16658 12680
rect 16508 12619 16658 12624
rect 16574 12615 16658 12619
rect 16748 12627 16900 12660
rect 16960 12627 17112 12660
rect 16748 12618 17112 12627
rect 16748 12616 16837 12618
rect 16748 12552 16792 12616
rect 16893 12562 17112 12618
rect 16856 12553 17112 12562
rect 17879 12616 18011 12619
rect 18274 12616 18406 12619
rect 17879 12614 18406 12616
rect 17879 12558 17917 12614
rect 17973 12558 18312 12614
rect 18368 12558 18406 12614
rect 17879 12556 18406 12558
rect 17879 12553 18011 12556
rect 18274 12553 18406 12556
rect 16856 12552 16900 12553
rect 16748 12508 16900 12552
rect 16960 12508 17112 12553
rect 17384 12404 19656 12448
rect 17384 12381 18064 12404
rect 17333 12340 18064 12381
rect 18128 12340 19656 12404
rect 17333 12307 19656 12340
rect 17384 12296 19656 12307
rect 17384 12236 17536 12296
rect 19504 12236 19656 12296
rect 17384 12192 18596 12236
rect 17384 12128 18488 12192
rect 18552 12128 18596 12192
rect 17384 12084 18596 12128
rect 19504 12084 20716 12236
rect 24592 12192 28984 12236
rect 24592 12128 24636 12192
rect 24700 12128 26332 12192
rect 26396 12128 28984 12192
rect 24592 12084 28984 12128
rect 27136 11872 27500 12084
rect 28832 12024 28984 12084
rect 30316 12024 30680 12236
rect 31800 12024 32164 12236
rect 33496 12084 38312 12236
rect 33496 12024 33648 12084
rect 28832 11872 33648 12024
rect 34980 11872 35344 12084
rect 36464 11872 36828 12084
rect 38160 12024 38312 12084
rect 39644 12024 40008 12236
rect 41128 12024 41492 12236
rect 42824 12084 44672 12236
rect 42824 12024 42976 12084
rect 38160 11872 42976 12024
rect 44308 12024 44672 12084
rect 45792 12084 47640 12236
rect 45792 12024 46156 12084
rect 44308 11872 46156 12024
rect 47488 12024 47640 12084
rect 48972 12084 50820 12236
rect 48972 12024 49336 12084
rect 47488 11872 49336 12024
rect 50456 12024 50820 12084
rect 52152 12024 52304 12236
rect 53636 12084 56968 12236
rect 53636 12024 54000 12084
rect 50456 11872 54000 12024
rect 55120 11872 55484 12084
rect 56816 12024 56968 12084
rect 58300 12024 58664 12236
rect 59784 12024 60148 12236
rect 61480 12084 63328 12236
rect 61480 12024 61632 12084
rect 56816 11872 61632 12024
rect 62964 12024 63328 12084
rect 64448 12024 64812 12236
rect 66144 12024 66296 12236
rect 67628 12084 70960 12236
rect 67628 12024 67992 12084
rect 62964 11872 67992 12024
rect 69112 11872 69476 12084
rect 70808 12024 70960 12084
rect 72292 12084 75624 12236
rect 72292 12024 72656 12084
rect 70808 11872 72656 12024
rect 73988 11872 74140 12084
rect 75472 11980 75624 12084
rect 75472 11916 75516 11980
rect 75580 11916 75624 11980
rect 75472 11872 75624 11916
rect 18074 11712 18206 11715
rect 25058 11712 25190 11715
rect 18074 11710 25190 11712
rect 18074 11654 18112 11710
rect 18168 11654 25096 11710
rect 25152 11654 25190 11710
rect 18074 11652 25190 11654
rect 18074 11649 18206 11652
rect 25058 11649 25190 11652
rect 23956 11344 24744 11388
rect 23956 11280 24636 11344
rect 24700 11280 24744 11344
rect 23956 11236 24744 11280
rect 27136 11344 27500 11388
rect 27136 11280 27180 11344
rect 27244 11280 27500 11344
rect 23956 11132 24320 11236
rect 23956 11068 24212 11132
rect 24276 11068 24320 11132
rect 23956 11024 24320 11068
rect 27136 11132 27500 11280
rect 27136 11068 27392 11132
rect 27456 11068 27500 11132
rect 27136 11024 27500 11068
rect 28832 11132 28984 11388
rect 28832 11068 28876 11132
rect 28940 11068 28984 11132
rect 28832 11024 28984 11068
rect 30316 11176 30680 11388
rect 30316 11132 30816 11176
rect 31800 11132 32164 11388
rect 30316 11068 30784 11132
rect 30848 11068 30892 11132
rect 31800 11068 32056 11132
rect 32120 11068 32164 11132
rect 30316 11024 30816 11068
rect 31800 11024 32164 11068
rect 33496 11176 33648 11388
rect 33496 11132 33784 11176
rect 34980 11132 35344 11388
rect 33496 11068 33752 11132
rect 33816 11068 33860 11132
rect 34980 11068 35236 11132
rect 35300 11068 35344 11132
rect 33496 11024 33784 11068
rect 34980 11024 35344 11068
rect 36464 11132 36828 11388
rect 36464 11068 36720 11132
rect 36784 11068 36828 11132
rect 36464 11024 36828 11068
rect 38160 11176 38312 11388
rect 39644 11176 40008 11388
rect 41128 11176 41492 11388
rect 38160 11132 38448 11176
rect 39644 11132 41492 11176
rect 38160 11068 38416 11132
rect 38480 11068 38524 11132
rect 39644 11068 39900 11132
rect 39964 11068 41492 11132
rect 38160 11024 38448 11068
rect 39644 11024 41492 11068
rect 42824 11176 42976 11388
rect 42824 11132 43112 11176
rect 44308 11132 44672 11388
rect 45792 11176 46156 11388
rect 45656 11132 46156 11176
rect 42824 11068 43080 11132
rect 43144 11068 43188 11132
rect 44308 11068 44564 11132
rect 44628 11068 44672 11132
rect 45580 11068 45624 11132
rect 45688 11068 46156 11132
rect 42824 11024 43112 11068
rect 44308 11024 44672 11068
rect 45656 11024 46156 11068
rect 47488 11132 47640 11388
rect 48972 11176 49336 11388
rect 50456 11176 50820 11388
rect 48624 11132 49336 11176
rect 50320 11132 50820 11176
rect 47488 11068 47532 11132
rect 47596 11068 47640 11132
rect 48548 11068 48592 11132
rect 48656 11068 49336 11132
rect 50244 11068 50288 11132
rect 50352 11068 50820 11132
rect 47488 11024 47640 11068
rect 48624 11024 49336 11068
rect 50320 11024 50820 11068
rect 52152 11132 52304 11388
rect 52152 11068 52196 11132
rect 52260 11068 52304 11132
rect 52152 11024 52304 11068
rect 53636 11132 54000 11388
rect 55120 11176 55484 11388
rect 56816 11176 56968 11388
rect 54984 11132 55484 11176
rect 56468 11132 56968 11176
rect 53636 11068 53680 11132
rect 53744 11068 54000 11132
rect 54908 11068 54952 11132
rect 55016 11068 55484 11132
rect 56392 11068 56436 11132
rect 56500 11068 56968 11132
rect 53636 11024 54000 11068
rect 54984 11024 55484 11068
rect 56468 11024 56968 11068
rect 58300 11132 58664 11388
rect 59784 11176 60148 11388
rect 61480 11176 61632 11388
rect 62964 11176 63328 11388
rect 59648 11132 60148 11176
rect 61132 11132 61632 11176
rect 62828 11132 63328 11176
rect 58300 11068 58344 11132
rect 58408 11068 58664 11132
rect 59572 11068 59616 11132
rect 59680 11068 60148 11132
rect 61056 11068 61100 11132
rect 61164 11068 61632 11132
rect 62752 11068 62796 11132
rect 62860 11068 63328 11132
rect 58300 11024 58664 11068
rect 59648 11024 60148 11068
rect 61132 11024 61632 11068
rect 62828 11024 63328 11068
rect 64448 11132 64812 11388
rect 66144 11176 66296 11388
rect 67628 11176 67992 11388
rect 69112 11176 69476 11388
rect 65796 11132 66296 11176
rect 67492 11132 67992 11176
rect 68976 11132 69476 11176
rect 64448 11068 64492 11132
rect 64556 11068 64812 11132
rect 65720 11068 65764 11132
rect 65828 11068 66296 11132
rect 67416 11068 67460 11132
rect 67524 11068 67992 11132
rect 68900 11068 68944 11132
rect 69008 11068 69476 11132
rect 64448 11024 64812 11068
rect 65796 11024 66296 11068
rect 67492 11024 67992 11068
rect 68976 11024 69476 11068
rect 70808 11132 70960 11388
rect 70808 11068 70852 11132
rect 70916 11068 70960 11132
rect 70808 11024 70960 11068
rect 72292 11132 72656 11388
rect 72292 11068 72336 11132
rect 72400 11068 72656 11132
rect 72292 11024 72656 11068
rect 73988 11132 74140 11388
rect 75472 11176 75624 11388
rect 75124 11132 77956 11176
rect 73988 11068 74032 11132
rect 74096 11068 74140 11132
rect 75048 11068 75092 11132
rect 75156 11068 77848 11132
rect 77912 11068 77956 11132
rect 73988 11024 74140 11068
rect 75124 11024 77956 11068
rect 18444 10920 76472 10964
rect 18444 10856 18488 10920
rect 18552 10856 75516 10920
rect 75580 10856 76472 10920
rect 18074 10776 18206 10779
rect 18444 10776 76472 10856
rect 76654 10776 76786 10779
rect 18074 10774 76786 10776
rect 18074 10718 18112 10774
rect 18168 10718 76692 10774
rect 76748 10718 76786 10774
rect 18074 10716 76786 10718
rect 18074 10713 18206 10716
rect 18444 10600 26440 10716
rect 26712 10712 27076 10716
rect 26712 10656 26909 10712
rect 26965 10708 27076 10712
rect 26965 10656 26968 10708
rect 26712 10647 26968 10656
rect 26712 10600 26864 10647
rect 26924 10644 26968 10647
rect 27032 10644 27076 10708
rect 26924 10600 27076 10644
rect 27136 10712 27288 10716
rect 27136 10708 27181 10712
rect 27237 10708 27288 10712
rect 27136 10644 27180 10708
rect 27244 10644 27288 10708
rect 27136 10600 27288 10644
rect 27348 10600 28136 10716
rect 28408 10712 28560 10716
rect 28408 10708 28465 10712
rect 28408 10644 28452 10708
rect 28521 10656 28560 10712
rect 28516 10644 28560 10656
rect 28408 10600 28560 10644
rect 28620 10712 28984 10716
rect 28620 10708 28737 10712
rect 28620 10644 28664 10708
rect 28728 10656 28737 10708
rect 28793 10656 28984 10712
rect 28728 10647 28984 10656
rect 28728 10644 28772 10647
rect 28620 10600 28772 10644
rect 28832 10600 28984 10647
rect 29044 10600 29620 10716
rect 29892 10712 30468 10716
rect 29892 10708 30021 10712
rect 29892 10644 29936 10708
rect 30000 10656 30021 10708
rect 30077 10656 30293 10712
rect 30349 10708 30468 10712
rect 30349 10656 30360 10708
rect 30000 10647 30360 10656
rect 30000 10644 30044 10647
rect 29892 10600 30044 10644
rect 30104 10600 30256 10647
rect 30316 10644 30360 10647
rect 30424 10644 30468 10708
rect 30316 10600 30468 10644
rect 30740 10600 31104 10716
rect 31376 10712 31740 10716
rect 31376 10656 31577 10712
rect 31633 10708 31740 10712
rect 31376 10647 31632 10656
rect 31376 10600 31528 10647
rect 31588 10644 31632 10647
rect 31696 10644 31740 10708
rect 31588 10600 31740 10644
rect 31800 10712 31952 10716
rect 31800 10708 31849 10712
rect 31905 10708 31952 10712
rect 31800 10644 31844 10708
rect 31908 10644 31952 10708
rect 31800 10600 31952 10644
rect 32012 10600 33012 10716
rect 33072 10712 33648 10716
rect 33072 10656 33133 10712
rect 33189 10708 33405 10712
rect 33189 10656 33328 10708
rect 33072 10644 33328 10656
rect 33392 10656 33405 10708
rect 33461 10708 33648 10712
rect 33461 10656 33540 10708
rect 33392 10647 33540 10656
rect 33392 10644 33436 10647
rect 33072 10600 33436 10644
rect 33496 10644 33540 10647
rect 33604 10644 33648 10708
rect 33496 10600 33648 10644
rect 33708 10600 34284 10716
rect 34556 10712 34920 10716
rect 34556 10708 34689 10712
rect 34556 10644 34600 10708
rect 34664 10656 34689 10708
rect 34745 10656 34920 10712
rect 34664 10647 34920 10656
rect 34923 10712 35132 10716
rect 34923 10656 34961 10712
rect 35017 10708 35132 10712
rect 35017 10656 35024 10708
rect 34923 10647 35024 10656
rect 34664 10644 34708 10647
rect 34556 10600 34708 10644
rect 34768 10600 34920 10647
rect 34980 10644 35024 10647
rect 35088 10644 35132 10708
rect 34980 10600 35132 10644
rect 35192 10600 35980 10716
rect 36040 10712 36404 10716
rect 36040 10708 36245 10712
rect 36040 10644 36084 10708
rect 36148 10656 36245 10708
rect 36301 10656 36404 10712
rect 36148 10647 36404 10656
rect 36148 10644 36192 10647
rect 36040 10600 36192 10644
rect 36252 10600 36404 10647
rect 36464 10712 36616 10716
rect 36464 10708 36517 10712
rect 36464 10644 36508 10708
rect 36573 10656 36616 10712
rect 36572 10644 36616 10656
rect 36464 10600 36616 10644
rect 36676 10600 37676 10716
rect 37736 10712 38312 10716
rect 37736 10656 37801 10712
rect 37857 10708 38073 10712
rect 37857 10656 37992 10708
rect 37736 10644 37992 10656
rect 38056 10656 38073 10708
rect 38129 10708 38312 10712
rect 38129 10656 38204 10708
rect 38056 10647 38204 10656
rect 38056 10644 38100 10647
rect 37736 10600 38100 10644
rect 38160 10644 38204 10647
rect 38268 10644 38312 10708
rect 38160 10600 38312 10644
rect 38372 10600 38948 10716
rect 39220 10712 39584 10716
rect 39220 10656 39357 10712
rect 39413 10708 39584 10712
rect 39413 10656 39476 10708
rect 39220 10647 39476 10656
rect 39220 10600 39372 10647
rect 39432 10644 39476 10647
rect 39540 10644 39584 10708
rect 39591 10712 39796 10716
rect 39591 10656 39629 10712
rect 39685 10708 39796 10712
rect 39685 10656 39688 10708
rect 39591 10647 39688 10656
rect 39432 10600 39584 10644
rect 39644 10644 39688 10647
rect 39752 10644 39796 10708
rect 39644 10600 39796 10644
rect 39856 10600 40432 10716
rect 40704 10712 41068 10716
rect 40704 10708 40913 10712
rect 40704 10644 40748 10708
rect 40812 10656 40913 10708
rect 40969 10656 41068 10712
rect 40812 10647 41068 10656
rect 40812 10644 40856 10647
rect 40704 10600 40856 10644
rect 40916 10600 41068 10647
rect 41128 10712 41280 10716
rect 41128 10708 41185 10712
rect 41128 10644 41172 10708
rect 41241 10656 41280 10712
rect 41236 10644 41280 10656
rect 41128 10600 41280 10644
rect 41340 10600 42128 10716
rect 42400 10712 42563 10716
rect 42400 10708 42469 10712
rect 42400 10644 42444 10708
rect 42525 10656 42563 10712
rect 42508 10647 42563 10656
rect 42612 10712 42976 10716
rect 42612 10708 42741 10712
rect 42508 10644 42552 10647
rect 42400 10600 42552 10644
rect 42612 10644 42656 10708
rect 42720 10656 42741 10708
rect 42797 10656 42976 10712
rect 42720 10647 42976 10656
rect 42720 10644 42764 10647
rect 42612 10600 42764 10644
rect 42824 10600 42976 10647
rect 43036 10600 43612 10716
rect 43884 10712 44248 10716
rect 43884 10656 44025 10712
rect 44081 10708 44248 10712
rect 44081 10656 44140 10708
rect 43884 10647 44140 10656
rect 43884 10600 44036 10647
rect 44096 10644 44140 10647
rect 44204 10644 44248 10708
rect 44259 10712 44460 10716
rect 44259 10656 44297 10712
rect 44353 10708 44460 10712
rect 44259 10647 44352 10656
rect 44096 10600 44248 10644
rect 44308 10644 44352 10647
rect 44416 10644 44460 10708
rect 44308 10600 44460 10644
rect 44520 10600 45096 10716
rect 45368 10712 45732 10716
rect 45368 10708 45581 10712
rect 45368 10644 45412 10708
rect 45476 10656 45581 10708
rect 45637 10656 45732 10712
rect 45476 10647 45732 10656
rect 45476 10644 45520 10647
rect 45368 10600 45520 10644
rect 45580 10600 45732 10647
rect 45792 10712 46156 10716
rect 45792 10656 45853 10712
rect 45909 10708 46156 10712
rect 45909 10656 46048 10708
rect 45792 10647 46048 10656
rect 45792 10600 45944 10647
rect 46004 10644 46048 10647
rect 46112 10644 46156 10708
rect 46004 10600 46156 10644
rect 46428 10600 46792 10716
rect 47064 10712 47231 10716
rect 47064 10708 47137 10712
rect 47064 10644 47108 10708
rect 47193 10656 47231 10712
rect 47172 10647 47231 10656
rect 47276 10712 47640 10716
rect 47276 10708 47409 10712
rect 47172 10644 47216 10647
rect 47064 10600 47216 10644
rect 47276 10644 47320 10708
rect 47384 10656 47409 10708
rect 47465 10656 47640 10712
rect 47384 10647 47640 10656
rect 47384 10644 47428 10647
rect 47276 10600 47428 10644
rect 47488 10600 47640 10647
rect 47700 10600 48276 10716
rect 48548 10712 48912 10716
rect 48548 10656 48693 10712
rect 48749 10708 48912 10712
rect 48749 10656 48804 10708
rect 48548 10647 48804 10656
rect 48548 10600 48700 10647
rect 48760 10644 48804 10647
rect 48868 10644 48912 10708
rect 48927 10712 49124 10716
rect 48927 10656 48965 10712
rect 49021 10708 49124 10712
rect 48927 10647 49016 10656
rect 48760 10600 48912 10644
rect 48972 10644 49016 10647
rect 49080 10644 49124 10708
rect 48972 10600 49124 10644
rect 49184 10600 49760 10716
rect 50032 10712 50396 10716
rect 50032 10708 50249 10712
rect 50032 10644 50076 10708
rect 50140 10656 50249 10708
rect 50305 10656 50396 10712
rect 50140 10647 50396 10656
rect 50140 10644 50184 10647
rect 50032 10600 50184 10644
rect 50244 10600 50396 10647
rect 50456 10712 50820 10716
rect 50456 10708 50521 10712
rect 50456 10644 50500 10708
rect 50577 10656 50820 10712
rect 50564 10647 50820 10656
rect 50564 10644 50608 10647
rect 50456 10600 50608 10644
rect 50668 10600 50820 10647
rect 51092 10708 76472 10716
rect 76654 10713 76786 10716
rect 51092 10644 76364 10708
rect 76428 10644 76472 10708
rect 51092 10600 76472 10644
rect 23956 10328 24320 10540
rect 23956 10176 26864 10328
rect 18074 10037 18206 10040
rect 26180 10037 26312 10040
rect 18074 10035 26312 10037
rect 18074 9979 18112 10035
rect 18168 9979 26218 10035
rect 26274 9979 26312 10035
rect 18074 9977 26312 9979
rect 18074 9974 18206 9977
rect 26180 9974 26312 9977
rect 26712 9904 26864 10176
rect 27136 9964 28348 10116
rect 27136 9904 27288 9964
rect 28196 9904 28348 9964
rect 28408 10072 28984 10116
rect 28408 10008 28876 10072
rect 28940 10008 28984 10072
rect 28408 9964 28984 10008
rect 29892 10072 30892 10116
rect 29892 10008 30784 10072
rect 30848 10008 30892 10072
rect 29892 9964 30892 10008
rect 31588 10072 32164 10116
rect 31588 10008 32056 10072
rect 32120 10008 32164 10072
rect 31588 9964 32164 10008
rect 33284 9964 34708 10116
rect 28408 9904 28560 9964
rect 29892 9904 30044 9964
rect 31588 9904 31740 9964
rect 33284 9904 33436 9964
rect 34556 9904 34708 9964
rect 36464 9964 37676 10116
rect 36464 9904 36616 9964
rect 37524 9904 37676 9964
rect 37948 9964 39372 10116
rect 37948 9904 38100 9964
rect 39220 9904 39372 9964
rect 39644 9964 40856 10116
rect 39644 9904 39796 9964
rect 40704 9904 40856 9964
rect 42400 10072 43188 10116
rect 42400 10008 43080 10072
rect 43144 10008 43188 10072
rect 42400 9964 43188 10008
rect 44096 9964 45520 10116
rect 42400 9904 42552 9964
rect 44096 9904 44248 9964
rect 45368 9904 45520 9964
rect 47276 9964 48700 10116
rect 47276 9904 47428 9964
rect 48548 9904 48700 9964
rect 51940 9964 53364 10116
rect 51940 9904 52092 9964
rect 53212 9904 53364 9964
rect 64236 9964 65660 10116
rect 64236 9904 64388 9964
rect 65508 9904 65660 9964
rect 73776 9964 74988 10116
rect 73776 9904 73928 9964
rect 74836 9904 74988 9964
rect 26712 9860 27500 9904
rect 26712 9796 27392 9860
rect 27456 9796 27500 9860
rect 26712 9752 27500 9796
rect 28196 9860 33860 9904
rect 28196 9796 33752 9860
rect 33816 9796 33860 9860
rect 28196 9752 33860 9796
rect 34556 9860 36828 9904
rect 34556 9796 36720 9860
rect 36784 9796 36828 9860
rect 34556 9752 36828 9796
rect 37524 9860 38524 9904
rect 37524 9796 38416 9860
rect 38480 9796 38524 9860
rect 37524 9752 38524 9796
rect 39220 9860 40008 9904
rect 39220 9796 39900 9860
rect 39964 9796 40008 9860
rect 39220 9752 40008 9796
rect 40704 9860 44672 9904
rect 40704 9796 44564 9860
rect 44628 9796 44672 9860
rect 40704 9752 44672 9796
rect 45368 9860 47640 9904
rect 45368 9796 45624 9860
rect 45688 9796 47532 9860
rect 47596 9796 47640 9860
rect 45368 9752 47640 9796
rect 48548 9860 52304 9904
rect 48548 9796 48592 9860
rect 48656 9796 50288 9860
rect 50352 9796 52196 9860
rect 52260 9796 52304 9860
rect 48548 9752 52304 9796
rect 53212 9860 74140 9904
rect 53212 9796 53680 9860
rect 53744 9796 54952 9860
rect 55016 9796 56436 9860
rect 56500 9796 58344 9860
rect 58408 9796 59616 9860
rect 59680 9796 61100 9860
rect 61164 9796 62796 9860
rect 62860 9796 64492 9860
rect 64556 9796 65764 9860
rect 65828 9796 67460 9860
rect 67524 9796 68944 9860
rect 69008 9796 70852 9860
rect 70916 9796 72336 9860
rect 72400 9796 74032 9860
rect 74096 9796 74140 9860
rect 53212 9752 74140 9796
rect 74836 9860 75624 9904
rect 74836 9796 75092 9860
rect 75156 9796 75624 9860
rect 74836 9752 75624 9796
rect 34556 9692 34708 9752
rect 44308 9692 44460 9752
rect 45368 9692 45520 9752
rect 23956 9648 24320 9692
rect 23956 9584 24212 9648
rect 24276 9584 24320 9648
rect 23956 9328 24320 9584
rect 34556 9648 35344 9692
rect 34556 9584 35236 9648
rect 35300 9584 35344 9648
rect 34556 9540 35344 9584
rect 44308 9540 45520 9692
rect 27136 8376 79016 8420
rect 27136 8312 76364 8376
rect 76428 8312 78908 8376
rect 78972 8312 79016 8376
rect 27136 8268 79016 8312
rect 2544 7952 2696 7996
rect 2544 7888 2588 7952
rect 2652 7888 2696 7952
rect 2544 7844 2696 7888
rect 2546 7825 2678 7844
rect 2753 7644 2885 7653
rect 2753 7588 2791 7644
rect 2847 7588 2885 7644
rect 2753 7579 2885 7588
rect 2968 7429 6512 7572
rect 2968 7420 6313 7429
rect 2968 7360 3120 7420
rect 0 7208 3120 7360
rect 6148 7373 6313 7420
rect 6369 7373 6512 7429
rect 6148 7208 6512 7373
rect 2546 6936 2678 7061
rect 1908 6892 2696 6936
rect 1908 6828 1952 6892
rect 2016 6828 2696 6892
rect 1908 6784 2696 6828
rect 2753 6460 2885 6469
rect 2753 6404 2791 6460
rect 2847 6404 2885 6460
rect 2753 6395 2885 6404
rect 26712 6300 26864 6512
rect 27348 6300 27712 6512
rect 28196 6300 28560 6512
rect 29044 6300 29196 6512
rect 29680 6360 32376 6512
rect 29680 6300 30044 6360
rect 848 6256 2696 6300
rect 848 6192 892 6256
rect 956 6192 2588 6256
rect 2652 6192 2696 6256
rect 848 6148 2696 6192
rect 26712 6148 30044 6300
rect 30528 6148 30892 6360
rect 31376 6148 31528 6360
rect 32012 6300 32376 6360
rect 32860 6360 33860 6512
rect 32860 6300 33224 6360
rect 32012 6148 33224 6300
rect 33708 6300 33860 6360
rect 34344 6360 35556 6512
rect 34344 6300 34708 6360
rect 33708 6148 34708 6300
rect 35192 6300 35556 6360
rect 36040 6300 36192 6512
rect 36676 6300 37040 6512
rect 37524 6300 37888 6512
rect 38372 6300 38524 6512
rect 39008 6360 40856 6512
rect 39008 6300 39372 6360
rect 35192 6148 39372 6300
rect 39856 6148 40220 6360
rect 40704 6300 40856 6360
rect 41340 6300 41704 6512
rect 42188 6360 43188 6512
rect 42188 6300 42552 6360
rect 40704 6148 42552 6300
rect 43036 6300 43188 6360
rect 43672 6300 44036 6512
rect 44520 6300 44884 6512
rect 45368 6300 45520 6512
rect 46004 6300 46368 6512
rect 46852 6300 47216 6512
rect 47700 6360 49548 6512
rect 47700 6300 47852 6360
rect 43036 6148 47852 6300
rect 48336 6348 48614 6360
rect 48336 6148 48488 6348
rect 49184 6300 49548 6360
rect 50032 6360 51032 6512
rect 50032 6300 50184 6360
rect 49184 6148 50184 6300
rect 50880 6300 51032 6360
rect 51516 6360 53364 6512
rect 51516 6300 51880 6360
rect 50880 6148 51880 6300
rect 52364 6148 52516 6360
rect 53212 6300 53364 6360
rect 53848 6300 54212 6512
rect 54696 6300 54848 6512
rect 55544 6300 55696 6512
rect 56180 6300 56544 6512
rect 57028 6300 57180 6512
rect 57876 6360 58876 6512
rect 57876 6300 58028 6360
rect 53212 6148 58028 6300
rect 58512 6300 58876 6360
rect 59360 6300 59512 6512
rect 60208 6360 61844 6512
rect 60208 6300 60360 6360
rect 58512 6148 60360 6300
rect 60844 6148 61208 6360
rect 61692 6300 61844 6360
rect 62540 6360 63540 6512
rect 62540 6300 62692 6360
rect 61692 6148 62692 6300
rect 63176 6300 63540 6360
rect 64024 6300 64176 6512
rect 64872 6300 65024 6512
rect 65508 6360 66720 6512
rect 65508 6300 65872 6360
rect 66442 6348 66720 6360
rect 63176 6148 65872 6300
rect 66568 6300 66720 6348
rect 67204 6300 67356 6512
rect 67840 6360 69688 6512
rect 67840 6300 68204 6360
rect 66568 6148 68204 6300
rect 68688 6148 69052 6360
rect 69536 6300 69688 6360
rect 70172 6360 71384 6512
rect 70172 6300 70536 6360
rect 69536 6148 70536 6300
rect 71020 6300 71384 6360
rect 71868 6300 72020 6512
rect 72504 6300 72868 6512
rect 73352 6360 74352 6512
rect 73352 6300 73716 6360
rect 71020 6148 73716 6300
rect 74200 6300 74352 6360
rect 74836 6360 76048 6512
rect 74836 6300 75200 6360
rect 74200 6148 75200 6300
rect 75684 6300 76048 6360
rect 76532 6468 77956 6512
rect 76532 6404 77848 6468
rect 77912 6404 77956 6468
rect 76532 6360 77956 6404
rect 76532 6300 76684 6360
rect 75684 6148 76684 6300
rect 20140 3544 20504 3756
rect 21624 3544 21988 3756
rect 23108 3544 23472 3756
rect 24592 3604 27924 3756
rect 24592 3544 24956 3604
rect 20140 3500 24956 3544
rect 20140 3436 21880 3500
rect 21944 3436 24956 3500
rect 20140 3392 24956 3436
rect 26076 3392 26440 3604
rect 27560 3392 27924 3604
rect 29044 3544 29408 3756
rect 30528 3544 30892 3756
rect 32012 3544 32376 3756
rect 29044 3500 32376 3544
rect 29044 3436 29300 3500
rect 29364 3436 32376 3500
rect 29044 3392 32376 3436
rect 33496 3604 35344 3756
rect 33496 3500 33860 3604
rect 33496 3436 33752 3500
rect 33816 3436 33860 3500
rect 33496 3392 33860 3436
rect 34980 3392 35344 3604
rect 36464 3544 36828 3756
rect 37948 3544 38312 3756
rect 39432 3544 39796 3756
rect 36464 3500 39796 3544
rect 36464 3436 36720 3500
rect 36784 3436 39796 3500
rect 36464 3392 39796 3436
rect 40916 3544 41280 3756
rect 42400 3604 45732 3756
rect 42400 3544 42764 3604
rect 40916 3392 42764 3544
rect 43884 3392 44248 3604
rect 45368 3500 45732 3604
rect 45368 3436 45624 3500
rect 45688 3436 45732 3500
rect 45368 3392 45732 3436
rect 46852 3604 48700 3756
rect 46852 3392 47216 3604
rect 48336 3544 48700 3604
rect 49820 3604 51668 3756
rect 49820 3544 50184 3604
rect 48336 3500 50184 3544
rect 48336 3436 48592 3500
rect 48656 3436 50184 3500
rect 48336 3392 50184 3436
rect 51304 3392 51668 3604
rect 52788 3544 53152 3756
rect 54272 3544 54636 3756
rect 52788 3500 54636 3544
rect 52788 3436 54316 3500
rect 54380 3436 54636 3500
rect 52788 3392 54636 3436
rect 55756 3604 57604 3756
rect 55756 3392 56120 3604
rect 57240 3544 57604 3604
rect 58724 3604 60572 3756
rect 58724 3544 59088 3604
rect 57240 3500 59088 3544
rect 57240 3436 57496 3500
rect 57560 3436 59088 3500
rect 57240 3392 59088 3436
rect 60208 3544 60572 3604
rect 61692 3544 62056 3756
rect 60208 3392 62056 3544
rect 63176 3544 63540 3756
rect 64660 3604 67992 3756
rect 64660 3544 65024 3604
rect 63176 3392 65024 3544
rect 66144 3392 66508 3604
rect 67628 3500 67992 3604
rect 67628 3436 67672 3500
rect 67736 3436 67992 3500
rect 67628 3392 67992 3436
rect 16508 3104 16640 3107
rect 19716 3104 19868 3120
rect 19928 3104 20080 3120
rect 21200 3104 21352 3120
rect 21412 3104 21564 3120
rect 22684 3104 22836 3120
rect 22896 3104 23048 3120
rect 24168 3104 24320 3120
rect 24380 3104 24532 3120
rect 25652 3104 25804 3120
rect 25864 3104 26016 3120
rect 27136 3104 27288 3120
rect 27348 3104 27500 3120
rect 28620 3104 28772 3120
rect 28832 3104 28984 3120
rect 30104 3104 30256 3120
rect 30316 3104 30468 3120
rect 31588 3104 31740 3120
rect 31800 3104 31952 3120
rect 33072 3104 33224 3120
rect 33284 3104 33436 3120
rect 34556 3104 34708 3120
rect 34768 3104 34920 3120
rect 36040 3104 36192 3120
rect 36252 3104 36404 3120
rect 37524 3104 37676 3120
rect 37736 3104 37888 3120
rect 39008 3104 39160 3120
rect 39220 3104 39372 3120
rect 40492 3104 40644 3120
rect 41976 3104 42128 3120
rect 43460 3104 43612 3120
rect 16508 3102 44816 3104
rect 16508 3046 16546 3102
rect 16602 3076 44816 3102
rect 16602 3046 19760 3076
rect 16508 3044 19760 3046
rect 16508 3041 16640 3044
rect 19716 3012 19760 3044
rect 19824 3044 21244 3076
rect 19824 3040 20080 3044
rect 19716 2984 19801 3012
rect 19857 2984 20080 3040
rect 19716 2975 20080 2984
rect 19716 2968 19868 2975
rect 19928 2968 20080 2975
rect 21200 3012 21244 3044
rect 21308 3044 22728 3076
rect 21308 3040 21564 3044
rect 21200 2984 21283 3012
rect 21339 2984 21564 3040
rect 21200 2975 21564 2984
rect 21200 2968 21352 2975
rect 21412 2968 21564 2975
rect 22684 3012 22728 3044
rect 22792 3044 24212 3076
rect 22792 3040 23048 3044
rect 22684 2984 22765 3012
rect 22821 2984 23048 3040
rect 22684 2975 23048 2984
rect 22684 2968 22836 2975
rect 22896 2968 23048 2975
rect 24168 3012 24212 3044
rect 24276 3044 25696 3076
rect 24276 3040 24532 3044
rect 24168 2984 24247 3012
rect 24303 2984 24532 3040
rect 24168 2975 24532 2984
rect 24168 2968 24320 2975
rect 24380 2968 24532 2975
rect 25652 3012 25696 3044
rect 25760 3044 27392 3076
rect 25760 3040 26016 3044
rect 25652 2984 25729 3012
rect 25785 2984 26016 3040
rect 25652 2975 26016 2984
rect 25652 2968 25804 2975
rect 25864 2968 26016 2975
rect 27136 3040 27392 3044
rect 27136 2984 27211 3040
rect 27267 3012 27392 3040
rect 27456 3044 28876 3076
rect 27456 3012 27500 3044
rect 27267 2984 27500 3012
rect 27136 2975 27500 2984
rect 27136 2968 27288 2975
rect 27348 2968 27500 2975
rect 28620 3040 28876 3044
rect 28620 2984 28693 3040
rect 28749 3012 28876 3040
rect 28940 3044 30148 3076
rect 28940 3012 28984 3044
rect 28749 2984 28984 3012
rect 28620 2975 28984 2984
rect 28620 2968 28772 2975
rect 28832 2968 28984 2975
rect 30104 3012 30148 3044
rect 30212 3044 31844 3076
rect 30212 3040 30468 3044
rect 30104 2984 30175 3012
rect 30231 2984 30468 3040
rect 30104 2975 30468 2984
rect 30104 2968 30256 2975
rect 30316 2968 30468 2975
rect 31588 3040 31844 3044
rect 31588 2984 31657 3040
rect 31713 3012 31844 3040
rect 31908 3044 33116 3076
rect 31908 3012 31952 3044
rect 31713 2984 31952 3012
rect 31588 2975 31952 2984
rect 31588 2968 31740 2975
rect 31800 2968 31952 2975
rect 33072 3012 33116 3044
rect 33180 3044 34812 3076
rect 33180 3040 33436 3044
rect 33072 2984 33139 3012
rect 33195 2984 33436 3040
rect 33072 2975 33436 2984
rect 33072 2968 33224 2975
rect 33284 2968 33436 2975
rect 34556 3040 34812 3044
rect 34556 2984 34621 3040
rect 34677 3012 34812 3040
rect 34876 3044 36296 3076
rect 34876 3012 34920 3044
rect 34677 2984 34920 3012
rect 34556 2975 34920 2984
rect 34556 2968 34708 2975
rect 34768 2968 34920 2975
rect 36040 3040 36296 3044
rect 36040 2984 36103 3040
rect 36159 3012 36296 3040
rect 36360 3044 37780 3076
rect 36360 3012 36404 3044
rect 36159 2984 36404 3012
rect 36040 2975 36404 2984
rect 36040 2968 36192 2975
rect 36252 2968 36404 2975
rect 37524 3040 37780 3044
rect 37524 2984 37585 3040
rect 37641 3012 37780 3040
rect 37844 3044 39264 3076
rect 37844 3012 37888 3044
rect 37641 2984 37888 3012
rect 37524 2975 37888 2984
rect 37524 2968 37676 2975
rect 37736 2968 37888 2975
rect 39008 3040 39264 3044
rect 39008 2984 39067 3040
rect 39123 3012 39264 3040
rect 39328 3044 40536 3076
rect 39328 3012 39372 3044
rect 39123 2984 39372 3012
rect 39008 2975 39372 2984
rect 39008 2968 39160 2975
rect 39220 2968 39372 2975
rect 40492 3012 40536 3044
rect 40600 3044 42020 3076
rect 40600 3040 40644 3044
rect 40492 2984 40549 3012
rect 40605 2984 40644 3040
rect 40492 2968 40644 2984
rect 41976 3012 42020 3044
rect 42084 3044 43504 3076
rect 42084 3040 42128 3044
rect 41976 2984 42031 3012
rect 42087 2984 42128 3040
rect 41976 2968 42128 2984
rect 43460 3012 43504 3044
rect 43568 3044 44816 3076
rect 44944 3076 45096 3120
rect 43568 3040 43612 3044
rect 43460 2984 43513 3012
rect 43569 2984 43612 3040
rect 43460 2968 43612 2984
rect 44944 3012 44988 3076
rect 45052 3012 45096 3076
rect 44944 2984 44995 3012
rect 45051 2984 45096 3012
rect 44944 2968 45096 2984
rect 46428 3076 46580 3120
rect 46428 3012 46472 3076
rect 46536 3012 46580 3076
rect 46428 2984 46477 3012
rect 46533 2984 46580 3012
rect 46428 2968 46580 2984
rect 47912 3076 48064 3120
rect 47912 3012 47956 3076
rect 48020 3012 48064 3076
rect 47912 2984 47959 3012
rect 48015 2984 48064 3012
rect 47912 2968 48064 2984
rect 49396 3076 49548 3120
rect 49396 3012 49440 3076
rect 49504 3012 49548 3076
rect 49396 2984 49441 3012
rect 49497 2984 49548 3012
rect 49396 2968 49548 2984
rect 50880 3076 51032 3120
rect 50880 3040 50924 3076
rect 50880 2984 50923 3040
rect 50988 3012 51032 3076
rect 50979 2984 51032 3012
rect 50880 2968 51032 2984
rect 52364 3076 52516 3120
rect 52364 3040 52408 3076
rect 52364 2984 52405 3040
rect 52472 3012 52516 3076
rect 52461 2984 52516 3012
rect 52364 2968 52516 2984
rect 53848 3076 54000 3120
rect 53848 3040 53892 3076
rect 53848 2984 53887 3040
rect 53956 3012 54000 3076
rect 53943 2984 54000 3012
rect 53848 2968 54000 2984
rect 55120 3049 55272 3120
rect 55332 3076 55484 3120
rect 55332 3049 55376 3076
rect 55120 3040 55376 3049
rect 55120 2984 55369 3040
rect 55440 3012 55484 3076
rect 55425 2984 55484 3012
rect 55120 2975 55484 2984
rect 55120 2968 55272 2975
rect 55332 2968 55484 2975
rect 56604 3049 56756 3120
rect 56816 3076 56968 3120
rect 56816 3049 56860 3076
rect 56604 3040 56860 3049
rect 56604 2984 56851 3040
rect 56924 3012 56968 3076
rect 56907 2984 56968 3012
rect 56604 2975 56968 2984
rect 56604 2968 56756 2975
rect 56816 2968 56968 2975
rect 58088 3076 58240 3120
rect 58088 3012 58132 3076
rect 58196 3049 58240 3076
rect 58300 3049 58452 3120
rect 58196 3040 58452 3049
rect 58196 3012 58333 3040
rect 58088 2984 58333 3012
rect 58389 2984 58452 3040
rect 58088 2975 58452 2984
rect 58088 2968 58240 2975
rect 58300 2968 58452 2975
rect 59572 3049 59724 3120
rect 59784 3076 59936 3120
rect 59784 3049 59828 3076
rect 59572 3040 59828 3049
rect 59572 2984 59815 3040
rect 59892 3012 59936 3076
rect 59871 2984 59936 3012
rect 59572 2975 59936 2984
rect 59572 2968 59724 2975
rect 59784 2968 59936 2975
rect 61056 3049 61208 3120
rect 61268 3076 61420 3120
rect 61268 3049 61312 3076
rect 61056 3040 61312 3049
rect 61056 2984 61297 3040
rect 61376 3012 61420 3076
rect 61353 2984 61420 3012
rect 61056 2975 61420 2984
rect 61056 2968 61208 2975
rect 61268 2968 61420 2975
rect 62540 3076 62692 3120
rect 62540 3012 62584 3076
rect 62648 3049 62692 3076
rect 62752 3049 62904 3120
rect 62648 3040 62904 3049
rect 62648 3012 62779 3040
rect 62540 2984 62779 3012
rect 62835 2984 62904 3040
rect 62540 2975 62904 2984
rect 62540 2968 62692 2975
rect 62752 2968 62904 2975
rect 64024 3049 64176 3120
rect 64236 3076 64388 3120
rect 64236 3049 64280 3076
rect 64024 3040 64280 3049
rect 64024 2984 64261 3040
rect 64344 3012 64388 3076
rect 64317 2984 64388 3012
rect 64024 2975 64388 2984
rect 64024 2968 64176 2975
rect 64236 2968 64388 2975
rect 65508 3049 65660 3120
rect 65720 3076 65872 3120
rect 65720 3049 65764 3076
rect 65508 3040 65764 3049
rect 65508 2984 65743 3040
rect 65828 3012 65872 3076
rect 65799 2984 65872 3012
rect 65508 2975 65872 2984
rect 65508 2968 65660 2975
rect 65720 2968 65872 2975
rect 66992 3049 67144 3120
rect 67204 3076 67356 3120
rect 67204 3049 67248 3076
rect 66992 3040 67248 3049
rect 66992 2984 67225 3040
rect 67312 3012 67356 3076
rect 67281 2984 67356 3012
rect 66992 2975 67356 2984
rect 66992 2968 67144 2975
rect 67204 2968 67356 2975
rect 20140 2756 23472 2908
rect 20140 2544 20504 2756
rect 21624 2544 21988 2756
rect 23108 2696 23472 2756
rect 24592 2696 24956 2908
rect 26076 2696 26440 2908
rect 27560 2696 27924 2908
rect 29044 2864 32588 2908
rect 29044 2800 32480 2864
rect 32544 2800 32588 2864
rect 29044 2756 32588 2800
rect 29044 2696 29408 2756
rect 23108 2544 29408 2696
rect 30528 2544 30892 2756
rect 32012 2696 32376 2756
rect 33496 2696 33860 2908
rect 34980 2756 36828 2908
rect 34980 2696 35344 2756
rect 32012 2544 35344 2696
rect 36464 2696 36828 2756
rect 37948 2756 41280 2908
rect 37948 2696 38312 2756
rect 36464 2544 38312 2696
rect 39432 2544 39796 2756
rect 40916 2696 41280 2756
rect 42400 2696 42764 2908
rect 43884 2696 44248 2908
rect 45368 2756 47216 2908
rect 45368 2696 45732 2756
rect 40916 2544 45732 2696
rect 46852 2696 47216 2756
rect 48336 2696 48700 2908
rect 49820 2696 50184 2908
rect 51304 2756 53152 2908
rect 51304 2696 51668 2756
rect 46852 2544 51668 2696
rect 52788 2696 53152 2756
rect 54272 2756 56120 2908
rect 54272 2696 54636 2756
rect 52788 2544 54636 2696
rect 55756 2696 56120 2756
rect 57240 2756 59088 2908
rect 57240 2696 57604 2756
rect 55756 2544 57604 2696
rect 58724 2696 59088 2756
rect 60208 2756 65024 2908
rect 60208 2696 60572 2756
rect 58724 2544 60572 2696
rect 61692 2544 62056 2756
rect 63176 2544 63540 2756
rect 64660 2696 65024 2756
rect 66144 2696 66508 2908
rect 67628 2696 67992 2908
rect 64660 2544 67992 2696
rect 1484 2016 78380 2060
rect 1484 1952 1528 2016
rect 1592 1952 1740 2016
rect 1804 1952 1952 2016
rect 2016 1952 21880 2016
rect 21944 1952 29300 2016
rect 29364 1952 33752 2016
rect 33816 1952 36720 2016
rect 36784 1952 45624 2016
rect 45688 1952 48592 2016
rect 48656 1952 54316 2016
rect 54380 1952 57496 2016
rect 57560 1952 67672 2016
rect 67736 1952 77848 2016
rect 77912 1952 78060 2016
rect 78124 1952 78272 2016
rect 78336 1952 78380 2016
rect 1484 1804 78380 1952
rect 1484 1740 1528 1804
rect 1592 1740 1740 1804
rect 1804 1740 1952 1804
rect 2016 1740 77848 1804
rect 77912 1740 78060 1804
rect 78124 1740 78272 1804
rect 78336 1740 78380 1804
rect 1484 1592 78380 1740
rect 1484 1528 1528 1592
rect 1592 1528 1740 1592
rect 1804 1528 1952 1592
rect 2016 1528 77848 1592
rect 77912 1528 78060 1592
rect 78124 1528 78272 1592
rect 78336 1528 78380 1592
rect 1484 1484 78380 1528
rect 424 956 79440 1000
rect 424 892 468 956
rect 532 892 680 956
rect 744 892 892 956
rect 956 892 32480 956
rect 32544 892 78908 956
rect 78972 892 79120 956
rect 79184 892 79332 956
rect 79396 892 79440 956
rect 424 744 79440 892
rect 424 680 468 744
rect 532 680 680 744
rect 744 680 892 744
rect 956 680 78908 744
rect 78972 680 79120 744
rect 79184 680 79332 744
rect 79396 680 79440 744
rect 424 532 79440 680
rect 424 468 468 532
rect 532 468 680 532
rect 744 468 892 532
rect 956 468 78908 532
rect 78972 468 79120 532
rect 79184 468 79332 532
rect 79396 468 79440 532
rect 424 424 79440 468
<< via3 >>
rect 468 112828 532 112892
rect 680 112828 744 112892
rect 892 112828 956 112892
rect 78908 112828 78972 112892
rect 79120 112828 79184 112892
rect 79332 112828 79396 112892
rect 468 112616 532 112680
rect 680 112616 744 112680
rect 892 112616 956 112680
rect 78908 112616 78972 112680
rect 79120 112616 79184 112680
rect 79332 112616 79396 112680
rect 468 112404 532 112468
rect 680 112404 744 112468
rect 892 112404 956 112468
rect 26332 112404 26396 112468
rect 78908 112404 78972 112468
rect 79120 112404 79184 112468
rect 79332 112404 79396 112468
rect 1528 111768 1592 111832
rect 1740 111768 1804 111832
rect 1952 111768 2016 111832
rect 77848 111768 77912 111832
rect 78060 111768 78124 111832
rect 78272 111768 78336 111832
rect 1528 111556 1592 111620
rect 1740 111556 1804 111620
rect 1952 111556 2016 111620
rect 77848 111556 77912 111620
rect 78060 111556 78124 111620
rect 78272 111556 78336 111620
rect 1528 111344 1592 111408
rect 1740 111344 1804 111408
rect 1952 111344 2016 111408
rect 24636 111344 24700 111408
rect 77848 111344 77912 111408
rect 78060 111344 78124 111408
rect 78272 111344 78336 111408
rect 26332 110708 26396 110772
rect 24848 110496 24912 110560
rect 24636 109012 24700 109076
rect 26332 109012 26396 109076
rect 24848 107528 24912 107592
rect 26544 107528 26608 107592
rect 26332 106044 26396 106108
rect 26120 105832 26184 105896
rect 26544 104560 26608 104624
rect 24848 104348 24912 104412
rect 24636 102864 24700 102928
rect 26120 102864 26184 102928
rect 24848 101380 24912 101444
rect 26120 101380 26184 101444
rect 24636 99896 24700 99960
rect 24636 99684 24700 99748
rect 26120 98412 26184 98476
rect 24424 98200 24488 98264
rect 24636 96716 24700 96780
rect 24848 96716 24912 96780
rect 24424 95232 24488 95296
rect 26332 95232 26396 95296
rect 24848 93748 24912 93812
rect 26120 93536 26184 93600
rect 26332 92264 26396 92328
rect 24636 90568 24700 90632
rect 26120 90568 26184 90632
rect 26332 88872 26396 88936
rect 24636 87600 24700 87664
rect 26120 87388 26184 87452
rect 26332 86116 26396 86180
rect 24848 85904 24912 85968
rect 26120 84420 26184 84484
rect 26332 84420 26396 84484
rect 24848 82936 24912 83000
rect 26120 82724 26184 82788
rect 26332 81452 26396 81516
rect 26332 81240 26396 81304
rect 26120 79968 26184 80032
rect 26544 79756 26608 79820
rect 26120 78272 26184 78336
rect 26332 78272 26396 78336
rect 26544 76788 26608 76852
rect 24848 76576 24912 76640
rect 26120 75304 26184 75368
rect 24636 75092 24700 75156
rect 24848 73820 24912 73884
rect 24848 73608 24912 73672
rect 24636 72124 24700 72188
rect 26120 72124 26184 72188
rect 24848 70640 24912 70704
rect 26332 70428 26396 70492
rect 26120 69156 26184 69220
rect 26120 68944 26184 69008
rect 26332 67672 26396 67736
rect 26544 67460 26608 67524
rect 26120 65976 26184 66040
rect 26332 65976 26396 66040
rect 26544 64492 26608 64556
rect 26120 64280 26184 64344
rect 26332 63008 26396 63072
rect 26332 62796 26396 62860
rect 26120 61524 26184 61588
rect 24848 61312 24912 61376
rect 26120 59828 26184 59892
rect 26332 59828 26396 59892
rect 24848 58344 24912 58408
rect 24848 58132 24912 58196
rect 26120 56860 26184 56924
rect 26120 56648 26184 56712
rect 24848 55376 24912 55440
rect 24636 55164 24700 55228
rect 26120 53680 26184 53744
rect 26332 53680 26396 53744
rect 24636 52196 24700 52260
rect 26544 51984 26608 52048
rect 26332 50712 26396 50776
rect 26120 50500 26184 50564
rect 20184 49016 20248 49080
rect 26544 49228 26608 49292
rect 24848 49016 24912 49080
rect 19336 47532 19400 47596
rect 24636 47532 24700 47596
rect 26120 47532 26184 47596
rect 20184 46048 20248 46112
rect 24848 46048 24912 46112
rect 20396 45836 20460 45900
rect 24848 45836 24912 45900
rect 19336 44564 19400 44628
rect 20608 44352 20672 44416
rect 24636 44564 24700 44628
rect 26120 44352 26184 44416
rect 20396 43080 20460 43144
rect 20396 42868 20460 42932
rect 24848 42868 24912 42932
rect 24848 42656 24912 42720
rect 19336 41384 19400 41448
rect 20608 41384 20672 41448
rect 24636 41384 24700 41448
rect 26120 41384 26184 41448
rect 20396 40112 20460 40176
rect 20608 39688 20672 39752
rect 24848 39900 24912 39964
rect 26332 39688 26396 39752
rect 19336 38416 19400 38480
rect 24636 38416 24700 38480
rect 24848 38204 24912 38268
rect 20608 36932 20672 36996
rect 20396 36720 20460 36784
rect 26120 36720 26184 36784
rect 26332 36720 26396 36784
rect 24848 35236 24912 35300
rect 20396 33752 20460 33816
rect 20184 33540 20248 33604
rect 26120 33752 26184 33816
rect 26332 33540 26396 33604
rect 20396 32056 20460 32120
rect 24636 32056 24700 32120
rect 20184 30784 20248 30848
rect 20820 30572 20884 30636
rect 26120 30572 26184 30636
rect 26332 30572 26396 30636
rect 20396 29088 20460 29152
rect 20608 29088 20672 29152
rect 24636 29088 24700 29152
rect 24848 29088 24912 29152
rect 20820 27604 20884 27668
rect 20396 27392 20460 27456
rect 26120 27604 26184 27668
rect 24636 27392 24700 27456
rect 20608 26120 20672 26184
rect 20184 25908 20248 25972
rect 24848 26120 24912 26184
rect 26120 25908 26184 25972
rect 19972 24424 20036 24488
rect 20396 24424 20460 24488
rect 24636 24424 24700 24488
rect 26544 24424 26608 24488
rect 19336 22940 19400 23004
rect 20184 22940 20248 23004
rect 26120 22940 26184 23004
rect 26332 22940 26396 23004
rect 19972 21244 20036 21308
rect 26544 21456 26608 21520
rect 24848 21244 24912 21308
rect 17216 20608 17280 20672
rect 19336 19972 19400 20036
rect 26332 19972 26396 20036
rect 17428 19760 17492 19824
rect 24636 19760 24700 19824
rect 17216 19124 17280 19188
rect 17640 18912 17704 18976
rect 24848 18488 24912 18552
rect 17428 18276 17492 18340
rect 19548 18276 19612 18340
rect 24848 18276 24912 18340
rect 17216 18064 17280 18128
rect 17428 17852 17492 17916
rect 19548 17852 19612 17916
rect 17428 17428 17492 17492
rect 17640 17428 17704 17492
rect 17428 17216 17492 17280
rect 24636 16792 24700 16856
rect 26120 16792 26184 16856
rect 17216 16580 17280 16644
rect 17004 16368 17068 16432
rect 16368 15944 16432 16008
rect 17640 15944 17704 16008
rect 17428 15732 17492 15796
rect 17852 15732 17916 15796
rect 17216 15308 17280 15372
rect 17640 15096 17704 15160
rect 24848 15308 24912 15372
rect 26332 15096 26396 15160
rect 17004 14884 17068 14948
rect 17640 14672 17704 14736
rect 18064 14460 18128 14524
rect 16580 14248 16644 14312
rect 17852 14036 17916 14100
rect 17004 13612 17068 13676
rect 26120 13824 26184 13888
rect 27180 13612 27244 13676
rect 17640 13188 17704 13252
rect 16792 12562 16837 12616
rect 16837 12562 16856 12616
rect 16792 12552 16856 12562
rect 18064 12340 18128 12404
rect 18488 12128 18552 12192
rect 24636 12128 24700 12192
rect 26332 12128 26396 12192
rect 75516 11916 75580 11980
rect 24636 11280 24700 11344
rect 27180 11280 27244 11344
rect 24212 11068 24276 11132
rect 27392 11068 27456 11132
rect 28876 11068 28940 11132
rect 30784 11068 30848 11132
rect 32056 11068 32120 11132
rect 33752 11068 33816 11132
rect 35236 11068 35300 11132
rect 36720 11068 36784 11132
rect 38416 11068 38480 11132
rect 39900 11068 39964 11132
rect 43080 11068 43144 11132
rect 44564 11068 44628 11132
rect 45624 11068 45688 11132
rect 47532 11068 47596 11132
rect 48592 11068 48656 11132
rect 50288 11068 50352 11132
rect 52196 11068 52260 11132
rect 53680 11068 53744 11132
rect 54952 11068 55016 11132
rect 56436 11068 56500 11132
rect 58344 11068 58408 11132
rect 59616 11068 59680 11132
rect 61100 11068 61164 11132
rect 62796 11068 62860 11132
rect 64492 11068 64556 11132
rect 65764 11068 65828 11132
rect 67460 11068 67524 11132
rect 68944 11068 69008 11132
rect 70852 11068 70916 11132
rect 72336 11068 72400 11132
rect 74032 11068 74096 11132
rect 75092 11068 75156 11132
rect 77848 11068 77912 11132
rect 18488 10856 18552 10920
rect 75516 10856 75580 10920
rect 26968 10644 27032 10708
rect 27180 10656 27181 10708
rect 27181 10656 27237 10708
rect 27237 10656 27244 10708
rect 27180 10644 27244 10656
rect 28452 10656 28465 10708
rect 28465 10656 28516 10708
rect 28452 10644 28516 10656
rect 28664 10644 28728 10708
rect 29936 10644 30000 10708
rect 30360 10644 30424 10708
rect 31632 10656 31633 10708
rect 31633 10656 31696 10708
rect 31632 10644 31696 10656
rect 31844 10656 31849 10708
rect 31849 10656 31905 10708
rect 31905 10656 31908 10708
rect 31844 10644 31908 10656
rect 33328 10644 33392 10708
rect 33540 10644 33604 10708
rect 34600 10644 34664 10708
rect 35024 10644 35088 10708
rect 36084 10644 36148 10708
rect 36508 10656 36517 10708
rect 36517 10656 36572 10708
rect 36508 10644 36572 10656
rect 37992 10644 38056 10708
rect 38204 10644 38268 10708
rect 39476 10644 39540 10708
rect 39688 10644 39752 10708
rect 40748 10644 40812 10708
rect 41172 10656 41185 10708
rect 41185 10656 41236 10708
rect 41172 10644 41236 10656
rect 42444 10656 42469 10708
rect 42469 10656 42508 10708
rect 42444 10644 42508 10656
rect 42656 10644 42720 10708
rect 44140 10644 44204 10708
rect 44352 10656 44353 10708
rect 44353 10656 44416 10708
rect 44352 10644 44416 10656
rect 45412 10644 45476 10708
rect 46048 10644 46112 10708
rect 47108 10656 47137 10708
rect 47137 10656 47172 10708
rect 47108 10644 47172 10656
rect 47320 10644 47384 10708
rect 48804 10644 48868 10708
rect 49016 10656 49021 10708
rect 49021 10656 49080 10708
rect 49016 10644 49080 10656
rect 50076 10644 50140 10708
rect 50500 10656 50521 10708
rect 50521 10656 50564 10708
rect 50500 10644 50564 10656
rect 76364 10644 76428 10708
rect 28876 10008 28940 10072
rect 30784 10008 30848 10072
rect 32056 10008 32120 10072
rect 43080 10008 43144 10072
rect 27392 9796 27456 9860
rect 33752 9796 33816 9860
rect 36720 9796 36784 9860
rect 38416 9796 38480 9860
rect 39900 9796 39964 9860
rect 44564 9796 44628 9860
rect 45624 9796 45688 9860
rect 47532 9796 47596 9860
rect 48592 9796 48656 9860
rect 50288 9796 50352 9860
rect 52196 9796 52260 9860
rect 53680 9796 53744 9860
rect 54952 9796 55016 9860
rect 56436 9796 56500 9860
rect 58344 9796 58408 9860
rect 59616 9796 59680 9860
rect 61100 9796 61164 9860
rect 62796 9796 62860 9860
rect 64492 9796 64556 9860
rect 65764 9796 65828 9860
rect 67460 9796 67524 9860
rect 68944 9796 69008 9860
rect 70852 9796 70916 9860
rect 72336 9796 72400 9860
rect 74032 9796 74096 9860
rect 75092 9796 75156 9860
rect 24212 9584 24276 9648
rect 35236 9584 35300 9648
rect 76364 8312 76428 8376
rect 78908 8312 78972 8376
rect 2588 7888 2652 7952
rect 1952 6828 2016 6892
rect 892 6192 956 6256
rect 2588 6192 2652 6256
rect 77848 6404 77912 6468
rect 21880 3436 21944 3500
rect 29300 3436 29364 3500
rect 33752 3436 33816 3500
rect 36720 3436 36784 3500
rect 45624 3436 45688 3500
rect 48592 3436 48656 3500
rect 54316 3436 54380 3500
rect 57496 3436 57560 3500
rect 67672 3436 67736 3500
rect 19760 3040 19824 3076
rect 19760 3012 19801 3040
rect 19801 3012 19824 3040
rect 21244 3040 21308 3076
rect 21244 3012 21283 3040
rect 21283 3012 21308 3040
rect 22728 3040 22792 3076
rect 22728 3012 22765 3040
rect 22765 3012 22792 3040
rect 24212 3040 24276 3076
rect 24212 3012 24247 3040
rect 24247 3012 24276 3040
rect 25696 3040 25760 3076
rect 25696 3012 25729 3040
rect 25729 3012 25760 3040
rect 27392 3012 27456 3076
rect 28876 3012 28940 3076
rect 30148 3040 30212 3076
rect 30148 3012 30175 3040
rect 30175 3012 30212 3040
rect 31844 3012 31908 3076
rect 33116 3040 33180 3076
rect 33116 3012 33139 3040
rect 33139 3012 33180 3040
rect 34812 3012 34876 3076
rect 36296 3012 36360 3076
rect 37780 3012 37844 3076
rect 39264 3012 39328 3076
rect 40536 3040 40600 3076
rect 40536 3012 40549 3040
rect 40549 3012 40600 3040
rect 42020 3040 42084 3076
rect 42020 3012 42031 3040
rect 42031 3012 42084 3040
rect 43504 3040 43568 3076
rect 43504 3012 43513 3040
rect 43513 3012 43568 3040
rect 44988 3040 45052 3076
rect 44988 3012 44995 3040
rect 44995 3012 45051 3040
rect 45051 3012 45052 3040
rect 46472 3040 46536 3076
rect 46472 3012 46477 3040
rect 46477 3012 46533 3040
rect 46533 3012 46536 3040
rect 47956 3040 48020 3076
rect 47956 3012 47959 3040
rect 47959 3012 48015 3040
rect 48015 3012 48020 3040
rect 49440 3040 49504 3076
rect 49440 3012 49441 3040
rect 49441 3012 49497 3040
rect 49497 3012 49504 3040
rect 50924 3040 50988 3076
rect 50924 3012 50979 3040
rect 50979 3012 50988 3040
rect 52408 3040 52472 3076
rect 52408 3012 52461 3040
rect 52461 3012 52472 3040
rect 53892 3040 53956 3076
rect 53892 3012 53943 3040
rect 53943 3012 53956 3040
rect 55376 3040 55440 3076
rect 55376 3012 55425 3040
rect 55425 3012 55440 3040
rect 56860 3040 56924 3076
rect 56860 3012 56907 3040
rect 56907 3012 56924 3040
rect 58132 3012 58196 3076
rect 59828 3040 59892 3076
rect 59828 3012 59871 3040
rect 59871 3012 59892 3040
rect 61312 3040 61376 3076
rect 61312 3012 61353 3040
rect 61353 3012 61376 3040
rect 62584 3012 62648 3076
rect 64280 3040 64344 3076
rect 64280 3012 64317 3040
rect 64317 3012 64344 3040
rect 65764 3040 65828 3076
rect 65764 3012 65799 3040
rect 65799 3012 65828 3040
rect 67248 3040 67312 3076
rect 67248 3012 67281 3040
rect 67281 3012 67312 3040
rect 32480 2800 32544 2864
rect 1528 1952 1592 2016
rect 1740 1952 1804 2016
rect 1952 1952 2016 2016
rect 21880 1952 21944 2016
rect 29300 1952 29364 2016
rect 33752 1952 33816 2016
rect 36720 1952 36784 2016
rect 45624 1952 45688 2016
rect 48592 1952 48656 2016
rect 54316 1952 54380 2016
rect 57496 1952 57560 2016
rect 67672 1952 67736 2016
rect 77848 1952 77912 2016
rect 78060 1952 78124 2016
rect 78272 1952 78336 2016
rect 1528 1740 1592 1804
rect 1740 1740 1804 1804
rect 1952 1740 2016 1804
rect 77848 1740 77912 1804
rect 78060 1740 78124 1804
rect 78272 1740 78336 1804
rect 1528 1528 1592 1592
rect 1740 1528 1804 1592
rect 1952 1528 2016 1592
rect 77848 1528 77912 1592
rect 78060 1528 78124 1592
rect 78272 1528 78336 1592
rect 468 892 532 956
rect 680 892 744 956
rect 892 892 956 956
rect 32480 892 32544 956
rect 78908 892 78972 956
rect 79120 892 79184 956
rect 79332 892 79396 956
rect 468 680 532 744
rect 680 680 744 744
rect 892 680 956 744
rect 78908 680 78972 744
rect 79120 680 79184 744
rect 79332 680 79396 744
rect 468 468 532 532
rect 680 468 744 532
rect 892 468 956 532
rect 78908 468 78972 532
rect 79120 468 79184 532
rect 79332 468 79396 532
<< metal4 >>
rect 424 112892 1000 112936
rect 424 112828 468 112892
rect 532 112828 680 112892
rect 744 112828 892 112892
rect 956 112828 1000 112892
rect 424 112680 1000 112828
rect 424 112616 468 112680
rect 532 112616 680 112680
rect 744 112616 892 112680
rect 956 112616 1000 112680
rect 424 112468 1000 112616
rect 78864 112892 79440 112936
rect 78864 112828 78908 112892
rect 78972 112828 79120 112892
rect 79184 112828 79332 112892
rect 79396 112828 79440 112892
rect 78864 112680 79440 112828
rect 78864 112616 78908 112680
rect 78972 112616 79120 112680
rect 79184 112616 79332 112680
rect 79396 112616 79440 112680
rect 424 112404 468 112468
rect 532 112404 680 112468
rect 744 112404 892 112468
rect 956 112404 1000 112468
rect 424 6256 1000 112404
rect 26288 112468 26440 112512
rect 26288 112404 26332 112468
rect 26396 112404 26440 112468
rect 424 6192 892 6256
rect 956 6192 1000 6256
rect 424 956 1000 6192
rect 1484 111832 2060 111876
rect 1484 111768 1528 111832
rect 1592 111768 1740 111832
rect 1804 111768 1952 111832
rect 2016 111768 2060 111832
rect 1484 111620 2060 111768
rect 1484 111556 1528 111620
rect 1592 111556 1740 111620
rect 1804 111556 1952 111620
rect 2016 111556 2060 111620
rect 1484 111408 2060 111556
rect 1484 111344 1528 111408
rect 1592 111344 1740 111408
rect 1804 111344 1952 111408
rect 2016 111344 2060 111408
rect 1484 6892 2060 111344
rect 24592 111408 24744 111452
rect 24592 111344 24636 111408
rect 24700 111344 24744 111408
rect 24592 109076 24744 111344
rect 26288 110772 26440 112404
rect 78864 112468 79440 112616
rect 78864 112404 78908 112468
rect 78972 112404 79120 112468
rect 79184 112404 79332 112468
rect 79396 112404 79440 112468
rect 26288 110740 26332 110772
rect 26318 110708 26332 110740
rect 26396 110740 26440 110772
rect 77804 111832 78380 111876
rect 77804 111768 77848 111832
rect 77912 111768 78060 111832
rect 78124 111768 78272 111832
rect 78336 111768 78380 111832
rect 77804 111620 78380 111768
rect 77804 111556 77848 111620
rect 77912 111556 78060 111620
rect 78124 111556 78272 111620
rect 78336 111556 78380 111620
rect 77804 111408 78380 111556
rect 77804 111344 77848 111408
rect 77912 111344 78060 111408
rect 78124 111344 78272 111408
rect 78336 111344 78380 111408
rect 26396 110708 26410 110740
rect 26318 110694 26410 110708
rect 24592 109044 24636 109076
rect 24622 109012 24636 109044
rect 24700 109044 24744 109076
rect 24804 110560 24956 110604
rect 24804 110496 24848 110560
rect 24912 110496 24956 110560
rect 24700 109012 24714 109044
rect 24622 108998 24714 109012
rect 24804 107592 24956 110496
rect 26318 109076 26410 109090
rect 26318 109044 26332 109076
rect 24804 107560 24848 107592
rect 24834 107528 24848 107560
rect 24912 107560 24956 107592
rect 26288 109012 26332 109044
rect 26396 109044 26410 109076
rect 26396 109012 26440 109044
rect 24912 107528 24926 107560
rect 24834 107514 24926 107528
rect 26288 106108 26440 109012
rect 26288 106044 26332 106108
rect 26396 106044 26440 106108
rect 26288 106000 26440 106044
rect 26500 107592 26652 107636
rect 26500 107528 26544 107592
rect 26608 107528 26652 107592
rect 26076 105896 26228 105940
rect 26076 105832 26120 105896
rect 26184 105832 26228 105896
rect 24804 104412 24956 104456
rect 24804 104348 24848 104412
rect 24912 104348 24956 104412
rect 24592 102928 24744 102972
rect 24592 102864 24636 102928
rect 24700 102864 24744 102928
rect 24592 99960 24744 102864
rect 24804 101444 24956 104348
rect 26076 102928 26228 105832
rect 26500 104624 26652 107528
rect 26500 104592 26544 104624
rect 26530 104560 26544 104592
rect 26608 104592 26652 104624
rect 26608 104560 26622 104592
rect 26530 104546 26622 104560
rect 26076 102896 26120 102928
rect 26106 102864 26120 102896
rect 26184 102896 26228 102928
rect 26184 102864 26198 102896
rect 26106 102850 26198 102864
rect 24804 101412 24848 101444
rect 24834 101380 24848 101412
rect 24912 101412 24956 101444
rect 26106 101444 26198 101458
rect 26106 101412 26120 101444
rect 24912 101380 24926 101412
rect 24834 101366 24926 101380
rect 26076 101380 26120 101412
rect 26184 101412 26198 101444
rect 26184 101380 26228 101412
rect 24592 99928 24636 99960
rect 24622 99896 24636 99928
rect 24700 99928 24744 99960
rect 24700 99896 24714 99928
rect 24622 99882 24714 99896
rect 24592 99748 24744 99792
rect 24592 99684 24636 99748
rect 24700 99684 24744 99748
rect 24410 98264 24502 98278
rect 24410 98232 24424 98264
rect 24380 98200 24424 98232
rect 24488 98232 24502 98264
rect 24488 98200 24532 98232
rect 24380 95296 24532 98200
rect 24592 96780 24744 99684
rect 26076 98476 26228 101380
rect 26076 98412 26120 98476
rect 26184 98412 26228 98476
rect 26076 98368 26228 98412
rect 24592 96748 24636 96780
rect 24622 96716 24636 96748
rect 24700 96748 24744 96780
rect 24834 96780 24926 96794
rect 24834 96748 24848 96780
rect 24700 96716 24714 96748
rect 24622 96702 24714 96716
rect 24804 96716 24848 96748
rect 24912 96748 24926 96780
rect 24912 96716 24956 96748
rect 24380 95232 24424 95296
rect 24488 95232 24532 95296
rect 24380 95188 24532 95232
rect 24804 93812 24956 96716
rect 24804 93748 24848 93812
rect 24912 93748 24956 93812
rect 24804 93704 24956 93748
rect 26288 95296 26440 95340
rect 26288 95232 26332 95296
rect 26396 95232 26440 95296
rect 26106 93600 26198 93614
rect 26106 93568 26120 93600
rect 26076 93536 26120 93568
rect 26184 93568 26198 93600
rect 26184 93536 26228 93568
rect 24622 90632 24714 90646
rect 24622 90600 24636 90632
rect 24592 90568 24636 90600
rect 24700 90600 24714 90632
rect 26076 90632 26228 93536
rect 26288 92328 26440 95232
rect 26288 92296 26332 92328
rect 26318 92264 26332 92296
rect 26396 92296 26440 92328
rect 26396 92264 26410 92296
rect 26318 92250 26410 92264
rect 24700 90568 24744 90600
rect 24592 87664 24744 90568
rect 26076 90568 26120 90632
rect 26184 90568 26228 90632
rect 26076 90524 26228 90568
rect 26318 88936 26410 88950
rect 26318 88904 26332 88936
rect 24592 87600 24636 87664
rect 24700 87600 24744 87664
rect 24592 87556 24744 87600
rect 26288 88872 26332 88904
rect 26396 88904 26410 88936
rect 26396 88872 26440 88904
rect 26076 87452 26228 87496
rect 26076 87388 26120 87452
rect 26184 87388 26228 87452
rect 24834 85968 24926 85982
rect 24834 85936 24848 85968
rect 24804 85904 24848 85936
rect 24912 85936 24926 85968
rect 24912 85904 24956 85936
rect 24804 83000 24956 85904
rect 26076 84484 26228 87388
rect 26288 86180 26440 88872
rect 26288 86116 26332 86180
rect 26396 86116 26440 86180
rect 26288 86072 26440 86116
rect 26076 84452 26120 84484
rect 26106 84420 26120 84452
rect 26184 84452 26228 84484
rect 26318 84484 26410 84498
rect 26318 84452 26332 84484
rect 26184 84420 26198 84452
rect 26106 84406 26198 84420
rect 26288 84420 26332 84452
rect 26396 84452 26410 84484
rect 26396 84420 26440 84452
rect 24804 82936 24848 83000
rect 24912 82936 24956 83000
rect 24804 82892 24956 82936
rect 26106 82788 26198 82802
rect 26106 82756 26120 82788
rect 26076 82724 26120 82756
rect 26184 82756 26198 82788
rect 26184 82724 26228 82756
rect 26076 80032 26228 82724
rect 26288 81516 26440 84420
rect 26288 81452 26332 81516
rect 26396 81452 26440 81516
rect 26288 81408 26440 81452
rect 26076 79968 26120 80032
rect 26184 79968 26228 80032
rect 26076 79924 26228 79968
rect 26288 81304 26440 81348
rect 26288 81240 26332 81304
rect 26396 81240 26440 81304
rect 26106 78336 26198 78350
rect 26106 78304 26120 78336
rect 26076 78272 26120 78304
rect 26184 78304 26198 78336
rect 26288 78336 26440 81240
rect 26288 78304 26332 78336
rect 26184 78272 26228 78304
rect 24804 76640 24956 76684
rect 24804 76576 24848 76640
rect 24912 76576 24956 76640
rect 24622 75156 24714 75170
rect 24622 75124 24636 75156
rect 24592 75092 24636 75124
rect 24700 75124 24714 75156
rect 24700 75092 24744 75124
rect 24592 72188 24744 75092
rect 24804 73884 24956 76576
rect 26076 75368 26228 78272
rect 26318 78272 26332 78304
rect 26396 78304 26440 78336
rect 26500 79820 26652 79864
rect 26500 79756 26544 79820
rect 26608 79756 26652 79820
rect 26396 78272 26410 78304
rect 26318 78258 26410 78272
rect 26500 76852 26652 79756
rect 26500 76820 26544 76852
rect 26530 76788 26544 76820
rect 26608 76820 26652 76852
rect 26608 76788 26622 76820
rect 26530 76774 26622 76788
rect 26076 75304 26120 75368
rect 26184 75304 26228 75368
rect 26076 75260 26228 75304
rect 24804 73852 24848 73884
rect 24834 73820 24848 73852
rect 24912 73852 24956 73884
rect 24912 73820 24926 73852
rect 24834 73806 24926 73820
rect 24834 73672 24926 73686
rect 24834 73640 24848 73672
rect 24592 72124 24636 72188
rect 24700 72124 24744 72188
rect 24592 72080 24744 72124
rect 24804 73608 24848 73640
rect 24912 73640 24926 73672
rect 24912 73608 24956 73640
rect 24804 70704 24956 73608
rect 26106 72188 26198 72202
rect 26106 72156 26120 72188
rect 24804 70640 24848 70704
rect 24912 70640 24956 70704
rect 24804 70596 24956 70640
rect 26076 72124 26120 72156
rect 26184 72156 26198 72188
rect 26184 72124 26228 72156
rect 26076 69220 26228 72124
rect 26318 70492 26410 70506
rect 26318 70460 26332 70492
rect 26076 69156 26120 69220
rect 26184 69156 26228 69220
rect 26076 69112 26228 69156
rect 26288 70428 26332 70460
rect 26396 70460 26410 70492
rect 26396 70428 26440 70460
rect 26076 69008 26228 69052
rect 26076 68944 26120 69008
rect 26184 68944 26228 69008
rect 26076 66040 26228 68944
rect 26288 67736 26440 70428
rect 26288 67672 26332 67736
rect 26396 67672 26440 67736
rect 26288 67628 26440 67672
rect 26530 67524 26622 67538
rect 26530 67492 26544 67524
rect 26500 67460 26544 67492
rect 26608 67492 26622 67524
rect 26608 67460 26652 67492
rect 26076 66008 26120 66040
rect 26106 65976 26120 66008
rect 26184 66008 26228 66040
rect 26318 66040 26410 66054
rect 26318 66008 26332 66040
rect 26184 65976 26198 66008
rect 26106 65962 26198 65976
rect 26288 65976 26332 66008
rect 26396 66008 26410 66040
rect 26396 65976 26440 66008
rect 26076 64344 26228 64388
rect 26076 64280 26120 64344
rect 26184 64280 26228 64344
rect 26076 61588 26228 64280
rect 26288 63072 26440 65976
rect 26500 64556 26652 67460
rect 26500 64492 26544 64556
rect 26608 64492 26652 64556
rect 26500 64448 26652 64492
rect 26288 63008 26332 63072
rect 26396 63008 26440 63072
rect 26288 62964 26440 63008
rect 26076 61556 26120 61588
rect 26106 61524 26120 61556
rect 26184 61556 26228 61588
rect 26288 62860 26440 62904
rect 26288 62796 26332 62860
rect 26396 62796 26440 62860
rect 26184 61524 26198 61556
rect 26106 61510 26198 61524
rect 24804 61376 24956 61420
rect 24804 61312 24848 61376
rect 24912 61312 24956 61376
rect 24804 58408 24956 61312
rect 24804 58376 24848 58408
rect 24834 58344 24848 58376
rect 24912 58376 24956 58408
rect 26076 59892 26228 59936
rect 26076 59828 26120 59892
rect 26184 59828 26228 59892
rect 26288 59892 26440 62796
rect 26288 59860 26332 59892
rect 24912 58344 24926 58376
rect 24834 58330 24926 58344
rect 24804 58196 24956 58240
rect 24804 58132 24848 58196
rect 24912 58132 24956 58196
rect 24804 55440 24956 58132
rect 26076 56924 26228 59828
rect 26318 59828 26332 59860
rect 26396 59860 26440 59892
rect 26396 59828 26410 59860
rect 26318 59814 26410 59828
rect 26076 56892 26120 56924
rect 26106 56860 26120 56892
rect 26184 56892 26228 56924
rect 26184 56860 26198 56892
rect 26106 56846 26198 56860
rect 24804 55408 24848 55440
rect 24834 55376 24848 55408
rect 24912 55408 24956 55440
rect 26076 56712 26228 56756
rect 26076 56648 26120 56712
rect 26184 56648 26228 56712
rect 24912 55376 24926 55408
rect 24834 55362 24926 55376
rect 24592 55228 24744 55272
rect 24592 55164 24636 55228
rect 24700 55164 24744 55228
rect 24592 52260 24744 55164
rect 26076 53744 26228 56648
rect 26076 53712 26120 53744
rect 26106 53680 26120 53712
rect 26184 53712 26228 53744
rect 26318 53744 26410 53758
rect 26318 53712 26332 53744
rect 26184 53680 26198 53712
rect 26106 53666 26198 53680
rect 26288 53680 26332 53712
rect 26396 53712 26410 53744
rect 26396 53680 26440 53712
rect 24592 52228 24636 52260
rect 24622 52196 24636 52228
rect 24700 52228 24744 52260
rect 24700 52196 24714 52228
rect 24622 52182 24714 52196
rect 26288 50776 26440 53680
rect 26530 52048 26622 52062
rect 26530 52016 26544 52048
rect 26288 50712 26332 50776
rect 26396 50712 26440 50776
rect 26288 50668 26440 50712
rect 26500 51984 26544 52016
rect 26608 52016 26622 52048
rect 26608 51984 26652 52016
rect 26076 50564 26228 50608
rect 26076 50500 26120 50564
rect 26184 50500 26228 50564
rect 20140 49080 20292 49124
rect 20140 49016 20184 49080
rect 20248 49016 20292 49080
rect 19322 47596 19414 47610
rect 19322 47564 19336 47596
rect 19292 47532 19336 47564
rect 19400 47564 19414 47596
rect 19400 47532 19444 47564
rect 19292 44628 19444 47532
rect 20140 46112 20292 49016
rect 24804 49080 24956 49124
rect 24804 49016 24848 49080
rect 24912 49016 24956 49080
rect 20140 46080 20184 46112
rect 20170 46048 20184 46080
rect 20248 46080 20292 46112
rect 24592 47596 24744 47640
rect 24592 47532 24636 47596
rect 24700 47532 24744 47596
rect 20248 46048 20262 46080
rect 20170 46034 20262 46048
rect 20382 45900 20474 45914
rect 20382 45868 20396 45900
rect 19292 44564 19336 44628
rect 19400 44564 19444 44628
rect 19292 44520 19444 44564
rect 20352 45836 20396 45868
rect 20460 45868 20474 45900
rect 20460 45836 20504 45868
rect 20352 43144 20504 45836
rect 24592 44628 24744 47532
rect 24804 46112 24956 49016
rect 26076 47596 26228 50500
rect 26500 49292 26652 51984
rect 26500 49228 26544 49292
rect 26608 49228 26652 49292
rect 26500 49184 26652 49228
rect 26076 47564 26120 47596
rect 26106 47532 26120 47564
rect 26184 47564 26228 47596
rect 26184 47532 26198 47564
rect 26106 47518 26198 47532
rect 24804 46080 24848 46112
rect 24834 46048 24848 46080
rect 24912 46080 24956 46112
rect 24912 46048 24926 46080
rect 24834 46034 24926 46048
rect 24834 45900 24926 45914
rect 24834 45868 24848 45900
rect 24592 44596 24636 44628
rect 24622 44564 24636 44596
rect 24700 44596 24744 44628
rect 24804 45836 24848 45868
rect 24912 45868 24926 45900
rect 24912 45836 24956 45868
rect 24700 44564 24714 44596
rect 24622 44550 24714 44564
rect 20594 44416 20686 44430
rect 20594 44384 20608 44416
rect 20352 43080 20396 43144
rect 20460 43080 20504 43144
rect 20352 43036 20504 43080
rect 20564 44352 20608 44384
rect 20672 44384 20686 44416
rect 20672 44352 20716 44384
rect 20352 42932 20504 42976
rect 20352 42868 20396 42932
rect 20460 42868 20504 42932
rect 19292 41448 19444 41492
rect 19292 41384 19336 41448
rect 19400 41384 19444 41448
rect 19292 38480 19444 41384
rect 20352 40176 20504 42868
rect 20564 41448 20716 44352
rect 24804 42932 24956 45836
rect 26106 44416 26198 44430
rect 26106 44384 26120 44416
rect 24804 42868 24848 42932
rect 24912 42868 24956 42932
rect 24804 42824 24956 42868
rect 26076 44352 26120 44384
rect 26184 44384 26198 44416
rect 26184 44352 26228 44384
rect 24804 42720 24956 42764
rect 24804 42656 24848 42720
rect 24912 42656 24956 42720
rect 20564 41384 20608 41448
rect 20672 41384 20716 41448
rect 24622 41448 24714 41462
rect 24622 41416 24636 41448
rect 20564 41340 20716 41384
rect 24592 41384 24636 41416
rect 24700 41416 24714 41448
rect 24700 41384 24744 41416
rect 20352 40144 20396 40176
rect 20382 40112 20396 40144
rect 20460 40144 20504 40176
rect 20460 40112 20474 40144
rect 20382 40098 20474 40112
rect 20594 39752 20686 39766
rect 20594 39720 20608 39752
rect 19292 38448 19336 38480
rect 19322 38416 19336 38448
rect 19400 38448 19444 38480
rect 20564 39688 20608 39720
rect 20672 39720 20686 39752
rect 20672 39688 20716 39720
rect 19400 38416 19414 38448
rect 19322 38402 19414 38416
rect 20564 36996 20716 39688
rect 24592 38480 24744 41384
rect 24804 39964 24956 42656
rect 26076 41448 26228 44352
rect 26076 41384 26120 41448
rect 26184 41384 26228 41448
rect 26076 41340 26228 41384
rect 24804 39932 24848 39964
rect 24834 39900 24848 39932
rect 24912 39932 24956 39964
rect 24912 39900 24926 39932
rect 24834 39886 24926 39900
rect 24592 38416 24636 38480
rect 24700 38416 24744 38480
rect 24592 38372 24744 38416
rect 26288 39752 26440 39796
rect 26288 39688 26332 39752
rect 26396 39688 26440 39752
rect 20564 36932 20608 36996
rect 20672 36932 20716 36996
rect 20564 36888 20716 36932
rect 24804 38268 24956 38312
rect 24804 38204 24848 38268
rect 24912 38204 24956 38268
rect 20382 36784 20474 36798
rect 20382 36752 20396 36784
rect 20352 36720 20396 36752
rect 20460 36752 20474 36784
rect 20460 36720 20504 36752
rect 20352 33816 20504 36720
rect 24804 35300 24956 38204
rect 26106 36784 26198 36798
rect 26106 36752 26120 36784
rect 24804 35268 24848 35300
rect 24834 35236 24848 35268
rect 24912 35268 24956 35300
rect 26076 36720 26120 36752
rect 26184 36752 26198 36784
rect 26288 36784 26440 39688
rect 26288 36752 26332 36784
rect 26184 36720 26228 36752
rect 24912 35236 24926 35268
rect 24834 35222 24926 35236
rect 20352 33752 20396 33816
rect 20460 33752 20504 33816
rect 20352 33708 20504 33752
rect 26076 33816 26228 36720
rect 26318 36720 26332 36752
rect 26396 36752 26440 36784
rect 26396 36720 26410 36752
rect 26318 36706 26410 36720
rect 26076 33752 26120 33816
rect 26184 33752 26228 33816
rect 26076 33708 26228 33752
rect 20170 33604 20262 33618
rect 20170 33572 20184 33604
rect 20140 33540 20184 33572
rect 20248 33572 20262 33604
rect 26288 33604 26440 33648
rect 20248 33540 20292 33572
rect 20140 30848 20292 33540
rect 26288 33540 26332 33604
rect 26396 33540 26440 33604
rect 20140 30784 20184 30848
rect 20248 30784 20292 30848
rect 20140 30740 20292 30784
rect 20352 32120 20504 32164
rect 20352 32056 20396 32120
rect 20460 32056 20504 32120
rect 24622 32120 24714 32134
rect 24622 32088 24636 32120
rect 20352 29152 20504 32056
rect 24592 32056 24636 32088
rect 24700 32088 24714 32120
rect 24700 32056 24744 32088
rect 20806 30636 20898 30650
rect 20806 30604 20820 30636
rect 20776 30572 20820 30604
rect 20884 30604 20898 30636
rect 20884 30572 20928 30604
rect 20352 29120 20396 29152
rect 20382 29088 20396 29120
rect 20460 29120 20504 29152
rect 20594 29152 20686 29166
rect 20594 29120 20608 29152
rect 20460 29088 20474 29120
rect 20382 29074 20474 29088
rect 20564 29088 20608 29120
rect 20672 29120 20686 29152
rect 20672 29088 20716 29120
rect 20352 27456 20504 27500
rect 20352 27392 20396 27456
rect 20460 27392 20504 27456
rect 20140 25972 20292 26016
rect 20140 25908 20184 25972
rect 20248 25908 20292 25972
rect 19958 24488 20050 24502
rect 19958 24456 19972 24488
rect 19928 24424 19972 24456
rect 20036 24456 20050 24488
rect 20036 24424 20080 24456
rect 19292 23004 19444 23048
rect 19292 22940 19336 23004
rect 19400 22940 19444 23004
rect 17202 20672 17294 20686
rect 17202 20640 17216 20672
rect 17172 20608 17216 20640
rect 17280 20640 17294 20672
rect 17280 20608 17324 20640
rect 17172 19188 17324 20608
rect 19292 20036 19444 22940
rect 19928 21308 20080 24424
rect 20140 23004 20292 25908
rect 20352 24488 20504 27392
rect 20564 26184 20716 29088
rect 20776 27668 20928 30572
rect 24592 29152 24744 32056
rect 26076 30636 26228 30680
rect 26076 30572 26120 30636
rect 26184 30572 26228 30636
rect 26288 30636 26440 33540
rect 26288 30604 26332 30636
rect 24592 29088 24636 29152
rect 24700 29088 24744 29152
rect 24834 29152 24926 29166
rect 24834 29120 24848 29152
rect 24592 29044 24744 29088
rect 24804 29088 24848 29120
rect 24912 29120 24926 29152
rect 24912 29088 24956 29120
rect 20776 27604 20820 27668
rect 20884 27604 20928 27668
rect 20776 27560 20928 27604
rect 24622 27456 24714 27470
rect 24622 27424 24636 27456
rect 20564 26120 20608 26184
rect 20672 26120 20716 26184
rect 20564 26076 20716 26120
rect 24592 27392 24636 27424
rect 24700 27424 24714 27456
rect 24700 27392 24744 27424
rect 20352 24456 20396 24488
rect 20382 24424 20396 24456
rect 20460 24456 20504 24488
rect 24592 24488 24744 27392
rect 24804 26184 24956 29088
rect 26076 27668 26228 30572
rect 26318 30572 26332 30604
rect 26396 30604 26440 30636
rect 26396 30572 26410 30604
rect 26318 30558 26410 30572
rect 26076 27636 26120 27668
rect 26106 27604 26120 27636
rect 26184 27636 26228 27668
rect 26184 27604 26198 27636
rect 26106 27590 26198 27604
rect 24804 26120 24848 26184
rect 24912 26120 24956 26184
rect 24804 26076 24956 26120
rect 26106 25972 26198 25986
rect 26106 25940 26120 25972
rect 20460 24424 20474 24456
rect 20382 24410 20474 24424
rect 24592 24424 24636 24488
rect 24700 24424 24744 24488
rect 24592 24380 24744 24424
rect 26076 25908 26120 25940
rect 26184 25940 26198 25972
rect 26184 25908 26228 25940
rect 20140 22972 20184 23004
rect 20170 22940 20184 22972
rect 20248 22972 20292 23004
rect 26076 23004 26228 25908
rect 26500 24488 26652 24532
rect 26500 24424 26544 24488
rect 26608 24424 26652 24488
rect 20248 22940 20262 22972
rect 20170 22926 20262 22940
rect 26076 22940 26120 23004
rect 26184 22940 26228 23004
rect 26076 22896 26228 22940
rect 26288 23004 26440 23048
rect 26288 22940 26332 23004
rect 26396 22940 26440 23004
rect 19928 21244 19972 21308
rect 20036 21244 20080 21308
rect 19928 21200 20080 21244
rect 24804 21308 24956 21352
rect 24804 21244 24848 21308
rect 24912 21244 24956 21308
rect 19292 20004 19336 20036
rect 19322 19972 19336 20004
rect 19400 20004 19444 20036
rect 19400 19972 19414 20004
rect 19322 19958 19414 19972
rect 17414 19824 17506 19838
rect 17414 19792 17428 19824
rect 17172 19124 17216 19188
rect 17280 19124 17324 19188
rect 17172 19080 17324 19124
rect 17384 19760 17428 19792
rect 17492 19792 17506 19824
rect 24622 19824 24714 19838
rect 24622 19792 24636 19824
rect 17492 19760 17536 19792
rect 17384 18340 17536 19760
rect 24592 19760 24636 19792
rect 24700 19792 24714 19824
rect 24700 19760 24744 19792
rect 17384 18276 17428 18340
rect 17492 18276 17536 18340
rect 17384 18232 17536 18276
rect 17596 18976 17748 19020
rect 17596 18912 17640 18976
rect 17704 18912 17748 18976
rect 17172 18128 17324 18172
rect 17172 18064 17216 18128
rect 17280 18064 17324 18128
rect 17172 16644 17324 18064
rect 17384 17916 17536 17960
rect 17384 17852 17428 17916
rect 17492 17852 17536 17916
rect 17384 17492 17536 17852
rect 17384 17460 17428 17492
rect 17414 17428 17428 17460
rect 17492 17460 17536 17492
rect 17596 17492 17748 18912
rect 19504 18340 19656 18384
rect 19504 18276 19548 18340
rect 19612 18276 19656 18340
rect 19504 17916 19656 18276
rect 19504 17884 19548 17916
rect 19534 17852 19548 17884
rect 19612 17884 19656 17916
rect 19612 17852 19626 17884
rect 19534 17838 19626 17852
rect 17596 17460 17640 17492
rect 17492 17428 17506 17460
rect 17414 17414 17506 17428
rect 17626 17428 17640 17460
rect 17704 17460 17748 17492
rect 17704 17428 17718 17460
rect 17626 17414 17718 17428
rect 17414 17280 17506 17294
rect 17414 17248 17428 17280
rect 17172 16612 17216 16644
rect 17202 16580 17216 16612
rect 17280 16612 17324 16644
rect 17384 17216 17428 17248
rect 17492 17248 17506 17280
rect 17492 17216 17536 17248
rect 17280 16580 17294 16612
rect 17202 16566 17294 16580
rect 16990 16432 17082 16446
rect 16990 16400 17004 16432
rect 16960 16368 17004 16400
rect 17068 16400 17082 16432
rect 17068 16368 17112 16400
rect 16354 16008 16446 16022
rect 16354 15976 16368 16008
rect 16324 15944 16368 15976
rect 16432 15976 16446 16008
rect 16432 15944 16476 15976
rect 2574 7952 2666 7966
rect 2574 7920 2588 7952
rect 1484 6828 1952 6892
rect 2016 6828 2060 6892
rect 1484 2016 2060 6828
rect 2544 7888 2588 7920
rect 2652 7920 2666 7952
rect 2652 7888 2696 7920
rect 2544 6256 2696 7888
rect 2544 6192 2588 6256
rect 2652 6192 2696 6256
rect 2544 6148 2696 6192
rect 1484 1952 1528 2016
rect 1592 1952 1740 2016
rect 1804 1952 1952 2016
rect 2016 1952 2060 2016
rect 1484 1804 2060 1952
rect 1484 1740 1528 1804
rect 1592 1740 1740 1804
rect 1804 1740 1952 1804
rect 2016 1740 2060 1804
rect 1484 1592 2060 1740
rect 1484 1528 1528 1592
rect 1592 1528 1740 1592
rect 1804 1528 1952 1592
rect 2016 1528 2060 1592
rect 1484 1484 2060 1528
rect 424 892 468 956
rect 532 892 680 956
rect 744 892 892 956
rect 956 892 1000 956
rect 424 744 1000 892
rect 424 680 468 744
rect 532 680 680 744
rect 744 680 892 744
rect 956 680 1000 744
rect 424 532 1000 680
rect 424 468 468 532
rect 532 468 680 532
rect 744 468 892 532
rect 956 468 1000 532
rect 424 424 1000 468
rect 16324 0 16476 15944
rect 16960 14948 17112 16368
rect 17384 15796 17536 17216
rect 24592 16856 24744 19760
rect 24804 18552 24956 21244
rect 26288 20036 26440 22940
rect 26500 21520 26652 24424
rect 26500 21488 26544 21520
rect 26530 21456 26544 21488
rect 26608 21488 26652 21520
rect 26608 21456 26622 21488
rect 26530 21442 26622 21456
rect 26288 20004 26332 20036
rect 26318 19972 26332 20004
rect 26396 20004 26440 20036
rect 26396 19972 26410 20004
rect 26318 19958 26410 19972
rect 24804 18520 24848 18552
rect 24834 18488 24848 18520
rect 24912 18520 24956 18552
rect 24912 18488 24926 18520
rect 24834 18474 24926 18488
rect 24834 18340 24926 18354
rect 24834 18308 24848 18340
rect 24592 16792 24636 16856
rect 24700 16792 24744 16856
rect 24592 16748 24744 16792
rect 24804 18276 24848 18308
rect 24912 18308 24926 18340
rect 24912 18276 24956 18308
rect 17626 16008 17718 16022
rect 17626 15976 17640 16008
rect 17384 15732 17428 15796
rect 17492 15732 17536 15796
rect 17384 15688 17536 15732
rect 17596 15944 17640 15976
rect 17704 15976 17718 16008
rect 17704 15944 17748 15976
rect 17202 15372 17294 15386
rect 17202 15340 17216 15372
rect 16960 14884 17004 14948
rect 17068 14884 17112 14948
rect 16960 14840 17112 14884
rect 17172 15308 17216 15340
rect 17280 15340 17294 15372
rect 17280 15308 17324 15340
rect 16566 14312 16658 14326
rect 16566 14280 16580 14312
rect 16536 14248 16580 14280
rect 16644 14280 16658 14312
rect 16644 14248 16688 14280
rect 16536 0 16688 14248
rect 16990 13676 17082 13690
rect 16990 13644 17004 13676
rect 16960 13612 17004 13644
rect 17068 13644 17082 13676
rect 17068 13612 17112 13644
rect 16778 12616 16870 12630
rect 16778 12584 16792 12616
rect 16748 12552 16792 12584
rect 16856 12584 16870 12616
rect 16856 12552 16900 12584
rect 16748 0 16900 12552
rect 16960 0 17112 13612
rect 17172 0 17324 15308
rect 17596 15160 17748 15944
rect 17838 15796 17930 15810
rect 17838 15764 17852 15796
rect 17596 15096 17640 15160
rect 17704 15096 17748 15160
rect 17596 15052 17748 15096
rect 17808 15732 17852 15764
rect 17916 15764 17930 15796
rect 17916 15732 17960 15764
rect 17626 14736 17718 14750
rect 17626 14704 17640 14736
rect 17596 14672 17640 14704
rect 17704 14704 17718 14736
rect 17704 14672 17748 14704
rect 17596 13252 17748 14672
rect 17808 14100 17960 15732
rect 24804 15372 24956 18276
rect 26106 16856 26198 16870
rect 26106 16824 26120 16856
rect 24804 15308 24848 15372
rect 24912 15308 24956 15372
rect 24804 15264 24956 15308
rect 26076 16792 26120 16824
rect 26184 16824 26198 16856
rect 26184 16792 26228 16824
rect 17808 14036 17852 14100
rect 17916 14036 17960 14100
rect 17808 13992 17960 14036
rect 18020 14524 18172 14568
rect 18020 14460 18064 14524
rect 18128 14460 18172 14524
rect 17596 13188 17640 13252
rect 17704 13188 17748 13252
rect 17596 13144 17748 13188
rect 18020 12404 18172 14460
rect 26076 13888 26228 16792
rect 26076 13824 26120 13888
rect 26184 13824 26228 13888
rect 26076 13780 26228 13824
rect 26288 15160 26440 15204
rect 26288 15096 26332 15160
rect 26396 15096 26440 15160
rect 18020 12372 18064 12404
rect 18050 12340 18064 12372
rect 18128 12372 18172 12404
rect 18128 12340 18142 12372
rect 18050 12326 18142 12340
rect 18474 12192 18566 12206
rect 18474 12160 18488 12192
rect 18444 12128 18488 12160
rect 18552 12160 18566 12192
rect 24592 12192 24744 12236
rect 18552 12128 18596 12160
rect 18444 10920 18596 12128
rect 24592 12128 24636 12192
rect 24700 12128 24744 12192
rect 26288 12192 26440 15096
rect 27166 13676 27258 13690
rect 27166 13644 27180 13676
rect 26288 12160 26332 12192
rect 24592 11344 24744 12128
rect 26318 12128 26332 12160
rect 26396 12160 26440 12192
rect 27136 13612 27180 13644
rect 27244 13644 27258 13676
rect 27244 13612 27288 13644
rect 26396 12128 26410 12160
rect 26318 12114 26410 12128
rect 24592 11312 24636 11344
rect 24622 11280 24636 11312
rect 24700 11312 24744 11344
rect 27136 11344 27288 13612
rect 24700 11280 24714 11312
rect 24622 11266 24714 11280
rect 27136 11280 27180 11344
rect 27244 11280 27288 11344
rect 27136 11236 27288 11280
rect 75472 11980 75624 12024
rect 75472 11916 75516 11980
rect 75580 11916 75624 11980
rect 24198 11132 24290 11146
rect 24198 11100 24212 11132
rect 18444 10856 18488 10920
rect 18552 10856 18596 10920
rect 18444 10812 18596 10856
rect 24168 11068 24212 11100
rect 24276 11100 24290 11132
rect 27348 11132 27500 11176
rect 24276 11068 24320 11100
rect 24168 9648 24320 11068
rect 27348 11068 27392 11132
rect 27456 11068 27500 11132
rect 26954 10708 27046 10722
rect 26954 10676 26968 10708
rect 24168 9584 24212 9648
rect 24276 9584 24320 9648
rect 24168 9540 24320 9584
rect 26924 10644 26968 10676
rect 27032 10676 27046 10708
rect 27166 10708 27258 10722
rect 27166 10676 27180 10708
rect 27032 10644 27076 10676
rect 21866 3500 21958 3514
rect 21866 3468 21880 3500
rect 21836 3436 21880 3468
rect 21944 3468 21958 3500
rect 21944 3436 21988 3468
rect 19746 3076 19838 3090
rect 19746 3044 19760 3076
rect 19716 3012 19760 3044
rect 19824 3044 19838 3076
rect 21230 3076 21322 3090
rect 21230 3044 21244 3076
rect 19824 3012 19868 3044
rect 19716 0 19868 3012
rect 21200 3012 21244 3044
rect 21308 3044 21322 3076
rect 21308 3012 21352 3044
rect 21200 0 21352 3012
rect 21836 2016 21988 3436
rect 22714 3076 22806 3090
rect 22714 3044 22728 3076
rect 21836 1952 21880 2016
rect 21944 1952 21988 2016
rect 21836 1908 21988 1952
rect 22684 3012 22728 3044
rect 22792 3044 22806 3076
rect 24198 3076 24290 3090
rect 24198 3044 24212 3076
rect 22792 3012 22836 3044
rect 22684 0 22836 3012
rect 24168 3012 24212 3044
rect 24276 3044 24290 3076
rect 25682 3076 25774 3090
rect 25682 3044 25696 3076
rect 24276 3012 24320 3044
rect 24168 0 24320 3012
rect 25652 3012 25696 3044
rect 25760 3044 25774 3076
rect 25760 3012 25804 3044
rect 25652 0 25804 3012
rect 26924 0 27076 10644
rect 27136 10644 27180 10676
rect 27244 10676 27258 10708
rect 27244 10644 27288 10676
rect 27136 0 27288 10644
rect 27348 9860 27500 11068
rect 28832 11132 28984 11176
rect 28832 11068 28876 11132
rect 28940 11068 28984 11132
rect 28438 10708 28530 10722
rect 28438 10676 28452 10708
rect 27348 9828 27392 9860
rect 27378 9796 27392 9828
rect 27456 9828 27500 9860
rect 28408 10644 28452 10676
rect 28516 10676 28530 10708
rect 28650 10708 28742 10722
rect 28650 10676 28664 10708
rect 28516 10644 28560 10676
rect 27456 9796 27470 9828
rect 27378 9782 27470 9796
rect 27378 3076 27470 3090
rect 27378 3044 27392 3076
rect 27348 3012 27392 3044
rect 27456 3044 27470 3076
rect 27456 3012 27500 3044
rect 27348 0 27500 3012
rect 28408 0 28560 10644
rect 28620 10644 28664 10676
rect 28728 10676 28742 10708
rect 28728 10644 28772 10676
rect 28620 0 28772 10644
rect 28832 10072 28984 11068
rect 30740 11132 30892 11176
rect 30740 11068 30784 11132
rect 30848 11068 30892 11132
rect 29922 10708 30014 10722
rect 29922 10676 29936 10708
rect 28832 10040 28876 10072
rect 28862 10008 28876 10040
rect 28940 10040 28984 10072
rect 29892 10644 29936 10676
rect 30000 10676 30014 10708
rect 30346 10708 30438 10722
rect 30346 10676 30360 10708
rect 30000 10644 30044 10676
rect 28940 10008 28954 10040
rect 28862 9994 28954 10008
rect 29286 3500 29378 3514
rect 29286 3468 29300 3500
rect 29256 3436 29300 3468
rect 29364 3468 29378 3500
rect 29364 3436 29408 3468
rect 28862 3076 28954 3090
rect 28862 3044 28876 3076
rect 28832 3012 28876 3044
rect 28940 3044 28954 3076
rect 28940 3012 28984 3044
rect 28832 0 28984 3012
rect 29256 2016 29408 3436
rect 29256 1952 29300 2016
rect 29364 1952 29408 2016
rect 29256 1908 29408 1952
rect 29892 0 30044 10644
rect 30316 10644 30360 10676
rect 30424 10676 30438 10708
rect 30424 10644 30468 10676
rect 30134 3076 30226 3090
rect 30134 3044 30148 3076
rect 30104 3012 30148 3044
rect 30212 3044 30226 3076
rect 30212 3012 30256 3044
rect 30104 0 30256 3012
rect 30316 0 30468 10644
rect 30740 10072 30892 11068
rect 32012 11132 32164 11176
rect 32012 11068 32056 11132
rect 32120 11068 32164 11132
rect 31618 10708 31710 10722
rect 31618 10676 31632 10708
rect 30740 10040 30784 10072
rect 30770 10008 30784 10040
rect 30848 10040 30892 10072
rect 31588 10644 31632 10676
rect 31696 10676 31710 10708
rect 31830 10708 31922 10722
rect 31830 10676 31844 10708
rect 31696 10644 31740 10676
rect 30848 10008 30862 10040
rect 30770 9994 30862 10008
rect 31588 0 31740 10644
rect 31800 10644 31844 10676
rect 31908 10676 31922 10708
rect 31908 10644 31952 10676
rect 31800 3332 31952 10644
rect 32012 10072 32164 11068
rect 33708 11132 33860 11176
rect 33708 11068 33752 11132
rect 33816 11068 33860 11132
rect 33314 10708 33406 10722
rect 33314 10676 33328 10708
rect 32012 10040 32056 10072
rect 32042 10008 32056 10040
rect 32120 10040 32164 10072
rect 33284 10644 33328 10676
rect 33392 10676 33406 10708
rect 33526 10708 33618 10722
rect 33526 10676 33540 10708
rect 33392 10644 33436 10676
rect 32120 10008 32134 10040
rect 32042 9994 32134 10008
rect 31800 3180 32164 3332
rect 31830 3076 31922 3090
rect 31830 3044 31844 3076
rect 31800 3012 31844 3044
rect 31908 3044 31922 3076
rect 31908 3012 31952 3044
rect 31800 0 31952 3012
rect 32012 0 32164 3180
rect 33102 3076 33194 3090
rect 33102 3044 33116 3076
rect 33072 3012 33116 3044
rect 33180 3044 33194 3076
rect 33180 3012 33224 3044
rect 32466 2864 32558 2878
rect 32466 2832 32480 2864
rect 32436 2800 32480 2832
rect 32544 2832 32558 2864
rect 32544 2800 32588 2832
rect 32436 956 32588 2800
rect 32436 892 32480 956
rect 32544 892 32588 956
rect 32436 848 32588 892
rect 33072 0 33224 3012
rect 33284 0 33436 10644
rect 33496 10644 33540 10676
rect 33604 10676 33618 10708
rect 33604 10644 33648 10676
rect 33496 0 33648 10644
rect 33708 9860 33860 11068
rect 35192 11132 35344 11176
rect 35192 11068 35236 11132
rect 35300 11068 35344 11132
rect 34586 10708 34678 10722
rect 34586 10676 34600 10708
rect 33708 9828 33752 9860
rect 33738 9796 33752 9828
rect 33816 9828 33860 9860
rect 34556 10644 34600 10676
rect 34664 10676 34678 10708
rect 35010 10708 35102 10722
rect 35010 10676 35024 10708
rect 34664 10644 34708 10676
rect 33816 9796 33830 9828
rect 33738 9782 33830 9796
rect 33738 3500 33830 3514
rect 33738 3468 33752 3500
rect 33708 3436 33752 3468
rect 33816 3468 33830 3500
rect 33816 3436 33860 3468
rect 33708 2016 33860 3436
rect 33708 1952 33752 2016
rect 33816 1952 33860 2016
rect 33708 1908 33860 1952
rect 34556 0 34708 10644
rect 34980 10644 35024 10676
rect 35088 10676 35102 10708
rect 35088 10644 35132 10676
rect 34798 3076 34890 3090
rect 34798 3044 34812 3076
rect 34768 3012 34812 3044
rect 34876 3044 34890 3076
rect 34876 3012 34920 3044
rect 34768 0 34920 3012
rect 34980 0 35132 10644
rect 35192 9648 35344 11068
rect 36676 11132 36828 11176
rect 36676 11068 36720 11132
rect 36784 11068 36828 11132
rect 36070 10708 36162 10722
rect 36070 10676 36084 10708
rect 35192 9616 35236 9648
rect 35222 9584 35236 9616
rect 35300 9616 35344 9648
rect 36040 10644 36084 10676
rect 36148 10676 36162 10708
rect 36494 10708 36586 10722
rect 36494 10676 36508 10708
rect 36148 10644 36192 10676
rect 35300 9584 35314 9616
rect 35222 9570 35314 9584
rect 36040 0 36192 10644
rect 36464 10644 36508 10676
rect 36572 10676 36586 10708
rect 36572 10644 36616 10676
rect 36282 3076 36374 3090
rect 36282 3044 36296 3076
rect 36252 3012 36296 3044
rect 36360 3044 36374 3076
rect 36360 3012 36404 3044
rect 36252 0 36404 3012
rect 36464 0 36616 10644
rect 36676 9860 36828 11068
rect 38372 11132 38524 11176
rect 38372 11068 38416 11132
rect 38480 11068 38524 11132
rect 37978 10708 38070 10722
rect 37978 10676 37992 10708
rect 36676 9828 36720 9860
rect 36706 9796 36720 9828
rect 36784 9828 36828 9860
rect 37948 10644 37992 10676
rect 38056 10676 38070 10708
rect 38190 10708 38282 10722
rect 38190 10676 38204 10708
rect 38056 10644 38100 10676
rect 36784 9796 36798 9828
rect 36706 9782 36798 9796
rect 36706 3500 36798 3514
rect 36706 3468 36720 3500
rect 36676 3436 36720 3468
rect 36784 3468 36798 3500
rect 36784 3436 36828 3468
rect 36676 2016 36828 3436
rect 37766 3076 37858 3090
rect 37766 3044 37780 3076
rect 36676 1952 36720 2016
rect 36784 1952 36828 2016
rect 36676 1908 36828 1952
rect 37736 3012 37780 3044
rect 37844 3044 37858 3076
rect 37844 3012 37888 3044
rect 37736 0 37888 3012
rect 37948 0 38100 10644
rect 38160 10644 38204 10676
rect 38268 10676 38282 10708
rect 38268 10644 38312 10676
rect 38160 0 38312 10644
rect 38372 9860 38524 11068
rect 39856 11132 40008 11176
rect 39856 11068 39900 11132
rect 39964 11068 40008 11132
rect 39462 10708 39554 10722
rect 39462 10676 39476 10708
rect 38372 9828 38416 9860
rect 38402 9796 38416 9828
rect 38480 9828 38524 9860
rect 39432 10644 39476 10676
rect 39540 10676 39554 10708
rect 39674 10708 39766 10722
rect 39674 10676 39688 10708
rect 39540 10644 39584 10676
rect 38480 9796 38494 9828
rect 38402 9782 38494 9796
rect 39250 3076 39342 3090
rect 39250 3044 39264 3076
rect 39220 3012 39264 3044
rect 39328 3044 39342 3076
rect 39328 3012 39372 3044
rect 39220 0 39372 3012
rect 39432 0 39584 10644
rect 39644 10644 39688 10676
rect 39752 10676 39766 10708
rect 39752 10644 39796 10676
rect 39644 0 39796 10644
rect 39856 9860 40008 11068
rect 43036 11132 43188 11176
rect 43036 11068 43080 11132
rect 43144 11068 43188 11132
rect 40734 10708 40826 10722
rect 40734 10676 40748 10708
rect 39856 9828 39900 9860
rect 39886 9796 39900 9828
rect 39964 9828 40008 9860
rect 40704 10644 40748 10676
rect 40812 10676 40826 10708
rect 41158 10708 41250 10722
rect 41158 10676 41172 10708
rect 40812 10644 40856 10676
rect 39964 9796 39978 9828
rect 39886 9782 39978 9796
rect 40522 3076 40614 3090
rect 40522 3044 40536 3076
rect 40492 3012 40536 3044
rect 40600 3044 40614 3076
rect 40600 3012 40644 3044
rect 40492 0 40644 3012
rect 40704 0 40856 10644
rect 41128 10644 41172 10676
rect 41236 10676 41250 10708
rect 42430 10708 42522 10722
rect 42430 10676 42444 10708
rect 41236 10644 41280 10676
rect 41128 0 41280 10644
rect 42400 10644 42444 10676
rect 42508 10676 42522 10708
rect 42642 10708 42734 10722
rect 42642 10676 42656 10708
rect 42508 10644 42552 10676
rect 42006 3076 42098 3090
rect 42006 3044 42020 3076
rect 41976 3012 42020 3044
rect 42084 3044 42098 3076
rect 42084 3012 42128 3044
rect 41976 0 42128 3012
rect 42400 0 42552 10644
rect 42612 10644 42656 10676
rect 42720 10676 42734 10708
rect 42720 10644 42764 10676
rect 42612 0 42764 10644
rect 43036 10072 43188 11068
rect 44520 11132 44672 11176
rect 44520 11068 44564 11132
rect 44628 11068 44672 11132
rect 44126 10708 44218 10722
rect 44126 10676 44140 10708
rect 43036 10040 43080 10072
rect 43066 10008 43080 10040
rect 43144 10040 43188 10072
rect 44096 10644 44140 10676
rect 44204 10676 44218 10708
rect 44338 10708 44430 10722
rect 44338 10676 44352 10708
rect 44204 10644 44248 10676
rect 43144 10008 43158 10040
rect 43066 9994 43158 10008
rect 43490 3076 43582 3090
rect 43490 3044 43504 3076
rect 43460 3012 43504 3044
rect 43568 3044 43582 3076
rect 43568 3012 43612 3044
rect 43460 0 43612 3012
rect 44096 0 44248 10644
rect 44308 10644 44352 10676
rect 44416 10676 44430 10708
rect 44416 10644 44460 10676
rect 44308 0 44460 10644
rect 44520 9860 44672 11068
rect 45580 11132 45732 11176
rect 45580 11068 45624 11132
rect 45688 11068 45732 11132
rect 45398 10708 45490 10722
rect 45398 10676 45412 10708
rect 44520 9828 44564 9860
rect 44550 9796 44564 9828
rect 44628 9828 44672 9860
rect 45368 10644 45412 10676
rect 45476 10676 45490 10708
rect 45476 10644 45520 10676
rect 44628 9796 44642 9828
rect 44550 9782 44642 9796
rect 44974 3076 45066 3090
rect 44974 3044 44988 3076
rect 44944 3012 44988 3044
rect 45052 3044 45066 3076
rect 45052 3012 45096 3044
rect 44944 0 45096 3012
rect 45368 0 45520 10644
rect 45580 9860 45732 11068
rect 47488 11132 47640 11176
rect 47488 11068 47532 11132
rect 47596 11068 47640 11132
rect 46034 10708 46126 10722
rect 46034 10676 46048 10708
rect 45580 9828 45624 9860
rect 45610 9796 45624 9828
rect 45688 9828 45732 9860
rect 46004 10644 46048 10676
rect 46112 10676 46126 10708
rect 47094 10708 47186 10722
rect 47094 10676 47108 10708
rect 46112 10644 46156 10676
rect 45688 9796 45702 9828
rect 45610 9782 45702 9796
rect 45610 3500 45702 3514
rect 45610 3468 45624 3500
rect 45580 3436 45624 3468
rect 45688 3468 45702 3500
rect 45688 3436 45732 3468
rect 45580 2016 45732 3436
rect 45580 1952 45624 2016
rect 45688 1952 45732 2016
rect 45580 1908 45732 1952
rect 46004 0 46156 10644
rect 47064 10644 47108 10676
rect 47172 10676 47186 10708
rect 47306 10708 47398 10722
rect 47306 10676 47320 10708
rect 47172 10644 47216 10676
rect 46458 3076 46550 3090
rect 46458 3044 46472 3076
rect 46428 3012 46472 3044
rect 46536 3044 46550 3076
rect 46536 3012 46580 3044
rect 46428 0 46580 3012
rect 47064 0 47216 10644
rect 47276 10644 47320 10676
rect 47384 10676 47398 10708
rect 47384 10644 47428 10676
rect 47276 0 47428 10644
rect 47488 9860 47640 11068
rect 47488 9828 47532 9860
rect 47518 9796 47532 9828
rect 47596 9828 47640 9860
rect 48548 11132 48700 11176
rect 48548 11068 48592 11132
rect 48656 11068 48700 11132
rect 48548 9860 48700 11068
rect 50244 11132 50396 11176
rect 50244 11068 50288 11132
rect 50352 11068 50396 11132
rect 48790 10708 48882 10722
rect 48790 10676 48804 10708
rect 48548 9828 48592 9860
rect 47596 9796 47610 9828
rect 47518 9782 47610 9796
rect 48578 9796 48592 9828
rect 48656 9828 48700 9860
rect 48760 10644 48804 10676
rect 48868 10676 48882 10708
rect 49002 10708 49094 10722
rect 49002 10676 49016 10708
rect 48868 10644 48912 10676
rect 48656 9796 48670 9828
rect 48578 9782 48670 9796
rect 48578 3500 48670 3514
rect 48578 3468 48592 3500
rect 48548 3436 48592 3468
rect 48656 3468 48670 3500
rect 48656 3436 48700 3468
rect 47942 3076 48034 3090
rect 47942 3044 47956 3076
rect 47912 3012 47956 3044
rect 48020 3044 48034 3076
rect 48020 3012 48064 3044
rect 47912 0 48064 3012
rect 48548 2016 48700 3436
rect 48548 1952 48592 2016
rect 48656 1952 48700 2016
rect 48548 1908 48700 1952
rect 48760 0 48912 10644
rect 48972 10644 49016 10676
rect 49080 10676 49094 10708
rect 50062 10708 50154 10722
rect 50062 10676 50076 10708
rect 49080 10644 49124 10676
rect 48972 0 49124 10644
rect 50032 10644 50076 10676
rect 50140 10676 50154 10708
rect 50140 10644 50184 10676
rect 49426 3076 49518 3090
rect 49426 3044 49440 3076
rect 49396 3012 49440 3044
rect 49504 3044 49518 3076
rect 49504 3012 49548 3044
rect 49396 0 49548 3012
rect 50032 0 50184 10644
rect 50244 9860 50396 11068
rect 52152 11132 52304 11176
rect 52152 11068 52196 11132
rect 52260 11068 52304 11132
rect 50486 10708 50578 10722
rect 50486 10676 50500 10708
rect 50244 9828 50288 9860
rect 50274 9796 50288 9828
rect 50352 9828 50396 9860
rect 50456 10644 50500 10676
rect 50564 10676 50578 10708
rect 50564 10644 50608 10676
rect 50352 9796 50366 9828
rect 50274 9782 50366 9796
rect 50456 0 50608 10644
rect 52152 9860 52304 11068
rect 52152 9828 52196 9860
rect 52182 9796 52196 9828
rect 52260 9828 52304 9860
rect 53636 11132 53788 11176
rect 53636 11068 53680 11132
rect 53744 11068 53788 11132
rect 53636 9860 53788 11068
rect 53636 9828 53680 9860
rect 52260 9796 52274 9828
rect 52182 9782 52274 9796
rect 53666 9796 53680 9828
rect 53744 9828 53788 9860
rect 54908 11132 55060 11176
rect 54908 11068 54952 11132
rect 55016 11068 55060 11132
rect 54908 9860 55060 11068
rect 54908 9828 54952 9860
rect 53744 9796 53758 9828
rect 53666 9782 53758 9796
rect 54938 9796 54952 9828
rect 55016 9828 55060 9860
rect 56392 11132 56544 11176
rect 56392 11068 56436 11132
rect 56500 11068 56544 11132
rect 56392 9860 56544 11068
rect 56392 9828 56436 9860
rect 55016 9796 55030 9828
rect 54938 9782 55030 9796
rect 56422 9796 56436 9828
rect 56500 9828 56544 9860
rect 58300 11132 58452 11176
rect 58300 11068 58344 11132
rect 58408 11068 58452 11132
rect 58300 9860 58452 11068
rect 58300 9828 58344 9860
rect 56500 9796 56514 9828
rect 56422 9782 56514 9796
rect 58330 9796 58344 9828
rect 58408 9828 58452 9860
rect 59572 11132 59724 11176
rect 59572 11068 59616 11132
rect 59680 11068 59724 11132
rect 59572 9860 59724 11068
rect 59572 9828 59616 9860
rect 58408 9796 58422 9828
rect 58330 9782 58422 9796
rect 59602 9796 59616 9828
rect 59680 9828 59724 9860
rect 61056 11132 61208 11176
rect 61056 11068 61100 11132
rect 61164 11068 61208 11132
rect 61056 9860 61208 11068
rect 61056 9828 61100 9860
rect 59680 9796 59694 9828
rect 59602 9782 59694 9796
rect 61086 9796 61100 9828
rect 61164 9828 61208 9860
rect 62752 11132 62904 11176
rect 62752 11068 62796 11132
rect 62860 11068 62904 11132
rect 62752 9860 62904 11068
rect 62752 9828 62796 9860
rect 61164 9796 61178 9828
rect 61086 9782 61178 9796
rect 62782 9796 62796 9828
rect 62860 9828 62904 9860
rect 64448 11132 64600 11176
rect 64448 11068 64492 11132
rect 64556 11068 64600 11132
rect 64448 9860 64600 11068
rect 64448 9828 64492 9860
rect 62860 9796 62874 9828
rect 62782 9782 62874 9796
rect 64478 9796 64492 9828
rect 64556 9828 64600 9860
rect 65720 11132 65872 11176
rect 65720 11068 65764 11132
rect 65828 11068 65872 11132
rect 65720 9860 65872 11068
rect 65720 9828 65764 9860
rect 64556 9796 64570 9828
rect 64478 9782 64570 9796
rect 65750 9796 65764 9828
rect 65828 9828 65872 9860
rect 67416 11132 67568 11176
rect 67416 11068 67460 11132
rect 67524 11068 67568 11132
rect 67416 9860 67568 11068
rect 67416 9828 67460 9860
rect 65828 9796 65842 9828
rect 65750 9782 65842 9796
rect 67446 9796 67460 9828
rect 67524 9828 67568 9860
rect 68900 11132 69052 11176
rect 68900 11068 68944 11132
rect 69008 11068 69052 11132
rect 68900 9860 69052 11068
rect 68900 9828 68944 9860
rect 67524 9796 67538 9828
rect 67446 9782 67538 9796
rect 68930 9796 68944 9828
rect 69008 9828 69052 9860
rect 70808 11132 70960 11176
rect 70808 11068 70852 11132
rect 70916 11068 70960 11132
rect 70808 9860 70960 11068
rect 70808 9828 70852 9860
rect 69008 9796 69022 9828
rect 68930 9782 69022 9796
rect 70838 9796 70852 9828
rect 70916 9828 70960 9860
rect 72292 11132 72444 11176
rect 72292 11068 72336 11132
rect 72400 11068 72444 11132
rect 72292 9860 72444 11068
rect 72292 9828 72336 9860
rect 70916 9796 70930 9828
rect 70838 9782 70930 9796
rect 72322 9796 72336 9828
rect 72400 9828 72444 9860
rect 73988 11132 74140 11176
rect 73988 11068 74032 11132
rect 74096 11068 74140 11132
rect 73988 9860 74140 11068
rect 73988 9828 74032 9860
rect 72400 9796 72414 9828
rect 72322 9782 72414 9796
rect 74018 9796 74032 9828
rect 74096 9828 74140 9860
rect 75048 11132 75200 11176
rect 75048 11068 75092 11132
rect 75156 11068 75200 11132
rect 75048 9860 75200 11068
rect 75472 10920 75624 11916
rect 75472 10888 75516 10920
rect 75502 10856 75516 10888
rect 75580 10888 75624 10920
rect 77804 11132 78380 111344
rect 77804 11068 77848 11132
rect 77912 11068 78380 11132
rect 75580 10856 75594 10888
rect 75502 10842 75594 10856
rect 76350 10708 76442 10722
rect 76350 10676 76364 10708
rect 75048 9828 75092 9860
rect 74096 9796 74110 9828
rect 74018 9782 74110 9796
rect 75078 9796 75092 9828
rect 75156 9828 75200 9860
rect 76320 10644 76364 10676
rect 76428 10676 76442 10708
rect 76428 10644 76472 10676
rect 75156 9796 75170 9828
rect 75078 9782 75170 9796
rect 76320 8376 76472 10644
rect 76320 8312 76364 8376
rect 76428 8312 76472 8376
rect 76320 8268 76472 8312
rect 77804 6468 78380 11068
rect 77804 6404 77848 6468
rect 77912 6404 78380 6468
rect 54302 3500 54394 3514
rect 54302 3468 54316 3500
rect 54272 3436 54316 3468
rect 54380 3468 54394 3500
rect 57482 3500 57574 3514
rect 57482 3468 57496 3500
rect 54380 3436 54424 3468
rect 50910 3076 51002 3090
rect 50910 3044 50924 3076
rect 50880 3012 50924 3044
rect 50988 3044 51002 3076
rect 52394 3076 52486 3090
rect 52394 3044 52408 3076
rect 50988 3012 51032 3044
rect 50880 0 51032 3012
rect 52364 3012 52408 3044
rect 52472 3044 52486 3076
rect 53878 3076 53970 3090
rect 53878 3044 53892 3076
rect 52472 3012 52516 3044
rect 52364 0 52516 3012
rect 53848 3012 53892 3044
rect 53956 3044 53970 3076
rect 53956 3012 54000 3044
rect 53848 0 54000 3012
rect 54272 2016 54424 3436
rect 57452 3436 57496 3468
rect 57560 3468 57574 3500
rect 67658 3500 67750 3514
rect 67658 3468 67672 3500
rect 57560 3436 57604 3468
rect 55362 3076 55454 3090
rect 55362 3044 55376 3076
rect 54272 1952 54316 2016
rect 54380 1952 54424 2016
rect 54272 1908 54424 1952
rect 55332 3012 55376 3044
rect 55440 3044 55454 3076
rect 56846 3076 56938 3090
rect 56846 3044 56860 3076
rect 55440 3012 55484 3044
rect 55332 0 55484 3012
rect 56816 3012 56860 3044
rect 56924 3044 56938 3076
rect 56924 3012 56968 3044
rect 56816 0 56968 3012
rect 57452 2016 57604 3436
rect 67628 3436 67672 3468
rect 67736 3468 67750 3500
rect 67736 3436 67780 3468
rect 58118 3076 58210 3090
rect 58118 3044 58132 3076
rect 57452 1952 57496 2016
rect 57560 1952 57604 2016
rect 57452 1908 57604 1952
rect 58088 3012 58132 3044
rect 58196 3044 58210 3076
rect 59814 3076 59906 3090
rect 59814 3044 59828 3076
rect 58196 3012 58240 3044
rect 58088 0 58240 3012
rect 59784 3012 59828 3044
rect 59892 3044 59906 3076
rect 61298 3076 61390 3090
rect 61298 3044 61312 3076
rect 59892 3012 59936 3044
rect 59784 0 59936 3012
rect 61268 3012 61312 3044
rect 61376 3044 61390 3076
rect 62570 3076 62662 3090
rect 62570 3044 62584 3076
rect 61376 3012 61420 3044
rect 61268 0 61420 3012
rect 62540 3012 62584 3044
rect 62648 3044 62662 3076
rect 64266 3076 64358 3090
rect 64266 3044 64280 3076
rect 62648 3012 62692 3044
rect 62540 0 62692 3012
rect 64236 3012 64280 3044
rect 64344 3044 64358 3076
rect 65750 3076 65842 3090
rect 65750 3044 65764 3076
rect 64344 3012 64388 3044
rect 64236 0 64388 3012
rect 65720 3012 65764 3044
rect 65828 3044 65842 3076
rect 67234 3076 67326 3090
rect 67234 3044 67248 3076
rect 65828 3012 65872 3044
rect 65720 0 65872 3012
rect 67204 3012 67248 3044
rect 67312 3044 67326 3076
rect 67312 3012 67356 3044
rect 67204 0 67356 3012
rect 67628 2016 67780 3436
rect 67628 1952 67672 2016
rect 67736 1952 67780 2016
rect 67628 1908 67780 1952
rect 77804 2016 78380 6404
rect 77804 1952 77848 2016
rect 77912 1952 78060 2016
rect 78124 1952 78272 2016
rect 78336 1952 78380 2016
rect 77804 1804 78380 1952
rect 77804 1740 77848 1804
rect 77912 1740 78060 1804
rect 78124 1740 78272 1804
rect 78336 1740 78380 1804
rect 77804 1592 78380 1740
rect 77804 1528 77848 1592
rect 77912 1528 78060 1592
rect 78124 1528 78272 1592
rect 78336 1528 78380 1592
rect 77804 1484 78380 1528
rect 78864 8376 79440 112404
rect 78864 8312 78908 8376
rect 78972 8312 79440 8376
rect 78864 956 79440 8312
rect 78864 892 78908 956
rect 78972 892 79120 956
rect 79184 892 79332 956
rect 79396 892 79440 956
rect 78864 744 79440 892
rect 78864 680 78908 744
rect 78972 680 79120 744
rect 79184 680 79332 744
rect 79396 680 79440 744
rect 78864 532 79440 680
rect 78864 468 78908 532
rect 78972 468 79120 532
rect 79184 468 79332 532
rect 79396 468 79440 532
rect 78864 424 79440 468
use contact_32  contact_32_0
timestamp 1644969367
transform 1 0 78864 0 1 8298
box 0 0 1 1
use contact_32  contact_32_1
timestamp 1644969367
transform 1 0 32436 0 1 878
box 0 0 1 1
use contact_32  contact_32_2
timestamp 1644969367
transform 1 0 32436 0 1 2786
box 0 0 1 1
use contact_32  contact_32_3
timestamp 1644969367
transform 1 0 26076 0 1 64266
box 0 0 1 1
use contact_32  contact_32_4
timestamp 1644969367
transform 1 0 26076 0 1 61510
box 0 0 1 1
use contact_32  contact_32_5
timestamp 1644969367
transform 1 0 26288 0 1 15082
box 0 0 1 1
use contact_32  contact_32_6
timestamp 1644969367
transform 1 0 26288 0 1 12114
box 0 0 1 1
use contact_32  contact_32_7
timestamp 1644969367
transform 1 0 26500 0 1 49214
box 0 0 1 1
use contact_32  contact_32_8
timestamp 1644969367
transform 1 0 26500 0 1 51970
box 0 0 1 1
use contact_32  contact_32_9
timestamp 1644969367
transform 1 0 26500 0 1 64478
box 0 0 1 1
use contact_32  contact_32_10
timestamp 1644969367
transform 1 0 26500 0 1 67446
box 0 0 1 1
use contact_32  contact_32_11
timestamp 1644969367
transform 1 0 26288 0 1 39674
box 0 0 1 1
use contact_32  contact_32_12
timestamp 1644969367
transform 1 0 26288 0 1 36706
box 0 0 1 1
use contact_32  contact_32_13
timestamp 1644969367
transform 1 0 26076 0 1 33738
box 0 0 1 1
use contact_32  contact_32_14
timestamp 1644969367
transform 1 0 26076 0 1 36706
box 0 0 1 1
use contact_32  contact_32_15
timestamp 1644969367
transform 1 0 26076 0 1 98398
box 0 0 1 1
use contact_32  contact_32_16
timestamp 1644969367
transform 1 0 26076 0 1 101366
box 0 0 1 1
use contact_32  contact_32_17
timestamp 1644969367
transform 1 0 26288 0 1 33526
box 0 0 1 1
use contact_32  contact_32_18
timestamp 1644969367
transform 1 0 26288 0 1 30558
box 0 0 1 1
use contact_32  contact_32_19
timestamp 1644969367
transform 1 0 26500 0 1 107514
box 0 0 1 1
use contact_32  contact_32_20
timestamp 1644969367
transform 1 0 26500 0 1 104546
box 0 0 1 1
use contact_32  contact_32_21
timestamp 1644969367
transform 1 0 26076 0 1 79954
box 0 0 1 1
use contact_32  contact_32_22
timestamp 1644969367
transform 1 0 26076 0 1 82710
box 0 0 1 1
use contact_32  contact_32_23
timestamp 1644969367
transform 1 0 26500 0 1 24410
box 0 0 1 1
use contact_32  contact_32_24
timestamp 1644969367
transform 1 0 26500 0 1 21442
box 0 0 1 1
use contact_32  contact_32_25
timestamp 1644969367
transform 1 0 26288 0 1 112390
box 0 0 1 1
use contact_32  contact_32_26
timestamp 1644969367
transform 1 0 26288 0 1 110694
box 0 0 1 1
use contact_32  contact_32_27
timestamp 1644969367
transform 1 0 26076 0 1 30558
box 0 0 1 1
use contact_32  contact_32_28
timestamp 1644969367
transform 1 0 26076 0 1 27590
box 0 0 1 1
use contact_32  contact_32_29
timestamp 1644969367
transform 1 0 26288 0 1 67658
box 0 0 1 1
use contact_32  contact_32_30
timestamp 1644969367
transform 1 0 26288 0 1 70414
box 0 0 1 1
use contact_32  contact_32_31
timestamp 1644969367
transform 1 0 26500 0 1 79742
box 0 0 1 1
use contact_32  contact_32_32
timestamp 1644969367
transform 1 0 26500 0 1 76774
box 0 0 1 1
use contact_32  contact_32_33
timestamp 1644969367
transform 1 0 26288 0 1 95218
box 0 0 1 1
use contact_32  contact_32_34
timestamp 1644969367
transform 1 0 26288 0 1 92250
box 0 0 1 1
use contact_32  contact_32_35
timestamp 1644969367
transform 1 0 26288 0 1 86102
box 0 0 1 1
use contact_32  contact_32_36
timestamp 1644969367
transform 1 0 26288 0 1 88858
box 0 0 1 1
use contact_32  contact_32_37
timestamp 1644969367
transform 1 0 24804 0 1 61298
box 0 0 1 1
use contact_32  contact_32_38
timestamp 1644969367
transform 1 0 24804 0 1 58330
box 0 0 1 1
use contact_32  contact_32_39
timestamp 1644969367
transform 1 0 24804 0 1 110482
box 0 0 1 1
use contact_32  contact_32_40
timestamp 1644969367
transform 1 0 24804 0 1 107514
box 0 0 1 1
use contact_32  contact_32_41
timestamp 1644969367
transform 1 0 24804 0 1 82922
box 0 0 1 1
use contact_32  contact_32_42
timestamp 1644969367
transform 1 0 24804 0 1 85890
box 0 0 1 1
use contact_32  contact_32_43
timestamp 1644969367
transform 1 0 24804 0 1 58118
box 0 0 1 1
use contact_32  contact_32_44
timestamp 1644969367
transform 1 0 24804 0 1 55362
box 0 0 1 1
use contact_32  contact_32_45
timestamp 1644969367
transform 1 0 24804 0 1 21230
box 0 0 1 1
use contact_32  contact_32_46
timestamp 1644969367
transform 1 0 24804 0 1 18474
box 0 0 1 1
use contact_32  contact_32_47
timestamp 1644969367
transform 1 0 24804 0 1 15294
box 0 0 1 1
use contact_32  contact_32_48
timestamp 1644969367
transform 1 0 24804 0 1 18262
box 0 0 1 1
use contact_32  contact_32_49
timestamp 1644969367
transform 1 0 24804 0 1 70626
box 0 0 1 1
use contact_32  contact_32_50
timestamp 1644969367
transform 1 0 24804 0 1 73594
box 0 0 1 1
use contact_32  contact_32_51
timestamp 1644969367
transform 1 0 24804 0 1 76562
box 0 0 1 1
use contact_32  contact_32_52
timestamp 1644969367
transform 1 0 24804 0 1 73806
box 0 0 1 1
use contact_32  contact_32_53
timestamp 1644969367
transform 1 0 24592 0 1 24410
box 0 0 1 1
use contact_32  contact_32_54
timestamp 1644969367
transform 1 0 24592 0 1 27378
box 0 0 1 1
use contact_32  contact_32_55
timestamp 1644969367
transform 1 0 24592 0 1 55150
box 0 0 1 1
use contact_32  contact_32_56
timestamp 1644969367
transform 1 0 24592 0 1 52182
box 0 0 1 1
use contact_32  contact_32_57
timestamp 1644969367
transform 1 0 24380 0 1 95218
box 0 0 1 1
use contact_32  contact_32_58
timestamp 1644969367
transform 1 0 24380 0 1 98186
box 0 0 1 1
use contact_32  contact_32_59
timestamp 1644969367
transform 1 0 24804 0 1 104334
box 0 0 1 1
use contact_32  contact_32_60
timestamp 1644969367
transform 1 0 24804 0 1 101366
box 0 0 1 1
use contact_32  contact_32_61
timestamp 1644969367
transform 1 0 24804 0 1 42642
box 0 0 1 1
use contact_32  contact_32_62
timestamp 1644969367
transform 1 0 24804 0 1 39886
box 0 0 1 1
use contact_32  contact_32_63
timestamp 1644969367
transform 1 0 24804 0 1 42854
box 0 0 1 1
use contact_32  contact_32_64
timestamp 1644969367
transform 1 0 24804 0 1 45822
box 0 0 1 1
use contact_32  contact_32_65
timestamp 1644969367
transform 1 0 24804 0 1 49002
box 0 0 1 1
use contact_32  contact_32_66
timestamp 1644969367
transform 1 0 24804 0 1 46034
box 0 0 1 1
use contact_32  contact_32_67
timestamp 1644969367
transform 1 0 24592 0 1 12114
box 0 0 1 1
use contact_32  contact_32_68
timestamp 1644969367
transform 1 0 24592 0 1 11266
box 0 0 1 1
use contact_32  contact_32_69
timestamp 1644969367
transform 1 0 24168 0 1 9570
box 0 0 1 1
use contact_32  contact_32_70
timestamp 1644969367
transform 1 0 24168 0 1 11054
box 0 0 1 1
use contact_32  contact_32_71
timestamp 1644969367
transform 1 0 20352 0 1 27378
box 0 0 1 1
use contact_32  contact_32_72
timestamp 1644969367
transform 1 0 20352 0 1 24410
box 0 0 1 1
use contact_32  contact_32_73
timestamp 1644969367
transform 1 0 20776 0 1 27590
box 0 0 1 1
use contact_32  contact_32_74
timestamp 1644969367
transform 1 0 20776 0 1 30558
box 0 0 1 1
use contact_32  contact_32_75
timestamp 1644969367
transform 1 0 20352 0 1 33738
box 0 0 1 1
use contact_32  contact_32_76
timestamp 1644969367
transform 1 0 20352 0 1 36706
box 0 0 1 1
use contact_32  contact_32_77
timestamp 1644969367
transform 1 0 20564 0 1 36918
box 0 0 1 1
use contact_32  contact_32_78
timestamp 1644969367
transform 1 0 20564 0 1 39674
box 0 0 1 1
use contact_32  contact_32_79
timestamp 1644969367
transform 1 0 19928 0 1 21230
box 0 0 1 1
use contact_32  contact_32_80
timestamp 1644969367
transform 1 0 19928 0 1 24410
box 0 0 1 1
use contact_32  contact_32_81
timestamp 1644969367
transform 1 0 20352 0 1 42854
box 0 0 1 1
use contact_32  contact_32_82
timestamp 1644969367
transform 1 0 20352 0 1 40098
box 0 0 1 1
use contact_32  contact_32_83
timestamp 1644969367
transform 1 0 20140 0 1 30770
box 0 0 1 1
use contact_32  contact_32_84
timestamp 1644969367
transform 1 0 20140 0 1 33526
box 0 0 1 1
use contact_32  contact_32_85
timestamp 1644969367
transform 1 0 20352 0 1 43066
box 0 0 1 1
use contact_32  contact_32_86
timestamp 1644969367
transform 1 0 20352 0 1 45822
box 0 0 1 1
use contact_32  contact_32_87
timestamp 1644969367
transform 1 0 20140 0 1 49002
box 0 0 1 1
use contact_32  contact_32_88
timestamp 1644969367
transform 1 0 20140 0 1 46034
box 0 0 1 1
use contact_32  contact_32_89
timestamp 1644969367
transform 1 0 76320 0 1 8298
box 0 0 1 1
use contact_32  contact_32_90
timestamp 1644969367
transform 1 0 76320 0 1 10630
box 0 0 1 1
use contact_32  contact_32_91
timestamp 1644969367
transform 1 0 75472 0 1 11902
box 0 0 1 1
use contact_32  contact_32_92
timestamp 1644969367
transform 1 0 75472 0 1 10842
box 0 0 1 1
use contact_32  contact_32_93
timestamp 1644969367
transform 1 0 18444 0 1 10842
box 0 0 1 1
use contact_32  contact_32_94
timestamp 1644969367
transform 1 0 18444 0 1 12114
box 0 0 1 1
use contact_32  contact_32_95
timestamp 1644969367
transform 1 0 18020 0 1 14446
box 0 0 1 1
use contact_32  contact_32_96
timestamp 1644969367
transform 1 0 18020 0 1 12326
box 0 0 1 1
use contact_32  contact_32_97
timestamp 1644969367
transform 1 0 17172 0 1 19110
box 0 0 1 1
use contact_32  contact_32_98
timestamp 1644969367
transform 1 0 17172 0 1 20594
box 0 0 1 1
use contact_32  contact_32_99
timestamp 1644969367
transform 1 0 17596 0 1 15082
box 0 0 1 1
use contact_32  contact_32_100
timestamp 1644969367
transform 1 0 17596 0 1 15930
box 0 0 1 1
use contact_32  contact_32_101
timestamp 1644969367
transform 1 0 17808 0 1 14022
box 0 0 1 1
use contact_32  contact_32_102
timestamp 1644969367
transform 1 0 17808 0 1 15718
box 0 0 1 1
use contact_32  contact_32_103
timestamp 1644969367
transform 1 0 19504 0 1 18262
box 0 0 1 1
use contact_32  contact_32_104
timestamp 1644969367
transform 1 0 19504 0 1 17838
box 0 0 1 1
use contact_32  contact_32_105
timestamp 1644969367
transform 1 0 17384 0 1 17838
box 0 0 1 1
use contact_32  contact_32_106
timestamp 1644969367
transform 1 0 17384 0 1 17414
box 0 0 1 1
use contact_32  contact_32_107
timestamp 1644969367
transform 1 0 17596 0 1 18898
box 0 0 1 1
use contact_32  contact_32_108
timestamp 1644969367
transform 1 0 17596 0 1 17414
box 0 0 1 1
use contact_32  contact_32_109
timestamp 1644969367
transform 1 0 17384 0 1 15718
box 0 0 1 1
use contact_32  contact_32_110
timestamp 1644969367
transform 1 0 17384 0 1 17202
box 0 0 1 1
use contact_32  contact_32_111
timestamp 1644969367
transform 1 0 848 0 1 6178
box 0 0 1 1
use contact_32  contact_32_112
timestamp 1644969367
transform 1 0 2544 0 1 6178
box 0 0 1 1
use contact_32  contact_32_113
timestamp 1644969367
transform 1 0 2544 0 1 7874
box 0 0 1 1
use contact_32  contact_32_114
timestamp 1644969367
transform 1 0 77804 0 1 6390
box 0 0 1 1
use contact_32  contact_32_115
timestamp 1644969367
transform 1 0 77804 0 1 11054
box 0 0 1 1
use contact_32  contact_32_116
timestamp 1644969367
transform 1 0 75048 0 1 11054
box 0 0 1 1
use contact_32  contact_32_117
timestamp 1644969367
transform 1 0 75048 0 1 9782
box 0 0 1 1
use contact_32  contact_32_118
timestamp 1644969367
transform 1 0 73988 0 1 11054
box 0 0 1 1
use contact_32  contact_32_119
timestamp 1644969367
transform 1 0 73988 0 1 9782
box 0 0 1 1
use contact_32  contact_32_120
timestamp 1644969367
transform 1 0 72292 0 1 11054
box 0 0 1 1
use contact_32  contact_32_121
timestamp 1644969367
transform 1 0 72292 0 1 9782
box 0 0 1 1
use contact_32  contact_32_122
timestamp 1644969367
transform 1 0 70808 0 1 11054
box 0 0 1 1
use contact_32  contact_32_123
timestamp 1644969367
transform 1 0 70808 0 1 9782
box 0 0 1 1
use contact_32  contact_32_124
timestamp 1644969367
transform 1 0 68900 0 1 11054
box 0 0 1 1
use contact_32  contact_32_125
timestamp 1644969367
transform 1 0 68900 0 1 9782
box 0 0 1 1
use contact_32  contact_32_126
timestamp 1644969367
transform 1 0 67628 0 1 1938
box 0 0 1 1
use contact_32  contact_32_127
timestamp 1644969367
transform 1 0 67628 0 1 3422
box 0 0 1 1
use contact_32  contact_32_128
timestamp 1644969367
transform 1 0 67416 0 1 11054
box 0 0 1 1
use contact_32  contact_32_129
timestamp 1644969367
transform 1 0 67416 0 1 9782
box 0 0 1 1
use contact_32  contact_32_130
timestamp 1644969367
transform 1 0 65720 0 1 11054
box 0 0 1 1
use contact_32  contact_32_131
timestamp 1644969367
transform 1 0 65720 0 1 9782
box 0 0 1 1
use contact_32  contact_32_132
timestamp 1644969367
transform 1 0 64448 0 1 11054
box 0 0 1 1
use contact_32  contact_32_133
timestamp 1644969367
transform 1 0 64448 0 1 9782
box 0 0 1 1
use contact_32  contact_32_134
timestamp 1644969367
transform 1 0 62752 0 1 11054
box 0 0 1 1
use contact_32  contact_32_135
timestamp 1644969367
transform 1 0 62752 0 1 9782
box 0 0 1 1
use contact_32  contact_32_136
timestamp 1644969367
transform 1 0 61056 0 1 11054
box 0 0 1 1
use contact_32  contact_32_137
timestamp 1644969367
transform 1 0 61056 0 1 9782
box 0 0 1 1
use contact_32  contact_32_138
timestamp 1644969367
transform 1 0 59572 0 1 11054
box 0 0 1 1
use contact_32  contact_32_139
timestamp 1644969367
transform 1 0 59572 0 1 9782
box 0 0 1 1
use contact_32  contact_32_140
timestamp 1644969367
transform 1 0 58300 0 1 11054
box 0 0 1 1
use contact_32  contact_32_141
timestamp 1644969367
transform 1 0 58300 0 1 9782
box 0 0 1 1
use contact_32  contact_32_142
timestamp 1644969367
transform 1 0 57452 0 1 1938
box 0 0 1 1
use contact_32  contact_32_143
timestamp 1644969367
transform 1 0 57452 0 1 3422
box 0 0 1 1
use contact_32  contact_32_144
timestamp 1644969367
transform 1 0 56392 0 1 11054
box 0 0 1 1
use contact_32  contact_32_145
timestamp 1644969367
transform 1 0 56392 0 1 9782
box 0 0 1 1
use contact_32  contact_32_146
timestamp 1644969367
transform 1 0 54908 0 1 11054
box 0 0 1 1
use contact_32  contact_32_147
timestamp 1644969367
transform 1 0 54908 0 1 9782
box 0 0 1 1
use contact_32  contact_32_148
timestamp 1644969367
transform 1 0 54272 0 1 1938
box 0 0 1 1
use contact_32  contact_32_149
timestamp 1644969367
transform 1 0 54272 0 1 3422
box 0 0 1 1
use contact_32  contact_32_150
timestamp 1644969367
transform 1 0 53636 0 1 11054
box 0 0 1 1
use contact_32  contact_32_151
timestamp 1644969367
transform 1 0 53636 0 1 9782
box 0 0 1 1
use contact_32  contact_32_152
timestamp 1644969367
transform 1 0 52152 0 1 11054
box 0 0 1 1
use contact_32  contact_32_153
timestamp 1644969367
transform 1 0 52152 0 1 9782
box 0 0 1 1
use contact_32  contact_32_154
timestamp 1644969367
transform 1 0 50244 0 1 11054
box 0 0 1 1
use contact_32  contact_32_155
timestamp 1644969367
transform 1 0 50244 0 1 9782
box 0 0 1 1
use contact_32  contact_32_156
timestamp 1644969367
transform 1 0 48548 0 1 11054
box 0 0 1 1
use contact_32  contact_32_157
timestamp 1644969367
transform 1 0 48548 0 1 9782
box 0 0 1 1
use contact_32  contact_32_158
timestamp 1644969367
transform 1 0 48548 0 1 1938
box 0 0 1 1
use contact_32  contact_32_159
timestamp 1644969367
transform 1 0 48548 0 1 3422
box 0 0 1 1
use contact_32  contact_32_160
timestamp 1644969367
transform 1 0 47488 0 1 11054
box 0 0 1 1
use contact_32  contact_32_161
timestamp 1644969367
transform 1 0 47488 0 1 9782
box 0 0 1 1
use contact_32  contact_32_162
timestamp 1644969367
transform 1 0 45580 0 1 11054
box 0 0 1 1
use contact_32  contact_32_163
timestamp 1644969367
transform 1 0 45580 0 1 9782
box 0 0 1 1
use contact_32  contact_32_164
timestamp 1644969367
transform 1 0 45580 0 1 1938
box 0 0 1 1
use contact_32  contact_32_165
timestamp 1644969367
transform 1 0 45580 0 1 3422
box 0 0 1 1
use contact_32  contact_32_166
timestamp 1644969367
transform 1 0 44520 0 1 11054
box 0 0 1 1
use contact_32  contact_32_167
timestamp 1644969367
transform 1 0 44520 0 1 9782
box 0 0 1 1
use contact_32  contact_32_168
timestamp 1644969367
transform 1 0 43036 0 1 11054
box 0 0 1 1
use contact_32  contact_32_169
timestamp 1644969367
transform 1 0 43036 0 1 9994
box 0 0 1 1
use contact_32  contact_32_170
timestamp 1644969367
transform 1 0 39856 0 1 11054
box 0 0 1 1
use contact_32  contact_32_171
timestamp 1644969367
transform 1 0 39856 0 1 9782
box 0 0 1 1
use contact_32  contact_32_172
timestamp 1644969367
transform 1 0 38372 0 1 11054
box 0 0 1 1
use contact_32  contact_32_173
timestamp 1644969367
transform 1 0 38372 0 1 9782
box 0 0 1 1
use contact_32  contact_32_174
timestamp 1644969367
transform 1 0 36676 0 1 1938
box 0 0 1 1
use contact_32  contact_32_175
timestamp 1644969367
transform 1 0 36676 0 1 3422
box 0 0 1 1
use contact_32  contact_32_176
timestamp 1644969367
transform 1 0 36676 0 1 11054
box 0 0 1 1
use contact_32  contact_32_177
timestamp 1644969367
transform 1 0 36676 0 1 9782
box 0 0 1 1
use contact_32  contact_32_178
timestamp 1644969367
transform 1 0 35192 0 1 11054
box 0 0 1 1
use contact_32  contact_32_179
timestamp 1644969367
transform 1 0 35192 0 1 9570
box 0 0 1 1
use contact_32  contact_32_180
timestamp 1644969367
transform 1 0 33708 0 1 1938
box 0 0 1 1
use contact_32  contact_32_181
timestamp 1644969367
transform 1 0 33708 0 1 3422
box 0 0 1 1
use contact_32  contact_32_182
timestamp 1644969367
transform 1 0 33708 0 1 11054
box 0 0 1 1
use contact_32  contact_32_183
timestamp 1644969367
transform 1 0 33708 0 1 9782
box 0 0 1 1
use contact_32  contact_32_184
timestamp 1644969367
transform 1 0 32012 0 1 11054
box 0 0 1 1
use contact_32  contact_32_185
timestamp 1644969367
transform 1 0 32012 0 1 9994
box 0 0 1 1
use contact_32  contact_32_186
timestamp 1644969367
transform 1 0 30740 0 1 11054
box 0 0 1 1
use contact_32  contact_32_187
timestamp 1644969367
transform 1 0 30740 0 1 9994
box 0 0 1 1
use contact_32  contact_32_188
timestamp 1644969367
transform 1 0 29256 0 1 1938
box 0 0 1 1
use contact_32  contact_32_189
timestamp 1644969367
transform 1 0 29256 0 1 3422
box 0 0 1 1
use contact_32  contact_32_190
timestamp 1644969367
transform 1 0 28832 0 1 11054
box 0 0 1 1
use contact_32  contact_32_191
timestamp 1644969367
transform 1 0 28832 0 1 9994
box 0 0 1 1
use contact_32  contact_32_192
timestamp 1644969367
transform 1 0 27348 0 1 11054
box 0 0 1 1
use contact_32  contact_32_193
timestamp 1644969367
transform 1 0 27348 0 1 9782
box 0 0 1 1
use contact_32  contact_32_194
timestamp 1644969367
transform 1 0 27136 0 1 11266
box 0 0 1 1
use contact_32  contact_32_195
timestamp 1644969367
transform 1 0 27136 0 1 13598
box 0 0 1 1
use contact_32  contact_32_196
timestamp 1644969367
transform 1 0 26288 0 1 62782
box 0 0 1 1
use contact_32  contact_32_197
timestamp 1644969367
transform 1 0 26288 0 1 59814
box 0 0 1 1
use contact_32  contact_32_198
timestamp 1644969367
transform 1 0 26076 0 1 41370
box 0 0 1 1
use contact_32  contact_32_199
timestamp 1644969367
transform 1 0 26076 0 1 44338
box 0 0 1 1
use contact_32  contact_32_200
timestamp 1644969367
transform 1 0 26076 0 1 69142
box 0 0 1 1
use contact_32  contact_32_201
timestamp 1644969367
transform 1 0 26076 0 1 72110
box 0 0 1 1
use contact_32  contact_32_202
timestamp 1644969367
transform 1 0 26076 0 1 105818
box 0 0 1 1
use contact_32  contact_32_203
timestamp 1644969367
transform 1 0 26076 0 1 102850
box 0 0 1 1
use contact_32  contact_32_204
timestamp 1644969367
transform 1 0 26076 0 1 59814
box 0 0 1 1
use contact_32  contact_32_205
timestamp 1644969367
transform 1 0 26076 0 1 56846
box 0 0 1 1
use contact_32  contact_32_206
timestamp 1644969367
transform 1 0 26288 0 1 81226
box 0 0 1 1
use contact_32  contact_32_207
timestamp 1644969367
transform 1 0 26288 0 1 78258
box 0 0 1 1
use contact_32  contact_32_208
timestamp 1644969367
transform 1 0 26076 0 1 75290
box 0 0 1 1
use contact_32  contact_32_209
timestamp 1644969367
transform 1 0 26076 0 1 78258
box 0 0 1 1
use contact_32  contact_32_210
timestamp 1644969367
transform 1 0 26076 0 1 13810
box 0 0 1 1
use contact_32  contact_32_211
timestamp 1644969367
transform 1 0 26076 0 1 16778
box 0 0 1 1
use contact_32  contact_32_212
timestamp 1644969367
transform 1 0 26076 0 1 50486
box 0 0 1 1
use contact_32  contact_32_213
timestamp 1644969367
transform 1 0 26076 0 1 47518
box 0 0 1 1
use contact_32  contact_32_214
timestamp 1644969367
transform 1 0 26288 0 1 50698
box 0 0 1 1
use contact_32  contact_32_215
timestamp 1644969367
transform 1 0 26288 0 1 53666
box 0 0 1 1
use contact_32  contact_32_216
timestamp 1644969367
transform 1 0 26076 0 1 56634
box 0 0 1 1
use contact_32  contact_32_217
timestamp 1644969367
transform 1 0 26076 0 1 53666
box 0 0 1 1
use contact_32  contact_32_218
timestamp 1644969367
transform 1 0 26288 0 1 62994
box 0 0 1 1
use contact_32  contact_32_219
timestamp 1644969367
transform 1 0 26288 0 1 65962
box 0 0 1 1
use contact_32  contact_32_220
timestamp 1644969367
transform 1 0 26076 0 1 68930
box 0 0 1 1
use contact_32  contact_32_221
timestamp 1644969367
transform 1 0 26076 0 1 65962
box 0 0 1 1
use contact_32  contact_32_222
timestamp 1644969367
transform 1 0 26076 0 1 90554
box 0 0 1 1
use contact_32  contact_32_223
timestamp 1644969367
transform 1 0 26076 0 1 93522
box 0 0 1 1
use contact_32  contact_32_224
timestamp 1644969367
transform 1 0 26288 0 1 106030
box 0 0 1 1
use contact_32  contact_32_225
timestamp 1644969367
transform 1 0 26288 0 1 108998
box 0 0 1 1
use contact_32  contact_32_226
timestamp 1644969367
transform 1 0 26288 0 1 81438
box 0 0 1 1
use contact_32  contact_32_227
timestamp 1644969367
transform 1 0 26288 0 1 84406
box 0 0 1 1
use contact_32  contact_32_228
timestamp 1644969367
transform 1 0 26076 0 1 87374
box 0 0 1 1
use contact_32  contact_32_229
timestamp 1644969367
transform 1 0 26076 0 1 84406
box 0 0 1 1
use contact_32  contact_32_230
timestamp 1644969367
transform 1 0 26288 0 1 22926
box 0 0 1 1
use contact_32  contact_32_231
timestamp 1644969367
transform 1 0 26288 0 1 19958
box 0 0 1 1
use contact_32  contact_32_232
timestamp 1644969367
transform 1 0 26076 0 1 22926
box 0 0 1 1
use contact_32  contact_32_233
timestamp 1644969367
transform 1 0 26076 0 1 25894
box 0 0 1 1
use contact_32  contact_32_234
timestamp 1644969367
transform 1 0 24592 0 1 102850
box 0 0 1 1
use contact_32  contact_32_235
timestamp 1644969367
transform 1 0 24592 0 1 99882
box 0 0 1 1
use contact_32  contact_32_236
timestamp 1644969367
transform 1 0 24592 0 1 111330
box 0 0 1 1
use contact_32  contact_32_237
timestamp 1644969367
transform 1 0 24592 0 1 108998
box 0 0 1 1
use contact_32  contact_32_238
timestamp 1644969367
transform 1 0 24804 0 1 26106
box 0 0 1 1
use contact_32  contact_32_239
timestamp 1644969367
transform 1 0 24804 0 1 29074
box 0 0 1 1
use contact_32  contact_32_240
timestamp 1644969367
transform 1 0 24592 0 1 87586
box 0 0 1 1
use contact_32  contact_32_241
timestamp 1644969367
transform 1 0 24592 0 1 90554
box 0 0 1 1
use contact_32  contact_32_242
timestamp 1644969367
transform 1 0 24804 0 1 93734
box 0 0 1 1
use contact_32  contact_32_243
timestamp 1644969367
transform 1 0 24804 0 1 96702
box 0 0 1 1
use contact_32  contact_32_244
timestamp 1644969367
transform 1 0 24592 0 1 99670
box 0 0 1 1
use contact_32  contact_32_245
timestamp 1644969367
transform 1 0 24592 0 1 96702
box 0 0 1 1
use contact_32  contact_32_246
timestamp 1644969367
transform 1 0 24592 0 1 72110
box 0 0 1 1
use contact_32  contact_32_247
timestamp 1644969367
transform 1 0 24592 0 1 75078
box 0 0 1 1
use contact_32  contact_32_248
timestamp 1644969367
transform 1 0 24592 0 1 38402
box 0 0 1 1
use contact_32  contact_32_249
timestamp 1644969367
transform 1 0 24592 0 1 41370
box 0 0 1 1
use contact_32  contact_32_250
timestamp 1644969367
transform 1 0 24592 0 1 16778
box 0 0 1 1
use contact_32  contact_32_251
timestamp 1644969367
transform 1 0 24592 0 1 19746
box 0 0 1 1
use contact_32  contact_32_252
timestamp 1644969367
transform 1 0 24804 0 1 38190
box 0 0 1 1
use contact_32  contact_32_253
timestamp 1644969367
transform 1 0 24804 0 1 35222
box 0 0 1 1
use contact_32  contact_32_254
timestamp 1644969367
transform 1 0 24592 0 1 29074
box 0 0 1 1
use contact_32  contact_32_255
timestamp 1644969367
transform 1 0 24592 0 1 32042
box 0 0 1 1
use contact_32  contact_32_256
timestamp 1644969367
transform 1 0 24592 0 1 47518
box 0 0 1 1
use contact_32  contact_32_257
timestamp 1644969367
transform 1 0 24592 0 1 44550
box 0 0 1 1
use contact_32  contact_32_258
timestamp 1644969367
transform 1 0 21836 0 1 1938
box 0 0 1 1
use contact_32  contact_32_259
timestamp 1644969367
transform 1 0 21836 0 1 3422
box 0 0 1 1
use contact_32  contact_32_260
timestamp 1644969367
transform 1 0 20352 0 1 32042
box 0 0 1 1
use contact_32  contact_32_261
timestamp 1644969367
transform 1 0 20352 0 1 29074
box 0 0 1 1
use contact_32  contact_32_262
timestamp 1644969367
transform 1 0 20564 0 1 26106
box 0 0 1 1
use contact_32  contact_32_263
timestamp 1644969367
transform 1 0 20564 0 1 29074
box 0 0 1 1
use contact_32  contact_32_264
timestamp 1644969367
transform 1 0 20564 0 1 41370
box 0 0 1 1
use contact_32  contact_32_265
timestamp 1644969367
transform 1 0 20564 0 1 44338
box 0 0 1 1
use contact_32  contact_32_266
timestamp 1644969367
transform 1 0 20140 0 1 25894
box 0 0 1 1
use contact_32  contact_32_267
timestamp 1644969367
transform 1 0 20140 0 1 22926
box 0 0 1 1
use contact_32  contact_32_268
timestamp 1644969367
transform 1 0 19292 0 1 44550
box 0 0 1 1
use contact_32  contact_32_269
timestamp 1644969367
transform 1 0 19292 0 1 47518
box 0 0 1 1
use contact_32  contact_32_270
timestamp 1644969367
transform 1 0 19292 0 1 41370
box 0 0 1 1
use contact_32  contact_32_271
timestamp 1644969367
transform 1 0 19292 0 1 38402
box 0 0 1 1
use contact_32  contact_32_272
timestamp 1644969367
transform 1 0 19292 0 1 22926
box 0 0 1 1
use contact_32  contact_32_273
timestamp 1644969367
transform 1 0 19292 0 1 19958
box 0 0 1 1
use contact_32  contact_32_274
timestamp 1644969367
transform 1 0 17384 0 1 18262
box 0 0 1 1
use contact_32  contact_32_275
timestamp 1644969367
transform 1 0 17384 0 1 19746
box 0 0 1 1
use contact_32  contact_32_276
timestamp 1644969367
transform 1 0 17596 0 1 13174
box 0 0 1 1
use contact_32  contact_32_277
timestamp 1644969367
transform 1 0 17596 0 1 14658
box 0 0 1 1
use contact_32  contact_32_278
timestamp 1644969367
transform 1 0 17172 0 1 18050
box 0 0 1 1
use contact_32  contact_32_279
timestamp 1644969367
transform 1 0 17172 0 1 16566
box 0 0 1 1
use contact_32  contact_32_280
timestamp 1644969367
transform 1 0 16960 0 1 14870
box 0 0 1 1
use contact_32  contact_32_281
timestamp 1644969367
transform 1 0 16960 0 1 16354
box 0 0 1 1
use contact_32  contact_32_282
timestamp 1644969367
transform 1 0 1908 0 1 6814
box 0 0 1 1
use contact_34  contact_34_0
timestamp 1644969367
transform 1 0 848 0 1 112602
box 0 0 1 1
use contact_34  contact_34_1
timestamp 1644969367
transform 1 0 848 0 1 666
box 0 0 1 1
use contact_34  contact_34_2
timestamp 1644969367
transform 1 0 79288 0 1 666
box 0 0 1 1
use contact_34  contact_34_3
timestamp 1644969367
transform 1 0 424 0 1 112602
box 0 0 1 1
use contact_34  contact_34_4
timestamp 1644969367
transform 1 0 424 0 1 666
box 0 0 1 1
use contact_34  contact_34_5
timestamp 1644969367
transform 1 0 78864 0 1 878
box 0 0 1 1
use contact_34  contact_34_6
timestamp 1644969367
transform 1 0 78864 0 1 112390
box 0 0 1 1
use contact_34  contact_34_7
timestamp 1644969367
transform 1 0 78864 0 1 454
box 0 0 1 1
use contact_34  contact_34_8
timestamp 1644969367
transform 1 0 636 0 1 112602
box 0 0 1 1
use contact_34  contact_34_9
timestamp 1644969367
transform 1 0 636 0 1 666
box 0 0 1 1
use contact_34  contact_34_10
timestamp 1644969367
transform 1 0 79288 0 1 112814
box 0 0 1 1
use contact_34  contact_34_11
timestamp 1644969367
transform 1 0 78864 0 1 112814
box 0 0 1 1
use contact_34  contact_34_12
timestamp 1644969367
transform 1 0 79076 0 1 112814
box 0 0 1 1
use contact_34  contact_34_13
timestamp 1644969367
transform 1 0 848 0 1 112814
box 0 0 1 1
use contact_34  contact_34_14
timestamp 1644969367
transform 1 0 79288 0 1 878
box 0 0 1 1
use contact_34  contact_34_15
timestamp 1644969367
transform 1 0 848 0 1 878
box 0 0 1 1
use contact_34  contact_34_16
timestamp 1644969367
transform 1 0 848 0 1 112390
box 0 0 1 1
use contact_34  contact_34_17
timestamp 1644969367
transform 1 0 79288 0 1 112390
box 0 0 1 1
use contact_34  contact_34_18
timestamp 1644969367
transform 1 0 636 0 1 112814
box 0 0 1 1
use contact_34  contact_34_19
timestamp 1644969367
transform 1 0 79288 0 1 454
box 0 0 1 1
use contact_34  contact_34_20
timestamp 1644969367
transform 1 0 78864 0 1 112602
box 0 0 1 1
use contact_34  contact_34_21
timestamp 1644969367
transform 1 0 636 0 1 112390
box 0 0 1 1
use contact_34  contact_34_22
timestamp 1644969367
transform 1 0 79076 0 1 112390
box 0 0 1 1
use contact_34  contact_34_23
timestamp 1644969367
transform 1 0 79076 0 1 454
box 0 0 1 1
use contact_34  contact_34_24
timestamp 1644969367
transform 1 0 79076 0 1 878
box 0 0 1 1
use contact_34  contact_34_25
timestamp 1644969367
transform 1 0 424 0 1 112814
box 0 0 1 1
use contact_34  contact_34_26
timestamp 1644969367
transform 1 0 424 0 1 878
box 0 0 1 1
use contact_34  contact_34_27
timestamp 1644969367
transform 1 0 424 0 1 112390
box 0 0 1 1
use contact_34  contact_34_28
timestamp 1644969367
transform 1 0 848 0 1 454
box 0 0 1 1
use contact_34  contact_34_29
timestamp 1644969367
transform 1 0 78864 0 1 666
box 0 0 1 1
use contact_34  contact_34_30
timestamp 1644969367
transform 1 0 636 0 1 878
box 0 0 1 1
use contact_34  contact_34_31
timestamp 1644969367
transform 1 0 636 0 1 454
box 0 0 1 1
use contact_34  contact_34_32
timestamp 1644969367
transform 1 0 424 0 1 454
box 0 0 1 1
use contact_34  contact_34_33
timestamp 1644969367
transform 1 0 79288 0 1 112602
box 0 0 1 1
use contact_34  contact_34_34
timestamp 1644969367
transform 1 0 79076 0 1 112602
box 0 0 1 1
use contact_34  contact_34_35
timestamp 1644969367
transform 1 0 79076 0 1 666
box 0 0 1 1
use contact_34  contact_34_36
timestamp 1644969367
transform 1 0 78228 0 1 111330
box 0 0 1 1
use contact_34  contact_34_37
timestamp 1644969367
transform 1 0 77804 0 1 1514
box 0 0 1 1
use contact_34  contact_34_38
timestamp 1644969367
transform 1 0 78016 0 1 111542
box 0 0 1 1
use contact_34  contact_34_39
timestamp 1644969367
transform 1 0 1696 0 1 1938
box 0 0 1 1
use contact_34  contact_34_40
timestamp 1644969367
transform 1 0 1484 0 1 111542
box 0 0 1 1
use contact_34  contact_34_41
timestamp 1644969367
transform 1 0 1696 0 1 1514
box 0 0 1 1
use contact_34  contact_34_42
timestamp 1644969367
transform 1 0 1484 0 1 1938
box 0 0 1 1
use contact_34  contact_34_43
timestamp 1644969367
transform 1 0 78228 0 1 1726
box 0 0 1 1
use contact_34  contact_34_44
timestamp 1644969367
transform 1 0 77804 0 1 111754
box 0 0 1 1
use contact_34  contact_34_45
timestamp 1644969367
transform 1 0 1484 0 1 1514
box 0 0 1 1
use contact_34  contact_34_46
timestamp 1644969367
transform 1 0 78016 0 1 1938
box 0 0 1 1
use contact_34  contact_34_47
timestamp 1644969367
transform 1 0 1908 0 1 111542
box 0 0 1 1
use contact_34  contact_34_48
timestamp 1644969367
transform 1 0 1908 0 1 1938
box 0 0 1 1
use contact_34  contact_34_49
timestamp 1644969367
transform 1 0 77804 0 1 111330
box 0 0 1 1
use contact_34  contact_34_50
timestamp 1644969367
transform 1 0 1696 0 1 111754
box 0 0 1 1
use contact_34  contact_34_51
timestamp 1644969367
transform 1 0 77804 0 1 1726
box 0 0 1 1
use contact_34  contact_34_52
timestamp 1644969367
transform 1 0 1696 0 1 111330
box 0 0 1 1
use contact_34  contact_34_53
timestamp 1644969367
transform 1 0 1696 0 1 1726
box 0 0 1 1
use contact_34  contact_34_54
timestamp 1644969367
transform 1 0 78016 0 1 1514
box 0 0 1 1
use contact_34  contact_34_55
timestamp 1644969367
transform 1 0 1484 0 1 111754
box 0 0 1 1
use contact_34  contact_34_56
timestamp 1644969367
transform 1 0 78228 0 1 111542
box 0 0 1 1
use contact_34  contact_34_57
timestamp 1644969367
transform 1 0 1908 0 1 1514
box 0 0 1 1
use contact_34  contact_34_58
timestamp 1644969367
transform 1 0 1484 0 1 111330
box 0 0 1 1
use contact_34  contact_34_59
timestamp 1644969367
transform 1 0 78016 0 1 111754
box 0 0 1 1
use contact_34  contact_34_60
timestamp 1644969367
transform 1 0 78228 0 1 1514
box 0 0 1 1
use contact_34  contact_34_61
timestamp 1644969367
transform 1 0 1908 0 1 111754
box 0 0 1 1
use contact_34  contact_34_62
timestamp 1644969367
transform 1 0 78228 0 1 1938
box 0 0 1 1
use contact_34  contact_34_63
timestamp 1644969367
transform 1 0 77804 0 1 111542
box 0 0 1 1
use contact_34  contact_34_64
timestamp 1644969367
transform 1 0 78016 0 1 111330
box 0 0 1 1
use contact_34  contact_34_65
timestamp 1644969367
transform 1 0 78016 0 1 1726
box 0 0 1 1
use contact_34  contact_34_66
timestamp 1644969367
transform 1 0 1484 0 1 1726
box 0 0 1 1
use contact_34  contact_34_67
timestamp 1644969367
transform 1 0 1908 0 1 111330
box 0 0 1 1
use contact_34  contact_34_68
timestamp 1644969367
transform 1 0 1908 0 1 1726
box 0 0 1 1
use contact_34  contact_34_69
timestamp 1644969367
transform 1 0 77804 0 1 1938
box 0 0 1 1
use contact_34  contact_34_70
timestamp 1644969367
transform 1 0 1696 0 1 111542
box 0 0 1 1
use contact_34  contact_34_71
timestamp 1644969367
transform 1 0 78228 0 1 111754
box 0 0 1 1
use contact_32  contact_32_283
timestamp 1644969367
transform 1 0 16324 0 1 15930
box 0 0 1 1
use contact_32  contact_32_284
timestamp 1644969367
transform 1 0 17172 0 1 15294
box 0 0 1 1
use contact_32  contact_32_285
timestamp 1644969367
transform 1 0 16536 0 1 14234
box 0 0 1 1
use contact_32  contact_32_286
timestamp 1644969367
transform 1 0 16960 0 1 13598
box 0 0 1 1
use contact_32  contact_32_287
timestamp 1644969367
transform 1 0 16748 0 1 12538
box 0 0 1 1
use contact_32  contact_32_288
timestamp 1644969367
transform 1 0 50456 0 1 10630
box 0 0 1 1
use contact_32  contact_32_289
timestamp 1644969367
transform 1 0 50032 0 1 10630
box 0 0 1 1
use contact_32  contact_32_290
timestamp 1644969367
transform 1 0 48972 0 1 10630
box 0 0 1 1
use contact_32  contact_32_291
timestamp 1644969367
transform 1 0 48760 0 1 10630
box 0 0 1 1
use contact_32  contact_32_292
timestamp 1644969367
transform 1 0 47276 0 1 10630
box 0 0 1 1
use contact_32  contact_32_293
timestamp 1644969367
transform 1 0 47064 0 1 10630
box 0 0 1 1
use contact_32  contact_32_294
timestamp 1644969367
transform 1 0 46004 0 1 10630
box 0 0 1 1
use contact_32  contact_32_295
timestamp 1644969367
transform 1 0 45368 0 1 10630
box 0 0 1 1
use contact_32  contact_32_296
timestamp 1644969367
transform 1 0 44308 0 1 10630
box 0 0 1 1
use contact_32  contact_32_297
timestamp 1644969367
transform 1 0 44096 0 1 10630
box 0 0 1 1
use contact_32  contact_32_298
timestamp 1644969367
transform 1 0 42612 0 1 10630
box 0 0 1 1
use contact_32  contact_32_299
timestamp 1644969367
transform 1 0 42400 0 1 10630
box 0 0 1 1
use contact_32  contact_32_300
timestamp 1644969367
transform 1 0 41128 0 1 10630
box 0 0 1 1
use contact_32  contact_32_301
timestamp 1644969367
transform 1 0 40704 0 1 10630
box 0 0 1 1
use contact_32  contact_32_302
timestamp 1644969367
transform 1 0 39644 0 1 10630
box 0 0 1 1
use contact_32  contact_32_303
timestamp 1644969367
transform 1 0 39432 0 1 10630
box 0 0 1 1
use contact_32  contact_32_304
timestamp 1644969367
transform 1 0 38160 0 1 10630
box 0 0 1 1
use contact_32  contact_32_305
timestamp 1644969367
transform 1 0 37948 0 1 10630
box 0 0 1 1
use contact_32  contact_32_306
timestamp 1644969367
transform 1 0 36464 0 1 10630
box 0 0 1 1
use contact_32  contact_32_307
timestamp 1644969367
transform 1 0 36040 0 1 10630
box 0 0 1 1
use contact_32  contact_32_308
timestamp 1644969367
transform 1 0 34980 0 1 10630
box 0 0 1 1
use contact_32  contact_32_309
timestamp 1644969367
transform 1 0 34556 0 1 10630
box 0 0 1 1
use contact_32  contact_32_310
timestamp 1644969367
transform 1 0 33496 0 1 10630
box 0 0 1 1
use contact_32  contact_32_311
timestamp 1644969367
transform 1 0 33284 0 1 10630
box 0 0 1 1
use contact_32  contact_32_312
timestamp 1644969367
transform 1 0 31800 0 1 10630
box 0 0 1 1
use contact_32  contact_32_313
timestamp 1644969367
transform 1 0 31588 0 1 10630
box 0 0 1 1
use contact_32  contact_32_314
timestamp 1644969367
transform 1 0 30316 0 1 10630
box 0 0 1 1
use contact_32  contact_32_315
timestamp 1644969367
transform 1 0 29892 0 1 10630
box 0 0 1 1
use contact_32  contact_32_316
timestamp 1644969367
transform 1 0 28620 0 1 10630
box 0 0 1 1
use contact_32  contact_32_317
timestamp 1644969367
transform 1 0 28408 0 1 10630
box 0 0 1 1
use contact_32  contact_32_318
timestamp 1644969367
transform 1 0 27136 0 1 10630
box 0 0 1 1
use contact_32  contact_32_319
timestamp 1644969367
transform 1 0 26924 0 1 10630
box 0 0 1 1
use contact_32  contact_32_320
timestamp 1644969367
transform 1 0 19716 0 1 2998
box 0 0 1 1
use contact_32  contact_32_321
timestamp 1644969367
transform 1 0 67204 0 1 2998
box 0 0 1 1
use contact_32  contact_32_322
timestamp 1644969367
transform 1 0 65720 0 1 2998
box 0 0 1 1
use contact_32  contact_32_323
timestamp 1644969367
transform 1 0 64236 0 1 2998
box 0 0 1 1
use contact_32  contact_32_324
timestamp 1644969367
transform 1 0 62540 0 1 2998
box 0 0 1 1
use contact_32  contact_32_325
timestamp 1644969367
transform 1 0 61268 0 1 2998
box 0 0 1 1
use contact_32  contact_32_326
timestamp 1644969367
transform 1 0 59784 0 1 2998
box 0 0 1 1
use contact_32  contact_32_327
timestamp 1644969367
transform 1 0 58088 0 1 2998
box 0 0 1 1
use contact_32  contact_32_328
timestamp 1644969367
transform 1 0 56816 0 1 2998
box 0 0 1 1
use contact_32  contact_32_329
timestamp 1644969367
transform 1 0 55332 0 1 2998
box 0 0 1 1
use contact_32  contact_32_330
timestamp 1644969367
transform 1 0 53848 0 1 2998
box 0 0 1 1
use contact_32  contact_32_331
timestamp 1644969367
transform 1 0 52364 0 1 2998
box 0 0 1 1
use contact_32  contact_32_332
timestamp 1644969367
transform 1 0 50880 0 1 2998
box 0 0 1 1
use contact_32  contact_32_333
timestamp 1644969367
transform 1 0 49396 0 1 2998
box 0 0 1 1
use contact_32  contact_32_334
timestamp 1644969367
transform 1 0 47912 0 1 2998
box 0 0 1 1
use contact_32  contact_32_335
timestamp 1644969367
transform 1 0 46428 0 1 2998
box 0 0 1 1
use contact_32  contact_32_336
timestamp 1644969367
transform 1 0 44944 0 1 2998
box 0 0 1 1
use contact_32  contact_32_337
timestamp 1644969367
transform 1 0 43460 0 1 2998
box 0 0 1 1
use contact_32  contact_32_338
timestamp 1644969367
transform 1 0 41976 0 1 2998
box 0 0 1 1
use contact_32  contact_32_339
timestamp 1644969367
transform 1 0 40492 0 1 2998
box 0 0 1 1
use contact_32  contact_32_340
timestamp 1644969367
transform 1 0 39220 0 1 2998
box 0 0 1 1
use contact_32  contact_32_341
timestamp 1644969367
transform 1 0 37736 0 1 2998
box 0 0 1 1
use contact_32  contact_32_342
timestamp 1644969367
transform 1 0 36252 0 1 2998
box 0 0 1 1
use contact_32  contact_32_343
timestamp 1644969367
transform 1 0 34768 0 1 2998
box 0 0 1 1
use contact_32  contact_32_344
timestamp 1644969367
transform 1 0 33072 0 1 2998
box 0 0 1 1
use contact_32  contact_32_345
timestamp 1644969367
transform 1 0 31800 0 1 2998
box 0 0 1 1
use contact_32  contact_32_346
timestamp 1644969367
transform 1 0 30104 0 1 2998
box 0 0 1 1
use contact_32  contact_32_347
timestamp 1644969367
transform 1 0 28832 0 1 2998
box 0 0 1 1
use contact_32  contact_32_348
timestamp 1644969367
transform 1 0 27348 0 1 2998
box 0 0 1 1
use contact_32  contact_32_349
timestamp 1644969367
transform 1 0 25652 0 1 2998
box 0 0 1 1
use contact_32  contact_32_350
timestamp 1644969367
transform 1 0 24168 0 1 2998
box 0 0 1 1
use contact_32  contact_32_351
timestamp 1644969367
transform 1 0 22684 0 1 2998
box 0 0 1 1
use contact_32  contact_32_352
timestamp 1644969367
transform 1 0 21200 0 1 2998
box 0 0 1 1
use contact_18  contact_18_0
timestamp 1644969367
transform 1 0 16799 0 1 18765
box 0 0 1 1
use contact_18  contact_18_1
timestamp 1644969367
transform 1 0 16799 0 1 17581
box 0 0 1 1
use contact_18  contact_18_2
timestamp 1644969367
transform 1 0 16799 0 1 17089
box 0 0 1 1
use contact_18  contact_18_3
timestamp 1644969367
transform 1 0 16799 0 1 15905
box 0 0 1 1
use contact_18  contact_18_4
timestamp 1644969367
transform 1 0 16799 0 1 15413
box 0 0 1 1
use contact_18  contact_18_5
timestamp 1644969367
transform 1 0 16799 0 1 14229
box 0 0 1 1
use contact_18  contact_18_6
timestamp 1644969367
transform 1 0 16799 0 1 13737
box 0 0 1 1
use contact_18  contact_18_7
timestamp 1644969367
transform 1 0 16799 0 1 12553
box 0 0 1 1
use contact_18  contact_18_8
timestamp 1644969367
transform 1 0 19763 0 1 2975
box 0 0 1 1
use contact_18  contact_18_9
timestamp 1644969367
transform 1 0 50483 0 1 10647
box 0 0 1 1
use contact_18  contact_18_10
timestamp 1644969367
transform 1 0 50483 0 1 10647
box 0 0 1 1
use contact_18  contact_18_11
timestamp 1644969367
transform 1 0 50211 0 1 10647
box 0 0 1 1
use contact_18  contact_18_12
timestamp 1644969367
transform 1 0 50211 0 1 10647
box 0 0 1 1
use contact_18  contact_18_13
timestamp 1644969367
transform 1 0 48927 0 1 10647
box 0 0 1 1
use contact_18  contact_18_14
timestamp 1644969367
transform 1 0 48927 0 1 10647
box 0 0 1 1
use contact_18  contact_18_15
timestamp 1644969367
transform 1 0 48655 0 1 10647
box 0 0 1 1
use contact_18  contact_18_16
timestamp 1644969367
transform 1 0 48655 0 1 10647
box 0 0 1 1
use contact_18  contact_18_17
timestamp 1644969367
transform 1 0 47371 0 1 10647
box 0 0 1 1
use contact_18  contact_18_18
timestamp 1644969367
transform 1 0 47371 0 1 10647
box 0 0 1 1
use contact_18  contact_18_19
timestamp 1644969367
transform 1 0 47099 0 1 10647
box 0 0 1 1
use contact_18  contact_18_20
timestamp 1644969367
transform 1 0 47099 0 1 10647
box 0 0 1 1
use contact_18  contact_18_21
timestamp 1644969367
transform 1 0 45815 0 1 10647
box 0 0 1 1
use contact_18  contact_18_22
timestamp 1644969367
transform 1 0 45815 0 1 10647
box 0 0 1 1
use contact_18  contact_18_23
timestamp 1644969367
transform 1 0 45543 0 1 10647
box 0 0 1 1
use contact_18  contact_18_24
timestamp 1644969367
transform 1 0 45543 0 1 10647
box 0 0 1 1
use contact_18  contact_18_25
timestamp 1644969367
transform 1 0 44259 0 1 10647
box 0 0 1 1
use contact_18  contact_18_26
timestamp 1644969367
transform 1 0 44259 0 1 10647
box 0 0 1 1
use contact_18  contact_18_27
timestamp 1644969367
transform 1 0 43987 0 1 10647
box 0 0 1 1
use contact_18  contact_18_28
timestamp 1644969367
transform 1 0 43987 0 1 10647
box 0 0 1 1
use contact_18  contact_18_29
timestamp 1644969367
transform 1 0 42703 0 1 10647
box 0 0 1 1
use contact_18  contact_18_30
timestamp 1644969367
transform 1 0 42703 0 1 10647
box 0 0 1 1
use contact_18  contact_18_31
timestamp 1644969367
transform 1 0 42431 0 1 10647
box 0 0 1 1
use contact_18  contact_18_32
timestamp 1644969367
transform 1 0 42431 0 1 10647
box 0 0 1 1
use contact_18  contact_18_33
timestamp 1644969367
transform 1 0 41147 0 1 10647
box 0 0 1 1
use contact_18  contact_18_34
timestamp 1644969367
transform 1 0 41147 0 1 10647
box 0 0 1 1
use contact_18  contact_18_35
timestamp 1644969367
transform 1 0 40875 0 1 10647
box 0 0 1 1
use contact_18  contact_18_36
timestamp 1644969367
transform 1 0 40875 0 1 10647
box 0 0 1 1
use contact_18  contact_18_37
timestamp 1644969367
transform 1 0 39591 0 1 10647
box 0 0 1 1
use contact_18  contact_18_38
timestamp 1644969367
transform 1 0 39591 0 1 10647
box 0 0 1 1
use contact_18  contact_18_39
timestamp 1644969367
transform 1 0 39319 0 1 10647
box 0 0 1 1
use contact_18  contact_18_40
timestamp 1644969367
transform 1 0 39319 0 1 10647
box 0 0 1 1
use contact_18  contact_18_41
timestamp 1644969367
transform 1 0 38035 0 1 10647
box 0 0 1 1
use contact_18  contact_18_42
timestamp 1644969367
transform 1 0 38035 0 1 10647
box 0 0 1 1
use contact_18  contact_18_43
timestamp 1644969367
transform 1 0 37763 0 1 10647
box 0 0 1 1
use contact_18  contact_18_44
timestamp 1644969367
transform 1 0 37763 0 1 10647
box 0 0 1 1
use contact_18  contact_18_45
timestamp 1644969367
transform 1 0 36479 0 1 10647
box 0 0 1 1
use contact_18  contact_18_46
timestamp 1644969367
transform 1 0 36479 0 1 10647
box 0 0 1 1
use contact_18  contact_18_47
timestamp 1644969367
transform 1 0 36207 0 1 10647
box 0 0 1 1
use contact_18  contact_18_48
timestamp 1644969367
transform 1 0 36207 0 1 10647
box 0 0 1 1
use contact_18  contact_18_49
timestamp 1644969367
transform 1 0 34923 0 1 10647
box 0 0 1 1
use contact_18  contact_18_50
timestamp 1644969367
transform 1 0 34923 0 1 10647
box 0 0 1 1
use contact_18  contact_18_51
timestamp 1644969367
transform 1 0 34651 0 1 10647
box 0 0 1 1
use contact_18  contact_18_52
timestamp 1644969367
transform 1 0 34651 0 1 10647
box 0 0 1 1
use contact_18  contact_18_53
timestamp 1644969367
transform 1 0 33367 0 1 10647
box 0 0 1 1
use contact_18  contact_18_54
timestamp 1644969367
transform 1 0 33367 0 1 10647
box 0 0 1 1
use contact_18  contact_18_55
timestamp 1644969367
transform 1 0 33095 0 1 10647
box 0 0 1 1
use contact_18  contact_18_56
timestamp 1644969367
transform 1 0 33095 0 1 10647
box 0 0 1 1
use contact_18  contact_18_57
timestamp 1644969367
transform 1 0 31811 0 1 10647
box 0 0 1 1
use contact_18  contact_18_58
timestamp 1644969367
transform 1 0 31811 0 1 10647
box 0 0 1 1
use contact_18  contact_18_59
timestamp 1644969367
transform 1 0 31539 0 1 10647
box 0 0 1 1
use contact_18  contact_18_60
timestamp 1644969367
transform 1 0 31539 0 1 10647
box 0 0 1 1
use contact_18  contact_18_61
timestamp 1644969367
transform 1 0 30255 0 1 10647
box 0 0 1 1
use contact_18  contact_18_62
timestamp 1644969367
transform 1 0 30255 0 1 10647
box 0 0 1 1
use contact_18  contact_18_63
timestamp 1644969367
transform 1 0 29983 0 1 10647
box 0 0 1 1
use contact_18  contact_18_64
timestamp 1644969367
transform 1 0 29983 0 1 10647
box 0 0 1 1
use contact_18  contact_18_65
timestamp 1644969367
transform 1 0 28699 0 1 10647
box 0 0 1 1
use contact_18  contact_18_66
timestamp 1644969367
transform 1 0 28699 0 1 10647
box 0 0 1 1
use contact_18  contact_18_67
timestamp 1644969367
transform 1 0 28427 0 1 10647
box 0 0 1 1
use contact_18  contact_18_68
timestamp 1644969367
transform 1 0 28427 0 1 10647
box 0 0 1 1
use contact_18  contact_18_69
timestamp 1644969367
transform 1 0 27143 0 1 10647
box 0 0 1 1
use contact_18  contact_18_70
timestamp 1644969367
transform 1 0 27143 0 1 10647
box 0 0 1 1
use contact_18  contact_18_71
timestamp 1644969367
transform 1 0 26871 0 1 10647
box 0 0 1 1
use contact_18  contact_18_72
timestamp 1644969367
transform 1 0 26871 0 1 10647
box 0 0 1 1
use contact_18  contact_18_73
timestamp 1644969367
transform 1 0 67187 0 1 2975
box 0 0 1 1
use contact_18  contact_18_74
timestamp 1644969367
transform 1 0 65705 0 1 2975
box 0 0 1 1
use contact_18  contact_18_75
timestamp 1644969367
transform 1 0 64223 0 1 2975
box 0 0 1 1
use contact_18  contact_18_76
timestamp 1644969367
transform 1 0 62741 0 1 2975
box 0 0 1 1
use contact_18  contact_18_77
timestamp 1644969367
transform 1 0 61259 0 1 2975
box 0 0 1 1
use contact_18  contact_18_78
timestamp 1644969367
transform 1 0 59777 0 1 2975
box 0 0 1 1
use contact_18  contact_18_79
timestamp 1644969367
transform 1 0 58295 0 1 2975
box 0 0 1 1
use contact_18  contact_18_80
timestamp 1644969367
transform 1 0 56813 0 1 2975
box 0 0 1 1
use contact_18  contact_18_81
timestamp 1644969367
transform 1 0 55331 0 1 2975
box 0 0 1 1
use contact_18  contact_18_82
timestamp 1644969367
transform 1 0 53849 0 1 2975
box 0 0 1 1
use contact_18  contact_18_83
timestamp 1644969367
transform 1 0 52367 0 1 2975
box 0 0 1 1
use contact_18  contact_18_84
timestamp 1644969367
transform 1 0 50885 0 1 2975
box 0 0 1 1
use contact_18  contact_18_85
timestamp 1644969367
transform 1 0 49403 0 1 2975
box 0 0 1 1
use contact_18  contact_18_86
timestamp 1644969367
transform 1 0 47921 0 1 2975
box 0 0 1 1
use contact_18  contact_18_87
timestamp 1644969367
transform 1 0 46439 0 1 2975
box 0 0 1 1
use contact_18  contact_18_88
timestamp 1644969367
transform 1 0 44957 0 1 2975
box 0 0 1 1
use contact_18  contact_18_89
timestamp 1644969367
transform 1 0 43475 0 1 2975
box 0 0 1 1
use contact_18  contact_18_90
timestamp 1644969367
transform 1 0 41993 0 1 2975
box 0 0 1 1
use contact_18  contact_18_91
timestamp 1644969367
transform 1 0 40511 0 1 2975
box 0 0 1 1
use contact_18  contact_18_92
timestamp 1644969367
transform 1 0 39029 0 1 2975
box 0 0 1 1
use contact_18  contact_18_93
timestamp 1644969367
transform 1 0 37547 0 1 2975
box 0 0 1 1
use contact_18  contact_18_94
timestamp 1644969367
transform 1 0 36065 0 1 2975
box 0 0 1 1
use contact_18  contact_18_95
timestamp 1644969367
transform 1 0 34583 0 1 2975
box 0 0 1 1
use contact_18  contact_18_96
timestamp 1644969367
transform 1 0 33101 0 1 2975
box 0 0 1 1
use contact_18  contact_18_97
timestamp 1644969367
transform 1 0 31619 0 1 2975
box 0 0 1 1
use contact_18  contact_18_98
timestamp 1644969367
transform 1 0 30137 0 1 2975
box 0 0 1 1
use contact_18  contact_18_99
timestamp 1644969367
transform 1 0 28655 0 1 2975
box 0 0 1 1
use contact_18  contact_18_100
timestamp 1644969367
transform 1 0 27173 0 1 2975
box 0 0 1 1
use contact_18  contact_18_101
timestamp 1644969367
transform 1 0 25691 0 1 2975
box 0 0 1 1
use contact_18  contact_18_102
timestamp 1644969367
transform 1 0 24209 0 1 2975
box 0 0 1 1
use contact_18  contact_18_103
timestamp 1644969367
transform 1 0 22727 0 1 2975
box 0 0 1 1
use contact_18  contact_18_104
timestamp 1644969367
transform 1 0 21245 0 1 2975
box 0 0 1 1
use contact_18  contact_18_105
timestamp 1644969367
transform 1 0 6275 0 1 7364
box 0 0 1 1
use contact_18  contact_18_106
timestamp 1644969367
transform 1 0 2753 0 1 7579
box 0 0 1 1
use contact_18  contact_18_107
timestamp 1644969367
transform 1 0 2753 0 1 6395
box 0 0 1 1
use contact_18  contact_18_108
timestamp 1644969367
transform 1 0 18862 0 1 18769
box 0 0 1 1
use contact_18  contact_18_109
timestamp 1644969367
transform 1 0 17879 0 1 18769
box 0 0 1 1
use contact_18  contact_18_110
timestamp 1644969367
transform 1 0 18778 0 1 17577
box 0 0 1 1
use contact_18  contact_18_111
timestamp 1644969367
transform 1 0 17879 0 1 17577
box 0 0 1 1
use contact_18  contact_18_112
timestamp 1644969367
transform 1 0 18694 0 1 17093
box 0 0 1 1
use contact_18  contact_18_113
timestamp 1644969367
transform 1 0 17879 0 1 17093
box 0 0 1 1
use contact_18  contact_18_114
timestamp 1644969367
transform 1 0 18610 0 1 15901
box 0 0 1 1
use contact_18  contact_18_115
timestamp 1644969367
transform 1 0 17879 0 1 15901
box 0 0 1 1
use contact_18  contact_18_116
timestamp 1644969367
transform 1 0 18526 0 1 15417
box 0 0 1 1
use contact_18  contact_18_117
timestamp 1644969367
transform 1 0 17879 0 1 15417
box 0 0 1 1
use contact_18  contact_18_118
timestamp 1644969367
transform 1 0 18442 0 1 14225
box 0 0 1 1
use contact_18  contact_18_119
timestamp 1644969367
transform 1 0 17879 0 1 14225
box 0 0 1 1
use contact_18  contact_18_120
timestamp 1644969367
transform 1 0 18358 0 1 13741
box 0 0 1 1
use contact_18  contact_18_121
timestamp 1644969367
transform 1 0 17879 0 1 13741
box 0 0 1 1
use contact_18  contact_18_122
timestamp 1644969367
transform 1 0 18274 0 1 12549
box 0 0 1 1
use contact_18  contact_18_123
timestamp 1644969367
transform 1 0 17879 0 1 12549
box 0 0 1 1
use contact_18  contact_18_124
timestamp 1644969367
transform 1 0 25058 0 1 11645
box 0 0 1 1
use contact_18  contact_18_125
timestamp 1644969367
transform 1 0 18074 0 1 11645
box 0 0 1 1
use contact_18  contact_18_126
timestamp 1644969367
transform 1 0 76654 0 1 10709
box 0 0 1 1
use contact_18  contact_18_127
timestamp 1644969367
transform 1 0 18074 0 1 10709
box 0 0 1 1
use contact_18  contact_18_128
timestamp 1644969367
transform 1 0 26180 0 1 9970
box 0 0 1 1
use contact_18  contact_18_129
timestamp 1644969367
transform 1 0 18074 0 1 9970
box 0 0 1 1
use contact_30  contact_30_0
timestamp 1644969367
transform 1 0 16508 0 1 3037
box 0 0 1 1
use contact_30  contact_30_1
timestamp 1644969367
transform 1 0 16508 0 1 3037
box 0 0 1 1
use contact_30  contact_30_2
timestamp 1644969367
transform 1 0 16508 0 1 12615
box 0 0 1 1
use data_dff  data_dff_0
timestamp 1644969367
transform 1 0 21104 0 1 2766
box -39 -42 47424 916
use col_addr_dff  col_addr_dff_0
timestamp 1644969367
transform 1 0 19622 0 1 2766
box -39 -42 1482 916
use row_addr_dff  row_addr_dff_0
timestamp 1644969367
transform 1 0 16658 0 1 12344
box -39 -42 1482 8422
use control_logic_multiport  control_logic_multiport_0
timestamp 1644969367
transform 1 0 2612 0 1 6186
box -66 -42 15528 5906
use bank  bank_0
timestamp 1644969367
transform 1 0 18308 0 1 5800
box 0 0 58866 105020
<< labels >>
rlabel metal3 s 2752 6394 2884 6468 4 web
rlabel metal3 s 2752 7578 2884 7652 4 csb
rlabel metal3 s 0 7208 364 7360 4 clk
rlabel metal4 s 21200 0 21352 364 4 din0[0]
rlabel metal4 s 22684 0 22836 364 4 din0[1]
rlabel metal4 s 24168 0 24320 364 4 din0[2]
rlabel metal4 s 25652 0 25804 364 4 din0[3]
rlabel metal4 s 27348 0 27500 364 4 din0[4]
rlabel metal4 s 28832 0 28984 364 4 din0[5]
rlabel metal4 s 30104 0 30256 364 4 din0[6]
rlabel metal4 s 31800 0 31952 364 4 din0[7]
rlabel metal4 s 33072 0 33224 364 4 din0[8]
rlabel metal4 s 34768 0 34920 364 4 din0[9]
rlabel metal4 s 36252 0 36404 364 4 din0[10]
rlabel metal4 s 37736 0 37888 364 4 din0[11]
rlabel metal4 s 39220 0 39372 364 4 din0[12]
rlabel metal4 s 40492 0 40644 364 4 din0[13]
rlabel metal4 s 41976 0 42128 364 4 din0[14]
rlabel metal4 s 43460 0 43612 364 4 din0[15]
rlabel metal4 s 44944 0 45096 364 4 din0[16]
rlabel metal4 s 46428 0 46580 364 4 din0[17]
rlabel metal4 s 47912 0 48064 364 4 din0[18]
rlabel metal4 s 49396 0 49548 364 4 din0[19]
rlabel metal4 s 50880 0 51032 364 4 din0[20]
rlabel metal4 s 52364 0 52516 364 4 din0[21]
rlabel metal4 s 53848 0 54000 364 4 din0[22]
rlabel metal4 s 55332 0 55484 364 4 din0[23]
rlabel metal4 s 56816 0 56968 364 4 din0[24]
rlabel metal4 s 58088 0 58240 364 4 din0[25]
rlabel metal4 s 59784 0 59936 364 4 din0[26]
rlabel metal4 s 61268 0 61420 364 4 din0[27]
rlabel metal4 s 62540 0 62692 364 4 din0[28]
rlabel metal4 s 64236 0 64388 364 4 din0[29]
rlabel metal4 s 65720 0 65872 364 4 din0[30]
rlabel metal4 s 67204 0 67356 364 4 din0[31]
rlabel metal4 s 26924 0 27076 364 4 dout0[0]
rlabel metal3 s 26870 10646 27002 10720 4 dout1[0]
rlabel metal4 s 27136 0 27288 364 4 dout0[1]
rlabel metal3 s 27142 10646 27274 10720 4 dout1[1]
rlabel metal4 s 28408 0 28560 364 4 dout0[2]
rlabel metal3 s 28426 10646 28558 10720 4 dout1[2]
rlabel metal4 s 28620 0 28772 364 4 dout0[3]
rlabel metal3 s 28698 10646 28830 10720 4 dout1[3]
rlabel metal4 s 29892 0 30044 364 4 dout0[4]
rlabel metal3 s 29982 10646 30114 10720 4 dout1[4]
rlabel metal4 s 30316 0 30468 364 4 dout0[5]
rlabel metal3 s 30254 10646 30386 10720 4 dout1[5]
rlabel metal4 s 31588 0 31740 364 4 dout0[6]
rlabel metal3 s 31538 10646 31670 10720 4 dout1[6]
rlabel metal4 s 32012 0 32164 364 4 dout0[7]
rlabel metal3 s 31810 10646 31942 10720 4 dout1[7]
rlabel metal4 s 33284 0 33436 364 4 dout0[8]
rlabel metal3 s 33094 10646 33226 10720 4 dout1[8]
rlabel metal4 s 33496 0 33648 364 4 dout0[9]
rlabel metal3 s 33366 10646 33498 10720 4 dout1[9]
rlabel metal4 s 34556 0 34708 364 4 dout0[10]
rlabel metal3 s 34650 10646 34782 10720 4 dout1[10]
rlabel metal4 s 34980 0 35132 364 4 dout0[11]
rlabel metal3 s 34922 10646 35054 10720 4 dout1[11]
rlabel metal4 s 36040 0 36192 364 4 dout0[12]
rlabel metal3 s 36206 10646 36338 10720 4 dout1[12]
rlabel metal4 s 36464 0 36616 364 4 dout0[13]
rlabel metal3 s 36478 10646 36610 10720 4 dout1[13]
rlabel metal4 s 37948 0 38100 364 4 dout0[14]
rlabel metal3 s 37762 10646 37894 10720 4 dout1[14]
rlabel metal4 s 38160 0 38312 364 4 dout0[15]
rlabel metal3 s 38034 10646 38166 10720 4 dout1[15]
rlabel metal4 s 39432 0 39584 364 4 dout0[16]
rlabel metal3 s 39318 10646 39450 10720 4 dout1[16]
rlabel metal4 s 39644 0 39796 364 4 dout0[17]
rlabel metal3 s 39590 10646 39722 10720 4 dout1[17]
rlabel metal4 s 40704 0 40856 364 4 dout0[18]
rlabel metal3 s 40874 10646 41006 10720 4 dout1[18]
rlabel metal4 s 41128 0 41280 364 4 dout0[19]
rlabel metal3 s 41146 10646 41278 10720 4 dout1[19]
rlabel metal4 s 42400 0 42552 364 4 dout0[20]
rlabel metal3 s 42430 10646 42562 10720 4 dout1[20]
rlabel metal4 s 42612 0 42764 364 4 dout0[21]
rlabel metal3 s 42702 10646 42834 10720 4 dout1[21]
rlabel metal4 s 44096 0 44248 364 4 dout0[22]
rlabel metal3 s 43986 10646 44118 10720 4 dout1[22]
rlabel metal4 s 44308 0 44460 364 4 dout0[23]
rlabel metal3 s 44258 10646 44390 10720 4 dout1[23]
rlabel metal4 s 45368 0 45520 364 4 dout0[24]
rlabel metal3 s 45542 10646 45674 10720 4 dout1[24]
rlabel metal4 s 46004 0 46156 364 4 dout0[25]
rlabel metal3 s 45814 10646 45946 10720 4 dout1[25]
rlabel metal4 s 47064 0 47216 364 4 dout0[26]
rlabel metal3 s 47098 10646 47230 10720 4 dout1[26]
rlabel metal4 s 47276 0 47428 364 4 dout0[27]
rlabel metal3 s 47370 10646 47502 10720 4 dout1[27]
rlabel metal4 s 48760 0 48912 364 4 dout0[28]
rlabel metal3 s 48654 10646 48786 10720 4 dout1[28]
rlabel metal4 s 48972 0 49124 364 4 dout0[29]
rlabel metal3 s 48926 10646 49058 10720 4 dout1[29]
rlabel metal4 s 50032 0 50184 364 4 dout0[30]
rlabel metal3 s 50210 10646 50342 10720 4 dout1[30]
rlabel metal4 s 50456 0 50608 364 4 dout0[31]
rlabel metal3 s 50482 10646 50614 10720 4 dout1[31]
rlabel metal4 s 19716 0 19868 364 4 addr0
rlabel metal4 s 16748 0 16900 364 4 addr1[1]
rlabel metal4 s 16960 0 17112 364 4 addr1[2]
rlabel metal4 s 16536 0 16688 364 4 addr1[3]
rlabel metal4 s 17172 0 17324 364 4 addr1[4]
rlabel metal4 s 16324 0 16476 364 4 addr1[5]
rlabel metal3 s 0 16960 364 17112 4 addr1[6]
rlabel metal3 s 0 17596 364 17748 4 addr1[7]
rlabel metal3 s 0 18656 364 18808 4 addr1[8]
rlabel metal3 s 1484 1484 78380 2060 4 vdd
rlabel metal4 s 77804 1484 78380 111876 4 vdd
rlabel metal3 s 1484 111300 78380 111876 4 vdd
rlabel metal4 s 1484 1484 2060 111876 4 vdd
rlabel metal3 s 424 424 79440 1000 4 gnd
rlabel metal4 s 424 424 1000 112936 4 gnd
rlabel metal3 s 424 112360 79440 112936 4 gnd
rlabel metal4 s 78864 424 79440 112936 4 gnd
<< properties >>
string FIXED_BBOX 0 0 79440 112936
string GDS_FILE sram_0rw2r1w_32_128_sky130A.gds
string GDS_END 298632
string GDS_START 128
<< end >>
