magic
tech sky130A
timestamp 1644922390
<< nwell >>
rect 0 523 602 808
<< nmos >>
rect 47 154 62 209
rect 95 154 110 209
rect 143 154 158 209
rect 191 154 206 209
rect 293 154 308 209
rect 341 154 356 209
rect 392 154 407 196
rect 492 154 507 196
rect 540 154 555 196
<< pmos >>
rect 47 541 62 583
rect 95 541 110 583
rect 143 541 158 583
rect 191 541 206 583
rect 293 541 308 583
rect 341 541 356 583
rect 392 541 407 676
rect 492 541 507 676
rect 540 541 555 676
<< ndiff >>
rect 18 191 47 209
rect 18 174 22 191
rect 39 174 47 191
rect 18 154 47 174
rect 62 154 95 209
rect 110 191 143 209
rect 110 174 118 191
rect 135 174 143 191
rect 110 154 143 174
rect 158 154 191 209
rect 206 191 235 209
rect 206 174 214 191
rect 231 174 235 191
rect 206 154 235 174
rect 264 191 293 209
rect 264 174 268 191
rect 285 174 293 191
rect 264 154 293 174
rect 308 154 341 209
rect 356 196 384 209
rect 356 191 392 196
rect 356 174 364 191
rect 381 174 392 191
rect 356 154 392 174
rect 407 184 436 196
rect 407 167 415 184
rect 432 167 436 184
rect 407 154 436 167
rect 463 184 492 196
rect 463 167 467 184
rect 484 167 492 184
rect 463 154 492 167
rect 507 184 540 196
rect 507 167 515 184
rect 532 167 540 184
rect 507 154 540 167
rect 555 184 584 196
rect 555 167 563 184
rect 580 167 584 184
rect 555 154 584 167
<< pdiff >>
rect 364 660 392 676
rect 364 643 368 660
rect 385 643 392 660
rect 364 618 392 643
rect 364 601 368 618
rect 385 601 392 618
rect 364 583 392 601
rect 18 570 47 583
rect 18 553 22 570
rect 39 553 47 570
rect 18 541 47 553
rect 62 570 95 583
rect 62 553 70 570
rect 87 553 95 570
rect 62 541 95 553
rect 110 570 143 583
rect 110 553 118 570
rect 135 553 143 570
rect 110 541 143 553
rect 158 570 191 583
rect 158 553 166 570
rect 183 553 191 570
rect 158 541 191 553
rect 206 570 235 583
rect 206 553 214 570
rect 231 553 235 570
rect 206 541 235 553
rect 264 570 293 583
rect 264 553 268 570
rect 285 553 293 570
rect 264 541 293 553
rect 308 569 341 583
rect 308 552 316 569
rect 333 552 341 569
rect 308 541 341 552
rect 356 569 392 583
rect 356 552 366 569
rect 383 552 392 569
rect 356 541 392 552
rect 407 660 436 676
rect 407 643 415 660
rect 432 643 436 660
rect 407 618 436 643
rect 407 601 415 618
rect 432 601 436 618
rect 407 575 436 601
rect 407 558 415 575
rect 432 558 436 575
rect 407 541 436 558
rect 463 660 492 676
rect 463 643 467 660
rect 484 643 492 660
rect 463 618 492 643
rect 463 601 467 618
rect 484 601 492 618
rect 463 575 492 601
rect 463 558 467 575
rect 484 558 492 575
rect 463 541 492 558
rect 507 660 540 676
rect 507 643 515 660
rect 532 643 540 660
rect 507 618 540 643
rect 507 601 515 618
rect 532 601 540 618
rect 507 575 540 601
rect 507 558 515 575
rect 532 558 540 575
rect 507 541 540 558
rect 555 660 584 676
rect 555 643 563 660
rect 580 643 584 660
rect 555 618 584 643
rect 555 601 563 618
rect 580 601 584 618
rect 555 575 584 601
rect 555 558 563 575
rect 580 558 584 575
rect 555 541 584 558
<< ndiffc >>
rect 22 174 39 191
rect 118 174 135 191
rect 214 174 231 191
rect 268 174 285 191
rect 364 174 381 191
rect 415 167 432 184
rect 467 167 484 184
rect 515 167 532 184
rect 563 167 580 184
<< pdiffc >>
rect 368 643 385 660
rect 368 601 385 618
rect 22 553 39 570
rect 70 553 87 570
rect 118 553 135 570
rect 166 553 183 570
rect 214 553 231 570
rect 268 553 285 570
rect 316 552 333 569
rect 366 552 383 569
rect 415 643 432 660
rect 415 601 432 618
rect 415 558 432 575
rect 467 643 484 660
rect 467 601 484 618
rect 467 558 484 575
rect 515 643 532 660
rect 515 601 532 618
rect 515 558 532 575
rect 563 643 580 660
rect 563 601 580 618
rect 563 558 580 575
<< psubdiff >>
rect 92 9 128 21
rect 92 -9 101 9
rect 119 -9 128 9
rect 92 -21 128 -9
rect 219 9 255 21
rect 219 -9 228 9
rect 246 -9 255 9
rect 219 -21 255 -9
rect 347 9 383 21
rect 347 -9 356 9
rect 374 -9 383 9
rect 347 -21 383 -9
rect 474 9 510 21
rect 474 -9 483 9
rect 500 -9 510 9
rect 474 -21 510 -9
<< nsubdiff >>
rect 92 778 128 790
rect 92 760 101 778
rect 119 760 128 778
rect 92 748 128 760
rect 219 778 255 790
rect 219 760 228 778
rect 246 760 255 778
rect 219 748 255 760
rect 347 778 383 790
rect 347 760 356 778
rect 374 760 383 778
rect 347 748 383 760
rect 474 778 510 790
rect 474 760 483 778
rect 501 760 510 778
rect 474 748 510 760
<< psubdiffcont >>
rect 101 -9 119 9
rect 228 -9 246 9
rect 356 -9 374 9
rect 483 -9 500 9
<< nsubdiffcont >>
rect 101 760 119 778
rect 228 760 246 778
rect 356 760 374 778
rect 483 760 501 778
<< poly >>
rect 392 676 407 689
rect 492 676 507 689
rect 540 676 555 689
rect 47 583 62 596
rect 95 583 110 596
rect 143 583 158 596
rect 191 583 206 596
rect 293 583 308 596
rect 341 583 356 596
rect 47 508 62 541
rect 35 500 62 508
rect 35 483 40 500
rect 57 483 62 500
rect 35 475 62 483
rect 47 209 62 475
rect 95 464 110 541
rect 83 456 110 464
rect 83 439 88 456
rect 105 439 110 456
rect 83 431 110 439
rect 95 209 110 431
rect 143 420 158 541
rect 131 412 158 420
rect 131 395 136 412
rect 153 395 158 412
rect 131 387 158 395
rect 143 209 158 387
rect 191 376 206 541
rect 179 368 206 376
rect 179 351 184 368
rect 201 351 206 368
rect 179 343 206 351
rect 191 209 206 343
rect 293 319 308 541
rect 281 311 308 319
rect 281 294 286 311
rect 303 294 308 311
rect 281 286 308 294
rect 293 209 308 286
rect 341 276 356 541
rect 392 350 407 541
rect 380 342 407 350
rect 380 325 385 342
rect 402 325 407 342
rect 380 317 407 325
rect 329 268 356 276
rect 329 251 334 268
rect 351 251 356 268
rect 329 243 356 251
rect 341 209 356 243
rect 392 196 407 317
rect 492 393 507 541
rect 540 457 555 541
rect 528 449 555 457
rect 528 432 533 449
rect 550 432 555 449
rect 528 424 555 432
rect 492 385 519 393
rect 492 368 497 385
rect 514 368 519 385
rect 492 360 519 368
rect 492 196 507 360
rect 540 196 555 424
rect 47 141 62 154
rect 95 141 110 154
rect 143 141 158 154
rect 191 141 206 154
rect 293 141 308 154
rect 341 141 356 154
rect 392 141 407 154
rect 492 141 507 154
rect 540 141 555 154
<< polycont >>
rect 40 483 57 500
rect 88 439 105 456
rect 136 395 153 412
rect 184 351 201 368
rect 286 294 303 311
rect 385 325 402 342
rect 334 251 351 268
rect 533 432 550 449
rect 497 368 514 385
<< locali >>
rect 22 778 580 786
rect 22 760 101 778
rect 119 760 228 778
rect 246 760 356 778
rect 374 760 483 778
rect 501 760 580 778
rect 22 752 580 760
rect 22 583 39 752
rect 118 583 135 752
rect 214 583 231 752
rect 268 583 285 752
rect 368 676 385 752
rect 515 676 532 752
rect 364 660 387 676
rect 364 643 368 660
rect 385 643 387 660
rect 364 618 387 643
rect 364 601 368 618
rect 385 601 387 618
rect 364 583 387 601
rect 18 570 42 583
rect 18 553 22 570
rect 39 553 42 570
rect 18 541 42 553
rect 67 570 90 583
rect 67 553 70 570
rect 87 553 90 570
rect 67 541 90 553
rect 115 570 138 583
rect 115 553 118 570
rect 135 553 138 570
rect 115 541 138 553
rect 163 570 186 583
rect 163 553 166 570
rect 183 553 186 570
rect 163 541 186 553
rect 211 570 235 583
rect 211 553 214 570
rect 231 553 235 570
rect 211 541 235 553
rect 264 570 288 583
rect 264 553 268 570
rect 285 553 288 570
rect 264 541 288 553
rect 313 569 336 583
rect 313 552 316 569
rect 333 552 336 569
rect 313 541 336 552
rect 361 569 387 583
rect 361 552 366 569
rect 383 552 387 569
rect 361 541 387 552
rect 412 660 436 676
rect 412 643 415 660
rect 432 643 436 660
rect 412 618 436 643
rect 412 601 415 618
rect 432 601 436 618
rect 412 575 436 601
rect 412 558 415 575
rect 432 558 436 575
rect 412 541 436 558
rect 40 500 57 508
rect 40 475 57 483
rect 88 456 105 464
rect 169 456 186 541
rect 169 439 255 456
rect 88 431 105 439
rect 136 412 153 420
rect 136 387 153 395
rect 184 368 201 376
rect 184 343 201 351
rect 218 323 235 396
rect 25 306 235 323
rect 25 209 42 306
rect 252 289 269 439
rect 316 376 333 541
rect 316 359 402 376
rect 380 342 402 359
rect 380 333 385 342
rect 218 272 269 289
rect 286 311 303 319
rect 385 317 402 325
rect 286 286 303 294
rect 419 298 436 541
rect 218 209 235 272
rect 334 268 351 276
rect 334 243 351 251
rect 18 191 42 209
rect 18 174 22 191
rect 39 174 42 191
rect 18 154 42 174
rect 115 191 138 209
rect 115 174 118 191
rect 135 174 138 191
rect 115 154 138 174
rect 211 191 235 209
rect 211 174 214 191
rect 231 174 235 191
rect 211 154 235 174
rect 264 191 288 209
rect 264 174 268 191
rect 285 174 288 191
rect 264 154 288 174
rect 361 191 384 209
rect 419 196 436 281
rect 361 174 364 191
rect 381 174 384 191
rect 361 154 384 174
rect 412 184 436 196
rect 412 167 415 184
rect 432 167 436 184
rect 412 154 436 167
rect 463 660 487 676
rect 463 643 467 660
rect 484 643 487 660
rect 463 618 487 643
rect 463 601 467 618
rect 484 601 487 618
rect 463 575 487 601
rect 463 558 467 575
rect 484 558 487 575
rect 463 541 487 558
rect 512 660 535 676
rect 512 643 515 660
rect 532 643 535 660
rect 512 618 535 643
rect 512 601 515 618
rect 532 601 535 618
rect 512 575 535 601
rect 512 558 515 575
rect 532 558 535 575
rect 512 541 535 558
rect 560 660 584 676
rect 560 643 563 660
rect 580 643 584 660
rect 560 618 584 643
rect 560 601 563 618
rect 580 601 584 618
rect 560 575 584 601
rect 560 558 563 575
rect 580 558 584 575
rect 560 541 584 558
rect 463 342 480 541
rect 533 449 550 457
rect 533 424 550 432
rect 567 439 584 541
rect 567 422 571 439
rect 497 385 514 393
rect 497 360 514 368
rect 463 196 480 325
rect 567 196 584 422
rect 463 184 487 196
rect 463 167 467 184
rect 484 167 487 184
rect 463 154 487 167
rect 512 184 535 196
rect 512 167 515 184
rect 532 167 535 184
rect 512 154 535 167
rect 560 184 584 196
rect 560 167 563 184
rect 580 167 584 184
rect 560 154 584 167
rect 118 17 135 154
rect 364 17 381 154
rect 515 17 532 154
rect 69 9 532 17
rect 69 -9 101 9
rect 119 -9 228 9
rect 246 -9 356 9
rect 374 -9 483 9
rect 500 -9 532 9
rect 69 -17 532 -9
<< viali >>
rect 101 760 119 778
rect 228 760 246 778
rect 356 760 374 778
rect 483 760 501 778
rect 70 553 87 570
rect 40 483 57 500
rect 88 439 105 456
rect 255 439 272 456
rect 136 395 153 412
rect 218 396 235 413
rect 184 351 201 368
rect 385 325 402 342
rect 286 294 303 311
rect 419 281 436 298
rect 334 251 351 268
rect 268 174 285 191
rect 533 432 550 449
rect 571 422 588 439
rect 497 368 514 385
rect 463 325 480 342
rect 101 -9 119 9
rect 228 -9 246 9
rect 356 -9 374 9
rect 483 -9 500 9
<< metal1 >>
rect 0 778 602 784
rect 0 760 101 778
rect 119 760 228 778
rect 246 760 356 778
rect 374 760 483 778
rect 501 760 602 778
rect 0 754 602 760
rect 67 570 90 576
rect 67 553 70 570
rect 87 561 90 570
rect 87 553 238 561
rect 67 547 238 553
rect 36 500 63 507
rect 36 490 40 500
rect 35 483 40 490
rect 57 483 63 500
rect 35 476 63 483
rect 84 456 111 463
rect 84 446 88 456
rect 83 439 88 446
rect 105 439 111 456
rect 83 432 111 439
rect 224 419 238 547
rect 252 456 275 462
rect 252 439 255 456
rect 272 447 275 456
rect 529 449 553 455
rect 529 447 533 449
rect 272 439 533 447
rect 252 433 533 439
rect 529 432 533 433
rect 550 432 553 449
rect 529 425 553 432
rect 568 439 591 446
rect 132 412 159 419
rect 132 402 136 412
rect 131 395 136 402
rect 153 395 159 412
rect 131 388 159 395
rect 215 413 238 419
rect 568 422 571 439
rect 588 438 591 439
rect 588 424 602 438
rect 588 422 591 424
rect 568 415 591 422
rect 215 396 218 413
rect 235 403 238 413
rect 235 396 517 403
rect 215 389 517 396
rect 494 385 517 389
rect 180 368 207 375
rect 180 358 184 368
rect 179 351 184 358
rect 201 351 207 368
rect 494 368 497 385
rect 514 368 517 385
rect 494 362 517 368
rect 179 344 207 351
rect 556 351 602 365
rect 371 342 406 349
rect 371 325 385 342
rect 402 325 406 342
rect 371 319 406 325
rect 460 343 483 348
rect 556 343 570 351
rect 460 342 570 343
rect 460 325 463 342
rect 480 329 570 342
rect 480 325 483 329
rect 460 319 483 325
rect 282 311 309 318
rect 282 301 286 311
rect 281 294 286 301
rect 303 294 309 311
rect 281 287 309 294
rect 330 268 357 275
rect 330 258 334 268
rect 329 251 334 258
rect 351 251 357 268
rect 329 244 357 251
rect 371 197 385 319
rect 416 298 602 304
rect 416 281 419 298
rect 436 290 602 298
rect 436 281 439 290
rect 416 275 439 281
rect 265 191 385 197
rect 265 174 268 191
rect 285 183 385 191
rect 285 174 288 183
rect 265 168 288 174
rect 0 9 602 15
rect 0 -9 101 9
rect 119 -9 228 9
rect 246 -9 356 9
rect 374 -9 483 9
rect 500 -9 602 9
rect 0 -15 602 -9
<< labels >>
flabel metal1 281 294 281 294 0 FreeSans 80 0 0 0 A2
port 5 nsew
flabel metal1 595 297 595 297 0 FreeSans 80 0 0 0 OUT2
port 9 nsew
flabel ndiff 78 178 78 178 0 FreeSans 80 0 0 0 net1
flabel metal1 229 478 229 478 0 FreeSans 80 0 0 0 net2
flabel ndiff 174 177 174 177 0 FreeSans 80 0 0 0 net3
flabel metal1 280 438 280 438 0 FreeSans 80 0 0 0 net4
flabel ndiff 326 174 326 174 0 FreeSans 80 0 0 0 net5
flabel metal1 378 281 378 281 0 FreeSans 80 0 0 0 net6
flabel metal1 298 764 298 764 0 FreeSans 80 0 0 0 vdd
port 10 nsew
flabel metal1 284 0 284 0 0 FreeSans 80 0 0 0 gnd
port 11 nsew
flabel metal1 596 431 596 431 0 FreeSans 80 0 0 0 OUT0
port 12 nsew
flabel metal1 594 357 594 357 0 FreeSans 80 0 0 0 OUT1
port 13 nsew
flabel metal1 35 482 35 482 0 FreeSans 80 0 0 0 A0
port 0 nsew
flabel metal1 83 438 83 438 0 FreeSans 80 0 0 0 B0
port 1 nsew
flabel metal1 131 393 131 393 0 FreeSans 80 0 0 0 A1
port 3 nsew
flabel metal1 179 350 179 350 0 FreeSans 80 0 0 0 B1
port 4 nsew
flabel metal1 329 250 329 250 0 FreeSans 80 0 0 0 B2
port 6 nsew
<< properties >>
string FIXED_BBOX 0 -21 602 769
<< end >>
