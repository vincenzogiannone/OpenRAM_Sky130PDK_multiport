magic
tech sky130A
magscale 1 2
timestamp 1643678851
<< checkpaint >>
rect -1271 -1302 6690 50504
<< viali >>
rect 2545 30047 2579 30081
rect 2545 28423 2579 28457
rect 2545 26967 2579 27001
rect 2545 25343 2579 25377
rect 2545 23887 2579 23921
rect 2545 22263 2579 22297
rect 2545 20807 2579 20841
rect 2545 19183 2579 19217
rect 2545 14651 2579 14685
rect 2545 13027 2579 13061
rect 2545 11571 2579 11605
rect 2545 9947 2579 9981
rect 2545 5415 2579 5449
rect 2545 3791 2579 3825
rect 2545 2335 2579 2369
rect 2545 711 2579 745
<< metal1 >>
rect 3692 47954 4844 47982
rect 3284 47898 4748 47926
rect 2944 47842 4652 47870
rect 4984 47840 5350 47868
rect 3692 47786 4448 47814
rect 3284 47730 4352 47758
rect 5066 47718 5350 47746
rect 2876 47674 4256 47702
rect 3692 47618 4160 47646
rect 3284 47562 4064 47590
rect 5274 47572 5350 47600
rect 2808 47506 3968 47534
rect 2876 46334 3968 46362
rect 3216 46278 4064 46306
rect 5274 46268 5350 46296
rect 3692 46222 4160 46250
rect 2944 46166 4256 46194
rect 3216 46110 4352 46138
rect 5066 46122 5350 46150
rect 3692 46054 4448 46082
rect 3012 45998 4652 46026
rect 4984 46000 5350 46028
rect 3216 45942 4748 45970
rect 3692 45886 4844 45914
rect 3692 44926 4844 44954
rect 3216 44870 4748 44898
rect 2808 44814 4652 44842
rect 4984 44812 5350 44840
rect 3692 44758 4448 44786
rect 3148 44702 4352 44730
rect 5066 44690 5350 44718
rect 3012 44646 4256 44674
rect 3692 44590 4160 44618
rect 3148 44534 4064 44562
rect 5274 44544 5350 44572
rect 2944 44478 3968 44506
rect 3012 43306 3968 43334
rect 3080 43250 4064 43278
rect 5274 43240 5350 43268
rect 3692 43194 4160 43222
rect 2808 43138 4256 43166
rect 3148 43082 4352 43110
rect 5066 43094 5350 43122
rect 3692 43026 4448 43054
rect 2876 42970 4652 42998
rect 4984 42972 5350 43000
rect 3148 42914 4748 42942
rect 3692 42858 4844 42886
rect 3692 41898 4844 41926
rect 3080 41842 4748 41870
rect 2944 41786 4652 41814
rect 4984 41784 5350 41812
rect 3692 41730 4448 41758
rect 3080 41674 4352 41702
rect 5066 41662 5350 41690
rect 2876 41618 4256 41646
rect 3692 41562 4160 41590
rect 3080 41506 4064 41534
rect 5274 41516 5350 41544
rect 2808 41450 3968 41478
rect 2876 40278 3968 40306
rect 3284 40222 4064 40250
rect 5274 40212 5350 40240
rect 3624 40166 4160 40194
rect 2944 40110 4256 40138
rect 3284 40054 4352 40082
rect 5066 40066 5350 40094
rect 3624 39998 4448 40026
rect 3012 39942 4652 39970
rect 4984 39944 5350 39972
rect 3284 39886 4748 39914
rect 3624 39830 4844 39858
rect 3624 38870 4844 38898
rect 3284 38814 4748 38842
rect 2808 38758 4652 38786
rect 4984 38756 5350 38784
rect 3624 38702 4448 38730
rect 3216 38646 4352 38674
rect 5066 38634 5350 38662
rect 3012 38590 4256 38618
rect 3624 38534 4160 38562
rect 3216 38478 4064 38506
rect 5274 38488 5350 38516
rect 2944 38422 3968 38450
rect 3012 37250 3968 37278
rect 3148 37194 4064 37222
rect 5274 37184 5350 37212
rect 3624 37138 4160 37166
rect 2808 37082 4256 37110
rect 3216 37026 4352 37054
rect 5066 37038 5350 37066
rect 3624 36970 4448 36998
rect 2876 36914 4652 36942
rect 4984 36916 5350 36944
rect 3216 36858 4748 36886
rect 3624 36802 4844 36830
rect 3624 35842 4844 35870
rect 3148 35786 4748 35814
rect 2944 35730 4652 35758
rect 4984 35728 5350 35756
rect 3624 35674 4448 35702
rect 3148 35618 4352 35646
rect 5066 35606 5350 35634
rect 2876 35562 4256 35590
rect 3624 35506 4160 35534
rect 3148 35450 4064 35478
rect 5274 35460 5350 35488
rect 2808 35394 3968 35422
rect 2876 34222 3968 34250
rect 3080 34166 4064 34194
rect 5274 34156 5350 34184
rect 3624 34110 4160 34138
rect 2944 34054 4256 34082
rect 3080 33998 4352 34026
rect 5066 34010 5350 34038
rect 3624 33942 4448 33970
rect 3012 33886 4652 33914
rect 4984 33888 5350 33916
rect 3080 33830 4748 33858
rect 3624 33774 4844 33802
rect 3624 32814 4844 32842
rect 3080 32758 4748 32786
rect 2808 32702 4652 32730
rect 4984 32700 5350 32728
rect 3556 32646 4448 32674
rect 3284 32590 4352 32618
rect 5066 32578 5350 32606
rect 3012 32534 4256 32562
rect 3556 32478 4160 32506
rect 3284 32422 4064 32450
rect 5274 32432 5350 32460
rect 2944 32366 3968 32394
rect 3012 31194 3968 31222
rect 3216 31138 4064 31166
rect 5274 31128 5350 31156
rect 3556 31082 4160 31110
rect 2808 31026 4256 31054
rect 3284 30970 4352 30998
rect 5066 30982 5350 31010
rect 3556 30914 4448 30942
rect 2876 30858 4652 30886
rect 4984 30860 5350 30888
rect 3284 30802 4748 30830
rect 3556 30746 4844 30774
rect 2533 30079 2536 30087
rect 2507 30049 2536 30079
rect 2533 30041 2536 30049
rect 2588 30079 2591 30087
rect 2588 30049 2618 30079
rect 2588 30041 2591 30049
rect 3556 29786 4844 29814
rect 3216 29730 4748 29758
rect 2944 29674 4652 29702
rect 4984 29672 5350 29700
rect 3556 29618 4448 29646
rect 3216 29562 4352 29590
rect 5066 29550 5350 29578
rect 2876 29506 4256 29534
rect 3556 29450 4160 29478
rect 3216 29394 4064 29422
rect 5274 29404 5350 29432
rect 2808 29338 3968 29366
rect 2533 28455 2536 28463
rect 2507 28425 2536 28455
rect 2533 28417 2536 28425
rect 2588 28455 2591 28463
rect 2588 28425 2618 28455
rect 2588 28417 2591 28425
rect 2876 28166 3968 28194
rect 3148 28110 4064 28138
rect 5274 28100 5350 28128
rect 3556 28054 4160 28082
rect 2944 27998 4256 28026
rect 3148 27942 4352 27970
rect 5066 27954 5350 27982
rect 3556 27886 4448 27914
rect 3012 27830 4652 27858
rect 4984 27832 5350 27860
rect 3148 27774 4748 27802
rect 3556 27718 4844 27746
rect 2533 26999 2536 27007
rect 2507 26969 2536 26999
rect 2533 26961 2536 26969
rect 2588 26999 2591 27007
rect 2588 26969 2618 26999
rect 2588 26961 2591 26969
rect 3556 26758 4844 26786
rect 3148 26702 4748 26730
rect 2808 26646 4652 26674
rect 4984 26644 5350 26672
rect 3556 26590 4448 26618
rect 3080 26534 4352 26562
rect 5066 26522 5350 26550
rect 3012 26478 4256 26506
rect 3556 26422 4160 26450
rect 3080 26366 4064 26394
rect 5274 26376 5350 26404
rect 2944 26310 3968 26338
rect 2533 25375 2536 25383
rect 2507 25345 2536 25375
rect 2533 25337 2536 25345
rect 2588 25375 2591 25383
rect 2588 25345 2618 25375
rect 2588 25337 2591 25345
rect 3012 25138 3968 25166
rect 3284 25082 4064 25110
rect 5274 25072 5350 25100
rect 3488 25026 4160 25054
rect 2808 24970 4256 24998
rect 3080 24914 4352 24942
rect 5066 24926 5350 24954
rect 3556 24858 4448 24886
rect 2876 24802 4652 24830
rect 4984 24804 5350 24832
rect 3080 24746 4748 24774
rect 3556 24690 4844 24718
rect 2533 23919 2536 23927
rect 2507 23889 2536 23919
rect 2533 23881 2536 23889
rect 2588 23919 2591 23927
rect 2588 23889 2618 23919
rect 2588 23881 2591 23889
rect 3488 23730 4844 23758
rect 3284 23674 4748 23702
rect 2944 23618 4652 23646
rect 4984 23616 5350 23644
rect 3488 23562 4448 23590
rect 3284 23506 4352 23534
rect 5066 23494 5350 23522
rect 2876 23450 4256 23478
rect 3488 23394 4160 23422
rect 3284 23338 4064 23366
rect 5274 23348 5350 23376
rect 2808 23282 3968 23310
rect 449 22266 697 22294
rect 2533 22295 2536 22303
rect 2507 22265 2536 22295
rect 2533 22257 2536 22265
rect 2588 22295 2591 22303
rect 2588 22265 2618 22295
rect 2588 22257 2591 22265
rect 2876 22110 3968 22138
rect 3216 22054 4064 22082
rect 5274 22044 5350 22072
rect 3488 21998 4160 22026
rect 2944 21942 4256 21970
rect 3216 21886 4352 21914
rect 5066 21898 5350 21926
rect 3488 21830 4448 21858
rect 3012 21774 4652 21802
rect 4984 21776 5350 21804
rect 3216 21718 4748 21746
rect 3488 21662 4844 21690
rect 381 20810 629 20838
rect 2533 20839 2536 20847
rect 2507 20809 2536 20839
rect 2533 20801 2536 20809
rect 2588 20839 2591 20847
rect 2588 20809 2618 20839
rect 2588 20801 2591 20809
rect 3488 20702 4844 20730
rect 3216 20646 4748 20674
rect 2808 20590 4652 20618
rect 4984 20588 5350 20616
rect 3488 20534 4448 20562
rect 3148 20478 4352 20506
rect 5066 20466 5350 20494
rect 3012 20422 4256 20450
rect 3488 20366 4160 20394
rect 3148 20310 4064 20338
rect 5274 20320 5350 20348
rect 2944 20254 3968 20282
rect 313 19186 561 19214
rect 2533 19215 2536 19223
rect 2507 19185 2536 19215
rect 2533 19177 2536 19185
rect 2588 19215 2591 19223
rect 2588 19185 2618 19215
rect 2588 19177 2591 19185
rect 3012 19082 3968 19110
rect 3080 19026 4064 19054
rect 5274 19016 5350 19044
rect 3488 18970 4160 18998
rect 2808 18914 4256 18942
rect 3148 18858 4352 18886
rect 5066 18870 5350 18898
rect 3488 18802 4448 18830
rect 2876 18746 4652 18774
rect 4984 18748 5350 18776
rect 3148 18690 4748 18718
rect 3488 18634 4844 18662
rect 3488 17674 4844 17702
rect 3080 17618 4748 17646
rect 2944 17562 4652 17590
rect 4984 17560 5350 17588
rect 3488 17506 4448 17534
rect 3080 17450 4352 17478
rect 5066 17438 5350 17466
rect 2876 17394 4256 17422
rect 3488 17338 4160 17366
rect 3080 17282 4064 17310
rect 5274 17292 5350 17320
rect 2808 17226 3968 17254
rect 2876 16054 3968 16082
rect 3284 15998 4064 16026
rect 5274 15988 5350 16016
rect 3420 15942 4160 15970
rect 2944 15886 4256 15914
rect 3284 15830 4352 15858
rect 5066 15842 5350 15870
rect 3420 15774 4448 15802
rect 3012 15718 4652 15746
rect 4984 15720 5350 15748
rect 3284 15662 4748 15690
rect 3420 15606 4844 15634
rect 2533 14683 2536 14691
rect 2507 14653 2536 14683
rect 2533 14645 2536 14653
rect 2588 14683 2591 14691
rect 2588 14653 2618 14683
rect 2588 14645 2591 14653
rect 3420 14646 4844 14674
rect 3284 14590 4748 14618
rect 2808 14534 4652 14562
rect 4984 14532 5350 14560
rect 3420 14478 4448 14506
rect 3216 14422 4352 14450
rect 5066 14410 5350 14438
rect 3012 14366 4256 14394
rect 3420 14310 4160 14338
rect 3216 14254 4064 14282
rect 5274 14264 5350 14292
rect 2944 14198 3968 14226
rect 2533 13059 2536 13067
rect 2507 13029 2536 13059
rect 2533 13021 2536 13029
rect 2588 13059 2591 13067
rect 2588 13029 2618 13059
rect 2588 13021 2591 13029
rect 3012 13026 3968 13054
rect 3148 12970 4064 12998
rect 5274 12960 5350 12988
rect 3420 12914 4160 12942
rect 2808 12858 4256 12886
rect 3216 12802 4352 12830
rect 5066 12814 5350 12842
rect 3420 12746 4448 12774
rect 2876 12690 4652 12718
rect 4984 12692 5350 12720
rect 3216 12634 4748 12662
rect 3420 12578 4844 12606
rect 245 11574 991 11602
rect 2533 11603 2536 11611
rect 2507 11573 2536 11603
rect 2533 11565 2536 11573
rect 2588 11603 2591 11611
rect 3420 11618 4844 11646
rect 2588 11573 2618 11603
rect 2588 11565 2591 11573
rect 3148 11562 4748 11590
rect 2944 11506 4652 11534
rect 4984 11504 5350 11532
rect 3420 11450 4448 11478
rect 3148 11394 4352 11422
rect 5066 11382 5350 11410
rect 2876 11338 4256 11366
rect 3420 11282 4160 11310
rect 3148 11226 4064 11254
rect 5274 11236 5350 11264
rect 2808 11170 3968 11198
rect 177 9950 923 9978
rect 2533 9979 2536 9987
rect 2507 9949 2536 9979
rect 2533 9941 2536 9949
rect 2588 9979 2591 9987
rect 2876 9998 3968 10026
rect 2588 9949 2618 9979
rect 2588 9941 2591 9949
rect 3080 9942 4064 9970
rect 5274 9932 5350 9960
rect 3420 9886 4160 9914
rect 2944 9830 4256 9858
rect 3080 9774 4352 9802
rect 5066 9786 5350 9814
rect 3420 9718 4448 9746
rect 3012 9662 4652 9690
rect 4984 9664 5350 9692
rect 3080 9606 4748 9634
rect 3420 9550 4844 9578
rect 3420 8590 4844 8618
rect 3080 8534 4748 8562
rect 2808 8478 4652 8506
rect 4984 8476 5350 8504
rect 3352 8422 4448 8450
rect 3284 8366 4352 8394
rect 5066 8354 5350 8382
rect 3012 8310 4256 8338
rect 3352 8254 4160 8282
rect 3284 8198 4064 8226
rect 5274 8208 5350 8236
rect 2944 8142 3968 8170
rect 3012 6970 3968 6998
rect 3216 6914 4064 6942
rect 5274 6904 5350 6932
rect 3352 6858 4160 6886
rect 2808 6802 4256 6830
rect 3284 6746 4352 6774
rect 5066 6758 5350 6786
rect 3352 6690 4448 6718
rect 2876 6634 4652 6662
rect 4984 6636 5350 6664
rect 3284 6578 4748 6606
rect 3352 6522 4844 6550
rect 3352 5562 4844 5590
rect 3216 5506 4748 5534
rect 2533 5447 2536 5455
rect 2507 5417 2536 5447
rect 2533 5409 2536 5417
rect 2588 5447 2591 5455
rect 2588 5417 2618 5447
rect 2944 5450 4652 5478
rect 4984 5448 5350 5476
rect 2588 5409 2591 5417
rect 3352 5394 4448 5422
rect 3216 5338 4352 5366
rect 5066 5326 5350 5354
rect 2876 5282 4256 5310
rect 3352 5226 4160 5254
rect 3216 5170 4064 5198
rect 5274 5180 5350 5208
rect 2808 5114 3968 5142
rect 2876 3942 3968 3970
rect 3148 3886 4064 3914
rect 5274 3876 5350 3904
rect 2533 3823 2536 3831
rect 2507 3793 2536 3823
rect 2533 3785 2536 3793
rect 2588 3823 2591 3831
rect 2588 3793 2618 3823
rect 3352 3830 4160 3858
rect 2588 3785 2591 3793
rect 2944 3774 4256 3802
rect 3148 3718 4352 3746
rect 5066 3730 5350 3758
rect 3352 3662 4448 3690
rect 3012 3606 4652 3634
rect 4984 3608 5350 3636
rect 3148 3550 4748 3578
rect 3352 3494 4844 3522
rect 3352 2534 4844 2562
rect 3148 2478 4748 2506
rect 2808 2422 4652 2450
rect 4984 2420 5350 2448
rect 109 2338 991 2366
rect 2533 2367 2536 2375
rect 2507 2337 2536 2367
rect 2533 2329 2536 2337
rect 2588 2367 2591 2375
rect 2588 2337 2618 2367
rect 3352 2366 4448 2394
rect 2588 2329 2591 2337
rect 3080 2310 4352 2338
rect 5066 2298 5350 2326
rect 3012 2254 4256 2282
rect 3352 2198 4160 2226
rect 3080 2142 4064 2170
rect 5274 2152 5350 2180
rect 2944 2086 3968 2114
rect 2784 914 2960 942
rect 2880 858 3232 886
rect 5274 848 5350 876
rect 2976 802 3640 830
rect 41 714 923 742
rect 2533 743 2536 751
rect 2507 713 2536 743
rect 2533 705 2536 713
rect 2588 743 2591 751
rect 2588 713 2618 743
rect 2808 746 4256 774
rect 2588 705 2591 713
rect 3080 690 4352 718
rect 5066 702 5350 730
rect 3352 634 4448 662
rect 2876 578 4652 606
rect 4984 580 5350 608
rect 3080 522 4748 550
rect 3352 466 4844 494
<< via1 >>
rect 5338 48422 5390 48474
rect 3640 47942 3692 47994
rect 3232 47886 3284 47938
rect 2892 47830 2944 47882
rect 3640 47774 3692 47826
rect 3232 47718 3284 47770
rect 2824 47662 2876 47714
rect 3640 47606 3692 47658
rect 3232 47550 3284 47602
rect 2756 47494 2808 47546
rect 5338 46908 5390 46960
rect 2824 46322 2876 46374
rect 3164 46266 3216 46318
rect 3640 46210 3692 46262
rect 2892 46154 2944 46206
rect 3164 46098 3216 46150
rect 3640 46042 3692 46094
rect 2960 45986 3012 46038
rect 3164 45930 3216 45982
rect 3640 45874 3692 45926
rect 5338 45394 5390 45446
rect 3640 44914 3692 44966
rect 3164 44858 3216 44910
rect 2756 44802 2808 44854
rect 3640 44746 3692 44798
rect 3096 44690 3148 44742
rect 2960 44634 3012 44686
rect 3640 44578 3692 44630
rect 3096 44522 3148 44574
rect 2892 44466 2944 44518
rect 5338 43880 5390 43932
rect 2960 43294 3012 43346
rect 3028 43238 3080 43290
rect 3640 43182 3692 43234
rect 2756 43126 2808 43178
rect 3096 43070 3148 43122
rect 3640 43014 3692 43066
rect 2824 42958 2876 43010
rect 3096 42902 3148 42954
rect 3640 42846 3692 42898
rect 5338 42366 5390 42418
rect 3640 41886 3692 41938
rect 3028 41830 3080 41882
rect 2892 41774 2944 41826
rect 3640 41718 3692 41770
rect 3028 41662 3080 41714
rect 2824 41606 2876 41658
rect 3640 41550 3692 41602
rect 3028 41494 3080 41546
rect 2756 41438 2808 41490
rect 5338 40852 5390 40904
rect 2824 40266 2876 40318
rect 3232 40210 3284 40262
rect 3572 40154 3624 40206
rect 2892 40098 2944 40150
rect 3232 40042 3284 40094
rect 3572 39986 3624 40038
rect 2960 39930 3012 39982
rect 3232 39874 3284 39926
rect 3572 39818 3624 39870
rect 5338 39338 5390 39390
rect 3572 38858 3624 38910
rect 3232 38802 3284 38854
rect 2756 38746 2808 38798
rect 3572 38690 3624 38742
rect 3164 38634 3216 38686
rect 2960 38578 3012 38630
rect 3572 38522 3624 38574
rect 3164 38466 3216 38518
rect 2892 38410 2944 38462
rect 5338 37824 5390 37876
rect 2960 37238 3012 37290
rect 3096 37182 3148 37234
rect 3572 37126 3624 37178
rect 2756 37070 2808 37122
rect 3164 37014 3216 37066
rect 3572 36958 3624 37010
rect 2824 36902 2876 36954
rect 3164 36846 3216 36898
rect 3572 36790 3624 36842
rect 5338 36310 5390 36362
rect 3572 35830 3624 35882
rect 3096 35774 3148 35826
rect 2892 35718 2944 35770
rect 3572 35662 3624 35714
rect 3096 35606 3148 35658
rect 2824 35550 2876 35602
rect 3572 35494 3624 35546
rect 3096 35438 3148 35490
rect 2756 35382 2808 35434
rect 5338 34796 5390 34848
rect 2824 34210 2876 34262
rect 3028 34154 3080 34206
rect 3572 34098 3624 34150
rect 2892 34042 2944 34094
rect 3028 33986 3080 34038
rect 3572 33930 3624 33982
rect 2960 33874 3012 33926
rect 3028 33818 3080 33870
rect 3572 33762 3624 33814
rect 5338 33282 5390 33334
rect 3572 32802 3624 32854
rect 3028 32746 3080 32798
rect 2756 32690 2808 32742
rect 3504 32634 3556 32686
rect 3232 32578 3284 32630
rect 2960 32522 3012 32574
rect 3504 32466 3556 32518
rect 3232 32410 3284 32462
rect 2892 32354 2944 32406
rect 5338 31768 5390 31820
rect 2960 31182 3012 31234
rect 3164 31126 3216 31178
rect 3504 31070 3556 31122
rect 2756 31014 2808 31066
rect 3232 30958 3284 31010
rect 3504 30902 3556 30954
rect 2824 30846 2876 30898
rect 3232 30790 3284 30842
rect 3504 30734 3556 30786
rect 5338 30254 5390 30306
rect 2536 30081 2588 30090
rect 2536 30047 2545 30081
rect 2545 30047 2579 30081
rect 2579 30047 2588 30081
rect 2536 30038 2588 30047
rect 3504 29774 3556 29826
rect 3164 29718 3216 29770
rect 2892 29662 2944 29714
rect 3504 29606 3556 29658
rect 3164 29550 3216 29602
rect 2824 29494 2876 29546
rect 3504 29438 3556 29490
rect 3164 29382 3216 29434
rect 2756 29326 2808 29378
rect 5338 28740 5390 28792
rect 2536 28457 2588 28466
rect 2536 28423 2545 28457
rect 2545 28423 2579 28457
rect 2579 28423 2588 28457
rect 2536 28414 2588 28423
rect 2824 28154 2876 28206
rect 3096 28098 3148 28150
rect 3504 28042 3556 28094
rect 2892 27986 2944 28038
rect 3096 27930 3148 27982
rect 3504 27874 3556 27926
rect 2960 27818 3012 27870
rect 3096 27762 3148 27814
rect 3504 27706 3556 27758
rect 5338 27226 5390 27278
rect 2536 27001 2588 27010
rect 2536 26967 2545 27001
rect 2545 26967 2579 27001
rect 2579 26967 2588 27001
rect 2536 26958 2588 26967
rect 3504 26746 3556 26798
rect 3096 26690 3148 26742
rect 2756 26634 2808 26686
rect 3504 26578 3556 26630
rect 3028 26522 3080 26574
rect 2960 26466 3012 26518
rect 3504 26410 3556 26462
rect 3028 26354 3080 26406
rect 2892 26298 2944 26350
rect 5338 25712 5390 25764
rect 2536 25377 2588 25386
rect 2536 25343 2545 25377
rect 2545 25343 2579 25377
rect 2579 25343 2588 25377
rect 2536 25334 2588 25343
rect 2960 25126 3012 25178
rect 3232 25070 3284 25122
rect 3436 25014 3488 25066
rect 2756 24958 2808 25010
rect 3028 24902 3080 24954
rect 3504 24846 3556 24898
rect 2824 24790 2876 24842
rect 3028 24734 3080 24786
rect 3504 24678 3556 24730
rect 5338 24198 5390 24250
rect 2536 23921 2588 23930
rect 2536 23887 2545 23921
rect 2545 23887 2579 23921
rect 2579 23887 2588 23921
rect 2536 23878 2588 23887
rect 3436 23718 3488 23770
rect 3232 23662 3284 23714
rect 2892 23606 2944 23658
rect 3436 23550 3488 23602
rect 3232 23494 3284 23546
rect 2824 23438 2876 23490
rect 3436 23382 3488 23434
rect 3232 23326 3284 23378
rect 2756 23270 2808 23322
rect 5338 22684 5390 22736
rect 397 22254 449 22306
rect 697 22254 749 22306
rect 2536 22297 2588 22306
rect 2536 22263 2545 22297
rect 2545 22263 2579 22297
rect 2579 22263 2588 22297
rect 2536 22254 2588 22263
rect 2824 22098 2876 22150
rect 3164 22042 3216 22094
rect 3436 21986 3488 22038
rect 2892 21930 2944 21982
rect 3164 21874 3216 21926
rect 3436 21818 3488 21870
rect 2960 21762 3012 21814
rect 3164 21706 3216 21758
rect 3436 21650 3488 21702
rect 5338 21170 5390 21222
rect 329 20798 381 20850
rect 629 20798 681 20850
rect 2536 20841 2588 20850
rect 2536 20807 2545 20841
rect 2545 20807 2579 20841
rect 2579 20807 2588 20841
rect 2536 20798 2588 20807
rect 3436 20690 3488 20742
rect 3164 20634 3216 20686
rect 2756 20578 2808 20630
rect 3436 20522 3488 20574
rect 3096 20466 3148 20518
rect 2960 20410 3012 20462
rect 3436 20354 3488 20406
rect 3096 20298 3148 20350
rect 2892 20242 2944 20294
rect 5338 19656 5390 19708
rect 261 19174 313 19226
rect 561 19174 613 19226
rect 2536 19217 2588 19226
rect 2536 19183 2545 19217
rect 2545 19183 2579 19217
rect 2579 19183 2588 19217
rect 2536 19174 2588 19183
rect 2960 19070 3012 19122
rect 3028 19014 3080 19066
rect 3436 18958 3488 19010
rect 2756 18902 2808 18954
rect 3096 18846 3148 18898
rect 3436 18790 3488 18842
rect 2824 18734 2876 18786
rect 3096 18678 3148 18730
rect 3436 18622 3488 18674
rect 5338 18142 5390 18194
rect 3436 17662 3488 17714
rect 3028 17606 3080 17658
rect 2892 17550 2944 17602
rect 3436 17494 3488 17546
rect 3028 17438 3080 17490
rect 2824 17382 2876 17434
rect 3436 17326 3488 17378
rect 3028 17270 3080 17322
rect 2756 17214 2808 17266
rect 5338 16628 5390 16680
rect 2824 16042 2876 16094
rect 3232 15986 3284 16038
rect 3368 15930 3420 15982
rect 2892 15874 2944 15926
rect 3232 15818 3284 15870
rect 3368 15762 3420 15814
rect 2960 15706 3012 15758
rect 3232 15650 3284 15702
rect 3368 15594 3420 15646
rect 5338 15114 5390 15166
rect 2536 14685 2588 14694
rect 2536 14651 2545 14685
rect 2545 14651 2579 14685
rect 2579 14651 2588 14685
rect 2536 14642 2588 14651
rect 3368 14634 3420 14686
rect 3232 14578 3284 14630
rect 2756 14522 2808 14574
rect 3368 14466 3420 14518
rect 3164 14410 3216 14462
rect 2960 14354 3012 14406
rect 3368 14298 3420 14350
rect 3164 14242 3216 14294
rect 2892 14186 2944 14238
rect 5338 13600 5390 13652
rect 2536 13061 2588 13070
rect 2536 13027 2545 13061
rect 2545 13027 2579 13061
rect 2579 13027 2588 13061
rect 2536 13018 2588 13027
rect 2960 13014 3012 13066
rect 3096 12958 3148 13010
rect 3368 12902 3420 12954
rect 2756 12846 2808 12898
rect 3164 12790 3216 12842
rect 3368 12734 3420 12786
rect 2824 12678 2876 12730
rect 3164 12622 3216 12674
rect 3368 12566 3420 12618
rect 5338 12086 5390 12138
rect 193 11562 245 11614
rect 991 11562 1043 11614
rect 2536 11605 2588 11614
rect 2536 11571 2545 11605
rect 2545 11571 2579 11605
rect 2579 11571 2588 11605
rect 3368 11606 3420 11658
rect 2536 11562 2588 11571
rect 3096 11550 3148 11602
rect 2892 11494 2944 11546
rect 3368 11438 3420 11490
rect 3096 11382 3148 11434
rect 2824 11326 2876 11378
rect 3368 11270 3420 11322
rect 3096 11214 3148 11266
rect 2756 11158 2808 11210
rect 5338 10572 5390 10624
rect 125 9938 177 9990
rect 923 9938 975 9990
rect 2536 9981 2588 9990
rect 2536 9947 2545 9981
rect 2545 9947 2579 9981
rect 2579 9947 2588 9981
rect 2824 9986 2876 10038
rect 2536 9938 2588 9947
rect 3028 9930 3080 9982
rect 3368 9874 3420 9926
rect 2892 9818 2944 9870
rect 3028 9762 3080 9814
rect 3368 9706 3420 9758
rect 2960 9650 3012 9702
rect 3028 9594 3080 9646
rect 3368 9538 3420 9590
rect 5338 9058 5390 9110
rect 3368 8578 3420 8630
rect 3028 8522 3080 8574
rect 2756 8466 2808 8518
rect 3300 8410 3352 8462
rect 3232 8354 3284 8406
rect 2960 8298 3012 8350
rect 3300 8242 3352 8294
rect 3232 8186 3284 8238
rect 2892 8130 2944 8182
rect 5338 7544 5390 7596
rect 2960 6958 3012 7010
rect 3164 6902 3216 6954
rect 3300 6846 3352 6898
rect 2756 6790 2808 6842
rect 3232 6734 3284 6786
rect 3300 6678 3352 6730
rect 2824 6622 2876 6674
rect 3232 6566 3284 6618
rect 3300 6510 3352 6562
rect 5338 6030 5390 6082
rect 3300 5550 3352 5602
rect 3164 5494 3216 5546
rect 2536 5449 2588 5458
rect 2536 5415 2545 5449
rect 2545 5415 2579 5449
rect 2579 5415 2588 5449
rect 2892 5438 2944 5490
rect 2536 5406 2588 5415
rect 3300 5382 3352 5434
rect 3164 5326 3216 5378
rect 2824 5270 2876 5322
rect 3300 5214 3352 5266
rect 3164 5158 3216 5210
rect 2756 5102 2808 5154
rect 5338 4516 5390 4568
rect 2824 3930 2876 3982
rect 3096 3874 3148 3926
rect 2536 3825 2588 3834
rect 2536 3791 2545 3825
rect 2545 3791 2579 3825
rect 2579 3791 2588 3825
rect 3300 3818 3352 3870
rect 2536 3782 2588 3791
rect 2892 3762 2944 3814
rect 3096 3706 3148 3758
rect 3300 3650 3352 3702
rect 2960 3594 3012 3646
rect 3096 3538 3148 3590
rect 3300 3482 3352 3534
rect 5338 3002 5390 3054
rect 3300 2522 3352 2574
rect 3096 2466 3148 2518
rect 2756 2410 2808 2462
rect 57 2326 109 2378
rect 991 2326 1043 2378
rect 2536 2369 2588 2378
rect 2536 2335 2545 2369
rect 2545 2335 2579 2369
rect 2579 2335 2588 2369
rect 3300 2354 3352 2406
rect 2536 2326 2588 2335
rect 3028 2298 3080 2350
rect 2960 2242 3012 2294
rect 3300 2186 3352 2238
rect 3028 2130 3080 2182
rect 2892 2074 2944 2126
rect 5338 1488 5390 1540
rect 2960 902 3012 954
rect 3232 846 3284 898
rect 3640 790 3692 842
rect -11 702 41 754
rect 923 702 975 754
rect 2536 745 2588 754
rect 2536 711 2545 745
rect 2545 711 2579 745
rect 2579 711 2588 745
rect 2756 734 2808 786
rect 2536 702 2588 711
rect 3028 678 3080 730
rect 3300 622 3352 674
rect 2824 566 2876 618
rect 3028 510 3080 562
rect 3300 454 3352 506
rect 5338 -26 5390 26
<< metal2 >>
rect 2768 47546 2796 49244
rect 2836 47714 2864 49244
rect 2904 47882 2932 49244
rect 2768 44854 2796 47494
rect 2836 46374 2864 47662
rect 2768 43178 2796 44802
rect 2768 41490 2796 43126
rect 2836 43010 2864 46322
rect 2904 46206 2932 47830
rect 2904 44518 2932 46154
rect 2972 46038 3000 49244
rect 2972 44686 3000 45986
rect 2836 41658 2864 42958
rect 2904 41826 2932 44466
rect 2972 43346 3000 44634
rect 2768 38798 2796 41438
rect 2836 40318 2864 41606
rect 2768 37122 2796 38746
rect 2768 35434 2796 37070
rect 2836 36954 2864 40266
rect 2904 40150 2932 41774
rect 2904 38462 2932 40098
rect 2972 39982 3000 43294
rect 3040 43290 3068 49244
rect 3108 44742 3136 49244
rect 3176 46318 3204 49244
rect 3244 47938 3272 49244
rect 3244 47770 3272 47886
rect 3244 47602 3272 47718
rect 3176 46150 3204 46266
rect 3176 45982 3204 46098
rect 3176 44910 3204 45930
rect 3108 44574 3136 44690
rect 3040 41882 3068 43238
rect 3108 43122 3136 44522
rect 3108 42954 3136 43070
rect 3040 41714 3068 41830
rect 3040 41546 3068 41662
rect 2972 38630 3000 39930
rect 2836 35602 2864 36902
rect 2904 35770 2932 38410
rect 2972 37290 3000 38578
rect 2768 32742 2796 35382
rect 2836 34262 2864 35550
rect 2768 31066 2796 32690
rect 1 754 29 30792
rect 69 2378 97 30792
rect 137 9990 165 30792
rect 205 11614 233 30792
rect 273 19226 301 30792
rect 341 20850 369 30792
rect 409 22306 437 30792
rect 2542 30092 2582 30098
rect 2542 30030 2582 30036
rect 2768 29378 2796 31014
rect 2836 30898 2864 34210
rect 2904 34094 2932 35718
rect 2904 32406 2932 34042
rect 2972 33926 3000 37238
rect 3040 34206 3068 41494
rect 3108 37234 3136 42902
rect 3176 38686 3204 44858
rect 3244 40262 3272 47550
rect 3244 40094 3272 40210
rect 3244 39926 3272 40042
rect 3244 38854 3272 39874
rect 3176 38518 3204 38634
rect 3108 35826 3136 37182
rect 3176 37066 3204 38466
rect 3176 36898 3204 37014
rect 3108 35658 3136 35774
rect 3108 35490 3136 35606
rect 3040 34038 3068 34154
rect 2972 32574 3000 33874
rect 3040 33870 3068 33986
rect 3040 32798 3068 33818
rect 2836 29546 2864 30846
rect 2904 29714 2932 32354
rect 2972 31234 3000 32522
rect 2542 28468 2582 28474
rect 2542 28406 2582 28412
rect 2542 27012 2582 27018
rect 2542 26950 2582 26956
rect 2768 26686 2796 29326
rect 2836 28206 2864 29494
rect 2542 25388 2582 25394
rect 2542 25326 2582 25332
rect 2768 25010 2796 26634
rect 2542 23932 2582 23938
rect 2542 23870 2582 23876
rect 2768 23322 2796 24958
rect 2836 24842 2864 28154
rect 2904 28038 2932 29662
rect 2904 26350 2932 27986
rect 2972 27870 3000 31182
rect 2972 26518 3000 27818
rect 3040 26574 3068 32746
rect 3108 28150 3136 35438
rect 3176 31178 3204 36846
rect 3244 32630 3272 38802
rect 3244 32462 3272 32578
rect 3176 29770 3204 31126
rect 3244 31010 3272 32410
rect 3244 30842 3272 30958
rect 3176 29602 3204 29718
rect 3176 29434 3204 29550
rect 3108 27982 3136 28098
rect 3108 27814 3136 27930
rect 3108 26742 3136 27762
rect 2836 23490 2864 24790
rect 2904 23658 2932 26298
rect 2972 25178 3000 26466
rect 3040 26406 3068 26522
rect 2542 22308 2582 22314
rect 1 0 29 702
rect 69 0 97 2326
rect 137 0 165 9938
rect 205 0 233 11562
rect 273 0 301 19174
rect 341 0 369 20798
rect 409 0 437 22254
rect 2542 22246 2582 22252
rect 2542 20852 2582 20858
rect 2542 20790 2582 20796
rect 2768 20630 2796 23270
rect 2836 22150 2864 23438
rect 2542 19228 2582 19234
rect 2542 19166 2582 19172
rect 2768 18954 2796 20578
rect 2768 17266 2796 18902
rect 2836 18786 2864 22098
rect 2904 21982 2932 23606
rect 2904 20294 2932 21930
rect 2972 21814 3000 25126
rect 3040 24954 3068 26354
rect 3040 24786 3068 24902
rect 2972 20462 3000 21762
rect 2836 17434 2864 18734
rect 2904 17602 2932 20242
rect 2972 19122 3000 20410
rect 2542 14696 2582 14702
rect 2542 14634 2582 14640
rect 2768 14574 2796 17214
rect 2836 16094 2864 17382
rect 2542 13072 2582 13078
rect 2542 13010 2582 13016
rect 2768 12898 2796 14522
rect 2542 11616 2582 11622
rect 2542 11554 2582 11560
rect 2768 11210 2796 12846
rect 2836 12730 2864 16042
rect 2904 15926 2932 17550
rect 2904 14238 2932 15874
rect 2972 15758 3000 19070
rect 3040 19066 3068 24734
rect 3108 20518 3136 26690
rect 3176 22094 3204 29382
rect 3244 25122 3272 30790
rect 3244 23714 3272 25070
rect 3244 23546 3272 23662
rect 3244 23378 3272 23494
rect 3176 21926 3204 22042
rect 3176 21758 3204 21874
rect 3176 20686 3204 21706
rect 3108 20350 3136 20466
rect 3040 17658 3068 19014
rect 3108 18898 3136 20298
rect 3108 18730 3136 18846
rect 3040 17490 3068 17606
rect 3040 17322 3068 17438
rect 2972 14406 3000 15706
rect 2836 11378 2864 12678
rect 2904 11546 2932 14186
rect 2972 13066 3000 14354
rect 2542 9992 2582 9998
rect 2542 9930 2582 9936
rect 2768 8518 2796 11158
rect 2836 10038 2864 11326
rect 2768 6842 2796 8466
rect 2542 5460 2582 5466
rect 2542 5398 2582 5404
rect 2768 5154 2796 6790
rect 2836 6674 2864 9986
rect 2904 9870 2932 11494
rect 2904 8182 2932 9818
rect 2972 9702 3000 13014
rect 3040 9982 3068 17270
rect 3108 13010 3136 18678
rect 3176 14462 3204 20634
rect 3244 16038 3272 23326
rect 3312 18500 3340 49244
rect 3380 20040 3408 49244
rect 3448 25066 3476 49244
rect 3516 32686 3544 49244
rect 3584 40206 3612 49244
rect 3652 47994 3680 49244
rect 3652 47826 3680 47942
rect 3652 47658 3680 47774
rect 3652 46262 3680 47606
rect 3652 46094 3680 46210
rect 3652 45926 3680 46042
rect 3652 44966 3680 45874
rect 3652 44798 3680 44914
rect 3652 44630 3680 44746
rect 3652 43234 3680 44578
rect 3652 43066 3680 43182
rect 3652 42898 3680 43014
rect 3652 41938 3680 42846
rect 3652 41770 3680 41886
rect 3652 41602 3680 41718
rect 3584 40038 3612 40154
rect 3584 39870 3612 39986
rect 3584 38910 3612 39818
rect 3584 38742 3612 38858
rect 3584 38574 3612 38690
rect 3584 37178 3612 38522
rect 3584 37010 3612 37126
rect 3584 36842 3612 36958
rect 3584 35882 3612 36790
rect 3584 35714 3612 35830
rect 3584 35546 3612 35662
rect 3584 34150 3612 35494
rect 3584 33982 3612 34098
rect 3584 33814 3612 33930
rect 3584 32854 3612 33762
rect 3516 32518 3544 32634
rect 3516 31122 3544 32466
rect 3516 30954 3544 31070
rect 3516 30786 3544 30902
rect 3516 29826 3544 30734
rect 3516 29658 3544 29774
rect 3516 29490 3544 29606
rect 3516 28094 3544 29438
rect 3516 27926 3544 28042
rect 3516 27758 3544 27874
rect 3516 26798 3544 27706
rect 3516 26630 3544 26746
rect 3516 26462 3544 26578
rect 3448 23770 3476 25014
rect 3516 24898 3544 26410
rect 3516 24730 3544 24846
rect 3448 23602 3476 23718
rect 3448 23434 3476 23550
rect 3448 22167 3476 23382
rect 3516 23120 3544 24678
rect 3584 24660 3612 32802
rect 3652 26200 3680 41550
rect 3720 27740 3748 49244
rect 3788 29280 3816 49244
rect 5344 48476 5384 48482
rect 5344 48414 5384 48420
rect 5344 46962 5384 46968
rect 5344 46900 5384 46906
rect 5344 45448 5384 45454
rect 5344 45386 5384 45392
rect 5344 43934 5384 43940
rect 5344 43872 5384 43878
rect 5344 42420 5384 42426
rect 5344 42358 5384 42364
rect 5344 40906 5384 40912
rect 5344 40844 5384 40850
rect 5344 39392 5384 39398
rect 5344 39330 5384 39336
rect 5344 37878 5384 37884
rect 5344 37816 5384 37822
rect 5344 36364 5384 36370
rect 5344 36302 5384 36308
rect 5344 34850 5384 34856
rect 5344 34788 5384 34794
rect 5344 33336 5384 33342
rect 5344 33274 5384 33280
rect 5344 31822 5384 31828
rect 5344 31760 5384 31766
rect 5344 30308 5384 30314
rect 5344 30246 5384 30252
rect 3448 22038 3476 22111
rect 3448 21870 3476 21986
rect 3448 21702 3476 21818
rect 3448 20742 3476 21650
rect 3448 20574 3476 20690
rect 3448 20406 3476 20522
rect 3244 15870 3272 15986
rect 3244 15702 3272 15818
rect 3244 14630 3272 15650
rect 3176 14294 3204 14410
rect 3108 11602 3136 12958
rect 3176 12842 3204 14242
rect 3244 13884 3272 14578
rect 3176 12674 3204 12790
rect 3176 12344 3204 12622
rect 3108 11434 3136 11550
rect 3108 11266 3136 11382
rect 3108 10804 3136 11214
rect 3040 9814 3068 9930
rect 2972 8350 3000 9650
rect 3040 9646 3068 9762
rect 3040 9264 3068 9594
rect 3040 8574 3068 9208
rect 2836 5322 2864 6622
rect 2904 5490 2932 8130
rect 2972 7010 3000 8298
rect 2542 3836 2582 3842
rect 2542 3774 2582 3780
rect 2768 2462 2796 5102
rect 2836 3982 2864 5270
rect 2542 2380 2582 2386
rect 2542 2318 2582 2324
rect 2768 786 2796 2410
rect 2836 1568 2864 3930
rect 2904 3814 2932 5438
rect 2972 4648 3000 6958
rect 2904 3108 2932 3762
rect 2972 3646 3000 4592
rect 2904 2126 2932 3052
rect 2972 2294 3000 3594
rect 3040 2350 3068 8522
rect 3108 3926 3136 10748
rect 3176 6954 3204 12288
rect 3244 8406 3272 13828
rect 3312 8462 3340 18444
rect 3380 15982 3408 19984
rect 3448 19010 3476 20354
rect 3448 18842 3476 18958
rect 3448 18674 3476 18790
rect 3448 17714 3476 18622
rect 3448 17546 3476 17662
rect 3448 17378 3476 17494
rect 3380 15814 3408 15930
rect 3380 15646 3408 15762
rect 3380 14686 3408 15594
rect 3380 14518 3408 14634
rect 3380 14350 3408 14466
rect 3380 12954 3408 14298
rect 3380 12786 3408 12902
rect 3380 12618 3408 12734
rect 3380 11658 3408 12566
rect 3380 11490 3408 11606
rect 3380 11322 3408 11438
rect 3380 9926 3408 11270
rect 3380 9758 3408 9874
rect 3380 9590 3408 9706
rect 3380 8630 3408 9538
rect 3244 8238 3272 8354
rect 3312 8294 3340 8410
rect 3176 5546 3204 6902
rect 3244 6786 3272 8186
rect 3312 6898 3340 8242
rect 3244 6618 3272 6734
rect 3312 6730 3340 6846
rect 3176 5378 3204 5494
rect 3176 5210 3204 5326
rect 3108 3758 3136 3874
rect 3108 3590 3136 3706
rect 3108 2518 3136 3538
rect 2542 756 2582 762
rect 2542 694 2582 700
rect 2768 28 2796 734
rect 2836 618 2864 1512
rect 2836 0 2864 566
rect 2904 0 2932 2074
rect 2972 954 3000 2242
rect 3040 2182 3068 2298
rect 2972 0 3000 902
rect 3040 730 3068 2130
rect 3040 562 3068 678
rect 3040 0 3068 510
rect 3108 0 3136 2466
rect 3176 0 3204 5158
rect 3244 898 3272 6566
rect 3312 6562 3340 6678
rect 3312 5602 3340 6510
rect 3312 5434 3340 5550
rect 3312 5266 3340 5382
rect 3312 3870 3340 5214
rect 3312 3702 3340 3818
rect 3312 3534 3340 3650
rect 3312 2574 3340 3482
rect 3312 2406 3340 2522
rect 3312 2238 3340 2354
rect 3244 0 3272 846
rect 3312 674 3340 2186
rect 3312 506 3340 622
rect 3312 0 3340 454
rect 3380 0 3408 8578
rect 3448 0 3476 17326
rect 3516 0 3544 23064
rect 3584 0 3612 24604
rect 3652 842 3680 26144
rect 3652 0 3680 790
rect 3720 0 3748 27684
rect 3788 0 3816 29224
rect 5344 28794 5384 28800
rect 5344 28732 5384 28738
rect 5344 27280 5384 27286
rect 5344 27218 5384 27224
rect 5344 25766 5384 25772
rect 5344 25704 5384 25710
rect 5344 24252 5384 24258
rect 5344 24190 5384 24196
rect 5344 22738 5384 22744
rect 5344 22676 5384 22682
rect 5344 21224 5384 21230
rect 5344 21162 5384 21168
rect 5344 19710 5384 19716
rect 5344 19648 5384 19654
rect 5344 18196 5384 18202
rect 5344 18134 5384 18140
rect 5344 16682 5384 16688
rect 5344 16620 5384 16626
rect 5344 15168 5384 15174
rect 5344 15106 5384 15112
rect 5344 13654 5384 13660
rect 5344 13592 5384 13598
rect 5344 12140 5384 12146
rect 5344 12078 5384 12084
rect 5344 10626 5384 10632
rect 5344 10564 5384 10570
rect 5344 9112 5384 9118
rect 5344 9050 5384 9056
rect 5344 7598 5384 7604
rect 5344 7536 5384 7542
rect 5344 6084 5384 6090
rect 5344 6022 5384 6028
rect 5344 4570 5384 4576
rect 5344 4508 5384 4514
rect 5344 3056 5384 3062
rect 5344 2994 5384 3000
rect 5344 1542 5384 1548
rect 5344 1480 5384 1486
rect 5344 28 5384 34
rect 5344 -34 5384 -28
<< via2 >>
rect 2534 30090 2590 30092
rect 2534 30038 2536 30090
rect 2536 30038 2588 30090
rect 2588 30038 2590 30090
rect 2534 30036 2590 30038
rect 2534 28466 2590 28468
rect 2534 28414 2536 28466
rect 2536 28414 2588 28466
rect 2588 28414 2590 28466
rect 2534 28412 2590 28414
rect 2534 27010 2590 27012
rect 2534 26958 2536 27010
rect 2536 26958 2588 27010
rect 2588 26958 2590 27010
rect 2534 26956 2590 26958
rect 2534 25386 2590 25388
rect 2534 25334 2536 25386
rect 2536 25334 2588 25386
rect 2588 25334 2590 25386
rect 2534 25332 2590 25334
rect 2534 23930 2590 23932
rect 2534 23878 2536 23930
rect 2536 23878 2588 23930
rect 2588 23878 2590 23930
rect 2534 23876 2590 23878
rect 2534 22306 2590 22308
rect 2534 22254 2536 22306
rect 2536 22254 2588 22306
rect 2588 22254 2590 22306
rect 2534 22252 2590 22254
rect 2534 20850 2590 20852
rect 2534 20798 2536 20850
rect 2536 20798 2588 20850
rect 2588 20798 2590 20850
rect 2534 20796 2590 20798
rect 2534 19226 2590 19228
rect 2534 19174 2536 19226
rect 2536 19174 2588 19226
rect 2588 19174 2590 19226
rect 2534 19172 2590 19174
rect 2534 14694 2590 14696
rect 2534 14642 2536 14694
rect 2536 14642 2588 14694
rect 2588 14642 2590 14694
rect 2534 14640 2590 14642
rect 2534 13070 2590 13072
rect 2534 13018 2536 13070
rect 2536 13018 2588 13070
rect 2588 13018 2590 13070
rect 2534 13016 2590 13018
rect 2534 11614 2590 11616
rect 2534 11562 2536 11614
rect 2536 11562 2588 11614
rect 2588 11562 2590 11614
rect 2534 11560 2590 11562
rect 2534 9990 2590 9992
rect 2534 9938 2536 9990
rect 2536 9938 2588 9990
rect 2588 9938 2590 9990
rect 2534 9936 2590 9938
rect 2534 5458 2590 5460
rect 2534 5406 2536 5458
rect 2536 5406 2588 5458
rect 2588 5406 2590 5458
rect 2534 5404 2590 5406
rect 5336 48474 5392 48476
rect 5336 48422 5338 48474
rect 5338 48422 5390 48474
rect 5390 48422 5392 48474
rect 5336 48420 5392 48422
rect 5336 46960 5392 46962
rect 5336 46908 5338 46960
rect 5338 46908 5390 46960
rect 5390 46908 5392 46960
rect 5336 46906 5392 46908
rect 5336 45446 5392 45448
rect 5336 45394 5338 45446
rect 5338 45394 5390 45446
rect 5390 45394 5392 45446
rect 5336 45392 5392 45394
rect 5336 43932 5392 43934
rect 5336 43880 5338 43932
rect 5338 43880 5390 43932
rect 5390 43880 5392 43932
rect 5336 43878 5392 43880
rect 5336 42418 5392 42420
rect 5336 42366 5338 42418
rect 5338 42366 5390 42418
rect 5390 42366 5392 42418
rect 5336 42364 5392 42366
rect 5336 40904 5392 40906
rect 5336 40852 5338 40904
rect 5338 40852 5390 40904
rect 5390 40852 5392 40904
rect 5336 40850 5392 40852
rect 5336 39390 5392 39392
rect 5336 39338 5338 39390
rect 5338 39338 5390 39390
rect 5390 39338 5392 39390
rect 5336 39336 5392 39338
rect 5336 37876 5392 37878
rect 5336 37824 5338 37876
rect 5338 37824 5390 37876
rect 5390 37824 5392 37876
rect 5336 37822 5392 37824
rect 5336 36362 5392 36364
rect 5336 36310 5338 36362
rect 5338 36310 5390 36362
rect 5390 36310 5392 36362
rect 5336 36308 5392 36310
rect 5336 34848 5392 34850
rect 5336 34796 5338 34848
rect 5338 34796 5390 34848
rect 5390 34796 5392 34848
rect 5336 34794 5392 34796
rect 5336 33334 5392 33336
rect 5336 33282 5338 33334
rect 5338 33282 5390 33334
rect 5390 33282 5392 33334
rect 5336 33280 5392 33282
rect 5336 31820 5392 31822
rect 5336 31768 5338 31820
rect 5338 31768 5390 31820
rect 5390 31768 5392 31820
rect 5336 31766 5392 31768
rect 5336 30306 5392 30308
rect 5336 30254 5338 30306
rect 5338 30254 5390 30306
rect 5390 30254 5392 30306
rect 5336 30252 5392 30254
rect 3774 29224 3830 29280
rect 3706 27684 3762 27740
rect 3638 26144 3694 26200
rect 3570 24604 3626 24660
rect 3502 23064 3558 23120
rect 3434 22111 3490 22167
rect 3366 19984 3422 20040
rect 3298 18444 3354 18500
rect 3230 13828 3286 13884
rect 3162 12288 3218 12344
rect 3094 10748 3150 10804
rect 3026 9208 3082 9264
rect 2534 3834 2590 3836
rect 2534 3782 2536 3834
rect 2536 3782 2588 3834
rect 2588 3782 2590 3834
rect 2534 3780 2590 3782
rect 2534 2378 2590 2380
rect 2534 2326 2536 2378
rect 2536 2326 2588 2378
rect 2588 2326 2590 2378
rect 2534 2324 2590 2326
rect 2958 4592 3014 4648
rect 2890 3052 2946 3108
rect 2822 1512 2878 1568
rect 2534 754 2590 756
rect 2534 702 2536 754
rect 2536 702 2588 754
rect 2588 702 2590 754
rect 2534 700 2590 702
rect 2754 -28 2810 28
rect 5336 28792 5392 28794
rect 5336 28740 5338 28792
rect 5338 28740 5390 28792
rect 5390 28740 5392 28792
rect 5336 28738 5392 28740
rect 5336 27278 5392 27280
rect 5336 27226 5338 27278
rect 5338 27226 5390 27278
rect 5390 27226 5392 27278
rect 5336 27224 5392 27226
rect 5336 25764 5392 25766
rect 5336 25712 5338 25764
rect 5338 25712 5390 25764
rect 5390 25712 5392 25764
rect 5336 25710 5392 25712
rect 5336 24250 5392 24252
rect 5336 24198 5338 24250
rect 5338 24198 5390 24250
rect 5390 24198 5392 24250
rect 5336 24196 5392 24198
rect 5336 22736 5392 22738
rect 5336 22684 5338 22736
rect 5338 22684 5390 22736
rect 5390 22684 5392 22736
rect 5336 22682 5392 22684
rect 5336 21222 5392 21224
rect 5336 21170 5338 21222
rect 5338 21170 5390 21222
rect 5390 21170 5392 21222
rect 5336 21168 5392 21170
rect 5336 19708 5392 19710
rect 5336 19656 5338 19708
rect 5338 19656 5390 19708
rect 5390 19656 5392 19708
rect 5336 19654 5392 19656
rect 5336 18194 5392 18196
rect 5336 18142 5338 18194
rect 5338 18142 5390 18194
rect 5390 18142 5392 18194
rect 5336 18140 5392 18142
rect 5336 16680 5392 16682
rect 5336 16628 5338 16680
rect 5338 16628 5390 16680
rect 5390 16628 5392 16680
rect 5336 16626 5392 16628
rect 5336 15166 5392 15168
rect 5336 15114 5338 15166
rect 5338 15114 5390 15166
rect 5390 15114 5392 15166
rect 5336 15112 5392 15114
rect 5336 13652 5392 13654
rect 5336 13600 5338 13652
rect 5338 13600 5390 13652
rect 5390 13600 5392 13652
rect 5336 13598 5392 13600
rect 5336 12138 5392 12140
rect 5336 12086 5338 12138
rect 5338 12086 5390 12138
rect 5390 12086 5392 12138
rect 5336 12084 5392 12086
rect 5336 10624 5392 10626
rect 5336 10572 5338 10624
rect 5338 10572 5390 10624
rect 5390 10572 5392 10624
rect 5336 10570 5392 10572
rect 5336 9110 5392 9112
rect 5336 9058 5338 9110
rect 5338 9058 5390 9110
rect 5390 9058 5392 9110
rect 5336 9056 5392 9058
rect 5336 7596 5392 7598
rect 5336 7544 5338 7596
rect 5338 7544 5390 7596
rect 5390 7544 5392 7596
rect 5336 7542 5392 7544
rect 5336 6082 5392 6084
rect 5336 6030 5338 6082
rect 5338 6030 5390 6082
rect 5390 6030 5392 6082
rect 5336 6028 5392 6030
rect 5336 4568 5392 4570
rect 5336 4516 5338 4568
rect 5338 4516 5390 4568
rect 5390 4516 5392 4568
rect 5336 4514 5392 4516
rect 5336 3054 5392 3056
rect 5336 3002 5338 3054
rect 5338 3002 5390 3054
rect 5390 3002 5392 3054
rect 5336 3000 5392 3002
rect 5336 1540 5392 1542
rect 5336 1488 5338 1540
rect 5338 1488 5390 1540
rect 5390 1488 5392 1540
rect 5336 1486 5392 1488
rect 5336 26 5392 28
rect 5336 -26 5338 26
rect 5338 -26 5390 26
rect 5390 -26 5392 26
rect 5336 -28 5392 -26
<< metal3 >>
rect 5298 48476 5430 48481
rect 5298 48420 5336 48476
rect 5392 48420 5430 48476
rect 5298 48415 5430 48420
rect 5298 46962 5430 46967
rect 5298 46906 5336 46962
rect 5392 46906 5430 46962
rect 5298 46901 5430 46906
rect 5298 45448 5430 45453
rect 5298 45392 5336 45448
rect 5392 45392 5430 45448
rect 5298 45387 5430 45392
rect 5298 43934 5430 43939
rect 5298 43878 5336 43934
rect 5392 43878 5430 43934
rect 5298 43873 5430 43878
rect 5298 42420 5430 42425
rect 5298 42364 5336 42420
rect 5392 42364 5430 42420
rect 5298 42359 5430 42364
rect 5298 40906 5430 40911
rect 5298 40850 5336 40906
rect 5392 40850 5430 40906
rect 5298 40845 5430 40850
rect 5298 39392 5430 39397
rect 5298 39336 5336 39392
rect 5392 39336 5430 39392
rect 5298 39331 5430 39336
rect 5298 37878 5430 37883
rect 5298 37822 5336 37878
rect 5392 37822 5430 37878
rect 5298 37817 5430 37822
rect 5298 36364 5430 36369
rect 5298 36308 5336 36364
rect 5392 36308 5430 36364
rect 5298 36303 5430 36308
rect 5298 34850 5430 34855
rect 5298 34794 5336 34850
rect 5392 34794 5430 34850
rect 5298 34789 5430 34794
rect 5298 33336 5430 33341
rect 5298 33280 5336 33336
rect 5392 33280 5430 33336
rect 5298 33275 5430 33280
rect 5298 31822 5430 31827
rect 5298 31766 5336 31822
rect 5392 31766 5430 31822
rect 5298 31761 5430 31766
rect 751 30759 883 30825
rect 1646 30759 1778 30825
rect 5298 30308 5430 30313
rect 5298 30252 5336 30308
rect 5392 30252 5430 30308
rect 5298 30247 5430 30252
rect 2496 30092 2628 30097
rect 2496 30036 2534 30092
rect 2590 30036 2628 30092
rect 2496 30031 2628 30036
rect 751 29219 883 29285
rect 1646 29219 1778 29285
rect 2532 29282 2592 30031
rect 3736 29282 3868 29285
rect 2532 29280 3868 29282
rect 2532 29224 3774 29280
rect 3830 29224 3868 29280
rect 2532 29222 3868 29224
rect 3736 29219 3868 29222
rect 5298 28794 5430 28799
rect 5298 28738 5336 28794
rect 5392 28738 5430 28794
rect 5298 28733 5430 28738
rect 2496 28468 2628 28473
rect 2496 28412 2534 28468
rect 2590 28412 2628 28468
rect 2496 28407 2628 28412
rect 751 27679 883 27745
rect 1646 27679 1778 27745
rect 2532 27742 2592 28407
rect 3668 27742 3800 27745
rect 2532 27740 3800 27742
rect 2532 27684 3706 27740
rect 3762 27684 3800 27740
rect 2532 27682 3800 27684
rect 3668 27679 3800 27682
rect 5298 27280 5430 27285
rect 5298 27224 5336 27280
rect 5392 27224 5430 27280
rect 5298 27219 5430 27224
rect 2496 27012 2628 27017
rect 2496 26956 2534 27012
rect 2590 26956 2628 27012
rect 2496 26951 2628 26956
rect 751 26139 883 26205
rect 1646 26139 1778 26205
rect 2532 26202 2592 26951
rect 3600 26202 3732 26205
rect 2532 26200 3732 26202
rect 2532 26144 3638 26200
rect 3694 26144 3732 26200
rect 2532 26142 3732 26144
rect 3600 26139 3732 26142
rect 5298 25766 5430 25771
rect 5298 25710 5336 25766
rect 5392 25710 5430 25766
rect 5298 25705 5430 25710
rect 2496 25388 2628 25393
rect 2496 25332 2534 25388
rect 2590 25332 2628 25388
rect 2496 25327 2628 25332
rect 751 24599 883 24665
rect 1646 24599 1778 24665
rect 2532 24662 2592 25327
rect 3532 24662 3664 24665
rect 2532 24660 3664 24662
rect 2532 24604 3570 24660
rect 3626 24604 3664 24660
rect 2532 24602 3664 24604
rect 3532 24599 3664 24602
rect 5298 24252 5430 24257
rect 5298 24196 5336 24252
rect 5392 24196 5430 24252
rect 5298 24191 5430 24196
rect 2496 23932 2628 23937
rect 2496 23876 2534 23932
rect 2590 23876 2628 23932
rect 2496 23871 2628 23876
rect 751 23059 883 23125
rect 1646 23059 1778 23125
rect 2532 23122 2592 23871
rect 3464 23122 3596 23125
rect 2532 23120 3596 23122
rect 2532 23064 3502 23120
rect 3558 23064 3596 23120
rect 2532 23062 3596 23064
rect 3464 23059 3596 23062
rect 5298 22738 5430 22743
rect 5298 22682 5336 22738
rect 5392 22682 5430 22738
rect 5298 22677 5430 22682
rect 2496 22308 2628 22313
rect 2496 22252 2534 22308
rect 2590 22252 2628 22308
rect 2496 22247 2628 22252
rect 2532 22169 2592 22247
rect 3396 22169 3528 22172
rect 2532 22167 3528 22169
rect 2532 22111 3434 22167
rect 3490 22111 3528 22167
rect 2532 22109 3528 22111
rect 3396 22106 3528 22109
rect 751 21519 883 21585
rect 1646 21519 1778 21585
rect 5298 21224 5430 21229
rect 5298 21168 5336 21224
rect 5392 21168 5430 21224
rect 5298 21163 5430 21168
rect 2496 20852 2628 20857
rect 2496 20796 2534 20852
rect 2590 20796 2628 20852
rect 2496 20791 2628 20796
rect 751 19979 883 20045
rect 1646 19979 1778 20045
rect 2532 20042 2592 20791
rect 3328 20042 3460 20045
rect 2532 20040 3460 20042
rect 2532 19984 3366 20040
rect 3422 19984 3460 20040
rect 2532 19982 3460 19984
rect 3328 19979 3460 19982
rect 5298 19710 5430 19715
rect 5298 19654 5336 19710
rect 5392 19654 5430 19710
rect 5298 19649 5430 19654
rect 2496 19228 2628 19233
rect 2496 19172 2534 19228
rect 2590 19172 2628 19228
rect 2496 19167 2628 19172
rect 751 18439 883 18505
rect 1646 18439 1778 18505
rect 2532 18502 2592 19167
rect 3260 18502 3392 18505
rect 2532 18500 3392 18502
rect 2532 18444 3298 18500
rect 3354 18444 3392 18500
rect 2532 18442 3392 18444
rect 3260 18439 3392 18442
rect 5298 18196 5430 18201
rect 5298 18140 5336 18196
rect 5392 18140 5430 18196
rect 5298 18135 5430 18140
rect 5298 16682 5430 16687
rect 5298 16626 5336 16682
rect 5392 16626 5430 16682
rect 5298 16621 5430 16626
rect 1045 15363 1177 15429
rect 1804 15363 1936 15429
rect 5298 15168 5430 15173
rect 5298 15112 5336 15168
rect 5392 15112 5430 15168
rect 5298 15107 5430 15112
rect 2496 14696 2628 14701
rect 2496 14640 2534 14696
rect 2590 14640 2628 14696
rect 2496 14635 2628 14640
rect 1045 13823 1177 13889
rect 1804 13823 1936 13889
rect 2532 13886 2592 14635
rect 3192 13886 3324 13889
rect 2532 13884 3324 13886
rect 2532 13828 3230 13884
rect 3286 13828 3324 13884
rect 2532 13826 3324 13828
rect 3192 13823 3324 13826
rect 5298 13654 5430 13659
rect 5298 13598 5336 13654
rect 5392 13598 5430 13654
rect 5298 13593 5430 13598
rect 2496 13072 2628 13077
rect 2496 13016 2534 13072
rect 2590 13016 2628 13072
rect 2496 13011 2628 13016
rect 1045 12283 1177 12349
rect 1804 12283 1936 12349
rect 2532 12346 2592 13011
rect 3124 12346 3256 12349
rect 2532 12344 3256 12346
rect 2532 12288 3162 12344
rect 3218 12288 3256 12344
rect 2532 12286 3256 12288
rect 3124 12283 3256 12286
rect 5298 12140 5430 12145
rect 5298 12084 5336 12140
rect 5392 12084 5430 12140
rect 5298 12079 5430 12084
rect 2496 11616 2628 11621
rect 2496 11560 2534 11616
rect 2590 11560 2628 11616
rect 2496 11555 2628 11560
rect 1045 10743 1177 10809
rect 1804 10743 1936 10809
rect 2532 10806 2592 11555
rect 3056 10806 3188 10809
rect 2532 10804 3188 10806
rect 2532 10748 3094 10804
rect 3150 10748 3188 10804
rect 2532 10746 3188 10748
rect 3056 10743 3188 10746
rect 5298 10626 5430 10631
rect 5298 10570 5336 10626
rect 5392 10570 5430 10626
rect 5298 10565 5430 10570
rect 2496 9992 2628 9997
rect 2496 9936 2534 9992
rect 2590 9936 2628 9992
rect 2496 9931 2628 9936
rect 1045 9203 1177 9269
rect 1804 9203 1936 9269
rect 2532 9266 2592 9931
rect 2988 9266 3120 9269
rect 2532 9264 3120 9266
rect 2532 9208 3026 9264
rect 3082 9208 3120 9264
rect 2532 9206 3120 9208
rect 2988 9203 3120 9206
rect 5298 9112 5430 9117
rect 5298 9056 5336 9112
rect 5392 9056 5430 9112
rect 5298 9051 5430 9056
rect 5298 7598 5430 7603
rect 5298 7542 5336 7598
rect 5392 7542 5430 7598
rect 5298 7537 5430 7542
rect 1045 6127 1177 6193
rect 1804 6127 1936 6193
rect 5298 6084 5430 6089
rect 5298 6028 5336 6084
rect 5392 6028 5430 6084
rect 5298 6023 5430 6028
rect 2496 5460 2628 5465
rect 2496 5404 2534 5460
rect 2590 5404 2628 5460
rect 2496 5399 2628 5404
rect 1045 4587 1177 4653
rect 1804 4587 1936 4653
rect 2532 4650 2592 5399
rect 2920 4650 3052 4653
rect 2532 4648 3052 4650
rect 2532 4592 2958 4648
rect 3014 4592 3052 4648
rect 2532 4590 3052 4592
rect 2920 4587 3052 4590
rect 5298 4570 5430 4575
rect 5298 4514 5336 4570
rect 5392 4514 5430 4570
rect 5298 4509 5430 4514
rect 2496 3836 2628 3841
rect 2496 3780 2534 3836
rect 2590 3780 2628 3836
rect 2496 3775 2628 3780
rect 1045 3047 1177 3113
rect 1804 3047 1936 3113
rect 2532 3110 2592 3775
rect 2852 3110 2984 3113
rect 2532 3108 2984 3110
rect 2532 3052 2890 3108
rect 2946 3052 2984 3108
rect 2532 3050 2984 3052
rect 2852 3047 2984 3050
rect 5298 3056 5430 3061
rect 5298 3000 5336 3056
rect 5392 3000 5430 3056
rect 5298 2995 5430 3000
rect 2496 2380 2628 2385
rect 2496 2324 2534 2380
rect 2590 2324 2628 2380
rect 2496 2319 2628 2324
rect 1045 1507 1177 1573
rect 1804 1507 1936 1573
rect 2532 1570 2592 2319
rect 2784 1570 2916 1573
rect 2532 1568 2916 1570
rect 2532 1512 2822 1568
rect 2878 1512 2916 1568
rect 2532 1510 2916 1512
rect 2784 1507 2916 1510
rect 5298 1542 5430 1547
rect 5298 1486 5336 1542
rect 5392 1486 5430 1542
rect 5298 1481 5430 1486
rect 2496 756 2628 761
rect 2496 700 2534 756
rect 2590 700 2628 756
rect 2496 695 2628 700
rect 1045 -33 1177 33
rect 1804 -33 1936 33
rect 2532 30 2592 695
rect 2716 30 2848 33
rect 2532 28 2848 30
rect 2532 -28 2754 28
rect 2810 -28 2848 28
rect 2532 -30 2848 -28
rect 2716 -33 2848 -30
rect 5298 28 5430 33
rect 5298 -28 5336 28
rect 5392 -28 5430 28
rect 5298 -33 5430 -28
use contact_18  contact_18_0
timestamp 1643678851
transform 1 0 5298 0 1 -33
box 0 0 1 1
use contact_17  contact_17_0
timestamp 1643678851
transform 1 0 5349 0 1 -15
box 0 0 1 1
use contact_18  contact_18_1
timestamp 1643678851
transform 1 0 5298 0 1 1481
box 0 0 1 1
use contact_17  contact_17_1
timestamp 1643678851
transform 1 0 5349 0 1 1499
box 0 0 1 1
use contact_18  contact_18_2
timestamp 1643678851
transform 1 0 5298 0 1 -33
box 0 0 1 1
use contact_17  contact_17_2
timestamp 1643678851
transform 1 0 5349 0 1 -15
box 0 0 1 1
use contact_18  contact_18_3
timestamp 1643678851
transform 1 0 5298 0 1 1481
box 0 0 1 1
use contact_17  contact_17_3
timestamp 1643678851
transform 1 0 5349 0 1 1499
box 0 0 1 1
use contact_18  contact_18_4
timestamp 1643678851
transform 1 0 5298 0 1 -33
box 0 0 1 1
use contact_17  contact_17_4
timestamp 1643678851
transform 1 0 5349 0 1 -15
box 0 0 1 1
use contact_18  contact_18_5
timestamp 1643678851
transform 1 0 5298 0 1 1481
box 0 0 1 1
use contact_17  contact_17_5
timestamp 1643678851
transform 1 0 5349 0 1 1499
box 0 0 1 1
use contact_18  contact_18_6
timestamp 1643678851
transform 1 0 5298 0 1 -33
box 0 0 1 1
use contact_17  contact_17_6
timestamp 1643678851
transform 1 0 5349 0 1 -15
box 0 0 1 1
use contact_18  contact_18_7
timestamp 1643678851
transform 1 0 5298 0 1 1481
box 0 0 1 1
use contact_17  contact_17_7
timestamp 1643678851
transform 1 0 5349 0 1 1499
box 0 0 1 1
use contact_18  contact_18_8
timestamp 1643678851
transform 1 0 5298 0 1 -33
box 0 0 1 1
use contact_17  contact_17_8
timestamp 1643678851
transform 1 0 5349 0 1 -15
box 0 0 1 1
use contact_18  contact_18_9
timestamp 1643678851
transform 1 0 5298 0 1 1481
box 0 0 1 1
use contact_17  contact_17_9
timestamp 1643678851
transform 1 0 5349 0 1 1499
box 0 0 1 1
use contact_18  contact_18_10
timestamp 1643678851
transform 1 0 5298 0 1 -33
box 0 0 1 1
use contact_17  contact_17_10
timestamp 1643678851
transform 1 0 5349 0 1 -15
box 0 0 1 1
use contact_18  contact_18_11
timestamp 1643678851
transform 1 0 5298 0 1 1481
box 0 0 1 1
use contact_17  contact_17_11
timestamp 1643678851
transform 1 0 5349 0 1 1499
box 0 0 1 1
use contact_18  contact_18_12
timestamp 1643678851
transform 1 0 5298 0 1 -33
box 0 0 1 1
use contact_17  contact_17_12
timestamp 1643678851
transform 1 0 5349 0 1 -15
box 0 0 1 1
use contact_18  contact_18_13
timestamp 1643678851
transform 1 0 5298 0 1 1481
box 0 0 1 1
use contact_17  contact_17_13
timestamp 1643678851
transform 1 0 5349 0 1 1499
box 0 0 1 1
use contact_18  contact_18_14
timestamp 1643678851
transform 1 0 5298 0 1 -33
box 0 0 1 1
use contact_17  contact_17_14
timestamp 1643678851
transform 1 0 5349 0 1 -15
box 0 0 1 1
use contact_18  contact_18_15
timestamp 1643678851
transform 1 0 5298 0 1 1481
box 0 0 1 1
use contact_17  contact_17_15
timestamp 1643678851
transform 1 0 5349 0 1 1499
box 0 0 1 1
use contact_18  contact_18_16
timestamp 1643678851
transform 1 0 5298 0 1 -33
box 0 0 1 1
use contact_17  contact_17_16
timestamp 1643678851
transform 1 0 5349 0 1 -15
box 0 0 1 1
use contact_18  contact_18_17
timestamp 1643678851
transform 1 0 5298 0 1 1481
box 0 0 1 1
use contact_17  contact_17_17
timestamp 1643678851
transform 1 0 5349 0 1 1499
box 0 0 1 1
use contact_18  contact_18_18
timestamp 1643678851
transform 1 0 5298 0 1 -33
box 0 0 1 1
use contact_17  contact_17_18
timestamp 1643678851
transform 1 0 5349 0 1 -15
box 0 0 1 1
use contact_18  contact_18_19
timestamp 1643678851
transform 1 0 5298 0 1 1481
box 0 0 1 1
use contact_17  contact_17_19
timestamp 1643678851
transform 1 0 5349 0 1 1499
box 0 0 1 1
use contact_18  contact_18_20
timestamp 1643678851
transform 1 0 5298 0 1 -33
box 0 0 1 1
use contact_17  contact_17_20
timestamp 1643678851
transform 1 0 5349 0 1 -15
box 0 0 1 1
use contact_18  contact_18_21
timestamp 1643678851
transform 1 0 5298 0 1 1481
box 0 0 1 1
use contact_17  contact_17_21
timestamp 1643678851
transform 1 0 5349 0 1 1499
box 0 0 1 1
use contact_18  contact_18_22
timestamp 1643678851
transform 1 0 5298 0 1 -33
box 0 0 1 1
use contact_17  contact_17_22
timestamp 1643678851
transform 1 0 5349 0 1 -15
box 0 0 1 1
use contact_18  contact_18_23
timestamp 1643678851
transform 1 0 5298 0 1 1481
box 0 0 1 1
use contact_17  contact_17_23
timestamp 1643678851
transform 1 0 5349 0 1 1499
box 0 0 1 1
use contact_18  contact_18_24
timestamp 1643678851
transform 1 0 5298 0 1 -33
box 0 0 1 1
use contact_17  contact_17_24
timestamp 1643678851
transform 1 0 5349 0 1 -15
box 0 0 1 1
use contact_18  contact_18_25
timestamp 1643678851
transform 1 0 5298 0 1 1481
box 0 0 1 1
use contact_17  contact_17_25
timestamp 1643678851
transform 1 0 5349 0 1 1499
box 0 0 1 1
use contact_18  contact_18_26
timestamp 1643678851
transform 1 0 5298 0 1 -33
box 0 0 1 1
use contact_17  contact_17_26
timestamp 1643678851
transform 1 0 5349 0 1 -15
box 0 0 1 1
use contact_18  contact_18_27
timestamp 1643678851
transform 1 0 5298 0 1 1481
box 0 0 1 1
use contact_17  contact_17_27
timestamp 1643678851
transform 1 0 5349 0 1 1499
box 0 0 1 1
use contact_18  contact_18_28
timestamp 1643678851
transform 1 0 5298 0 1 -33
box 0 0 1 1
use contact_17  contact_17_28
timestamp 1643678851
transform 1 0 5349 0 1 -15
box 0 0 1 1
use contact_18  contact_18_29
timestamp 1643678851
transform 1 0 5298 0 1 1481
box 0 0 1 1
use contact_17  contact_17_29
timestamp 1643678851
transform 1 0 5349 0 1 1499
box 0 0 1 1
use contact_18  contact_18_30
timestamp 1643678851
transform 1 0 5298 0 1 -33
box 0 0 1 1
use contact_17  contact_17_30
timestamp 1643678851
transform 1 0 5349 0 1 -15
box 0 0 1 1
use contact_18  contact_18_31
timestamp 1643678851
transform 1 0 5298 0 1 1481
box 0 0 1 1
use contact_17  contact_17_31
timestamp 1643678851
transform 1 0 5349 0 1 1499
box 0 0 1 1
use contact_18  contact_18_32
timestamp 1643678851
transform 1 0 5298 0 1 -33
box 0 0 1 1
use contact_17  contact_17_32
timestamp 1643678851
transform 1 0 5349 0 1 -15
box 0 0 1 1
use contact_18  contact_18_33
timestamp 1643678851
transform 1 0 5298 0 1 1481
box 0 0 1 1
use contact_17  contact_17_33
timestamp 1643678851
transform 1 0 5349 0 1 1499
box 0 0 1 1
use contact_18  contact_18_34
timestamp 1643678851
transform 1 0 5298 0 1 -33
box 0 0 1 1
use contact_17  contact_17_34
timestamp 1643678851
transform 1 0 5349 0 1 -15
box 0 0 1 1
use contact_18  contact_18_35
timestamp 1643678851
transform 1 0 5298 0 1 1481
box 0 0 1 1
use contact_17  contact_17_35
timestamp 1643678851
transform 1 0 5349 0 1 1499
box 0 0 1 1
use contact_18  contact_18_36
timestamp 1643678851
transform 1 0 5298 0 1 -33
box 0 0 1 1
use contact_17  contact_17_36
timestamp 1643678851
transform 1 0 5349 0 1 -15
box 0 0 1 1
use contact_18  contact_18_37
timestamp 1643678851
transform 1 0 5298 0 1 1481
box 0 0 1 1
use contact_17  contact_17_37
timestamp 1643678851
transform 1 0 5349 0 1 1499
box 0 0 1 1
use contact_18  contact_18_38
timestamp 1643678851
transform 1 0 5298 0 1 -33
box 0 0 1 1
use contact_17  contact_17_38
timestamp 1643678851
transform 1 0 5349 0 1 -15
box 0 0 1 1
use contact_18  contact_18_39
timestamp 1643678851
transform 1 0 5298 0 1 1481
box 0 0 1 1
use contact_17  contact_17_39
timestamp 1643678851
transform 1 0 5349 0 1 1499
box 0 0 1 1
use contact_18  contact_18_40
timestamp 1643678851
transform 1 0 5298 0 1 -33
box 0 0 1 1
use contact_17  contact_17_40
timestamp 1643678851
transform 1 0 5349 0 1 -15
box 0 0 1 1
use contact_18  contact_18_41
timestamp 1643678851
transform 1 0 5298 0 1 1481
box 0 0 1 1
use contact_17  contact_17_41
timestamp 1643678851
transform 1 0 5349 0 1 1499
box 0 0 1 1
use contact_18  contact_18_42
timestamp 1643678851
transform 1 0 5298 0 1 -33
box 0 0 1 1
use contact_17  contact_17_42
timestamp 1643678851
transform 1 0 5349 0 1 -15
box 0 0 1 1
use contact_18  contact_18_43
timestamp 1643678851
transform 1 0 5298 0 1 1481
box 0 0 1 1
use contact_17  contact_17_43
timestamp 1643678851
transform 1 0 5349 0 1 1499
box 0 0 1 1
use contact_18  contact_18_44
timestamp 1643678851
transform 1 0 5298 0 1 -33
box 0 0 1 1
use contact_17  contact_17_44
timestamp 1643678851
transform 1 0 5349 0 1 -15
box 0 0 1 1
use contact_18  contact_18_45
timestamp 1643678851
transform 1 0 5298 0 1 1481
box 0 0 1 1
use contact_17  contact_17_45
timestamp 1643678851
transform 1 0 5349 0 1 1499
box 0 0 1 1
use contact_18  contact_18_46
timestamp 1643678851
transform 1 0 5298 0 1 -33
box 0 0 1 1
use contact_17  contact_17_46
timestamp 1643678851
transform 1 0 5349 0 1 -15
box 0 0 1 1
use contact_18  contact_18_47
timestamp 1643678851
transform 1 0 5298 0 1 1481
box 0 0 1 1
use contact_17  contact_17_47
timestamp 1643678851
transform 1 0 5349 0 1 1499
box 0 0 1 1
use contact_18  contact_18_48
timestamp 1643678851
transform 1 0 5298 0 1 -33
box 0 0 1 1
use contact_17  contact_17_48
timestamp 1643678851
transform 1 0 5349 0 1 -15
box 0 0 1 1
use contact_18  contact_18_49
timestamp 1643678851
transform 1 0 5298 0 1 1481
box 0 0 1 1
use contact_17  contact_17_49
timestamp 1643678851
transform 1 0 5349 0 1 1499
box 0 0 1 1
use contact_18  contact_18_50
timestamp 1643678851
transform 1 0 5298 0 1 -33
box 0 0 1 1
use contact_17  contact_17_50
timestamp 1643678851
transform 1 0 5349 0 1 -15
box 0 0 1 1
use contact_18  contact_18_51
timestamp 1643678851
transform 1 0 5298 0 1 1481
box 0 0 1 1
use contact_17  contact_17_51
timestamp 1643678851
transform 1 0 5349 0 1 1499
box 0 0 1 1
use contact_18  contact_18_52
timestamp 1643678851
transform 1 0 5298 0 1 -33
box 0 0 1 1
use contact_17  contact_17_52
timestamp 1643678851
transform 1 0 5349 0 1 -15
box 0 0 1 1
use contact_18  contact_18_53
timestamp 1643678851
transform 1 0 5298 0 1 1481
box 0 0 1 1
use contact_17  contact_17_53
timestamp 1643678851
transform 1 0 5349 0 1 1499
box 0 0 1 1
use contact_18  contact_18_54
timestamp 1643678851
transform 1 0 5298 0 1 -33
box 0 0 1 1
use contact_17  contact_17_54
timestamp 1643678851
transform 1 0 5349 0 1 -15
box 0 0 1 1
use contact_18  contact_18_55
timestamp 1643678851
transform 1 0 5298 0 1 1481
box 0 0 1 1
use contact_17  contact_17_55
timestamp 1643678851
transform 1 0 5349 0 1 1499
box 0 0 1 1
use contact_18  contact_18_56
timestamp 1643678851
transform 1 0 5298 0 1 -33
box 0 0 1 1
use contact_17  contact_17_56
timestamp 1643678851
transform 1 0 5349 0 1 -15
box 0 0 1 1
use contact_18  contact_18_57
timestamp 1643678851
transform 1 0 5298 0 1 1481
box 0 0 1 1
use contact_17  contact_17_57
timestamp 1643678851
transform 1 0 5349 0 1 1499
box 0 0 1 1
use contact_18  contact_18_58
timestamp 1643678851
transform 1 0 5298 0 1 -33
box 0 0 1 1
use contact_17  contact_17_58
timestamp 1643678851
transform 1 0 5349 0 1 -15
box 0 0 1 1
use contact_18  contact_18_59
timestamp 1643678851
transform 1 0 5298 0 1 1481
box 0 0 1 1
use contact_17  contact_17_59
timestamp 1643678851
transform 1 0 5349 0 1 1499
box 0 0 1 1
use contact_18  contact_18_60
timestamp 1643678851
transform 1 0 5298 0 1 -33
box 0 0 1 1
use contact_17  contact_17_60
timestamp 1643678851
transform 1 0 5349 0 1 -15
box 0 0 1 1
use contact_18  contact_18_61
timestamp 1643678851
transform 1 0 5298 0 1 1481
box 0 0 1 1
use contact_17  contact_17_61
timestamp 1643678851
transform 1 0 5349 0 1 1499
box 0 0 1 1
use contact_18  contact_18_62
timestamp 1643678851
transform 1 0 5298 0 1 -33
box 0 0 1 1
use contact_17  contact_17_62
timestamp 1643678851
transform 1 0 5349 0 1 -15
box 0 0 1 1
use contact_18  contact_18_63
timestamp 1643678851
transform 1 0 5298 0 1 1481
box 0 0 1 1
use contact_17  contact_17_63
timestamp 1643678851
transform 1 0 5349 0 1 1499
box 0 0 1 1
use contact_18  contact_18_64
timestamp 1643678851
transform 1 0 5298 0 1 -33
box 0 0 1 1
use contact_17  contact_17_64
timestamp 1643678851
transform 1 0 5349 0 1 -15
box 0 0 1 1
use contact_18  contact_18_65
timestamp 1643678851
transform 1 0 5298 0 1 1481
box 0 0 1 1
use contact_17  contact_17_65
timestamp 1643678851
transform 1 0 5349 0 1 1499
box 0 0 1 1
use contact_18  contact_18_66
timestamp 1643678851
transform 1 0 5298 0 1 -33
box 0 0 1 1
use contact_17  contact_17_66
timestamp 1643678851
transform 1 0 5349 0 1 -15
box 0 0 1 1
use contact_18  contact_18_67
timestamp 1643678851
transform 1 0 5298 0 1 1481
box 0 0 1 1
use contact_17  contact_17_67
timestamp 1643678851
transform 1 0 5349 0 1 1499
box 0 0 1 1
use contact_18  contact_18_68
timestamp 1643678851
transform 1 0 5298 0 1 -33
box 0 0 1 1
use contact_17  contact_17_68
timestamp 1643678851
transform 1 0 5349 0 1 -15
box 0 0 1 1
use contact_18  contact_18_69
timestamp 1643678851
transform 1 0 5298 0 1 1481
box 0 0 1 1
use contact_17  contact_17_69
timestamp 1643678851
transform 1 0 5349 0 1 1499
box 0 0 1 1
use contact_18  contact_18_70
timestamp 1643678851
transform 1 0 5298 0 1 -33
box 0 0 1 1
use contact_17  contact_17_70
timestamp 1643678851
transform 1 0 5349 0 1 -15
box 0 0 1 1
use contact_18  contact_18_71
timestamp 1643678851
transform 1 0 5298 0 1 1481
box 0 0 1 1
use contact_17  contact_17_71
timestamp 1643678851
transform 1 0 5349 0 1 1499
box 0 0 1 1
use contact_18  contact_18_72
timestamp 1643678851
transform 1 0 5298 0 1 -33
box 0 0 1 1
use contact_17  contact_17_72
timestamp 1643678851
transform 1 0 5349 0 1 -15
box 0 0 1 1
use contact_18  contact_18_73
timestamp 1643678851
transform 1 0 5298 0 1 1481
box 0 0 1 1
use contact_17  contact_17_73
timestamp 1643678851
transform 1 0 5349 0 1 1499
box 0 0 1 1
use contact_18  contact_18_74
timestamp 1643678851
transform 1 0 5298 0 1 -33
box 0 0 1 1
use contact_17  contact_17_74
timestamp 1643678851
transform 1 0 5349 0 1 -15
box 0 0 1 1
use contact_18  contact_18_75
timestamp 1643678851
transform 1 0 5298 0 1 1481
box 0 0 1 1
use contact_17  contact_17_75
timestamp 1643678851
transform 1 0 5349 0 1 1499
box 0 0 1 1
use contact_18  contact_18_76
timestamp 1643678851
transform 1 0 5298 0 1 -33
box 0 0 1 1
use contact_17  contact_17_76
timestamp 1643678851
transform 1 0 5349 0 1 -15
box 0 0 1 1
use contact_18  contact_18_77
timestamp 1643678851
transform 1 0 5298 0 1 1481
box 0 0 1 1
use contact_17  contact_17_77
timestamp 1643678851
transform 1 0 5349 0 1 1499
box 0 0 1 1
use contact_18  contact_18_78
timestamp 1643678851
transform 1 0 5298 0 1 -33
box 0 0 1 1
use contact_17  contact_17_78
timestamp 1643678851
transform 1 0 5349 0 1 -15
box 0 0 1 1
use contact_18  contact_18_79
timestamp 1643678851
transform 1 0 5298 0 1 1481
box 0 0 1 1
use contact_17  contact_17_79
timestamp 1643678851
transform 1 0 5349 0 1 1499
box 0 0 1 1
use contact_18  contact_18_80
timestamp 1643678851
transform 1 0 5298 0 1 -33
box 0 0 1 1
use contact_17  contact_17_80
timestamp 1643678851
transform 1 0 5349 0 1 -15
box 0 0 1 1
use contact_18  contact_18_81
timestamp 1643678851
transform 1 0 5298 0 1 1481
box 0 0 1 1
use contact_17  contact_17_81
timestamp 1643678851
transform 1 0 5349 0 1 1499
box 0 0 1 1
use contact_18  contact_18_82
timestamp 1643678851
transform 1 0 5298 0 1 -33
box 0 0 1 1
use contact_17  contact_17_82
timestamp 1643678851
transform 1 0 5349 0 1 -15
box 0 0 1 1
use contact_18  contact_18_83
timestamp 1643678851
transform 1 0 5298 0 1 1481
box 0 0 1 1
use contact_17  contact_17_83
timestamp 1643678851
transform 1 0 5349 0 1 1499
box 0 0 1 1
use contact_18  contact_18_84
timestamp 1643678851
transform 1 0 5298 0 1 -33
box 0 0 1 1
use contact_17  contact_17_84
timestamp 1643678851
transform 1 0 5349 0 1 -15
box 0 0 1 1
use contact_18  contact_18_85
timestamp 1643678851
transform 1 0 5298 0 1 1481
box 0 0 1 1
use contact_17  contact_17_85
timestamp 1643678851
transform 1 0 5349 0 1 1499
box 0 0 1 1
use contact_18  contact_18_86
timestamp 1643678851
transform 1 0 5298 0 1 -33
box 0 0 1 1
use contact_17  contact_17_86
timestamp 1643678851
transform 1 0 5349 0 1 -15
box 0 0 1 1
use contact_18  contact_18_87
timestamp 1643678851
transform 1 0 5298 0 1 1481
box 0 0 1 1
use contact_17  contact_17_87
timestamp 1643678851
transform 1 0 5349 0 1 1499
box 0 0 1 1
use contact_18  contact_18_88
timestamp 1643678851
transform 1 0 5298 0 1 -33
box 0 0 1 1
use contact_17  contact_17_88
timestamp 1643678851
transform 1 0 5349 0 1 -15
box 0 0 1 1
use contact_18  contact_18_89
timestamp 1643678851
transform 1 0 5298 0 1 1481
box 0 0 1 1
use contact_17  contact_17_89
timestamp 1643678851
transform 1 0 5349 0 1 1499
box 0 0 1 1
use contact_18  contact_18_90
timestamp 1643678851
transform 1 0 5298 0 1 -33
box 0 0 1 1
use contact_17  contact_17_90
timestamp 1643678851
transform 1 0 5349 0 1 -15
box 0 0 1 1
use contact_18  contact_18_91
timestamp 1643678851
transform 1 0 5298 0 1 1481
box 0 0 1 1
use contact_17  contact_17_91
timestamp 1643678851
transform 1 0 5349 0 1 1499
box 0 0 1 1
use contact_18  contact_18_92
timestamp 1643678851
transform 1 0 5298 0 1 -33
box 0 0 1 1
use contact_17  contact_17_92
timestamp 1643678851
transform 1 0 5349 0 1 -15
box 0 0 1 1
use contact_18  contact_18_93
timestamp 1643678851
transform 1 0 5298 0 1 1481
box 0 0 1 1
use contact_17  contact_17_93
timestamp 1643678851
transform 1 0 5349 0 1 1499
box 0 0 1 1
use contact_18  contact_18_94
timestamp 1643678851
transform 1 0 5298 0 1 -33
box 0 0 1 1
use contact_17  contact_17_94
timestamp 1643678851
transform 1 0 5349 0 1 -15
box 0 0 1 1
use contact_18  contact_18_95
timestamp 1643678851
transform 1 0 5298 0 1 1481
box 0 0 1 1
use contact_17  contact_17_95
timestamp 1643678851
transform 1 0 5349 0 1 1499
box 0 0 1 1
use contact_18  contact_18_96
timestamp 1643678851
transform 1 0 5298 0 1 -33
box 0 0 1 1
use contact_17  contact_17_96
timestamp 1643678851
transform 1 0 5349 0 1 -15
box 0 0 1 1
use contact_18  contact_18_97
timestamp 1643678851
transform 1 0 5298 0 1 1481
box 0 0 1 1
use contact_17  contact_17_97
timestamp 1643678851
transform 1 0 5349 0 1 1499
box 0 0 1 1
use contact_18  contact_18_98
timestamp 1643678851
transform 1 0 5298 0 1 -33
box 0 0 1 1
use contact_17  contact_17_98
timestamp 1643678851
transform 1 0 5349 0 1 -15
box 0 0 1 1
use contact_18  contact_18_99
timestamp 1643678851
transform 1 0 5298 0 1 1481
box 0 0 1 1
use contact_17  contact_17_99
timestamp 1643678851
transform 1 0 5349 0 1 1499
box 0 0 1 1
use contact_18  contact_18_100
timestamp 1643678851
transform 1 0 5298 0 1 -33
box 0 0 1 1
use contact_17  contact_17_100
timestamp 1643678851
transform 1 0 5349 0 1 -15
box 0 0 1 1
use contact_18  contact_18_101
timestamp 1643678851
transform 1 0 5298 0 1 1481
box 0 0 1 1
use contact_17  contact_17_101
timestamp 1643678851
transform 1 0 5349 0 1 1499
box 0 0 1 1
use contact_18  contact_18_102
timestamp 1643678851
transform 1 0 5298 0 1 -33
box 0 0 1 1
use contact_17  contact_17_102
timestamp 1643678851
transform 1 0 5349 0 1 -15
box 0 0 1 1
use contact_18  contact_18_103
timestamp 1643678851
transform 1 0 5298 0 1 1481
box 0 0 1 1
use contact_17  contact_17_103
timestamp 1643678851
transform 1 0 5349 0 1 1499
box 0 0 1 1
use contact_18  contact_18_104
timestamp 1643678851
transform 1 0 5298 0 1 -33
box 0 0 1 1
use contact_17  contact_17_104
timestamp 1643678851
transform 1 0 5349 0 1 -15
box 0 0 1 1
use contact_18  contact_18_105
timestamp 1643678851
transform 1 0 5298 0 1 1481
box 0 0 1 1
use contact_17  contact_17_105
timestamp 1643678851
transform 1 0 5349 0 1 1499
box 0 0 1 1
use contact_18  contact_18_106
timestamp 1643678851
transform 1 0 5298 0 1 -33
box 0 0 1 1
use contact_17  contact_17_106
timestamp 1643678851
transform 1 0 5349 0 1 -15
box 0 0 1 1
use contact_18  contact_18_107
timestamp 1643678851
transform 1 0 5298 0 1 1481
box 0 0 1 1
use contact_17  contact_17_107
timestamp 1643678851
transform 1 0 5349 0 1 1499
box 0 0 1 1
use contact_18  contact_18_108
timestamp 1643678851
transform 1 0 5298 0 1 -33
box 0 0 1 1
use contact_17  contact_17_108
timestamp 1643678851
transform 1 0 5349 0 1 -15
box 0 0 1 1
use contact_18  contact_18_109
timestamp 1643678851
transform 1 0 5298 0 1 1481
box 0 0 1 1
use contact_17  contact_17_109
timestamp 1643678851
transform 1 0 5349 0 1 1499
box 0 0 1 1
use contact_18  contact_18_110
timestamp 1643678851
transform 1 0 5298 0 1 -33
box 0 0 1 1
use contact_17  contact_17_110
timestamp 1643678851
transform 1 0 5349 0 1 -15
box 0 0 1 1
use contact_18  contact_18_111
timestamp 1643678851
transform 1 0 5298 0 1 1481
box 0 0 1 1
use contact_17  contact_17_111
timestamp 1643678851
transform 1 0 5349 0 1 1499
box 0 0 1 1
use contact_18  contact_18_112
timestamp 1643678851
transform 1 0 5298 0 1 -33
box 0 0 1 1
use contact_17  contact_17_112
timestamp 1643678851
transform 1 0 5349 0 1 -15
box 0 0 1 1
use contact_18  contact_18_113
timestamp 1643678851
transform 1 0 5298 0 1 1481
box 0 0 1 1
use contact_17  contact_17_113
timestamp 1643678851
transform 1 0 5349 0 1 1499
box 0 0 1 1
use contact_18  contact_18_114
timestamp 1643678851
transform 1 0 5298 0 1 -33
box 0 0 1 1
use contact_17  contact_17_114
timestamp 1643678851
transform 1 0 5349 0 1 -15
box 0 0 1 1
use contact_18  contact_18_115
timestamp 1643678851
transform 1 0 5298 0 1 1481
box 0 0 1 1
use contact_17  contact_17_115
timestamp 1643678851
transform 1 0 5349 0 1 1499
box 0 0 1 1
use contact_18  contact_18_116
timestamp 1643678851
transform 1 0 5298 0 1 -33
box 0 0 1 1
use contact_17  contact_17_116
timestamp 1643678851
transform 1 0 5349 0 1 -15
box 0 0 1 1
use contact_18  contact_18_117
timestamp 1643678851
transform 1 0 5298 0 1 1481
box 0 0 1 1
use contact_17  contact_17_117
timestamp 1643678851
transform 1 0 5349 0 1 1499
box 0 0 1 1
use contact_18  contact_18_118
timestamp 1643678851
transform 1 0 5298 0 1 -33
box 0 0 1 1
use contact_17  contact_17_118
timestamp 1643678851
transform 1 0 5349 0 1 -15
box 0 0 1 1
use contact_18  contact_18_119
timestamp 1643678851
transform 1 0 5298 0 1 1481
box 0 0 1 1
use contact_17  contact_17_119
timestamp 1643678851
transform 1 0 5349 0 1 1499
box 0 0 1 1
use contact_18  contact_18_120
timestamp 1643678851
transform 1 0 5298 0 1 -33
box 0 0 1 1
use contact_17  contact_17_120
timestamp 1643678851
transform 1 0 5349 0 1 -15
box 0 0 1 1
use contact_18  contact_18_121
timestamp 1643678851
transform 1 0 5298 0 1 1481
box 0 0 1 1
use contact_17  contact_17_121
timestamp 1643678851
transform 1 0 5349 0 1 1499
box 0 0 1 1
use contact_18  contact_18_122
timestamp 1643678851
transform 1 0 5298 0 1 -33
box 0 0 1 1
use contact_17  contact_17_122
timestamp 1643678851
transform 1 0 5349 0 1 -15
box 0 0 1 1
use contact_18  contact_18_123
timestamp 1643678851
transform 1 0 5298 0 1 1481
box 0 0 1 1
use contact_17  contact_17_123
timestamp 1643678851
transform 1 0 5349 0 1 1499
box 0 0 1 1
use contact_18  contact_18_124
timestamp 1643678851
transform 1 0 5298 0 1 -33
box 0 0 1 1
use contact_17  contact_17_124
timestamp 1643678851
transform 1 0 5349 0 1 -15
box 0 0 1 1
use contact_18  contact_18_125
timestamp 1643678851
transform 1 0 5298 0 1 1481
box 0 0 1 1
use contact_17  contact_17_125
timestamp 1643678851
transform 1 0 5349 0 1 1499
box 0 0 1 1
use contact_18  contact_18_126
timestamp 1643678851
transform 1 0 5298 0 1 -33
box 0 0 1 1
use contact_17  contact_17_126
timestamp 1643678851
transform 1 0 5349 0 1 -15
box 0 0 1 1
use contact_18  contact_18_127
timestamp 1643678851
transform 1 0 5298 0 1 1481
box 0 0 1 1
use contact_17  contact_17_127
timestamp 1643678851
transform 1 0 5349 0 1 1499
box 0 0 1 1
use contact_18  contact_18_128
timestamp 1643678851
transform 1 0 5298 0 1 48415
box 0 0 1 1
use contact_17  contact_17_128
timestamp 1643678851
transform 1 0 5349 0 1 48433
box 0 0 1 1
use contact_18  contact_18_129
timestamp 1643678851
transform 1 0 5298 0 1 46901
box 0 0 1 1
use contact_17  contact_17_129
timestamp 1643678851
transform 1 0 5349 0 1 46919
box 0 0 1 1
use contact_18  contact_18_130
timestamp 1643678851
transform 1 0 5298 0 1 45387
box 0 0 1 1
use contact_17  contact_17_130
timestamp 1643678851
transform 1 0 5349 0 1 45405
box 0 0 1 1
use contact_18  contact_18_131
timestamp 1643678851
transform 1 0 5298 0 1 46901
box 0 0 1 1
use contact_17  contact_17_131
timestamp 1643678851
transform 1 0 5349 0 1 46919
box 0 0 1 1
use contact_18  contact_18_132
timestamp 1643678851
transform 1 0 5298 0 1 45387
box 0 0 1 1
use contact_17  contact_17_132
timestamp 1643678851
transform 1 0 5349 0 1 45405
box 0 0 1 1
use contact_18  contact_18_133
timestamp 1643678851
transform 1 0 5298 0 1 43873
box 0 0 1 1
use contact_17  contact_17_133
timestamp 1643678851
transform 1 0 5349 0 1 43891
box 0 0 1 1
use contact_18  contact_18_134
timestamp 1643678851
transform 1 0 5298 0 1 42359
box 0 0 1 1
use contact_17  contact_17_134
timestamp 1643678851
transform 1 0 5349 0 1 42377
box 0 0 1 1
use contact_18  contact_18_135
timestamp 1643678851
transform 1 0 5298 0 1 43873
box 0 0 1 1
use contact_17  contact_17_135
timestamp 1643678851
transform 1 0 5349 0 1 43891
box 0 0 1 1
use contact_18  contact_18_136
timestamp 1643678851
transform 1 0 5298 0 1 42359
box 0 0 1 1
use contact_17  contact_17_136
timestamp 1643678851
transform 1 0 5349 0 1 42377
box 0 0 1 1
use contact_18  contact_18_137
timestamp 1643678851
transform 1 0 5298 0 1 40845
box 0 0 1 1
use contact_17  contact_17_137
timestamp 1643678851
transform 1 0 5349 0 1 40863
box 0 0 1 1
use contact_18  contact_18_138
timestamp 1643678851
transform 1 0 5298 0 1 39331
box 0 0 1 1
use contact_17  contact_17_138
timestamp 1643678851
transform 1 0 5349 0 1 39349
box 0 0 1 1
use contact_18  contact_18_139
timestamp 1643678851
transform 1 0 5298 0 1 40845
box 0 0 1 1
use contact_17  contact_17_139
timestamp 1643678851
transform 1 0 5349 0 1 40863
box 0 0 1 1
use contact_18  contact_18_140
timestamp 1643678851
transform 1 0 5298 0 1 39331
box 0 0 1 1
use contact_17  contact_17_140
timestamp 1643678851
transform 1 0 5349 0 1 39349
box 0 0 1 1
use contact_18  contact_18_141
timestamp 1643678851
transform 1 0 5298 0 1 37817
box 0 0 1 1
use contact_17  contact_17_141
timestamp 1643678851
transform 1 0 5349 0 1 37835
box 0 0 1 1
use contact_18  contact_18_142
timestamp 1643678851
transform 1 0 5298 0 1 36303
box 0 0 1 1
use contact_17  contact_17_142
timestamp 1643678851
transform 1 0 5349 0 1 36321
box 0 0 1 1
use contact_18  contact_18_143
timestamp 1643678851
transform 1 0 5298 0 1 37817
box 0 0 1 1
use contact_17  contact_17_143
timestamp 1643678851
transform 1 0 5349 0 1 37835
box 0 0 1 1
use contact_18  contact_18_144
timestamp 1643678851
transform 1 0 5298 0 1 36303
box 0 0 1 1
use contact_17  contact_17_144
timestamp 1643678851
transform 1 0 5349 0 1 36321
box 0 0 1 1
use contact_18  contact_18_145
timestamp 1643678851
transform 1 0 5298 0 1 34789
box 0 0 1 1
use contact_17  contact_17_145
timestamp 1643678851
transform 1 0 5349 0 1 34807
box 0 0 1 1
use contact_18  contact_18_146
timestamp 1643678851
transform 1 0 5298 0 1 33275
box 0 0 1 1
use contact_17  contact_17_146
timestamp 1643678851
transform 1 0 5349 0 1 33293
box 0 0 1 1
use contact_18  contact_18_147
timestamp 1643678851
transform 1 0 5298 0 1 34789
box 0 0 1 1
use contact_17  contact_17_147
timestamp 1643678851
transform 1 0 5349 0 1 34807
box 0 0 1 1
use contact_18  contact_18_148
timestamp 1643678851
transform 1 0 5298 0 1 33275
box 0 0 1 1
use contact_17  contact_17_148
timestamp 1643678851
transform 1 0 5349 0 1 33293
box 0 0 1 1
use contact_18  contact_18_149
timestamp 1643678851
transform 1 0 5298 0 1 31761
box 0 0 1 1
use contact_17  contact_17_149
timestamp 1643678851
transform 1 0 5349 0 1 31779
box 0 0 1 1
use contact_18  contact_18_150
timestamp 1643678851
transform 1 0 5298 0 1 30247
box 0 0 1 1
use contact_17  contact_17_150
timestamp 1643678851
transform 1 0 5349 0 1 30265
box 0 0 1 1
use contact_18  contact_18_151
timestamp 1643678851
transform 1 0 5298 0 1 31761
box 0 0 1 1
use contact_17  contact_17_151
timestamp 1643678851
transform 1 0 5349 0 1 31779
box 0 0 1 1
use contact_18  contact_18_152
timestamp 1643678851
transform 1 0 5298 0 1 30247
box 0 0 1 1
use contact_17  contact_17_152
timestamp 1643678851
transform 1 0 5349 0 1 30265
box 0 0 1 1
use contact_18  contact_18_153
timestamp 1643678851
transform 1 0 5298 0 1 28733
box 0 0 1 1
use contact_17  contact_17_153
timestamp 1643678851
transform 1 0 5349 0 1 28751
box 0 0 1 1
use contact_18  contact_18_154
timestamp 1643678851
transform 1 0 5298 0 1 27219
box 0 0 1 1
use contact_17  contact_17_154
timestamp 1643678851
transform 1 0 5349 0 1 27237
box 0 0 1 1
use contact_18  contact_18_155
timestamp 1643678851
transform 1 0 5298 0 1 28733
box 0 0 1 1
use contact_17  contact_17_155
timestamp 1643678851
transform 1 0 5349 0 1 28751
box 0 0 1 1
use contact_18  contact_18_156
timestamp 1643678851
transform 1 0 5298 0 1 27219
box 0 0 1 1
use contact_17  contact_17_156
timestamp 1643678851
transform 1 0 5349 0 1 27237
box 0 0 1 1
use contact_18  contact_18_157
timestamp 1643678851
transform 1 0 5298 0 1 25705
box 0 0 1 1
use contact_17  contact_17_157
timestamp 1643678851
transform 1 0 5349 0 1 25723
box 0 0 1 1
use contact_18  contact_18_158
timestamp 1643678851
transform 1 0 5298 0 1 24191
box 0 0 1 1
use contact_17  contact_17_158
timestamp 1643678851
transform 1 0 5349 0 1 24209
box 0 0 1 1
use contact_18  contact_18_159
timestamp 1643678851
transform 1 0 5298 0 1 25705
box 0 0 1 1
use contact_17  contact_17_159
timestamp 1643678851
transform 1 0 5349 0 1 25723
box 0 0 1 1
use contact_18  contact_18_160
timestamp 1643678851
transform 1 0 5298 0 1 24191
box 0 0 1 1
use contact_17  contact_17_160
timestamp 1643678851
transform 1 0 5349 0 1 24209
box 0 0 1 1
use contact_18  contact_18_161
timestamp 1643678851
transform 1 0 5298 0 1 22677
box 0 0 1 1
use contact_17  contact_17_161
timestamp 1643678851
transform 1 0 5349 0 1 22695
box 0 0 1 1
use contact_18  contact_18_162
timestamp 1643678851
transform 1 0 5298 0 1 21163
box 0 0 1 1
use contact_17  contact_17_162
timestamp 1643678851
transform 1 0 5349 0 1 21181
box 0 0 1 1
use contact_18  contact_18_163
timestamp 1643678851
transform 1 0 5298 0 1 22677
box 0 0 1 1
use contact_17  contact_17_163
timestamp 1643678851
transform 1 0 5349 0 1 22695
box 0 0 1 1
use contact_18  contact_18_164
timestamp 1643678851
transform 1 0 5298 0 1 21163
box 0 0 1 1
use contact_17  contact_17_164
timestamp 1643678851
transform 1 0 5349 0 1 21181
box 0 0 1 1
use contact_18  contact_18_165
timestamp 1643678851
transform 1 0 5298 0 1 19649
box 0 0 1 1
use contact_17  contact_17_165
timestamp 1643678851
transform 1 0 5349 0 1 19667
box 0 0 1 1
use contact_18  contact_18_166
timestamp 1643678851
transform 1 0 5298 0 1 18135
box 0 0 1 1
use contact_17  contact_17_166
timestamp 1643678851
transform 1 0 5349 0 1 18153
box 0 0 1 1
use contact_18  contact_18_167
timestamp 1643678851
transform 1 0 5298 0 1 19649
box 0 0 1 1
use contact_17  contact_17_167
timestamp 1643678851
transform 1 0 5349 0 1 19667
box 0 0 1 1
use contact_18  contact_18_168
timestamp 1643678851
transform 1 0 5298 0 1 18135
box 0 0 1 1
use contact_17  contact_17_168
timestamp 1643678851
transform 1 0 5349 0 1 18153
box 0 0 1 1
use contact_18  contact_18_169
timestamp 1643678851
transform 1 0 5298 0 1 16621
box 0 0 1 1
use contact_17  contact_17_169
timestamp 1643678851
transform 1 0 5349 0 1 16639
box 0 0 1 1
use contact_18  contact_18_170
timestamp 1643678851
transform 1 0 5298 0 1 15107
box 0 0 1 1
use contact_17  contact_17_170
timestamp 1643678851
transform 1 0 5349 0 1 15125
box 0 0 1 1
use contact_18  contact_18_171
timestamp 1643678851
transform 1 0 5298 0 1 16621
box 0 0 1 1
use contact_17  contact_17_171
timestamp 1643678851
transform 1 0 5349 0 1 16639
box 0 0 1 1
use contact_18  contact_18_172
timestamp 1643678851
transform 1 0 5298 0 1 15107
box 0 0 1 1
use contact_17  contact_17_172
timestamp 1643678851
transform 1 0 5349 0 1 15125
box 0 0 1 1
use contact_18  contact_18_173
timestamp 1643678851
transform 1 0 5298 0 1 13593
box 0 0 1 1
use contact_17  contact_17_173
timestamp 1643678851
transform 1 0 5349 0 1 13611
box 0 0 1 1
use contact_18  contact_18_174
timestamp 1643678851
transform 1 0 5298 0 1 12079
box 0 0 1 1
use contact_17  contact_17_174
timestamp 1643678851
transform 1 0 5349 0 1 12097
box 0 0 1 1
use contact_18  contact_18_175
timestamp 1643678851
transform 1 0 5298 0 1 13593
box 0 0 1 1
use contact_17  contact_17_175
timestamp 1643678851
transform 1 0 5349 0 1 13611
box 0 0 1 1
use contact_18  contact_18_176
timestamp 1643678851
transform 1 0 5298 0 1 12079
box 0 0 1 1
use contact_17  contact_17_176
timestamp 1643678851
transform 1 0 5349 0 1 12097
box 0 0 1 1
use contact_18  contact_18_177
timestamp 1643678851
transform 1 0 5298 0 1 10565
box 0 0 1 1
use contact_17  contact_17_177
timestamp 1643678851
transform 1 0 5349 0 1 10583
box 0 0 1 1
use contact_18  contact_18_178
timestamp 1643678851
transform 1 0 5298 0 1 9051
box 0 0 1 1
use contact_17  contact_17_178
timestamp 1643678851
transform 1 0 5349 0 1 9069
box 0 0 1 1
use contact_18  contact_18_179
timestamp 1643678851
transform 1 0 5298 0 1 10565
box 0 0 1 1
use contact_17  contact_17_179
timestamp 1643678851
transform 1 0 5349 0 1 10583
box 0 0 1 1
use contact_18  contact_18_180
timestamp 1643678851
transform 1 0 5298 0 1 9051
box 0 0 1 1
use contact_17  contact_17_180
timestamp 1643678851
transform 1 0 5349 0 1 9069
box 0 0 1 1
use contact_18  contact_18_181
timestamp 1643678851
transform 1 0 5298 0 1 7537
box 0 0 1 1
use contact_17  contact_17_181
timestamp 1643678851
transform 1 0 5349 0 1 7555
box 0 0 1 1
use contact_18  contact_18_182
timestamp 1643678851
transform 1 0 5298 0 1 6023
box 0 0 1 1
use contact_17  contact_17_182
timestamp 1643678851
transform 1 0 5349 0 1 6041
box 0 0 1 1
use contact_18  contact_18_183
timestamp 1643678851
transform 1 0 5298 0 1 7537
box 0 0 1 1
use contact_17  contact_17_183
timestamp 1643678851
transform 1 0 5349 0 1 7555
box 0 0 1 1
use contact_18  contact_18_184
timestamp 1643678851
transform 1 0 5298 0 1 6023
box 0 0 1 1
use contact_17  contact_17_184
timestamp 1643678851
transform 1 0 5349 0 1 6041
box 0 0 1 1
use contact_18  contact_18_185
timestamp 1643678851
transform 1 0 5298 0 1 4509
box 0 0 1 1
use contact_17  contact_17_185
timestamp 1643678851
transform 1 0 5349 0 1 4527
box 0 0 1 1
use contact_18  contact_18_186
timestamp 1643678851
transform 1 0 5298 0 1 2995
box 0 0 1 1
use contact_17  contact_17_186
timestamp 1643678851
transform 1 0 5349 0 1 3013
box 0 0 1 1
use contact_18  contact_18_187
timestamp 1643678851
transform 1 0 5298 0 1 4509
box 0 0 1 1
use contact_17  contact_17_187
timestamp 1643678851
transform 1 0 5349 0 1 4527
box 0 0 1 1
use contact_18  contact_18_188
timestamp 1643678851
transform 1 0 5298 0 1 2995
box 0 0 1 1
use contact_17  contact_17_188
timestamp 1643678851
transform 1 0 5349 0 1 3013
box 0 0 1 1
use contact_18  contact_18_189
timestamp 1643678851
transform 1 0 5298 0 1 1481
box 0 0 1 1
use contact_17  contact_17_189
timestamp 1643678851
transform 1 0 5349 0 1 1499
box 0 0 1 1
use contact_18  contact_18_190
timestamp 1643678851
transform 1 0 5298 0 1 -33
box 0 0 1 1
use contact_17  contact_17_190
timestamp 1643678851
transform 1 0 5349 0 1 -15
box 0 0 1 1
use contact_18  contact_18_191
timestamp 1643678851
transform 1 0 5298 0 1 1481
box 0 0 1 1
use contact_17  contact_17_191
timestamp 1643678851
transform 1 0 5349 0 1 1499
box 0 0 1 1
use contact_20  contact_20_0
timestamp 1643678851
transform 1 0 3736 0 1 29219
box 0 0 1 1
use contact_18  contact_18_192
timestamp 1643678851
transform 1 0 2496 0 1 30031
box 0 0 1 1
use contact_17  contact_17_192
timestamp 1643678851
transform 1 0 2547 0 1 30049
box 0 0 1 1
use contact_13  contact_13_0
timestamp 1643678851
transform 1 0 2533 0 1 30041
box 0 0 1 1
use contact_20  contact_20_1
timestamp 1643678851
transform 1 0 3668 0 1 27679
box 0 0 1 1
use contact_18  contact_18_193
timestamp 1643678851
transform 1 0 2496 0 1 28407
box 0 0 1 1
use contact_17  contact_17_193
timestamp 1643678851
transform 1 0 2547 0 1 28425
box 0 0 1 1
use contact_13  contact_13_1
timestamp 1643678851
transform 1 0 2533 0 1 28417
box 0 0 1 1
use contact_20  contact_20_2
timestamp 1643678851
transform 1 0 3600 0 1 26139
box 0 0 1 1
use contact_18  contact_18_194
timestamp 1643678851
transform 1 0 2496 0 1 26951
box 0 0 1 1
use contact_17  contact_17_194
timestamp 1643678851
transform 1 0 2547 0 1 26969
box 0 0 1 1
use contact_13  contact_13_2
timestamp 1643678851
transform 1 0 2533 0 1 26961
box 0 0 1 1
use contact_20  contact_20_3
timestamp 1643678851
transform 1 0 3532 0 1 24599
box 0 0 1 1
use contact_18  contact_18_195
timestamp 1643678851
transform 1 0 2496 0 1 25327
box 0 0 1 1
use contact_17  contact_17_195
timestamp 1643678851
transform 1 0 2547 0 1 25345
box 0 0 1 1
use contact_13  contact_13_3
timestamp 1643678851
transform 1 0 2533 0 1 25337
box 0 0 1 1
use contact_20  contact_20_4
timestamp 1643678851
transform 1 0 3464 0 1 23059
box 0 0 1 1
use contact_18  contact_18_196
timestamp 1643678851
transform 1 0 2496 0 1 23871
box 0 0 1 1
use contact_17  contact_17_196
timestamp 1643678851
transform 1 0 2547 0 1 23889
box 0 0 1 1
use contact_13  contact_13_4
timestamp 1643678851
transform 1 0 2533 0 1 23881
box 0 0 1 1
use contact_20  contact_20_5
timestamp 1643678851
transform 1 0 3396 0 1 22106
box 0 0 1 1
use contact_18  contact_18_197
timestamp 1643678851
transform 1 0 2496 0 1 22247
box 0 0 1 1
use contact_17  contact_17_197
timestamp 1643678851
transform 1 0 2547 0 1 22265
box 0 0 1 1
use contact_13  contact_13_5
timestamp 1643678851
transform 1 0 2533 0 1 22257
box 0 0 1 1
use contact_20  contact_20_6
timestamp 1643678851
transform 1 0 3328 0 1 19979
box 0 0 1 1
use contact_18  contact_18_198
timestamp 1643678851
transform 1 0 2496 0 1 20791
box 0 0 1 1
use contact_17  contact_17_198
timestamp 1643678851
transform 1 0 2547 0 1 20809
box 0 0 1 1
use contact_13  contact_13_6
timestamp 1643678851
transform 1 0 2533 0 1 20801
box 0 0 1 1
use contact_20  contact_20_7
timestamp 1643678851
transform 1 0 3260 0 1 18439
box 0 0 1 1
use contact_18  contact_18_199
timestamp 1643678851
transform 1 0 2496 0 1 19167
box 0 0 1 1
use contact_17  contact_17_199
timestamp 1643678851
transform 1 0 2547 0 1 19185
box 0 0 1 1
use contact_13  contact_13_7
timestamp 1643678851
transform 1 0 2533 0 1 19177
box 0 0 1 1
use contact_20  contact_20_8
timestamp 1643678851
transform 1 0 3192 0 1 13823
box 0 0 1 1
use contact_18  contact_18_200
timestamp 1643678851
transform 1 0 2496 0 1 14635
box 0 0 1 1
use contact_17  contact_17_200
timestamp 1643678851
transform 1 0 2547 0 1 14653
box 0 0 1 1
use contact_13  contact_13_8
timestamp 1643678851
transform 1 0 2533 0 1 14645
box 0 0 1 1
use contact_20  contact_20_9
timestamp 1643678851
transform 1 0 3124 0 1 12283
box 0 0 1 1
use contact_18  contact_18_201
timestamp 1643678851
transform 1 0 2496 0 1 13011
box 0 0 1 1
use contact_17  contact_17_201
timestamp 1643678851
transform 1 0 2547 0 1 13029
box 0 0 1 1
use contact_13  contact_13_9
timestamp 1643678851
transform 1 0 2533 0 1 13021
box 0 0 1 1
use contact_20  contact_20_10
timestamp 1643678851
transform 1 0 3056 0 1 10743
box 0 0 1 1
use contact_18  contact_18_202
timestamp 1643678851
transform 1 0 2496 0 1 11555
box 0 0 1 1
use contact_17  contact_17_202
timestamp 1643678851
transform 1 0 2547 0 1 11573
box 0 0 1 1
use contact_13  contact_13_10
timestamp 1643678851
transform 1 0 2533 0 1 11565
box 0 0 1 1
use contact_20  contact_20_11
timestamp 1643678851
transform 1 0 2988 0 1 9203
box 0 0 1 1
use contact_18  contact_18_203
timestamp 1643678851
transform 1 0 2496 0 1 9931
box 0 0 1 1
use contact_17  contact_17_203
timestamp 1643678851
transform 1 0 2547 0 1 9949
box 0 0 1 1
use contact_13  contact_13_11
timestamp 1643678851
transform 1 0 2533 0 1 9941
box 0 0 1 1
use contact_20  contact_20_12
timestamp 1643678851
transform 1 0 2920 0 1 4587
box 0 0 1 1
use contact_18  contact_18_204
timestamp 1643678851
transform 1 0 2496 0 1 5399
box 0 0 1 1
use contact_17  contact_17_204
timestamp 1643678851
transform 1 0 2547 0 1 5417
box 0 0 1 1
use contact_13  contact_13_12
timestamp 1643678851
transform 1 0 2533 0 1 5409
box 0 0 1 1
use contact_20  contact_20_13
timestamp 1643678851
transform 1 0 2852 0 1 3047
box 0 0 1 1
use contact_18  contact_18_205
timestamp 1643678851
transform 1 0 2496 0 1 3775
box 0 0 1 1
use contact_17  contact_17_205
timestamp 1643678851
transform 1 0 2547 0 1 3793
box 0 0 1 1
use contact_13  contact_13_13
timestamp 1643678851
transform 1 0 2533 0 1 3785
box 0 0 1 1
use contact_20  contact_20_14
timestamp 1643678851
transform 1 0 2784 0 1 1507
box 0 0 1 1
use contact_18  contact_18_206
timestamp 1643678851
transform 1 0 2496 0 1 2319
box 0 0 1 1
use contact_17  contact_17_206
timestamp 1643678851
transform 1 0 2547 0 1 2337
box 0 0 1 1
use contact_13  contact_13_14
timestamp 1643678851
transform 1 0 2533 0 1 2329
box 0 0 1 1
use contact_20  contact_20_15
timestamp 1643678851
transform 1 0 2716 0 1 -33
box 0 0 1 1
use contact_18  contact_18_207
timestamp 1643678851
transform 1 0 2496 0 1 695
box 0 0 1 1
use contact_17  contact_17_207
timestamp 1643678851
transform 1 0 2547 0 1 713
box 0 0 1 1
use contact_13  contact_13_15
timestamp 1643678851
transform 1 0 2533 0 1 705
box 0 0 1 1
use contact_14  contact_14_0
timestamp 1643678851
transform 1 0 3651 0 1 801
box 0 0 1 1
use contact_14  contact_14_1
timestamp 1643678851
transform 1 0 3243 0 1 857
box 0 0 1 1
use contact_14  contact_14_2
timestamp 1643678851
transform 1 0 2971 0 1 913
box 0 0 1 1
use contact_14  contact_14_3
timestamp 1643678851
transform 1 0 3651 0 1 47953
box 0 0 1 1
use contact_14  contact_14_4
timestamp 1643678851
transform 1 0 3243 0 1 47897
box 0 0 1 1
use contact_14  contact_14_5
timestamp 1643678851
transform 1 0 2903 0 1 47841
box 0 0 1 1
use contact_14  contact_14_6
timestamp 1643678851
transform 1 0 3651 0 1 47785
box 0 0 1 1
use contact_14  contact_14_7
timestamp 1643678851
transform 1 0 3243 0 1 47729
box 0 0 1 1
use contact_14  contact_14_8
timestamp 1643678851
transform 1 0 2835 0 1 47673
box 0 0 1 1
use contact_14  contact_14_9
timestamp 1643678851
transform 1 0 3651 0 1 47617
box 0 0 1 1
use contact_14  contact_14_10
timestamp 1643678851
transform 1 0 3243 0 1 47561
box 0 0 1 1
use contact_14  contact_14_11
timestamp 1643678851
transform 1 0 2767 0 1 47505
box 0 0 1 1
use contact_14  contact_14_12
timestamp 1643678851
transform 1 0 3651 0 1 45885
box 0 0 1 1
use contact_14  contact_14_13
timestamp 1643678851
transform 1 0 3175 0 1 45941
box 0 0 1 1
use contact_14  contact_14_14
timestamp 1643678851
transform 1 0 2971 0 1 45997
box 0 0 1 1
use contact_14  contact_14_15
timestamp 1643678851
transform 1 0 3651 0 1 46053
box 0 0 1 1
use contact_14  contact_14_16
timestamp 1643678851
transform 1 0 3175 0 1 46109
box 0 0 1 1
use contact_14  contact_14_17
timestamp 1643678851
transform 1 0 2903 0 1 46165
box 0 0 1 1
use contact_14  contact_14_18
timestamp 1643678851
transform 1 0 3651 0 1 46221
box 0 0 1 1
use contact_14  contact_14_19
timestamp 1643678851
transform 1 0 3175 0 1 46277
box 0 0 1 1
use contact_14  contact_14_20
timestamp 1643678851
transform 1 0 2835 0 1 46333
box 0 0 1 1
use contact_14  contact_14_21
timestamp 1643678851
transform 1 0 3651 0 1 44925
box 0 0 1 1
use contact_14  contact_14_22
timestamp 1643678851
transform 1 0 3175 0 1 44869
box 0 0 1 1
use contact_14  contact_14_23
timestamp 1643678851
transform 1 0 2767 0 1 44813
box 0 0 1 1
use contact_14  contact_14_24
timestamp 1643678851
transform 1 0 3651 0 1 44757
box 0 0 1 1
use contact_14  contact_14_25
timestamp 1643678851
transform 1 0 3107 0 1 44701
box 0 0 1 1
use contact_14  contact_14_26
timestamp 1643678851
transform 1 0 2971 0 1 44645
box 0 0 1 1
use contact_14  contact_14_27
timestamp 1643678851
transform 1 0 3651 0 1 44589
box 0 0 1 1
use contact_14  contact_14_28
timestamp 1643678851
transform 1 0 3107 0 1 44533
box 0 0 1 1
use contact_14  contact_14_29
timestamp 1643678851
transform 1 0 2903 0 1 44477
box 0 0 1 1
use contact_14  contact_14_30
timestamp 1643678851
transform 1 0 3651 0 1 42857
box 0 0 1 1
use contact_14  contact_14_31
timestamp 1643678851
transform 1 0 3107 0 1 42913
box 0 0 1 1
use contact_14  contact_14_32
timestamp 1643678851
transform 1 0 2835 0 1 42969
box 0 0 1 1
use contact_14  contact_14_33
timestamp 1643678851
transform 1 0 3651 0 1 43025
box 0 0 1 1
use contact_14  contact_14_34
timestamp 1643678851
transform 1 0 3107 0 1 43081
box 0 0 1 1
use contact_14  contact_14_35
timestamp 1643678851
transform 1 0 2767 0 1 43137
box 0 0 1 1
use contact_14  contact_14_36
timestamp 1643678851
transform 1 0 3651 0 1 43193
box 0 0 1 1
use contact_14  contact_14_37
timestamp 1643678851
transform 1 0 3039 0 1 43249
box 0 0 1 1
use contact_14  contact_14_38
timestamp 1643678851
transform 1 0 2971 0 1 43305
box 0 0 1 1
use contact_14  contact_14_39
timestamp 1643678851
transform 1 0 3651 0 1 41897
box 0 0 1 1
use contact_14  contact_14_40
timestamp 1643678851
transform 1 0 3039 0 1 41841
box 0 0 1 1
use contact_14  contact_14_41
timestamp 1643678851
transform 1 0 2903 0 1 41785
box 0 0 1 1
use contact_14  contact_14_42
timestamp 1643678851
transform 1 0 3651 0 1 41729
box 0 0 1 1
use contact_14  contact_14_43
timestamp 1643678851
transform 1 0 3039 0 1 41673
box 0 0 1 1
use contact_14  contact_14_44
timestamp 1643678851
transform 1 0 2835 0 1 41617
box 0 0 1 1
use contact_14  contact_14_45
timestamp 1643678851
transform 1 0 3651 0 1 41561
box 0 0 1 1
use contact_14  contact_14_46
timestamp 1643678851
transform 1 0 3039 0 1 41505
box 0 0 1 1
use contact_14  contact_14_47
timestamp 1643678851
transform 1 0 2767 0 1 41449
box 0 0 1 1
use contact_14  contact_14_48
timestamp 1643678851
transform 1 0 3583 0 1 39829
box 0 0 1 1
use contact_14  contact_14_49
timestamp 1643678851
transform 1 0 3243 0 1 39885
box 0 0 1 1
use contact_14  contact_14_50
timestamp 1643678851
transform 1 0 2971 0 1 39941
box 0 0 1 1
use contact_14  contact_14_51
timestamp 1643678851
transform 1 0 3583 0 1 39997
box 0 0 1 1
use contact_14  contact_14_52
timestamp 1643678851
transform 1 0 3243 0 1 40053
box 0 0 1 1
use contact_14  contact_14_53
timestamp 1643678851
transform 1 0 2903 0 1 40109
box 0 0 1 1
use contact_14  contact_14_54
timestamp 1643678851
transform 1 0 3583 0 1 40165
box 0 0 1 1
use contact_14  contact_14_55
timestamp 1643678851
transform 1 0 3243 0 1 40221
box 0 0 1 1
use contact_14  contact_14_56
timestamp 1643678851
transform 1 0 2835 0 1 40277
box 0 0 1 1
use contact_14  contact_14_57
timestamp 1643678851
transform 1 0 3583 0 1 38869
box 0 0 1 1
use contact_14  contact_14_58
timestamp 1643678851
transform 1 0 3243 0 1 38813
box 0 0 1 1
use contact_14  contact_14_59
timestamp 1643678851
transform 1 0 2767 0 1 38757
box 0 0 1 1
use contact_14  contact_14_60
timestamp 1643678851
transform 1 0 3583 0 1 38701
box 0 0 1 1
use contact_14  contact_14_61
timestamp 1643678851
transform 1 0 3175 0 1 38645
box 0 0 1 1
use contact_14  contact_14_62
timestamp 1643678851
transform 1 0 2971 0 1 38589
box 0 0 1 1
use contact_14  contact_14_63
timestamp 1643678851
transform 1 0 3583 0 1 38533
box 0 0 1 1
use contact_14  contact_14_64
timestamp 1643678851
transform 1 0 3175 0 1 38477
box 0 0 1 1
use contact_14  contact_14_65
timestamp 1643678851
transform 1 0 2903 0 1 38421
box 0 0 1 1
use contact_14  contact_14_66
timestamp 1643678851
transform 1 0 3583 0 1 36801
box 0 0 1 1
use contact_14  contact_14_67
timestamp 1643678851
transform 1 0 3175 0 1 36857
box 0 0 1 1
use contact_14  contact_14_68
timestamp 1643678851
transform 1 0 2835 0 1 36913
box 0 0 1 1
use contact_14  contact_14_69
timestamp 1643678851
transform 1 0 3583 0 1 36969
box 0 0 1 1
use contact_14  contact_14_70
timestamp 1643678851
transform 1 0 3175 0 1 37025
box 0 0 1 1
use contact_14  contact_14_71
timestamp 1643678851
transform 1 0 2767 0 1 37081
box 0 0 1 1
use contact_14  contact_14_72
timestamp 1643678851
transform 1 0 3583 0 1 37137
box 0 0 1 1
use contact_14  contact_14_73
timestamp 1643678851
transform 1 0 3107 0 1 37193
box 0 0 1 1
use contact_14  contact_14_74
timestamp 1643678851
transform 1 0 2971 0 1 37249
box 0 0 1 1
use contact_14  contact_14_75
timestamp 1643678851
transform 1 0 3583 0 1 35841
box 0 0 1 1
use contact_14  contact_14_76
timestamp 1643678851
transform 1 0 3107 0 1 35785
box 0 0 1 1
use contact_14  contact_14_77
timestamp 1643678851
transform 1 0 2903 0 1 35729
box 0 0 1 1
use contact_14  contact_14_78
timestamp 1643678851
transform 1 0 3583 0 1 35673
box 0 0 1 1
use contact_14  contact_14_79
timestamp 1643678851
transform 1 0 3107 0 1 35617
box 0 0 1 1
use contact_14  contact_14_80
timestamp 1643678851
transform 1 0 2835 0 1 35561
box 0 0 1 1
use contact_14  contact_14_81
timestamp 1643678851
transform 1 0 3583 0 1 35505
box 0 0 1 1
use contact_14  contact_14_82
timestamp 1643678851
transform 1 0 3107 0 1 35449
box 0 0 1 1
use contact_14  contact_14_83
timestamp 1643678851
transform 1 0 2767 0 1 35393
box 0 0 1 1
use contact_14  contact_14_84
timestamp 1643678851
transform 1 0 3583 0 1 33773
box 0 0 1 1
use contact_14  contact_14_85
timestamp 1643678851
transform 1 0 3039 0 1 33829
box 0 0 1 1
use contact_14  contact_14_86
timestamp 1643678851
transform 1 0 2971 0 1 33885
box 0 0 1 1
use contact_14  contact_14_87
timestamp 1643678851
transform 1 0 3583 0 1 33941
box 0 0 1 1
use contact_14  contact_14_88
timestamp 1643678851
transform 1 0 3039 0 1 33997
box 0 0 1 1
use contact_14  contact_14_89
timestamp 1643678851
transform 1 0 2903 0 1 34053
box 0 0 1 1
use contact_14  contact_14_90
timestamp 1643678851
transform 1 0 3583 0 1 34109
box 0 0 1 1
use contact_14  contact_14_91
timestamp 1643678851
transform 1 0 3039 0 1 34165
box 0 0 1 1
use contact_14  contact_14_92
timestamp 1643678851
transform 1 0 2835 0 1 34221
box 0 0 1 1
use contact_14  contact_14_93
timestamp 1643678851
transform 1 0 3583 0 1 32813
box 0 0 1 1
use contact_14  contact_14_94
timestamp 1643678851
transform 1 0 3039 0 1 32757
box 0 0 1 1
use contact_14  contact_14_95
timestamp 1643678851
transform 1 0 2767 0 1 32701
box 0 0 1 1
use contact_14  contact_14_96
timestamp 1643678851
transform 1 0 3515 0 1 32645
box 0 0 1 1
use contact_14  contact_14_97
timestamp 1643678851
transform 1 0 3243 0 1 32589
box 0 0 1 1
use contact_14  contact_14_98
timestamp 1643678851
transform 1 0 2971 0 1 32533
box 0 0 1 1
use contact_14  contact_14_99
timestamp 1643678851
transform 1 0 3515 0 1 32477
box 0 0 1 1
use contact_14  contact_14_100
timestamp 1643678851
transform 1 0 3243 0 1 32421
box 0 0 1 1
use contact_14  contact_14_101
timestamp 1643678851
transform 1 0 2903 0 1 32365
box 0 0 1 1
use contact_14  contact_14_102
timestamp 1643678851
transform 1 0 3515 0 1 30745
box 0 0 1 1
use contact_14  contact_14_103
timestamp 1643678851
transform 1 0 3243 0 1 30801
box 0 0 1 1
use contact_14  contact_14_104
timestamp 1643678851
transform 1 0 2835 0 1 30857
box 0 0 1 1
use contact_14  contact_14_105
timestamp 1643678851
transform 1 0 3515 0 1 30913
box 0 0 1 1
use contact_14  contact_14_106
timestamp 1643678851
transform 1 0 3243 0 1 30969
box 0 0 1 1
use contact_14  contact_14_107
timestamp 1643678851
transform 1 0 2767 0 1 31025
box 0 0 1 1
use contact_14  contact_14_108
timestamp 1643678851
transform 1 0 3515 0 1 31081
box 0 0 1 1
use contact_14  contact_14_109
timestamp 1643678851
transform 1 0 3175 0 1 31137
box 0 0 1 1
use contact_14  contact_14_110
timestamp 1643678851
transform 1 0 2971 0 1 31193
box 0 0 1 1
use contact_14  contact_14_111
timestamp 1643678851
transform 1 0 3515 0 1 29785
box 0 0 1 1
use contact_14  contact_14_112
timestamp 1643678851
transform 1 0 3175 0 1 29729
box 0 0 1 1
use contact_14  contact_14_113
timestamp 1643678851
transform 1 0 2903 0 1 29673
box 0 0 1 1
use contact_14  contact_14_114
timestamp 1643678851
transform 1 0 3515 0 1 29617
box 0 0 1 1
use contact_14  contact_14_115
timestamp 1643678851
transform 1 0 3175 0 1 29561
box 0 0 1 1
use contact_14  contact_14_116
timestamp 1643678851
transform 1 0 2835 0 1 29505
box 0 0 1 1
use contact_14  contact_14_117
timestamp 1643678851
transform 1 0 3515 0 1 29449
box 0 0 1 1
use contact_14  contact_14_118
timestamp 1643678851
transform 1 0 3175 0 1 29393
box 0 0 1 1
use contact_14  contact_14_119
timestamp 1643678851
transform 1 0 2767 0 1 29337
box 0 0 1 1
use contact_14  contact_14_120
timestamp 1643678851
transform 1 0 3515 0 1 27717
box 0 0 1 1
use contact_14  contact_14_121
timestamp 1643678851
transform 1 0 3107 0 1 27773
box 0 0 1 1
use contact_14  contact_14_122
timestamp 1643678851
transform 1 0 2971 0 1 27829
box 0 0 1 1
use contact_14  contact_14_123
timestamp 1643678851
transform 1 0 3515 0 1 27885
box 0 0 1 1
use contact_14  contact_14_124
timestamp 1643678851
transform 1 0 3107 0 1 27941
box 0 0 1 1
use contact_14  contact_14_125
timestamp 1643678851
transform 1 0 2903 0 1 27997
box 0 0 1 1
use contact_14  contact_14_126
timestamp 1643678851
transform 1 0 3515 0 1 28053
box 0 0 1 1
use contact_14  contact_14_127
timestamp 1643678851
transform 1 0 3107 0 1 28109
box 0 0 1 1
use contact_14  contact_14_128
timestamp 1643678851
transform 1 0 2835 0 1 28165
box 0 0 1 1
use contact_14  contact_14_129
timestamp 1643678851
transform 1 0 3515 0 1 26757
box 0 0 1 1
use contact_14  contact_14_130
timestamp 1643678851
transform 1 0 3107 0 1 26701
box 0 0 1 1
use contact_14  contact_14_131
timestamp 1643678851
transform 1 0 2767 0 1 26645
box 0 0 1 1
use contact_14  contact_14_132
timestamp 1643678851
transform 1 0 3515 0 1 26589
box 0 0 1 1
use contact_14  contact_14_133
timestamp 1643678851
transform 1 0 3039 0 1 26533
box 0 0 1 1
use contact_14  contact_14_134
timestamp 1643678851
transform 1 0 2971 0 1 26477
box 0 0 1 1
use contact_14  contact_14_135
timestamp 1643678851
transform 1 0 3515 0 1 26421
box 0 0 1 1
use contact_14  contact_14_136
timestamp 1643678851
transform 1 0 3039 0 1 26365
box 0 0 1 1
use contact_14  contact_14_137
timestamp 1643678851
transform 1 0 2903 0 1 26309
box 0 0 1 1
use contact_14  contact_14_138
timestamp 1643678851
transform 1 0 3515 0 1 24689
box 0 0 1 1
use contact_14  contact_14_139
timestamp 1643678851
transform 1 0 3039 0 1 24745
box 0 0 1 1
use contact_14  contact_14_140
timestamp 1643678851
transform 1 0 2835 0 1 24801
box 0 0 1 1
use contact_14  contact_14_141
timestamp 1643678851
transform 1 0 3515 0 1 24857
box 0 0 1 1
use contact_14  contact_14_142
timestamp 1643678851
transform 1 0 3039 0 1 24913
box 0 0 1 1
use contact_14  contact_14_143
timestamp 1643678851
transform 1 0 2767 0 1 24969
box 0 0 1 1
use contact_14  contact_14_144
timestamp 1643678851
transform 1 0 3447 0 1 25025
box 0 0 1 1
use contact_14  contact_14_145
timestamp 1643678851
transform 1 0 3243 0 1 25081
box 0 0 1 1
use contact_14  contact_14_146
timestamp 1643678851
transform 1 0 2971 0 1 25137
box 0 0 1 1
use contact_14  contact_14_147
timestamp 1643678851
transform 1 0 3447 0 1 23729
box 0 0 1 1
use contact_14  contact_14_148
timestamp 1643678851
transform 1 0 3243 0 1 23673
box 0 0 1 1
use contact_14  contact_14_149
timestamp 1643678851
transform 1 0 2903 0 1 23617
box 0 0 1 1
use contact_14  contact_14_150
timestamp 1643678851
transform 1 0 3447 0 1 23561
box 0 0 1 1
use contact_14  contact_14_151
timestamp 1643678851
transform 1 0 3243 0 1 23505
box 0 0 1 1
use contact_14  contact_14_152
timestamp 1643678851
transform 1 0 2835 0 1 23449
box 0 0 1 1
use contact_14  contact_14_153
timestamp 1643678851
transform 1 0 3447 0 1 23393
box 0 0 1 1
use contact_14  contact_14_154
timestamp 1643678851
transform 1 0 3243 0 1 23337
box 0 0 1 1
use contact_14  contact_14_155
timestamp 1643678851
transform 1 0 2767 0 1 23281
box 0 0 1 1
use contact_14  contact_14_156
timestamp 1643678851
transform 1 0 3447 0 1 21661
box 0 0 1 1
use contact_14  contact_14_157
timestamp 1643678851
transform 1 0 3175 0 1 21717
box 0 0 1 1
use contact_14  contact_14_158
timestamp 1643678851
transform 1 0 2971 0 1 21773
box 0 0 1 1
use contact_14  contact_14_159
timestamp 1643678851
transform 1 0 3447 0 1 21829
box 0 0 1 1
use contact_14  contact_14_160
timestamp 1643678851
transform 1 0 3175 0 1 21885
box 0 0 1 1
use contact_14  contact_14_161
timestamp 1643678851
transform 1 0 2903 0 1 21941
box 0 0 1 1
use contact_14  contact_14_162
timestamp 1643678851
transform 1 0 3447 0 1 21997
box 0 0 1 1
use contact_14  contact_14_163
timestamp 1643678851
transform 1 0 3175 0 1 22053
box 0 0 1 1
use contact_14  contact_14_164
timestamp 1643678851
transform 1 0 2835 0 1 22109
box 0 0 1 1
use contact_14  contact_14_165
timestamp 1643678851
transform 1 0 3447 0 1 20701
box 0 0 1 1
use contact_14  contact_14_166
timestamp 1643678851
transform 1 0 3175 0 1 20645
box 0 0 1 1
use contact_14  contact_14_167
timestamp 1643678851
transform 1 0 2767 0 1 20589
box 0 0 1 1
use contact_14  contact_14_168
timestamp 1643678851
transform 1 0 3447 0 1 20533
box 0 0 1 1
use contact_14  contact_14_169
timestamp 1643678851
transform 1 0 3107 0 1 20477
box 0 0 1 1
use contact_14  contact_14_170
timestamp 1643678851
transform 1 0 2971 0 1 20421
box 0 0 1 1
use contact_14  contact_14_171
timestamp 1643678851
transform 1 0 3447 0 1 20365
box 0 0 1 1
use contact_14  contact_14_172
timestamp 1643678851
transform 1 0 3107 0 1 20309
box 0 0 1 1
use contact_14  contact_14_173
timestamp 1643678851
transform 1 0 2903 0 1 20253
box 0 0 1 1
use contact_14  contact_14_174
timestamp 1643678851
transform 1 0 3447 0 1 18633
box 0 0 1 1
use contact_14  contact_14_175
timestamp 1643678851
transform 1 0 3107 0 1 18689
box 0 0 1 1
use contact_14  contact_14_176
timestamp 1643678851
transform 1 0 2835 0 1 18745
box 0 0 1 1
use contact_14  contact_14_177
timestamp 1643678851
transform 1 0 3447 0 1 18801
box 0 0 1 1
use contact_14  contact_14_178
timestamp 1643678851
transform 1 0 3107 0 1 18857
box 0 0 1 1
use contact_14  contact_14_179
timestamp 1643678851
transform 1 0 2767 0 1 18913
box 0 0 1 1
use contact_14  contact_14_180
timestamp 1643678851
transform 1 0 3447 0 1 18969
box 0 0 1 1
use contact_14  contact_14_181
timestamp 1643678851
transform 1 0 3039 0 1 19025
box 0 0 1 1
use contact_14  contact_14_182
timestamp 1643678851
transform 1 0 2971 0 1 19081
box 0 0 1 1
use contact_14  contact_14_183
timestamp 1643678851
transform 1 0 3447 0 1 17673
box 0 0 1 1
use contact_14  contact_14_184
timestamp 1643678851
transform 1 0 3039 0 1 17617
box 0 0 1 1
use contact_14  contact_14_185
timestamp 1643678851
transform 1 0 2903 0 1 17561
box 0 0 1 1
use contact_14  contact_14_186
timestamp 1643678851
transform 1 0 3447 0 1 17505
box 0 0 1 1
use contact_14  contact_14_187
timestamp 1643678851
transform 1 0 3039 0 1 17449
box 0 0 1 1
use contact_14  contact_14_188
timestamp 1643678851
transform 1 0 2835 0 1 17393
box 0 0 1 1
use contact_14  contact_14_189
timestamp 1643678851
transform 1 0 3447 0 1 17337
box 0 0 1 1
use contact_14  contact_14_190
timestamp 1643678851
transform 1 0 3039 0 1 17281
box 0 0 1 1
use contact_14  contact_14_191
timestamp 1643678851
transform 1 0 2767 0 1 17225
box 0 0 1 1
use contact_14  contact_14_192
timestamp 1643678851
transform 1 0 3379 0 1 15605
box 0 0 1 1
use contact_14  contact_14_193
timestamp 1643678851
transform 1 0 3243 0 1 15661
box 0 0 1 1
use contact_14  contact_14_194
timestamp 1643678851
transform 1 0 2971 0 1 15717
box 0 0 1 1
use contact_14  contact_14_195
timestamp 1643678851
transform 1 0 3379 0 1 15773
box 0 0 1 1
use contact_14  contact_14_196
timestamp 1643678851
transform 1 0 3243 0 1 15829
box 0 0 1 1
use contact_14  contact_14_197
timestamp 1643678851
transform 1 0 2903 0 1 15885
box 0 0 1 1
use contact_14  contact_14_198
timestamp 1643678851
transform 1 0 3379 0 1 15941
box 0 0 1 1
use contact_14  contact_14_199
timestamp 1643678851
transform 1 0 3243 0 1 15997
box 0 0 1 1
use contact_14  contact_14_200
timestamp 1643678851
transform 1 0 2835 0 1 16053
box 0 0 1 1
use contact_14  contact_14_201
timestamp 1643678851
transform 1 0 3379 0 1 14645
box 0 0 1 1
use contact_14  contact_14_202
timestamp 1643678851
transform 1 0 3243 0 1 14589
box 0 0 1 1
use contact_14  contact_14_203
timestamp 1643678851
transform 1 0 2767 0 1 14533
box 0 0 1 1
use contact_14  contact_14_204
timestamp 1643678851
transform 1 0 3379 0 1 14477
box 0 0 1 1
use contact_14  contact_14_205
timestamp 1643678851
transform 1 0 3175 0 1 14421
box 0 0 1 1
use contact_14  contact_14_206
timestamp 1643678851
transform 1 0 2971 0 1 14365
box 0 0 1 1
use contact_14  contact_14_207
timestamp 1643678851
transform 1 0 3379 0 1 14309
box 0 0 1 1
use contact_14  contact_14_208
timestamp 1643678851
transform 1 0 3175 0 1 14253
box 0 0 1 1
use contact_14  contact_14_209
timestamp 1643678851
transform 1 0 2903 0 1 14197
box 0 0 1 1
use contact_14  contact_14_210
timestamp 1643678851
transform 1 0 3379 0 1 12577
box 0 0 1 1
use contact_14  contact_14_211
timestamp 1643678851
transform 1 0 3175 0 1 12633
box 0 0 1 1
use contact_14  contact_14_212
timestamp 1643678851
transform 1 0 2835 0 1 12689
box 0 0 1 1
use contact_14  contact_14_213
timestamp 1643678851
transform 1 0 3379 0 1 12745
box 0 0 1 1
use contact_14  contact_14_214
timestamp 1643678851
transform 1 0 3175 0 1 12801
box 0 0 1 1
use contact_14  contact_14_215
timestamp 1643678851
transform 1 0 2767 0 1 12857
box 0 0 1 1
use contact_14  contact_14_216
timestamp 1643678851
transform 1 0 3379 0 1 12913
box 0 0 1 1
use contact_14  contact_14_217
timestamp 1643678851
transform 1 0 3107 0 1 12969
box 0 0 1 1
use contact_14  contact_14_218
timestamp 1643678851
transform 1 0 2971 0 1 13025
box 0 0 1 1
use contact_14  contact_14_219
timestamp 1643678851
transform 1 0 3379 0 1 11617
box 0 0 1 1
use contact_14  contact_14_220
timestamp 1643678851
transform 1 0 3107 0 1 11561
box 0 0 1 1
use contact_14  contact_14_221
timestamp 1643678851
transform 1 0 2903 0 1 11505
box 0 0 1 1
use contact_14  contact_14_222
timestamp 1643678851
transform 1 0 3379 0 1 11449
box 0 0 1 1
use contact_14  contact_14_223
timestamp 1643678851
transform 1 0 3107 0 1 11393
box 0 0 1 1
use contact_14  contact_14_224
timestamp 1643678851
transform 1 0 2835 0 1 11337
box 0 0 1 1
use contact_14  contact_14_225
timestamp 1643678851
transform 1 0 3379 0 1 11281
box 0 0 1 1
use contact_14  contact_14_226
timestamp 1643678851
transform 1 0 3107 0 1 11225
box 0 0 1 1
use contact_14  contact_14_227
timestamp 1643678851
transform 1 0 2767 0 1 11169
box 0 0 1 1
use contact_14  contact_14_228
timestamp 1643678851
transform 1 0 3379 0 1 9549
box 0 0 1 1
use contact_14  contact_14_229
timestamp 1643678851
transform 1 0 3039 0 1 9605
box 0 0 1 1
use contact_14  contact_14_230
timestamp 1643678851
transform 1 0 2971 0 1 9661
box 0 0 1 1
use contact_14  contact_14_231
timestamp 1643678851
transform 1 0 3379 0 1 9717
box 0 0 1 1
use contact_14  contact_14_232
timestamp 1643678851
transform 1 0 3039 0 1 9773
box 0 0 1 1
use contact_14  contact_14_233
timestamp 1643678851
transform 1 0 2903 0 1 9829
box 0 0 1 1
use contact_14  contact_14_234
timestamp 1643678851
transform 1 0 3379 0 1 9885
box 0 0 1 1
use contact_14  contact_14_235
timestamp 1643678851
transform 1 0 3039 0 1 9941
box 0 0 1 1
use contact_14  contact_14_236
timestamp 1643678851
transform 1 0 2835 0 1 9997
box 0 0 1 1
use contact_14  contact_14_237
timestamp 1643678851
transform 1 0 3379 0 1 8589
box 0 0 1 1
use contact_14  contact_14_238
timestamp 1643678851
transform 1 0 3039 0 1 8533
box 0 0 1 1
use contact_14  contact_14_239
timestamp 1643678851
transform 1 0 2767 0 1 8477
box 0 0 1 1
use contact_14  contact_14_240
timestamp 1643678851
transform 1 0 3311 0 1 8421
box 0 0 1 1
use contact_14  contact_14_241
timestamp 1643678851
transform 1 0 3243 0 1 8365
box 0 0 1 1
use contact_14  contact_14_242
timestamp 1643678851
transform 1 0 2971 0 1 8309
box 0 0 1 1
use contact_14  contact_14_243
timestamp 1643678851
transform 1 0 3311 0 1 8253
box 0 0 1 1
use contact_14  contact_14_244
timestamp 1643678851
transform 1 0 3243 0 1 8197
box 0 0 1 1
use contact_14  contact_14_245
timestamp 1643678851
transform 1 0 2903 0 1 8141
box 0 0 1 1
use contact_14  contact_14_246
timestamp 1643678851
transform 1 0 3311 0 1 6521
box 0 0 1 1
use contact_14  contact_14_247
timestamp 1643678851
transform 1 0 3243 0 1 6577
box 0 0 1 1
use contact_14  contact_14_248
timestamp 1643678851
transform 1 0 2835 0 1 6633
box 0 0 1 1
use contact_14  contact_14_249
timestamp 1643678851
transform 1 0 3311 0 1 6689
box 0 0 1 1
use contact_14  contact_14_250
timestamp 1643678851
transform 1 0 3243 0 1 6745
box 0 0 1 1
use contact_14  contact_14_251
timestamp 1643678851
transform 1 0 2767 0 1 6801
box 0 0 1 1
use contact_14  contact_14_252
timestamp 1643678851
transform 1 0 3311 0 1 6857
box 0 0 1 1
use contact_14  contact_14_253
timestamp 1643678851
transform 1 0 3175 0 1 6913
box 0 0 1 1
use contact_14  contact_14_254
timestamp 1643678851
transform 1 0 2971 0 1 6969
box 0 0 1 1
use contact_14  contact_14_255
timestamp 1643678851
transform 1 0 3311 0 1 5561
box 0 0 1 1
use contact_14  contact_14_256
timestamp 1643678851
transform 1 0 3175 0 1 5505
box 0 0 1 1
use contact_14  contact_14_257
timestamp 1643678851
transform 1 0 2903 0 1 5449
box 0 0 1 1
use contact_14  contact_14_258
timestamp 1643678851
transform 1 0 3311 0 1 5393
box 0 0 1 1
use contact_14  contact_14_259
timestamp 1643678851
transform 1 0 3175 0 1 5337
box 0 0 1 1
use contact_14  contact_14_260
timestamp 1643678851
transform 1 0 2835 0 1 5281
box 0 0 1 1
use contact_14  contact_14_261
timestamp 1643678851
transform 1 0 3311 0 1 5225
box 0 0 1 1
use contact_14  contact_14_262
timestamp 1643678851
transform 1 0 3175 0 1 5169
box 0 0 1 1
use contact_14  contact_14_263
timestamp 1643678851
transform 1 0 2767 0 1 5113
box 0 0 1 1
use contact_14  contact_14_264
timestamp 1643678851
transform 1 0 3311 0 1 3493
box 0 0 1 1
use contact_14  contact_14_265
timestamp 1643678851
transform 1 0 3107 0 1 3549
box 0 0 1 1
use contact_14  contact_14_266
timestamp 1643678851
transform 1 0 2971 0 1 3605
box 0 0 1 1
use contact_14  contact_14_267
timestamp 1643678851
transform 1 0 3311 0 1 3661
box 0 0 1 1
use contact_14  contact_14_268
timestamp 1643678851
transform 1 0 3107 0 1 3717
box 0 0 1 1
use contact_14  contact_14_269
timestamp 1643678851
transform 1 0 2903 0 1 3773
box 0 0 1 1
use contact_14  contact_14_270
timestamp 1643678851
transform 1 0 3311 0 1 3829
box 0 0 1 1
use contact_14  contact_14_271
timestamp 1643678851
transform 1 0 3107 0 1 3885
box 0 0 1 1
use contact_14  contact_14_272
timestamp 1643678851
transform 1 0 2835 0 1 3941
box 0 0 1 1
use contact_14  contact_14_273
timestamp 1643678851
transform 1 0 3311 0 1 2533
box 0 0 1 1
use contact_14  contact_14_274
timestamp 1643678851
transform 1 0 3107 0 1 2477
box 0 0 1 1
use contact_14  contact_14_275
timestamp 1643678851
transform 1 0 2767 0 1 2421
box 0 0 1 1
use contact_14  contact_14_276
timestamp 1643678851
transform 1 0 3311 0 1 2365
box 0 0 1 1
use contact_14  contact_14_277
timestamp 1643678851
transform 1 0 3039 0 1 2309
box 0 0 1 1
use contact_14  contact_14_278
timestamp 1643678851
transform 1 0 2971 0 1 2253
box 0 0 1 1
use contact_14  contact_14_279
timestamp 1643678851
transform 1 0 3311 0 1 2197
box 0 0 1 1
use contact_14  contact_14_280
timestamp 1643678851
transform 1 0 3039 0 1 2141
box 0 0 1 1
use contact_14  contact_14_281
timestamp 1643678851
transform 1 0 2903 0 1 2085
box 0 0 1 1
use contact_14  contact_14_282
timestamp 1643678851
transform 1 0 3311 0 1 465
box 0 0 1 1
use contact_14  contact_14_283
timestamp 1643678851
transform 1 0 3039 0 1 521
box 0 0 1 1
use contact_14  contact_14_284
timestamp 1643678851
transform 1 0 2835 0 1 577
box 0 0 1 1
use contact_14  contact_14_285
timestamp 1643678851
transform 1 0 3311 0 1 633
box 0 0 1 1
use contact_14  contact_14_286
timestamp 1643678851
transform 1 0 3039 0 1 689
box 0 0 1 1
use contact_14  contact_14_287
timestamp 1643678851
transform 1 0 2767 0 1 745
box 0 0 1 1
use contact_14  contact_14_288
timestamp 1643678851
transform 1 0 408 0 1 22265
box 0 0 1 1
use contact_17  contact_17_208
timestamp 1643678851
transform 1 0 708 0 1 22265
box 0 0 1 1
use contact_14  contact_14_289
timestamp 1643678851
transform 1 0 340 0 1 20809
box 0 0 1 1
use contact_17  contact_17_209
timestamp 1643678851
transform 1 0 640 0 1 20809
box 0 0 1 1
use contact_14  contact_14_290
timestamp 1643678851
transform 1 0 272 0 1 19185
box 0 0 1 1
use contact_17  contact_17_210
timestamp 1643678851
transform 1 0 572 0 1 19185
box 0 0 1 1
use contact_14  contact_14_291
timestamp 1643678851
transform 1 0 204 0 1 11573
box 0 0 1 1
use contact_17  contact_17_211
timestamp 1643678851
transform 1 0 1002 0 1 11573
box 0 0 1 1
use contact_14  contact_14_292
timestamp 1643678851
transform 1 0 136 0 1 9949
box 0 0 1 1
use contact_17  contact_17_212
timestamp 1643678851
transform 1 0 934 0 1 9949
box 0 0 1 1
use contact_14  contact_14_293
timestamp 1643678851
transform 1 0 68 0 1 2337
box 0 0 1 1
use contact_17  contact_17_213
timestamp 1643678851
transform 1 0 1002 0 1 2337
box 0 0 1 1
use contact_14  contact_14_294
timestamp 1643678851
transform 1 0 0 0 1 713
box 0 0 1 1
use contact_17  contact_17_214
timestamp 1643678851
transform 1 0 934 0 1 713
box 0 0 1 1
use dec_cell3_2r1w  dec_cell3_2r1w_0
timestamp 1643678851
transform 1 0 2700 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_1
timestamp 1643678851
transform 1 0 2700 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_2
timestamp 1643678851
transform 1 0 2700 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_3
timestamp 1643678851
transform 1 0 2700 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_4
timestamp 1643678851
transform 1 0 2700 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_5
timestamp 1643678851
transform 1 0 2700 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_6
timestamp 1643678851
transform 1 0 2700 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_7
timestamp 1643678851
transform 1 0 2700 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_8
timestamp 1643678851
transform 1 0 2700 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_9
timestamp 1643678851
transform 1 0 2700 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_10
timestamp 1643678851
transform 1 0 2700 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_11
timestamp 1643678851
transform 1 0 2700 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_12
timestamp 1643678851
transform 1 0 2700 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_13
timestamp 1643678851
transform 1 0 2700 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_14
timestamp 1643678851
transform 1 0 2700 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_15
timestamp 1643678851
transform 1 0 2700 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_16
timestamp 1643678851
transform 1 0 2700 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_17
timestamp 1643678851
transform 1 0 2700 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_18
timestamp 1643678851
transform 1 0 2700 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_19
timestamp 1643678851
transform 1 0 2700 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_20
timestamp 1643678851
transform 1 0 2700 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_21
timestamp 1643678851
transform 1 0 2700 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_22
timestamp 1643678851
transform 1 0 2700 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_23
timestamp 1643678851
transform 1 0 2700 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_24
timestamp 1643678851
transform 1 0 2700 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_25
timestamp 1643678851
transform 1 0 2700 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_26
timestamp 1643678851
transform 1 0 2700 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_27
timestamp 1643678851
transform 1 0 2700 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_28
timestamp 1643678851
transform 1 0 2700 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_29
timestamp 1643678851
transform 1 0 2700 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_30
timestamp 1643678851
transform 1 0 2700 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_31
timestamp 1643678851
transform 1 0 2700 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_32
timestamp 1643678851
transform 1 0 2700 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_33
timestamp 1643678851
transform 1 0 2700 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_34
timestamp 1643678851
transform 1 0 2700 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_35
timestamp 1643678851
transform 1 0 2700 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_36
timestamp 1643678851
transform 1 0 2700 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_37
timestamp 1643678851
transform 1 0 2700 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_38
timestamp 1643678851
transform 1 0 2700 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_39
timestamp 1643678851
transform 1 0 2700 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_40
timestamp 1643678851
transform 1 0 2700 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_41
timestamp 1643678851
transform 1 0 2700 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_42
timestamp 1643678851
transform 1 0 2700 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_43
timestamp 1643678851
transform 1 0 2700 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_44
timestamp 1643678851
transform 1 0 2700 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_45
timestamp 1643678851
transform 1 0 2700 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_46
timestamp 1643678851
transform 1 0 2700 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_47
timestamp 1643678851
transform 1 0 2700 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_48
timestamp 1643678851
transform 1 0 2700 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_49
timestamp 1643678851
transform 1 0 2700 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_50
timestamp 1643678851
transform 1 0 2700 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_51
timestamp 1643678851
transform 1 0 2700 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_52
timestamp 1643678851
transform 1 0 2700 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_53
timestamp 1643678851
transform 1 0 2700 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_54
timestamp 1643678851
transform 1 0 2700 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_55
timestamp 1643678851
transform 1 0 2700 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_56
timestamp 1643678851
transform 1 0 2700 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_57
timestamp 1643678851
transform 1 0 2700 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_58
timestamp 1643678851
transform 1 0 2700 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_59
timestamp 1643678851
transform 1 0 2700 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_60
timestamp 1643678851
transform 1 0 2700 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_61
timestamp 1643678851
transform 1 0 2700 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_62
timestamp 1643678851
transform 1 0 2700 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_63
timestamp 1643678851
transform 1 0 2700 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_64
timestamp 1643678851
transform 1 0 3856 0 -1 48448
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_65
timestamp 1643678851
transform 1 0 3856 0 1 45420
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_66
timestamp 1643678851
transform 1 0 3856 0 -1 45420
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_67
timestamp 1643678851
transform 1 0 3856 0 1 42392
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_68
timestamp 1643678851
transform 1 0 3856 0 -1 42392
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_69
timestamp 1643678851
transform 1 0 3856 0 1 39364
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_70
timestamp 1643678851
transform 1 0 3856 0 -1 39364
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_71
timestamp 1643678851
transform 1 0 3856 0 1 36336
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_72
timestamp 1643678851
transform 1 0 3856 0 -1 36336
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_73
timestamp 1643678851
transform 1 0 3856 0 1 33308
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_74
timestamp 1643678851
transform 1 0 3856 0 -1 33308
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_75
timestamp 1643678851
transform 1 0 3856 0 1 30280
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_76
timestamp 1643678851
transform 1 0 3856 0 -1 30280
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_77
timestamp 1643678851
transform 1 0 3856 0 1 27252
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_78
timestamp 1643678851
transform 1 0 3856 0 -1 27252
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_79
timestamp 1643678851
transform 1 0 3856 0 1 24224
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_80
timestamp 1643678851
transform 1 0 3856 0 -1 24224
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_81
timestamp 1643678851
transform 1 0 3856 0 1 21196
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_82
timestamp 1643678851
transform 1 0 3856 0 -1 21196
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_83
timestamp 1643678851
transform 1 0 3856 0 1 18168
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_84
timestamp 1643678851
transform 1 0 3856 0 -1 18168
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_85
timestamp 1643678851
transform 1 0 3856 0 1 15140
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_86
timestamp 1643678851
transform 1 0 3856 0 -1 15140
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_87
timestamp 1643678851
transform 1 0 3856 0 1 12112
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_88
timestamp 1643678851
transform 1 0 3856 0 -1 12112
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_89
timestamp 1643678851
transform 1 0 3856 0 1 9084
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_90
timestamp 1643678851
transform 1 0 3856 0 -1 9084
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_91
timestamp 1643678851
transform 1 0 3856 0 1 6056
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_92
timestamp 1643678851
transform 1 0 3856 0 -1 6056
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_93
timestamp 1643678851
transform 1 0 3856 0 1 3028
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_94
timestamp 1643678851
transform 1 0 3856 0 -1 3028
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_95
timestamp 1643678851
transform 1 0 3856 0 1 0
box 0 -42 1494 1616
use hierarchical_predecode3x8  hierarchical_predecode3x8_0
timestamp 1643678851
transform 1 0 505 0 1 18472
box 0 -34 2231 12354
use hierarchical_predecode2x4  hierarchical_predecode2x4_0
timestamp 1643678851
transform 1 0 867 0 1 9236
box 0 -34 1869 6194
use hierarchical_predecode2x4  hierarchical_predecode2x4_1
timestamp 1643678851
transform 1 0 867 0 1 0
box 0 -34 1869 6194
<< labels >>
rlabel metal2 s 1 0 29 30792 4 addr_0
rlabel metal2 s 69 0 97 30792 4 addr_1
rlabel metal2 s 137 0 165 30792 4 addr_2
rlabel metal2 s 205 0 233 30792 4 addr_3
rlabel metal2 s 273 0 301 30792 4 addr_4
rlabel metal2 s 341 0 369 30792 4 addr_5
rlabel metal2 s 409 0 437 30792 4 addr_6
rlabel metal1 s 5066 702 5350 730 4 decode0_0
rlabel metal1 s 5274 848 5350 876 4 decode1_0
rlabel metal1 s 4984 580 5350 608 4 decode2_0
rlabel metal1 s 5066 2298 5350 2326 4 decode0_1
rlabel metal1 s 5274 2152 5350 2180 4 decode1_1
rlabel metal1 s 4984 2420 5350 2448 4 decode2_1
rlabel metal1 s 5066 3730 5350 3758 4 decode0_2
rlabel metal1 s 5274 3876 5350 3904 4 decode1_2
rlabel metal1 s 4984 3608 5350 3636 4 decode2_2
rlabel metal1 s 5066 5326 5350 5354 4 decode0_3
rlabel metal1 s 5274 5180 5350 5208 4 decode1_3
rlabel metal1 s 4984 5448 5350 5476 4 decode2_3
rlabel metal1 s 5066 6758 5350 6786 4 decode0_4
rlabel metal1 s 5274 6904 5350 6932 4 decode1_4
rlabel metal1 s 4984 6636 5350 6664 4 decode2_4
rlabel metal1 s 5066 8354 5350 8382 4 decode0_5
rlabel metal1 s 5274 8208 5350 8236 4 decode1_5
rlabel metal1 s 4984 8476 5350 8504 4 decode2_5
rlabel metal1 s 5066 9786 5350 9814 4 decode0_6
rlabel metal1 s 5274 9932 5350 9960 4 decode1_6
rlabel metal1 s 4984 9664 5350 9692 4 decode2_6
rlabel metal1 s 5066 11382 5350 11410 4 decode0_7
rlabel metal1 s 5274 11236 5350 11264 4 decode1_7
rlabel metal1 s 4984 11504 5350 11532 4 decode2_7
rlabel metal1 s 5066 12814 5350 12842 4 decode0_8
rlabel metal1 s 5274 12960 5350 12988 4 decode1_8
rlabel metal1 s 4984 12692 5350 12720 4 decode2_8
rlabel metal1 s 5066 14410 5350 14438 4 decode0_9
rlabel metal1 s 5274 14264 5350 14292 4 decode1_9
rlabel metal1 s 4984 14532 5350 14560 4 decode2_9
rlabel metal1 s 5066 15842 5350 15870 4 decode0_10
rlabel metal1 s 5274 15988 5350 16016 4 decode1_10
rlabel metal1 s 4984 15720 5350 15748 4 decode2_10
rlabel metal1 s 5066 17438 5350 17466 4 decode0_11
rlabel metal1 s 5274 17292 5350 17320 4 decode1_11
rlabel metal1 s 4984 17560 5350 17588 4 decode2_11
rlabel metal1 s 5066 18870 5350 18898 4 decode0_12
rlabel metal1 s 5274 19016 5350 19044 4 decode1_12
rlabel metal1 s 4984 18748 5350 18776 4 decode2_12
rlabel metal1 s 5066 20466 5350 20494 4 decode0_13
rlabel metal1 s 5274 20320 5350 20348 4 decode1_13
rlabel metal1 s 4984 20588 5350 20616 4 decode2_13
rlabel metal1 s 5066 21898 5350 21926 4 decode0_14
rlabel metal1 s 5274 22044 5350 22072 4 decode1_14
rlabel metal1 s 4984 21776 5350 21804 4 decode2_14
rlabel metal1 s 5066 23494 5350 23522 4 decode0_15
rlabel metal1 s 5274 23348 5350 23376 4 decode1_15
rlabel metal1 s 4984 23616 5350 23644 4 decode2_15
rlabel metal1 s 5066 24926 5350 24954 4 decode0_16
rlabel metal1 s 5274 25072 5350 25100 4 decode1_16
rlabel metal1 s 4984 24804 5350 24832 4 decode2_16
rlabel metal1 s 5066 26522 5350 26550 4 decode0_17
rlabel metal1 s 5274 26376 5350 26404 4 decode1_17
rlabel metal1 s 4984 26644 5350 26672 4 decode2_17
rlabel metal1 s 5066 27954 5350 27982 4 decode0_18
rlabel metal1 s 5274 28100 5350 28128 4 decode1_18
rlabel metal1 s 4984 27832 5350 27860 4 decode2_18
rlabel metal1 s 5066 29550 5350 29578 4 decode0_19
rlabel metal1 s 5274 29404 5350 29432 4 decode1_19
rlabel metal1 s 4984 29672 5350 29700 4 decode2_19
rlabel metal1 s 5066 30982 5350 31010 4 decode0_20
rlabel metal1 s 5274 31128 5350 31156 4 decode1_20
rlabel metal1 s 4984 30860 5350 30888 4 decode2_20
rlabel metal1 s 5066 32578 5350 32606 4 decode0_21
rlabel metal1 s 5274 32432 5350 32460 4 decode1_21
rlabel metal1 s 4984 32700 5350 32728 4 decode2_21
rlabel metal1 s 5066 34010 5350 34038 4 decode0_22
rlabel metal1 s 5274 34156 5350 34184 4 decode1_22
rlabel metal1 s 4984 33888 5350 33916 4 decode2_22
rlabel metal1 s 5066 35606 5350 35634 4 decode0_23
rlabel metal1 s 5274 35460 5350 35488 4 decode1_23
rlabel metal1 s 4984 35728 5350 35756 4 decode2_23
rlabel metal1 s 5066 37038 5350 37066 4 decode0_24
rlabel metal1 s 5274 37184 5350 37212 4 decode1_24
rlabel metal1 s 4984 36916 5350 36944 4 decode2_24
rlabel metal1 s 5066 38634 5350 38662 4 decode0_25
rlabel metal1 s 5274 38488 5350 38516 4 decode1_25
rlabel metal1 s 4984 38756 5350 38784 4 decode2_25
rlabel metal1 s 5066 40066 5350 40094 4 decode0_26
rlabel metal1 s 5274 40212 5350 40240 4 decode1_26
rlabel metal1 s 4984 39944 5350 39972 4 decode2_26
rlabel metal1 s 5066 41662 5350 41690 4 decode0_27
rlabel metal1 s 5274 41516 5350 41544 4 decode1_27
rlabel metal1 s 4984 41784 5350 41812 4 decode2_27
rlabel metal1 s 5066 43094 5350 43122 4 decode0_28
rlabel metal1 s 5274 43240 5350 43268 4 decode1_28
rlabel metal1 s 4984 42972 5350 43000 4 decode2_28
rlabel metal1 s 5066 44690 5350 44718 4 decode0_29
rlabel metal1 s 5274 44544 5350 44572 4 decode1_29
rlabel metal1 s 4984 44812 5350 44840 4 decode2_29
rlabel metal1 s 5066 46122 5350 46150 4 decode0_30
rlabel metal1 s 5274 46268 5350 46296 4 decode1_30
rlabel metal1 s 4984 46000 5350 46028 4 decode2_30
rlabel metal1 s 5066 47718 5350 47746 4 decode0_31
rlabel metal1 s 5274 47572 5350 47600 4 decode1_31
rlabel metal1 s 4984 47840 5350 47868 4 decode2_31
rlabel metal2 s 2768 0 2796 49244 4 predecode_0
rlabel metal2 s 2836 0 2864 49244 4 predecode_1
rlabel metal2 s 2904 0 2932 49244 4 predecode_2
rlabel metal2 s 2972 0 3000 49244 4 predecode_3
rlabel metal2 s 3040 0 3068 49244 4 predecode_4
rlabel metal2 s 3108 0 3136 49244 4 predecode_5
rlabel metal2 s 3176 0 3204 49244 4 predecode_6
rlabel metal2 s 3244 0 3272 49244 4 predecode_7
rlabel metal2 s 3312 0 3340 49244 4 predecode_8
rlabel metal2 s 3380 0 3408 49244 4 predecode_9
rlabel metal2 s 3448 0 3476 49244 4 predecode_10
rlabel metal2 s 3516 0 3544 49244 4 predecode_11
rlabel metal2 s 3584 0 3612 49244 4 predecode_12
rlabel metal2 s 3652 0 3680 49244 4 predecode_13
rlabel metal2 s 3720 0 3748 49244 4 predecode_14
rlabel metal2 s 3788 0 3816 49244 4 predecode_15
rlabel metal3 s 1045 10743 1177 10809 4 vdd
rlabel metal3 s 5298 10565 5430 10631 4 vdd
rlabel metal3 s 5298 43873 5430 43939 4 vdd
rlabel metal3 s 1804 4587 1936 4653 4 vdd
rlabel metal3 s 1045 4587 1177 4653 4 vdd
rlabel metal3 s 5298 34789 5430 34855 4 vdd
rlabel metal3 s 5364 34822 5364 34822 4 vdd
rlabel metal3 s 5298 40845 5430 40911 4 vdd
rlabel metal3 s 1045 1507 1177 1573 4 vdd
rlabel metal3 s 5364 40878 5364 40878 4 vdd
rlabel metal3 s 5298 4509 5430 4575 4 vdd
rlabel metal3 s 751 26139 883 26205 4 vdd
rlabel metal3 s 1646 23059 1778 23125 4 vdd
rlabel metal3 s 5298 7537 5430 7603 4 vdd
rlabel metal3 s 5298 13593 5430 13659 4 vdd
rlabel metal3 s 751 29219 883 29285 4 vdd
rlabel metal3 s 751 23059 883 23125 4 vdd
rlabel metal3 s 1045 13823 1177 13889 4 vdd
rlabel metal3 s 5298 37817 5430 37883 4 vdd
rlabel metal3 s 1804 1507 1936 1573 4 vdd
rlabel metal3 s 1804 10743 1936 10809 4 vdd
rlabel metal3 s 5298 19649 5430 19715 4 vdd
rlabel metal3 s 5298 1481 5430 1547 4 vdd
rlabel metal3 s 1646 19979 1778 20045 4 vdd
rlabel metal3 s 5298 46901 5430 46967 4 vdd
rlabel metal3 s 5298 16621 5430 16687 4 vdd
rlabel metal3 s 5298 31761 5430 31827 4 vdd
rlabel metal3 s 5364 46934 5364 46934 4 vdd
rlabel metal3 s 1646 26139 1778 26205 4 vdd
rlabel metal3 s 5298 28733 5430 28799 4 vdd
rlabel metal3 s 1646 29219 1778 29285 4 vdd
rlabel metal3 s 5364 28766 5364 28766 4 vdd
rlabel metal3 s 5298 22677 5430 22743 4 vdd
rlabel metal3 s 1804 13823 1936 13889 4 vdd
rlabel metal3 s 5298 25705 5430 25771 4 vdd
rlabel metal3 s 751 19979 883 20045 4 vdd
rlabel metal3 s 751 24599 883 24665 4 gnd
rlabel metal3 s 1045 3047 1177 3113 4 gnd
rlabel metal3 s 751 21519 883 21585 4 gnd
rlabel metal3 s 5298 6023 5430 6089 4 gnd
rlabel metal3 s 1804 3047 1936 3113 4 gnd
rlabel metal3 s 5298 42359 5430 42425 4 gnd
rlabel metal3 s 751 18439 883 18505 4 gnd
rlabel metal3 s 5298 18135 5430 18201 4 gnd
rlabel metal3 s 5298 -33 5430 33 4 gnd
rlabel metal3 s 5298 45387 5430 45453 4 gnd
rlabel metal3 s 1646 27679 1778 27745 4 gnd
rlabel metal3 s 1646 24599 1778 24665 4 gnd
rlabel metal3 s 1646 30759 1778 30825 4 gnd
rlabel metal3 s 1646 18439 1778 18505 4 gnd
rlabel metal3 s 1804 15363 1936 15429 4 gnd
rlabel metal3 s 5298 2995 5430 3061 4 gnd
rlabel metal3 s 5298 21163 5430 21229 4 gnd
rlabel metal3 s 1646 21519 1778 21585 4 gnd
rlabel metal3 s 1045 12283 1177 12349 4 gnd
rlabel metal3 s 5298 33275 5430 33341 4 gnd
rlabel metal3 s 5298 15107 5430 15173 4 gnd
rlabel metal3 s 751 30759 883 30825 4 gnd
rlabel metal3 s 1045 -33 1177 33 4 gnd
rlabel metal3 s 1045 15363 1177 15429 4 gnd
rlabel metal3 s 5298 12079 5430 12145 4 gnd
rlabel metal3 s 5298 30247 5430 30313 4 gnd
rlabel metal3 s 1045 9203 1177 9269 4 gnd
rlabel metal3 s 5298 48415 5430 48481 4 gnd
rlabel metal3 s 1804 12283 1936 12349 4 gnd
rlabel metal3 s 5298 39331 5430 39397 4 gnd
rlabel metal3 s 1045 6127 1177 6193 4 gnd
rlabel metal3 s 5298 27219 5430 27285 4 gnd
rlabel metal3 s 1804 6127 1936 6193 4 gnd
rlabel metal3 s 5298 36303 5430 36369 4 gnd
rlabel metal3 s 5298 24191 5430 24257 4 gnd
rlabel metal3 s 1804 9203 1936 9269 4 gnd
rlabel metal3 s 5298 9051 5430 9117 4 gnd
rlabel metal3 s 1804 -33 1936 33 4 gnd
rlabel metal3 s 751 27679 883 27745 4 gnd
<< properties >>
string FIXED_BBOX 5298 -33 5430 0
string GDS_FILE sram_0rw2r1w_16_128_sky130A.gds
string GDS_END 1837190
string GDS_START 1711144
<< end >>
