magic
tech sky130A
magscale 1 2
timestamp 1644969367
<< checkpaint >>
rect -1260 -770 51830 7492
<< metal1 >>
rect 0 5824 49323 5852
rect 0 3434 49792 3462
rect 0 3354 49792 3382
rect 0 1503 50570 1531
<< metal2 >>
rect 585 5908 639 5936
rect 2141 5908 2195 5936
rect 3697 5908 3751 5936
rect 5253 5908 5307 5936
rect 6809 5908 6863 5936
rect 8365 5908 8419 5936
rect 9921 5908 9975 5936
rect 11477 5908 11531 5936
rect 13033 5908 13087 5936
rect 14589 5908 14643 5936
rect 16145 5908 16199 5936
rect 17701 5908 17755 5936
rect 19257 5908 19311 5936
rect 20813 5908 20867 5936
rect 22369 5908 22423 5936
rect 23925 5908 23979 5936
rect 25481 5908 25535 5936
rect 27037 5908 27091 5936
rect 28593 5908 28647 5936
rect 30149 5908 30203 5936
rect 31705 5908 31759 5936
rect 33261 5908 33315 5936
rect 34817 5908 34871 5936
rect 36373 5908 36427 5936
rect 37929 5908 37983 5936
rect 39485 5908 39539 5936
rect 41041 5908 41095 5936
rect 42597 5908 42651 5936
rect 44153 5908 44207 5936
rect 45709 5908 45763 5936
rect 47265 5908 47319 5936
rect 48821 5908 48875 5936
rect 1019 5256 1047 5886
rect 2575 5256 2603 5886
rect 319 4764 347 5004
rect 591 4764 619 5004
rect 1875 4764 1903 5004
rect 2147 4764 2175 5004
rect 3431 4764 3459 5004
rect 3703 4764 3731 5004
rect 4987 4764 5015 5004
rect 5259 4764 5287 5004
rect 6543 4764 6571 5004
rect 6815 4764 6843 5004
rect 8099 4764 8127 5004
rect 8371 4764 8399 5004
rect 9655 4764 9683 5004
rect 9927 4764 9955 5004
rect 11211 4764 11239 5004
rect 11483 4764 11511 5004
rect 12767 4764 12795 5004
rect 13039 4764 13067 5004
rect 14323 4764 14351 5004
rect 14595 4764 14623 5004
rect 15879 4764 15907 5004
rect 16151 4764 16179 5004
rect 17435 4764 17463 5004
rect 17707 4764 17735 5004
rect 18991 4764 19019 5004
rect 19263 4764 19291 5004
rect 20547 4764 20575 5004
rect 20819 4764 20847 5004
rect 22103 4764 22131 5004
rect 22375 4764 22403 5004
rect 23659 4764 23687 5004
rect 23931 4764 23959 5004
rect 84 1724 112 1794
rect 70 1696 112 1724
rect 70 504 98 1696
rect 694 1640 722 1794
rect 862 1724 890 1794
rect 532 1612 722 1640
rect 848 1696 890 1724
rect 532 504 560 1612
rect 848 504 876 1696
rect 1472 1640 1500 1794
rect 1640 1724 1668 1794
rect 1310 1612 1500 1640
rect 1626 1696 1668 1724
rect 1310 504 1338 1612
rect 1626 504 1654 1696
rect 2250 1640 2278 1794
rect 2418 1724 2446 1794
rect 2088 1612 2278 1640
rect 2404 1696 2446 1724
rect 2088 504 2116 1612
rect 2404 504 2432 1696
rect 3028 1640 3056 1794
rect 3196 1724 3224 1794
rect 2866 1612 3056 1640
rect 3182 1696 3224 1724
rect 2866 504 2894 1612
rect 3182 504 3210 1696
rect 3806 1640 3834 1794
rect 3974 1724 4002 1794
rect 3644 1612 3834 1640
rect 3960 1696 4002 1724
rect 3644 504 3672 1612
rect 3960 504 3988 1696
rect 4584 1640 4612 1794
rect 4752 1724 4780 1794
rect 4422 1612 4612 1640
rect 4738 1696 4780 1724
rect 4422 504 4450 1612
rect 4738 504 4766 1696
rect 5362 1640 5390 1794
rect 5530 1724 5558 1794
rect 5200 1612 5390 1640
rect 5516 1696 5558 1724
rect 5200 504 5228 1612
rect 5516 504 5544 1696
rect 6140 1640 6168 1794
rect 6308 1724 6336 1794
rect 5978 1612 6168 1640
rect 6294 1696 6336 1724
rect 5978 504 6006 1612
rect 6294 504 6322 1696
rect 6918 1640 6946 1794
rect 7086 1724 7114 1794
rect 6756 1612 6946 1640
rect 7072 1696 7114 1724
rect 6756 504 6784 1612
rect 7072 504 7100 1696
rect 7696 1640 7724 1794
rect 7864 1724 7892 1794
rect 7534 1612 7724 1640
rect 7850 1696 7892 1724
rect 7534 504 7562 1612
rect 7850 504 7878 1696
rect 8474 1640 8502 1794
rect 8642 1724 8670 1794
rect 8312 1612 8502 1640
rect 8628 1696 8670 1724
rect 8312 504 8340 1612
rect 8628 504 8656 1696
rect 9252 1640 9280 1794
rect 9420 1724 9448 1794
rect 9090 1612 9280 1640
rect 9406 1696 9448 1724
rect 9090 504 9118 1612
rect 9406 504 9434 1696
rect 10030 1640 10058 1794
rect 10198 1724 10226 1794
rect 9868 1612 10058 1640
rect 10184 1696 10226 1724
rect 9868 504 9896 1612
rect 10184 504 10212 1696
rect 10808 1640 10836 1794
rect 10976 1724 11004 1794
rect 10646 1612 10836 1640
rect 10962 1696 11004 1724
rect 10646 504 10674 1612
rect 10962 504 10990 1696
rect 11586 1640 11614 1794
rect 11754 1724 11782 1794
rect 11424 1612 11614 1640
rect 11740 1696 11782 1724
rect 11424 504 11452 1612
rect 11740 504 11768 1696
rect 12364 1640 12392 1794
rect 12532 1724 12560 1794
rect 12202 1612 12392 1640
rect 12518 1696 12560 1724
rect 12202 504 12230 1612
rect 12518 504 12546 1696
rect 13142 1640 13170 1794
rect 13310 1724 13338 1794
rect 12980 1612 13170 1640
rect 13296 1696 13338 1724
rect 12980 504 13008 1612
rect 13296 504 13324 1696
rect 13920 1640 13948 1794
rect 14088 1724 14116 1794
rect 13758 1612 13948 1640
rect 14074 1696 14116 1724
rect 13758 504 13786 1612
rect 14074 504 14102 1696
rect 14698 1640 14726 1794
rect 14866 1724 14894 1794
rect 14536 1612 14726 1640
rect 14852 1696 14894 1724
rect 14536 504 14564 1612
rect 14852 504 14880 1696
rect 15476 1640 15504 1794
rect 15644 1724 15672 1794
rect 15314 1612 15504 1640
rect 15630 1696 15672 1724
rect 15314 504 15342 1612
rect 15630 504 15658 1696
rect 16254 1640 16282 1794
rect 16422 1724 16450 1794
rect 16092 1612 16282 1640
rect 16408 1696 16450 1724
rect 16092 504 16120 1612
rect 16408 504 16436 1696
rect 17032 1640 17060 1794
rect 17200 1724 17228 1794
rect 16870 1612 17060 1640
rect 17186 1696 17228 1724
rect 16870 504 16898 1612
rect 17186 504 17214 1696
rect 17810 1640 17838 1794
rect 17978 1724 18006 1794
rect 17648 1612 17838 1640
rect 17964 1696 18006 1724
rect 17648 504 17676 1612
rect 17964 504 17992 1696
rect 18588 1640 18616 1794
rect 18756 1724 18784 1794
rect 18426 1612 18616 1640
rect 18742 1696 18784 1724
rect 18426 504 18454 1612
rect 18742 504 18770 1696
rect 19366 1640 19394 1794
rect 19534 1724 19562 1794
rect 19204 1612 19394 1640
rect 19520 1696 19562 1724
rect 19204 504 19232 1612
rect 19520 504 19548 1696
rect 20144 1640 20172 1794
rect 20312 1724 20340 1794
rect 19982 1612 20172 1640
rect 20298 1696 20340 1724
rect 19982 504 20010 1612
rect 20298 504 20326 1696
rect 20922 1640 20950 1794
rect 21090 1724 21118 1794
rect 20760 1612 20950 1640
rect 21076 1696 21118 1724
rect 20760 504 20788 1612
rect 21076 504 21104 1696
rect 21700 1640 21728 1794
rect 21868 1724 21896 1794
rect 21538 1612 21728 1640
rect 21854 1696 21896 1724
rect 21538 504 21566 1612
rect 21854 504 21882 1696
rect 22478 1640 22506 1794
rect 22646 1724 22674 1794
rect 22316 1612 22506 1640
rect 22632 1696 22674 1724
rect 22316 504 22344 1612
rect 22632 504 22660 1696
rect 23256 1640 23284 1794
rect 23424 1724 23452 1794
rect 23094 1612 23284 1640
rect 23410 1696 23452 1724
rect 23094 504 23122 1612
rect 23410 504 23438 1696
rect 24034 1640 24062 1794
rect 24202 1724 24230 1794
rect 23872 1612 24062 1640
rect 24188 1696 24230 1724
rect 23872 504 23900 1612
rect 24188 504 24216 1696
rect 24812 1640 24840 1794
rect 24980 1724 25008 1794
rect 24650 1612 24840 1640
rect 24966 1696 25008 1724
rect 24650 504 24678 1612
rect 24966 504 24994 1696
rect 25590 1640 25618 1794
rect 25758 1724 25786 1794
rect 25428 1612 25618 1640
rect 25744 1696 25786 1724
rect 25428 504 25456 1612
rect 25744 504 25772 1696
rect 26368 1640 26396 1794
rect 26536 1724 26564 1794
rect 26206 1612 26396 1640
rect 26522 1696 26564 1724
rect 26206 504 26234 1612
rect 26522 504 26550 1696
rect 27146 1640 27174 1794
rect 27314 1724 27342 1794
rect 26984 1612 27174 1640
rect 27300 1696 27342 1724
rect 26984 504 27012 1612
rect 27300 504 27328 1696
rect 27924 1640 27952 1794
rect 28092 1724 28120 1794
rect 27762 1612 27952 1640
rect 28078 1696 28120 1724
rect 27762 504 27790 1612
rect 28078 504 28106 1696
rect 28702 1640 28730 1794
rect 28870 1724 28898 1794
rect 28540 1612 28730 1640
rect 28856 1696 28898 1724
rect 28540 504 28568 1612
rect 28856 504 28884 1696
rect 29480 1640 29508 1794
rect 29648 1724 29676 1794
rect 29318 1612 29508 1640
rect 29634 1696 29676 1724
rect 29318 504 29346 1612
rect 29634 504 29662 1696
rect 30258 1640 30286 1794
rect 30426 1724 30454 1794
rect 30096 1612 30286 1640
rect 30412 1696 30454 1724
rect 30096 504 30124 1612
rect 30412 504 30440 1696
rect 31036 1640 31064 1794
rect 31204 1724 31232 1794
rect 30874 1612 31064 1640
rect 31190 1696 31232 1724
rect 30874 504 30902 1612
rect 31190 504 31218 1696
rect 31814 1640 31842 1794
rect 31982 1724 32010 1794
rect 31652 1612 31842 1640
rect 31968 1696 32010 1724
rect 31652 504 31680 1612
rect 31968 504 31996 1696
rect 32592 1640 32620 1794
rect 32760 1724 32788 1794
rect 32430 1612 32620 1640
rect 32746 1696 32788 1724
rect 32430 504 32458 1612
rect 32746 504 32774 1696
rect 33370 1640 33398 1794
rect 33538 1724 33566 1794
rect 33208 1612 33398 1640
rect 33524 1696 33566 1724
rect 33208 504 33236 1612
rect 33524 504 33552 1696
rect 34148 1640 34176 1794
rect 34316 1724 34344 1794
rect 33986 1612 34176 1640
rect 34302 1696 34344 1724
rect 33986 504 34014 1612
rect 34302 504 34330 1696
rect 34926 1640 34954 1794
rect 35094 1724 35122 1794
rect 34764 1612 34954 1640
rect 35080 1696 35122 1724
rect 34764 504 34792 1612
rect 35080 504 35108 1696
rect 35704 1640 35732 1794
rect 35872 1724 35900 1794
rect 35542 1612 35732 1640
rect 35858 1696 35900 1724
rect 35542 504 35570 1612
rect 35858 504 35886 1696
rect 36482 1640 36510 1794
rect 36650 1724 36678 1794
rect 36320 1612 36510 1640
rect 36636 1696 36678 1724
rect 36320 504 36348 1612
rect 36636 504 36664 1696
rect 37260 1640 37288 1794
rect 37428 1724 37456 1794
rect 37098 1612 37288 1640
rect 37414 1696 37456 1724
rect 37098 504 37126 1612
rect 37414 504 37442 1696
rect 38038 1640 38066 1794
rect 38206 1724 38234 1794
rect 37876 1612 38066 1640
rect 38192 1696 38234 1724
rect 37876 504 37904 1612
rect 38192 504 38220 1696
rect 38816 1640 38844 1794
rect 38984 1724 39012 1794
rect 38654 1612 38844 1640
rect 38970 1696 39012 1724
rect 38654 504 38682 1612
rect 38970 504 38998 1696
rect 39594 1640 39622 1794
rect 39762 1724 39790 1794
rect 39432 1612 39622 1640
rect 39748 1696 39790 1724
rect 39432 504 39460 1612
rect 39748 504 39776 1696
rect 40372 1640 40400 1794
rect 40540 1724 40568 1794
rect 40210 1612 40400 1640
rect 40526 1696 40568 1724
rect 40210 504 40238 1612
rect 40526 504 40554 1696
rect 41150 1640 41178 1794
rect 41318 1724 41346 1794
rect 40988 1612 41178 1640
rect 41304 1696 41346 1724
rect 40988 504 41016 1612
rect 41304 504 41332 1696
rect 41928 1640 41956 1794
rect 42096 1724 42124 1794
rect 41766 1612 41956 1640
rect 42082 1696 42124 1724
rect 41766 504 41794 1612
rect 42082 504 42110 1696
rect 42706 1640 42734 1794
rect 42874 1724 42902 1794
rect 42544 1612 42734 1640
rect 42860 1696 42902 1724
rect 42544 504 42572 1612
rect 42860 504 42888 1696
rect 43484 1640 43512 1794
rect 43652 1724 43680 1794
rect 43322 1612 43512 1640
rect 43638 1696 43680 1724
rect 43322 504 43350 1612
rect 43638 504 43666 1696
rect 44262 1640 44290 1794
rect 44430 1724 44458 1794
rect 44100 1612 44290 1640
rect 44416 1696 44458 1724
rect 44100 504 44128 1612
rect 44416 504 44444 1696
rect 45040 1640 45068 1794
rect 45208 1724 45236 1794
rect 44878 1612 45068 1640
rect 45194 1696 45236 1724
rect 44878 504 44906 1612
rect 45194 504 45222 1696
rect 45818 1640 45846 1794
rect 45986 1724 46014 1794
rect 45656 1612 45846 1640
rect 45972 1696 46014 1724
rect 45656 504 45684 1612
rect 45972 504 46000 1696
rect 46596 1640 46624 1794
rect 46764 1724 46792 1794
rect 46434 1612 46624 1640
rect 46750 1696 46792 1724
rect 46434 504 46462 1612
rect 46750 504 46778 1696
rect 47374 1640 47402 1794
rect 47542 1724 47570 1794
rect 47212 1612 47402 1640
rect 47528 1696 47570 1724
rect 47212 504 47240 1612
rect 47528 504 47556 1696
rect 48152 1640 48180 1794
rect 48320 1724 48348 1794
rect 47990 1612 48180 1640
rect 48306 1696 48348 1724
rect 47990 504 48018 1612
rect 48306 504 48334 1696
rect 48930 1640 48958 1794
rect 49098 1724 49126 1794
rect 48768 1612 48958 1640
rect 49084 1696 49126 1724
rect 48768 504 48796 1612
rect 49084 504 49112 1696
rect 49708 1640 49736 1794
rect 49546 1612 49736 1640
rect 49546 504 49574 1612
<< metal3 >>
rect 705 6100 771 6232
rect 2261 6100 2327 6232
rect 3817 6100 3883 6232
rect 5373 6100 5439 6232
rect 6929 6100 6995 6232
rect 8485 6100 8551 6232
rect 10041 6100 10107 6232
rect 11597 6100 11663 6232
rect 13153 6100 13219 6232
rect 14709 6100 14775 6232
rect 16265 6100 16331 6232
rect 17821 6100 17887 6232
rect 19377 6100 19443 6232
rect 20933 6100 20999 6232
rect 22489 6100 22555 6232
rect 24045 6100 24111 6232
rect 25601 6100 25667 6232
rect 27157 6100 27223 6232
rect 28713 6100 28779 6232
rect 30269 6100 30335 6232
rect 31825 6100 31891 6232
rect 33381 6100 33447 6232
rect 34937 6100 35003 6232
rect 36493 6100 36559 6232
rect 38049 6100 38115 6232
rect 39605 6100 39671 6232
rect 41161 6100 41227 6232
rect 42717 6100 42783 6232
rect 44273 6100 44339 6232
rect 45829 6100 45895 6232
rect 47385 6100 47451 6232
rect 48941 6100 49007 6232
rect 705 5268 771 5400
rect 2261 5268 2327 5400
rect 3817 5268 3883 5400
rect 5373 5268 5439 5400
rect 6929 5268 6995 5400
rect 8485 5268 8551 5400
rect 10041 5268 10107 5400
rect 11597 5268 11663 5400
rect 13153 5268 13219 5400
rect 14709 5268 14775 5400
rect 16265 5268 16331 5400
rect 17821 5268 17887 5400
rect 19377 5268 19443 5400
rect 20933 5268 20999 5400
rect 22489 5268 22555 5400
rect 24045 5268 24111 5400
rect 25601 5268 25667 5400
rect 27157 5268 27223 5400
rect 28713 5268 28779 5400
rect 30269 5268 30335 5400
rect 31825 5268 31891 5400
rect 33381 5268 33447 5400
rect 34937 5268 35003 5400
rect 36493 5268 36559 5400
rect 38049 5268 38115 5400
rect 39605 5268 39671 5400
rect 41161 5268 41227 5400
rect 42717 5268 42783 5400
rect 44273 5268 44339 5400
rect 45829 5268 45895 5400
rect 47385 5268 47451 5400
rect 48941 5268 49007 5400
rect 187 4933 319 5007
rect 459 4933 591 5007
rect 1743 4933 1875 5007
rect 2015 4933 2147 5007
rect 3299 4933 3431 5007
rect 3571 4933 3703 5007
rect 4855 4933 4987 5007
rect 5127 4933 5259 5007
rect 6411 4933 6543 5007
rect 6683 4933 6815 5007
rect 7967 4933 8099 5007
rect 8239 4933 8371 5007
rect 9523 4933 9655 5007
rect 9795 4933 9927 5007
rect 11079 4933 11211 5007
rect 11351 4933 11483 5007
rect 12635 4933 12767 5007
rect 12907 4933 13039 5007
rect 14191 4933 14323 5007
rect 14463 4933 14595 5007
rect 15747 4933 15879 5007
rect 16019 4933 16151 5007
rect 17303 4933 17435 5007
rect 17575 4933 17707 5007
rect 18859 4933 18991 5007
rect 19131 4933 19263 5007
rect 20415 4933 20547 5007
rect 20687 4933 20819 5007
rect 21971 4933 22103 5007
rect 22243 4933 22375 5007
rect 23527 4933 23659 5007
rect 23799 4933 23931 5007
rect 25083 4933 25215 5007
rect 25355 4933 25487 5007
rect 26639 4933 26771 5007
rect 26911 4933 27043 5007
rect 28195 4933 28327 5007
rect 28467 4933 28599 5007
rect 29751 4933 29883 5007
rect 30023 4933 30155 5007
rect 31307 4933 31439 5007
rect 31579 4933 31711 5007
rect 32863 4933 32995 5007
rect 33135 4933 33267 5007
rect 34419 4933 34551 5007
rect 34691 4933 34823 5007
rect 35975 4933 36107 5007
rect 36247 4933 36379 5007
rect 37531 4933 37663 5007
rect 37803 4933 37935 5007
rect 39087 4933 39219 5007
rect 39359 4933 39491 5007
rect 40643 4933 40775 5007
rect 40915 4933 41047 5007
rect 42199 4933 42331 5007
rect 42471 4933 42603 5007
rect 43755 4933 43887 5007
rect 44027 4933 44159 5007
rect 45311 4933 45443 5007
rect 45583 4933 45715 5007
rect 46867 4933 46999 5007
rect 47139 4933 47271 5007
rect 48423 4933 48555 5007
rect 48695 4933 48827 5007
rect 187 3987 319 4061
rect 459 3987 591 4061
rect 1743 3987 1875 4061
rect 2015 3987 2147 4061
rect 3299 3987 3431 4061
rect 3571 3987 3703 4061
rect 4855 3987 4987 4061
rect 5127 3987 5259 4061
rect 6411 3987 6543 4061
rect 6683 3987 6815 4061
rect 7967 3987 8099 4061
rect 8239 3987 8371 4061
rect 9523 3987 9655 4061
rect 9795 3987 9927 4061
rect 11079 3987 11211 4061
rect 11351 3987 11483 4061
rect 12635 3987 12767 4061
rect 12907 3987 13039 4061
rect 14191 3987 14323 4061
rect 14463 3987 14595 4061
rect 15747 3987 15879 4061
rect 16019 3987 16151 4061
rect 17303 3987 17435 4061
rect 17575 3987 17707 4061
rect 18859 3987 18991 4061
rect 19131 3987 19263 4061
rect 20415 3987 20547 4061
rect 20687 3987 20819 4061
rect 21971 3987 22103 4061
rect 22243 3987 22375 4061
rect 23527 3987 23659 4061
rect 23799 3987 23931 4061
rect 25083 3987 25215 4061
rect 25355 3987 25487 4061
rect 26639 3987 26771 4061
rect 26911 3987 27043 4061
rect 28195 3987 28327 4061
rect 28467 3987 28599 4061
rect 29751 3987 29883 4061
rect 30023 3987 30155 4061
rect 31307 3987 31439 4061
rect 31579 3987 31711 4061
rect 32863 3987 32995 4061
rect 33135 3987 33267 4061
rect 34419 3987 34551 4061
rect 34691 3987 34823 4061
rect 35975 3987 36107 4061
rect 36247 3987 36379 4061
rect 37531 3987 37663 4061
rect 37803 3987 37935 4061
rect 39087 3987 39219 4061
rect 39359 3987 39491 4061
rect 40643 3987 40775 4061
rect 40915 3987 41047 4061
rect 42199 3987 42331 4061
rect 42471 3987 42603 4061
rect 43755 3987 43887 4061
rect 44027 3987 44159 4061
rect 45311 3987 45443 4061
rect 45583 3987 45715 4061
rect 46867 3987 46999 4061
rect 47139 3987 47271 4061
rect 48423 3987 48555 4061
rect 48695 3987 48827 4061
rect 712 2506 844 2580
rect 1490 2506 1622 2580
rect 2268 2506 2400 2580
rect 3046 2506 3178 2580
rect 3824 2506 3956 2580
rect 4602 2506 4734 2580
rect 5380 2506 5512 2580
rect 6158 2506 6290 2580
rect 6936 2506 7068 2580
rect 7714 2506 7846 2580
rect 8492 2506 8624 2580
rect 9270 2506 9402 2580
rect 10048 2506 10180 2580
rect 10826 2506 10958 2580
rect 11604 2506 11736 2580
rect 12382 2506 12514 2580
rect 13160 2506 13292 2580
rect 13938 2506 14070 2580
rect 14716 2506 14848 2580
rect 15494 2506 15626 2580
rect 16272 2506 16404 2580
rect 17050 2506 17182 2580
rect 17828 2506 17960 2580
rect 18606 2506 18738 2580
rect 19384 2506 19516 2580
rect 20162 2506 20294 2580
rect 20940 2506 21072 2580
rect 21718 2506 21850 2580
rect 22496 2506 22628 2580
rect 23274 2506 23406 2580
rect 24052 2506 24184 2580
rect 24830 2506 24962 2580
rect 25608 2506 25740 2580
rect 26386 2506 26518 2580
rect 27164 2506 27296 2580
rect 27942 2506 28074 2580
rect 28720 2506 28852 2580
rect 29498 2506 29630 2580
rect 30276 2506 30408 2580
rect 31054 2506 31186 2580
rect 31832 2506 31964 2580
rect 32610 2506 32742 2580
rect 33388 2506 33520 2580
rect 34166 2506 34298 2580
rect 34944 2506 35076 2580
rect 35722 2506 35854 2580
rect 36500 2506 36632 2580
rect 37278 2506 37410 2580
rect 38056 2506 38188 2580
rect 38834 2506 38966 2580
rect 39612 2506 39744 2580
rect 40390 2506 40522 2580
rect 41168 2506 41300 2580
rect 41946 2506 42078 2580
rect 42724 2506 42856 2580
rect 43502 2506 43634 2580
rect 44280 2506 44412 2580
rect 45058 2506 45190 2580
rect 45836 2506 45968 2580
rect 46614 2506 46746 2580
rect 47392 2506 47524 2580
rect 48170 2506 48302 2580
rect 48948 2506 49080 2580
rect 49726 2506 49858 2580
rect 160 548 226 680
rect 938 548 1004 680
rect 1716 548 1782 680
rect 2494 548 2560 680
rect 3272 548 3338 680
rect 4050 548 4116 680
rect 4828 548 4894 680
rect 5606 548 5672 680
rect 6384 548 6450 680
rect 7162 548 7228 680
rect 7940 548 8006 680
rect 8718 548 8784 680
rect 9496 548 9562 680
rect 10274 548 10340 680
rect 11052 548 11118 680
rect 11830 548 11896 680
rect 12608 548 12674 680
rect 13386 548 13452 680
rect 14164 548 14230 680
rect 14942 548 15008 680
rect 15720 548 15786 680
rect 16498 548 16564 680
rect 17276 548 17342 680
rect 18054 548 18120 680
rect 18832 548 18898 680
rect 19610 548 19676 680
rect 20388 548 20454 680
rect 21166 548 21232 680
rect 21944 548 22010 680
rect 22722 548 22788 680
rect 23500 548 23566 680
rect 24278 548 24344 680
rect 25056 548 25122 680
rect 25834 548 25900 680
rect 26612 548 26678 680
rect 27390 548 27456 680
rect 28168 548 28234 680
rect 28946 548 29012 680
rect 29724 548 29790 680
rect 30502 548 30568 680
rect 31280 548 31346 680
rect 32058 548 32124 680
rect 32836 548 32902 680
rect 33614 548 33680 680
rect 34392 548 34458 680
rect 35170 548 35236 680
rect 35948 548 36014 680
rect 36726 548 36792 680
rect 37504 548 37570 680
rect 38282 548 38348 680
rect 39060 548 39126 680
rect 39838 548 39904 680
rect 40616 548 40682 680
rect 41394 548 41460 680
rect 42172 548 42238 680
rect 42950 548 43016 680
rect 43728 548 43794 680
rect 44506 548 44572 680
rect 45284 548 45350 680
rect 46062 548 46128 680
rect 46840 548 46906 680
rect 47618 548 47684 680
rect 48396 548 48462 680
rect 49174 548 49240 680
rect 49952 548 50018 680
use column_mux_array_multiport  column_mux_array_multiport_0
timestamp 1644969367
transform 1 0 0 0 -1 3702
box 0 48 49858 1908
use write_driver_array  write_driver_array_0
timestamp 1644969367
transform 1 0 0 0 -1 6208
box 0 -24 49323 952
use sense_amp_array  sense_amp_array_0
timestamp 1644969367
transform 1 0 0 0 -1 5004
box 117 -3 48897 1050
use precharge_array_multiport  precharge_array_multiport_0
timestamp 1644969367
transform 1 0 0 0 -1 1542
box 0 -8 50570 1052
<< labels >>
rlabel metal2 s 584 5908 638 5936 4 din0_0
rlabel metal2 s 2140 5908 2194 5936 4 din0_1
rlabel metal2 s 3696 5908 3750 5936 4 din0_2
rlabel metal2 s 5252 5908 5306 5936 4 din0_3
rlabel metal2 s 6808 5908 6862 5936 4 din0_4
rlabel metal2 s 8364 5908 8418 5936 4 din0_5
rlabel metal2 s 9920 5908 9974 5936 4 din0_6
rlabel metal2 s 11476 5908 11530 5936 4 din0_7
rlabel metal2 s 13032 5908 13086 5936 4 din0_8
rlabel metal2 s 14588 5908 14642 5936 4 din0_9
rlabel metal2 s 16144 5908 16198 5936 4 din0_10
rlabel metal2 s 17700 5908 17754 5936 4 din0_11
rlabel metal2 s 19256 5908 19310 5936 4 din0_12
rlabel metal2 s 20812 5908 20866 5936 4 din0_13
rlabel metal2 s 22368 5908 22422 5936 4 din0_14
rlabel metal2 s 23924 5908 23978 5936 4 din0_15
rlabel metal2 s 25480 5908 25534 5936 4 din0_16
rlabel metal2 s 27036 5908 27090 5936 4 din0_17
rlabel metal2 s 28592 5908 28646 5936 4 din0_18
rlabel metal2 s 30148 5908 30202 5936 4 din0_19
rlabel metal2 s 31704 5908 31758 5936 4 din0_20
rlabel metal2 s 33260 5908 33314 5936 4 din0_21
rlabel metal2 s 34816 5908 34870 5936 4 din0_22
rlabel metal2 s 36372 5908 36426 5936 4 din0_23
rlabel metal2 s 37928 5908 37982 5936 4 din0_24
rlabel metal2 s 39484 5908 39538 5936 4 din0_25
rlabel metal2 s 41040 5908 41094 5936 4 din0_26
rlabel metal2 s 42596 5908 42650 5936 4 din0_27
rlabel metal2 s 44152 5908 44206 5936 4 din0_28
rlabel metal2 s 45708 5908 45762 5936 4 din0_29
rlabel metal2 s 47264 5908 47318 5936 4 din0_30
rlabel metal2 s 48820 5908 48874 5936 4 din0_31
rlabel metal2 s 318 4764 346 5004 4 dout0_0
rlabel metal2 s 333 4884 333 4884 4 dout1_0
rlabel metal2 s 590 4764 618 5004 4 dout0_1
rlabel metal2 s 605 4884 605 4884 4 dout1_1
rlabel metal2 s 1874 4764 1902 5004 4 dout0_2
rlabel metal2 s 1889 4884 1889 4884 4 dout1_2
rlabel metal2 s 2146 4764 2174 5004 4 dout0_3
rlabel metal2 s 2161 4884 2161 4884 4 dout1_3
rlabel metal2 s 3430 4764 3458 5004 4 dout0_4
rlabel metal2 s 3445 4884 3445 4884 4 dout1_4
rlabel metal2 s 3702 4764 3730 5004 4 dout0_5
rlabel metal2 s 3717 4884 3717 4884 4 dout1_5
rlabel metal2 s 4986 4764 5014 5004 4 dout0_6
rlabel metal2 s 5001 4884 5001 4884 4 dout1_6
rlabel metal2 s 5258 4764 5286 5004 4 dout0_7
rlabel metal2 s 5273 4884 5273 4884 4 dout1_7
rlabel metal2 s 6542 4764 6570 5004 4 dout0_8
rlabel metal2 s 6557 4884 6557 4884 4 dout1_8
rlabel metal2 s 6814 4764 6842 5004 4 dout0_9
rlabel metal2 s 6829 4884 6829 4884 4 dout1_9
rlabel metal2 s 8098 4764 8126 5004 4 dout0_10
rlabel metal2 s 8113 4884 8113 4884 4 dout1_10
rlabel metal2 s 8370 4764 8398 5004 4 dout0_11
rlabel metal2 s 8385 4884 8385 4884 4 dout1_11
rlabel metal2 s 9654 4764 9682 5004 4 dout0_12
rlabel metal2 s 9669 4884 9669 4884 4 dout1_12
rlabel metal2 s 9926 4764 9954 5004 4 dout0_13
rlabel metal2 s 9941 4884 9941 4884 4 dout1_13
rlabel metal2 s 11210 4764 11238 5004 4 dout0_14
rlabel metal2 s 11225 4884 11225 4884 4 dout1_14
rlabel metal2 s 11482 4764 11510 5004 4 dout0_15
rlabel metal2 s 11497 4884 11497 4884 4 dout1_15
rlabel metal2 s 12766 4764 12794 5004 4 dout0_16
rlabel metal2 s 12781 4884 12781 4884 4 dout1_16
rlabel metal2 s 13038 4764 13066 5004 4 dout0_17
rlabel metal2 s 13053 4884 13053 4884 4 dout1_17
rlabel metal2 s 14322 4764 14350 5004 4 dout0_18
rlabel metal2 s 14337 4884 14337 4884 4 dout1_18
rlabel metal2 s 14594 4764 14622 5004 4 dout0_19
rlabel metal2 s 14609 4884 14609 4884 4 dout1_19
rlabel metal2 s 15878 4764 15906 5004 4 dout0_20
rlabel metal2 s 15893 4884 15893 4884 4 dout1_20
rlabel metal2 s 16150 4764 16178 5004 4 dout0_21
rlabel metal2 s 16165 4884 16165 4884 4 dout1_21
rlabel metal2 s 17434 4764 17462 5004 4 dout0_22
rlabel metal2 s 17449 4884 17449 4884 4 dout1_22
rlabel metal2 s 17706 4764 17734 5004 4 dout0_23
rlabel metal2 s 17721 4884 17721 4884 4 dout1_23
rlabel metal2 s 18990 4764 19018 5004 4 dout0_24
rlabel metal2 s 19005 4884 19005 4884 4 dout1_24
rlabel metal2 s 19262 4764 19290 5004 4 dout0_25
rlabel metal2 s 19277 4884 19277 4884 4 dout1_25
rlabel metal2 s 20546 4764 20574 5004 4 dout0_26
rlabel metal2 s 20561 4884 20561 4884 4 dout1_26
rlabel metal2 s 20818 4764 20846 5004 4 dout0_27
rlabel metal2 s 20833 4884 20833 4884 4 dout1_27
rlabel metal2 s 22102 4764 22130 5004 4 dout0_28
rlabel metal2 s 22117 4884 22117 4884 4 dout1_28
rlabel metal2 s 22374 4764 22402 5004 4 dout0_29
rlabel metal2 s 22389 4884 22389 4884 4 dout1_29
rlabel metal2 s 23658 4764 23686 5004 4 dout0_30
rlabel metal2 s 23673 4884 23673 4884 4 dout1_30
rlabel metal2 s 23930 4764 23958 5004 4 dout0_31
rlabel metal2 s 23945 4884 23945 4884 4 dout1_31
rlabel metal2 s 70 504 98 1542 4 rbl0_0
rlabel metal2 s 532 504 560 1542 4 rbl1_0
rlabel metal2 s 848 504 876 1542 4 rbl0_1
rlabel metal2 s 1310 504 1338 1542 4 rbl1_1
rlabel metal2 s 1626 504 1654 1542 4 rbl0_2
rlabel metal2 s 2088 504 2116 1542 4 rbl1_2
rlabel metal2 s 2404 504 2432 1542 4 rbl0_3
rlabel metal2 s 2866 504 2894 1542 4 rbl1_3
rlabel metal2 s 3182 504 3210 1542 4 rbl0_4
rlabel metal2 s 3644 504 3672 1542 4 rbl1_4
rlabel metal2 s 3960 504 3988 1542 4 rbl0_5
rlabel metal2 s 4422 504 4450 1542 4 rbl1_5
rlabel metal2 s 4738 504 4766 1542 4 rbl0_6
rlabel metal2 s 5200 504 5228 1542 4 rbl1_6
rlabel metal2 s 5516 504 5544 1542 4 rbl0_7
rlabel metal2 s 5978 504 6006 1542 4 rbl1_7
rlabel metal2 s 6294 504 6322 1542 4 rbl0_8
rlabel metal2 s 6756 504 6784 1542 4 rbl1_8
rlabel metal2 s 7072 504 7100 1542 4 rbl0_9
rlabel metal2 s 7534 504 7562 1542 4 rbl1_9
rlabel metal2 s 7850 504 7878 1542 4 rbl0_10
rlabel metal2 s 8312 504 8340 1542 4 rbl1_10
rlabel metal2 s 8628 504 8656 1542 4 rbl0_11
rlabel metal2 s 9090 504 9118 1542 4 rbl1_11
rlabel metal2 s 9406 504 9434 1542 4 rbl0_12
rlabel metal2 s 9868 504 9896 1542 4 rbl1_12
rlabel metal2 s 10184 504 10212 1542 4 rbl0_13
rlabel metal2 s 10646 504 10674 1542 4 rbl1_13
rlabel metal2 s 10962 504 10990 1542 4 rbl0_14
rlabel metal2 s 11424 504 11452 1542 4 rbl1_14
rlabel metal2 s 11740 504 11768 1542 4 rbl0_15
rlabel metal2 s 12202 504 12230 1542 4 rbl1_15
rlabel metal2 s 12518 504 12546 1542 4 rbl0_16
rlabel metal2 s 12980 504 13008 1542 4 rbl1_16
rlabel metal2 s 13296 504 13324 1542 4 rbl0_17
rlabel metal2 s 13758 504 13786 1542 4 rbl1_17
rlabel metal2 s 14074 504 14102 1542 4 rbl0_18
rlabel metal2 s 14536 504 14564 1542 4 rbl1_18
rlabel metal2 s 14852 504 14880 1542 4 rbl0_19
rlabel metal2 s 15314 504 15342 1542 4 rbl1_19
rlabel metal2 s 15630 504 15658 1542 4 rbl0_20
rlabel metal2 s 16092 504 16120 1542 4 rbl1_20
rlabel metal2 s 16408 504 16436 1542 4 rbl0_21
rlabel metal2 s 16870 504 16898 1542 4 rbl1_21
rlabel metal2 s 17186 504 17214 1542 4 rbl0_22
rlabel metal2 s 17648 504 17676 1542 4 rbl1_22
rlabel metal2 s 17964 504 17992 1542 4 rbl0_23
rlabel metal2 s 18426 504 18454 1542 4 rbl1_23
rlabel metal2 s 18742 504 18770 1542 4 rbl0_24
rlabel metal2 s 19204 504 19232 1542 4 rbl1_24
rlabel metal2 s 19520 504 19548 1542 4 rbl0_25
rlabel metal2 s 19982 504 20010 1542 4 rbl1_25
rlabel metal2 s 20298 504 20326 1542 4 rbl0_26
rlabel metal2 s 20760 504 20788 1542 4 rbl1_26
rlabel metal2 s 21076 504 21104 1542 4 rbl0_27
rlabel metal2 s 21538 504 21566 1542 4 rbl1_27
rlabel metal2 s 21854 504 21882 1542 4 rbl0_28
rlabel metal2 s 22316 504 22344 1542 4 rbl1_28
rlabel metal2 s 22632 504 22660 1542 4 rbl0_29
rlabel metal2 s 23094 504 23122 1542 4 rbl1_29
rlabel metal2 s 23410 504 23438 1542 4 rbl0_30
rlabel metal2 s 23872 504 23900 1542 4 rbl1_30
rlabel metal2 s 24188 504 24216 1542 4 rbl0_31
rlabel metal2 s 24650 504 24678 1542 4 rbl1_31
rlabel metal2 s 24966 504 24994 1542 4 rbl0_32
rlabel metal2 s 25428 504 25456 1542 4 rbl1_32
rlabel metal2 s 25744 504 25772 1542 4 rbl0_33
rlabel metal2 s 26206 504 26234 1542 4 rbl1_33
rlabel metal2 s 26522 504 26550 1542 4 rbl0_34
rlabel metal2 s 26984 504 27012 1542 4 rbl1_34
rlabel metal2 s 27300 504 27328 1542 4 rbl0_35
rlabel metal2 s 27762 504 27790 1542 4 rbl1_35
rlabel metal2 s 28078 504 28106 1542 4 rbl0_36
rlabel metal2 s 28540 504 28568 1542 4 rbl1_36
rlabel metal2 s 28856 504 28884 1542 4 rbl0_37
rlabel metal2 s 29318 504 29346 1542 4 rbl1_37
rlabel metal2 s 29634 504 29662 1542 4 rbl0_38
rlabel metal2 s 30096 504 30124 1542 4 rbl1_38
rlabel metal2 s 30412 504 30440 1542 4 rbl0_39
rlabel metal2 s 30874 504 30902 1542 4 rbl1_39
rlabel metal2 s 31190 504 31218 1542 4 rbl0_40
rlabel metal2 s 31652 504 31680 1542 4 rbl1_40
rlabel metal2 s 31968 504 31996 1542 4 rbl0_41
rlabel metal2 s 32430 504 32458 1542 4 rbl1_41
rlabel metal2 s 32746 504 32774 1542 4 rbl0_42
rlabel metal2 s 33208 504 33236 1542 4 rbl1_42
rlabel metal2 s 33524 504 33552 1542 4 rbl0_43
rlabel metal2 s 33986 504 34014 1542 4 rbl1_43
rlabel metal2 s 34302 504 34330 1542 4 rbl0_44
rlabel metal2 s 34764 504 34792 1542 4 rbl1_44
rlabel metal2 s 35080 504 35108 1542 4 rbl0_45
rlabel metal2 s 35542 504 35570 1542 4 rbl1_45
rlabel metal2 s 35858 504 35886 1542 4 rbl0_46
rlabel metal2 s 36320 504 36348 1542 4 rbl1_46
rlabel metal2 s 36636 504 36664 1542 4 rbl0_47
rlabel metal2 s 37098 504 37126 1542 4 rbl1_47
rlabel metal2 s 37414 504 37442 1542 4 rbl0_48
rlabel metal2 s 37876 504 37904 1542 4 rbl1_48
rlabel metal2 s 38192 504 38220 1542 4 rbl0_49
rlabel metal2 s 38654 504 38682 1542 4 rbl1_49
rlabel metal2 s 38970 504 38998 1542 4 rbl0_50
rlabel metal2 s 39432 504 39460 1542 4 rbl1_50
rlabel metal2 s 39748 504 39776 1542 4 rbl0_51
rlabel metal2 s 40210 504 40238 1542 4 rbl1_51
rlabel metal2 s 40526 504 40554 1542 4 rbl0_52
rlabel metal2 s 40988 504 41016 1542 4 rbl1_52
rlabel metal2 s 41304 504 41332 1542 4 rbl0_53
rlabel metal2 s 41766 504 41794 1542 4 rbl1_53
rlabel metal2 s 42082 504 42110 1542 4 rbl0_54
rlabel metal2 s 42544 504 42572 1542 4 rbl1_54
rlabel metal2 s 42860 504 42888 1542 4 rbl0_55
rlabel metal2 s 43322 504 43350 1542 4 rbl1_55
rlabel metal2 s 43638 504 43666 1542 4 rbl0_56
rlabel metal2 s 44100 504 44128 1542 4 rbl1_56
rlabel metal2 s 44416 504 44444 1542 4 rbl0_57
rlabel metal2 s 44878 504 44906 1542 4 rbl1_57
rlabel metal2 s 45194 504 45222 1542 4 rbl0_58
rlabel metal2 s 45656 504 45684 1542 4 rbl1_58
rlabel metal2 s 45972 504 46000 1542 4 rbl0_59
rlabel metal2 s 46434 504 46462 1542 4 rbl1_59
rlabel metal2 s 46750 504 46778 1542 4 rbl0_60
rlabel metal2 s 47212 504 47240 1542 4 rbl1_60
rlabel metal2 s 47528 504 47556 1542 4 rbl0_61
rlabel metal2 s 47990 504 48018 1542 4 rbl1_61
rlabel metal2 s 48306 504 48334 1542 4 rbl0_62
rlabel metal2 s 48768 504 48796 1542 4 rbl1_62
rlabel metal2 s 49084 504 49112 1542 4 rbl0_63
rlabel metal2 s 49546 504 49574 1542 4 rbl1_63
rlabel metal2 s 1018 5256 1046 5886 4 wbl0_0
rlabel metal2 s 2574 5256 2602 5886 4 wbl0_1
rlabel metal1 s 0 1502 50570 1530 4 p_en_bar
rlabel metal1 s 0 3434 49792 3462 4 sel_0
rlabel metal1 s 0 3354 49792 3382 4 sel_1
rlabel metal1 s 0 5824 49322 5852 4 w_en
rlabel metal3 s 30022 3986 30154 4060 4 vdd
rlabel metal3 s 10274 548 10340 680 4 vdd
rlabel metal3 s 12634 3986 12766 4060 4 vdd
rlabel metal3 s 32862 3986 32994 4060 4 vdd
rlabel metal3 s 23526 3986 23658 4060 4 vdd
rlabel metal3 s 27390 548 27456 680 4 vdd
rlabel metal3 s 30268 5268 30334 5400 4 vdd
rlabel metal3 s 9522 3986 9654 4060 4 vdd
rlabel metal3 s 6682 3986 6814 4060 4 vdd
rlabel metal3 s 36492 5268 36558 5400 4 vdd
rlabel metal3 s 1716 548 1782 680 4 vdd
rlabel metal3 s 25082 3986 25214 4060 4 vdd
rlabel metal3 s 47384 5268 47450 5400 4 vdd
rlabel metal3 s 14190 3986 14322 4060 4 vdd
rlabel metal3 s 47138 3986 47270 4060 4 vdd
rlabel metal3 s 13152 5268 13218 5400 4 vdd
rlabel metal3 s 14942 548 15008 680 4 vdd
rlabel metal3 s 7162 548 7228 680 4 vdd
rlabel metal3 s 5606 548 5672 680 4 vdd
rlabel metal3 s 16264 5268 16330 5400 4 vdd
rlabel metal3 s 20932 5268 20998 5400 4 vdd
rlabel metal3 s 39060 548 39126 680 4 vdd
rlabel metal3 s 30502 548 30568 680 4 vdd
rlabel metal3 s 15720 548 15786 680 4 vdd
rlabel metal3 s 16018 3986 16150 4060 4 vdd
rlabel metal3 s 31824 5268 31890 5400 4 vdd
rlabel metal3 s 4050 548 4116 680 4 vdd
rlabel metal3 s 17276 548 17342 680 4 vdd
rlabel metal3 s 5372 5268 5438 5400 4 vdd
rlabel metal3 s 42198 3986 42330 4060 4 vdd
rlabel metal3 s 34936 5268 35002 5400 4 vdd
rlabel metal3 s 48940 5268 49006 5400 4 vdd
rlabel metal3 s 17302 3986 17434 4060 4 vdd
rlabel metal3 s 28466 3986 28598 4060 4 vdd
rlabel metal3 s 36246 3986 36378 4060 4 vdd
rlabel metal3 s 10040 5268 10106 5400 4 vdd
rlabel metal3 s 45582 3986 45714 4060 4 vdd
rlabel metal3 s 6384 548 6450 680 4 vdd
rlabel metal3 s 23500 548 23566 680 4 vdd
rlabel metal3 s 39358 3986 39490 4060 4 vdd
rlabel metal3 s 33134 3986 33266 4060 4 vdd
rlabel metal3 s 38048 5268 38114 5400 4 vdd
rlabel metal3 s 35974 3986 36106 4060 4 vdd
rlabel metal3 s 49952 548 50018 680 4 vdd
rlabel metal3 s 38282 548 38348 680 4 vdd
rlabel metal3 s 13386 548 13452 680 4 vdd
rlabel metal3 s 28194 3986 28326 4060 4 vdd
rlabel metal3 s 45310 3986 45442 4060 4 vdd
rlabel metal3 s 8718 548 8784 680 4 vdd
rlabel metal3 s 186 3986 318 4060 4 vdd
rlabel metal3 s 14462 3986 14594 4060 4 vdd
rlabel metal3 s 11830 548 11896 680 4 vdd
rlabel metal3 s 17820 5268 17886 5400 4 vdd
rlabel metal3 s 22242 3986 22374 4060 4 vdd
rlabel metal3 s 45828 5268 45894 5400 4 vdd
rlabel metal3 s 42716 5268 42782 5400 4 vdd
rlabel metal3 s 11596 5268 11662 5400 4 vdd
rlabel metal3 s 42470 3986 42602 4060 4 vdd
rlabel metal3 s 20388 548 20454 680 4 vdd
rlabel metal3 s 44026 3986 44158 4060 4 vdd
rlabel metal3 s 42950 548 43016 680 4 vdd
rlabel metal3 s 18832 548 18898 680 4 vdd
rlabel metal3 s 46866 3986 46998 4060 4 vdd
rlabel metal3 s 34392 548 34458 680 4 vdd
rlabel metal3 s 3272 548 3338 680 4 vdd
rlabel metal3 s 44272 5268 44338 5400 4 vdd
rlabel metal3 s 6928 5268 6994 5400 4 vdd
rlabel metal3 s 2260 5268 2326 5400 4 vdd
rlabel metal3 s 39838 548 39904 680 4 vdd
rlabel metal3 s 33380 5268 33446 5400 4 vdd
rlabel metal3 s 25354 3986 25486 4060 4 vdd
rlabel metal3 s 29750 3986 29882 4060 4 vdd
rlabel metal3 s 5126 3986 5258 4060 4 vdd
rlabel metal3 s 19376 5268 19442 5400 4 vdd
rlabel metal3 s 2494 548 2560 680 4 vdd
rlabel metal3 s 29724 548 29790 680 4 vdd
rlabel metal3 s 4854 3986 4986 4060 4 vdd
rlabel metal3 s 3816 5268 3882 5400 4 vdd
rlabel metal3 s 35948 548 36014 680 4 vdd
rlabel metal3 s 22722 548 22788 680 4 vdd
rlabel metal3 s 458 3986 590 4060 4 vdd
rlabel metal3 s 18858 3986 18990 4060 4 vdd
rlabel metal3 s 25834 548 25900 680 4 vdd
rlabel metal3 s 4828 548 4894 680 4 vdd
rlabel metal3 s 34690 3986 34822 4060 4 vdd
rlabel metal3 s 31306 3986 31438 4060 4 vdd
rlabel metal3 s 40642 3986 40774 4060 4 vdd
rlabel metal3 s 21944 548 22010 680 4 vdd
rlabel metal3 s 48694 3986 48826 4060 4 vdd
rlabel metal3 s 25600 5268 25666 5400 4 vdd
rlabel metal3 s 14164 548 14230 680 4 vdd
rlabel metal3 s 11052 548 11118 680 4 vdd
rlabel metal3 s 18054 548 18120 680 4 vdd
rlabel metal3 s 9794 3986 9926 4060 4 vdd
rlabel metal3 s 21970 3986 22102 4060 4 vdd
rlabel metal3 s 15746 3986 15878 4060 4 vdd
rlabel metal3 s 46062 548 46128 680 4 vdd
rlabel metal3 s 11350 3986 11482 4060 4 vdd
rlabel metal3 s 48422 3986 48554 4060 4 vdd
rlabel metal3 s 40616 548 40682 680 4 vdd
rlabel metal3 s 41160 5268 41226 5400 4 vdd
rlabel metal3 s 24044 5268 24110 5400 4 vdd
rlabel metal3 s 49174 548 49240 680 4 vdd
rlabel metal3 s 43754 3986 43886 4060 4 vdd
rlabel metal3 s 3570 3986 3702 4060 4 vdd
rlabel metal3 s 39086 3986 39218 4060 4 vdd
rlabel metal3 s 32058 548 32124 680 4 vdd
rlabel metal3 s 14708 5268 14774 5400 4 vdd
rlabel metal3 s 31280 548 31346 680 4 vdd
rlabel metal3 s 36726 548 36792 680 4 vdd
rlabel metal3 s 31578 3986 31710 4060 4 vdd
rlabel metal3 s 17574 3986 17706 4060 4 vdd
rlabel metal3 s 8484 5268 8550 5400 4 vdd
rlabel metal3 s 26910 3986 27042 4060 4 vdd
rlabel metal3 s 37530 3986 37662 4060 4 vdd
rlabel metal3 s 32836 548 32902 680 4 vdd
rlabel metal3 s 48396 548 48462 680 4 vdd
rlabel metal3 s 704 5268 770 5400 4 vdd
rlabel metal3 s 43728 548 43794 680 4 vdd
rlabel metal3 s 938 548 1004 680 4 vdd
rlabel metal3 s 25056 548 25122 680 4 vdd
rlabel metal3 s 26638 3986 26770 4060 4 vdd
rlabel metal3 s 6410 3986 6542 4060 4 vdd
rlabel metal3 s 19610 548 19676 680 4 vdd
rlabel metal3 s 44506 548 44572 680 4 vdd
rlabel metal3 s 47618 548 47684 680 4 vdd
rlabel metal3 s 39604 5268 39670 5400 4 vdd
rlabel metal3 s 28168 548 28234 680 4 vdd
rlabel metal3 s 20686 3986 20818 4060 4 vdd
rlabel metal3 s 41394 548 41460 680 4 vdd
rlabel metal3 s 33614 548 33680 680 4 vdd
rlabel metal3 s 2014 3986 2146 4060 4 vdd
rlabel metal3 s 27156 5268 27222 5400 4 vdd
rlabel metal3 s 7966 3986 8098 4060 4 vdd
rlabel metal3 s 24278 548 24344 680 4 vdd
rlabel metal3 s 7940 548 8006 680 4 vdd
rlabel metal3 s 8238 3986 8370 4060 4 vdd
rlabel metal3 s 11078 3986 11210 4060 4 vdd
rlabel metal3 s 20414 3986 20546 4060 4 vdd
rlabel metal3 s 160 548 226 680 4 vdd
rlabel metal3 s 21166 548 21232 680 4 vdd
rlabel metal3 s 23798 3986 23930 4060 4 vdd
rlabel metal3 s 28946 548 29012 680 4 vdd
rlabel metal3 s 42172 548 42238 680 4 vdd
rlabel metal3 s 37802 3986 37934 4060 4 vdd
rlabel metal3 s 28712 5268 28778 5400 4 vdd
rlabel metal3 s 12906 3986 13038 4060 4 vdd
rlabel metal3 s 45284 548 45350 680 4 vdd
rlabel metal3 s 26612 548 26678 680 4 vdd
rlabel metal3 s 22488 5268 22554 5400 4 vdd
rlabel metal3 s 35170 548 35236 680 4 vdd
rlabel metal3 s 34418 3986 34550 4060 4 vdd
rlabel metal3 s 19130 3986 19262 4060 4 vdd
rlabel metal3 s 12608 548 12674 680 4 vdd
rlabel metal3 s 16498 548 16564 680 4 vdd
rlabel metal3 s 9496 548 9562 680 4 vdd
rlabel metal3 s 40914 3986 41046 4060 4 vdd
rlabel metal3 s 3298 3986 3430 4060 4 vdd
rlabel metal3 s 1742 3986 1874 4060 4 vdd
rlabel metal3 s 46840 548 46906 680 4 vdd
rlabel metal3 s 37504 548 37570 680 4 vdd
rlabel metal3 s 48170 2506 48302 2580 4 gnd
rlabel metal3 s 34936 6100 35002 6232 4 gnd
rlabel metal3 s 33134 4932 33266 5006 4 gnd
rlabel metal3 s 8484 6100 8550 6232 4 gnd
rlabel metal3 s 35974 4932 36106 5006 4 gnd
rlabel metal3 s 13152 6100 13218 6232 4 gnd
rlabel metal3 s 6928 6100 6994 6232 4 gnd
rlabel metal3 s 15494 2506 15626 2580 4 gnd
rlabel metal3 s 29750 4932 29882 5006 4 gnd
rlabel metal3 s 47384 6100 47450 6232 4 gnd
rlabel metal3 s 40642 4932 40774 5006 4 gnd
rlabel metal3 s 22488 6100 22554 6232 4 gnd
rlabel metal3 s 20932 6100 20998 6232 4 gnd
rlabel metal3 s 46866 4932 46998 5006 4 gnd
rlabel metal3 s 712 2506 844 2580 4 gnd
rlabel metal3 s 27942 2506 28074 2580 4 gnd
rlabel metal3 s 11078 4932 11210 5006 4 gnd
rlabel metal3 s 30276 2506 30408 2580 4 gnd
rlabel metal3 s 27164 2506 27296 2580 4 gnd
rlabel metal3 s 45828 6100 45894 6232 4 gnd
rlabel metal3 s 47138 4932 47270 5006 4 gnd
rlabel metal3 s 5126 4932 5258 5006 4 gnd
rlabel metal3 s 12634 4932 12766 5006 4 gnd
rlabel metal3 s 15746 4932 15878 5006 4 gnd
rlabel metal3 s 3816 6100 3882 6232 4 gnd
rlabel metal3 s 20162 2506 20294 2580 4 gnd
rlabel metal3 s 8238 4932 8370 5006 4 gnd
rlabel metal3 s 186 4932 318 5006 4 gnd
rlabel metal3 s 14190 4932 14322 5006 4 gnd
rlabel metal3 s 6682 4932 6814 5006 4 gnd
rlabel metal3 s 1490 2506 1622 2580 4 gnd
rlabel metal3 s 31054 2506 31186 2580 4 gnd
rlabel metal3 s 4602 2506 4734 2580 4 gnd
rlabel metal3 s 21718 2506 21850 2580 4 gnd
rlabel metal3 s 29498 2506 29630 2580 4 gnd
rlabel metal3 s 32862 4932 32994 5006 4 gnd
rlabel metal3 s 42716 6100 42782 6232 4 gnd
rlabel metal3 s 8492 2506 8624 2580 4 gnd
rlabel metal3 s 48948 2506 49080 2580 4 gnd
rlabel metal3 s 34944 2506 35076 2580 4 gnd
rlabel metal3 s 39358 4932 39490 5006 4 gnd
rlabel metal3 s 13938 2506 14070 2580 4 gnd
rlabel metal3 s 23798 4932 23930 5006 4 gnd
rlabel metal3 s 44272 6100 44338 6232 4 gnd
rlabel metal3 s 26910 4932 27042 5006 4 gnd
rlabel metal3 s 25082 4932 25214 5006 4 gnd
rlabel metal3 s 2268 2506 2400 2580 4 gnd
rlabel metal3 s 37802 4932 37934 5006 4 gnd
rlabel metal3 s 32610 2506 32742 2580 4 gnd
rlabel metal3 s 42198 4932 42330 5006 4 gnd
rlabel metal3 s 39604 6100 39670 6232 4 gnd
rlabel metal3 s 41160 6100 41226 6232 4 gnd
rlabel metal3 s 16264 6100 16330 6232 4 gnd
rlabel metal3 s 16272 2506 16404 2580 4 gnd
rlabel metal3 s 9270 2506 9402 2580 4 gnd
rlabel metal3 s 42724 2506 42856 2580 4 gnd
rlabel metal3 s 37278 2506 37410 2580 4 gnd
rlabel metal3 s 43502 2506 43634 2580 4 gnd
rlabel metal3 s 45058 2506 45190 2580 4 gnd
rlabel metal3 s 43754 4932 43886 5006 4 gnd
rlabel metal3 s 34166 2506 34298 2580 4 gnd
rlabel metal3 s 17302 4932 17434 5006 4 gnd
rlabel metal3 s 10826 2506 10958 2580 4 gnd
rlabel metal3 s 30268 6100 30334 6232 4 gnd
rlabel metal3 s 6158 2506 6290 2580 4 gnd
rlabel metal3 s 6936 2506 7068 2580 4 gnd
rlabel metal3 s 16018 4932 16150 5006 4 gnd
rlabel metal3 s 24830 2506 24962 2580 4 gnd
rlabel metal3 s 44280 2506 44412 2580 4 gnd
rlabel metal3 s 41168 2506 41300 2580 4 gnd
rlabel metal3 s 2260 6100 2326 6232 4 gnd
rlabel metal3 s 45310 4932 45442 5006 4 gnd
rlabel metal3 s 22496 2506 22628 2580 4 gnd
rlabel metal3 s 40390 2506 40522 2580 4 gnd
rlabel metal3 s 20686 4932 20818 5006 4 gnd
rlabel metal3 s 45582 4932 45714 5006 4 gnd
rlabel metal3 s 38048 6100 38114 6232 4 gnd
rlabel metal3 s 23526 4932 23658 5006 4 gnd
rlabel metal3 s 47392 2506 47524 2580 4 gnd
rlabel metal3 s 28194 4932 28326 5006 4 gnd
rlabel metal3 s 11596 6100 11662 6232 4 gnd
rlabel metal3 s 36492 6100 36558 6232 4 gnd
rlabel metal3 s 20414 4932 20546 5006 4 gnd
rlabel metal3 s 28712 6100 28778 6232 4 gnd
rlabel metal3 s 17828 2506 17960 2580 4 gnd
rlabel metal3 s 45836 2506 45968 2580 4 gnd
rlabel metal3 s 28720 2506 28852 2580 4 gnd
rlabel metal3 s 5372 6100 5438 6232 4 gnd
rlabel metal3 s 5380 2506 5512 2580 4 gnd
rlabel metal3 s 27156 6100 27222 6232 4 gnd
rlabel metal3 s 30022 4932 30154 5006 4 gnd
rlabel metal3 s 49726 2506 49858 2580 4 gnd
rlabel metal3 s 34690 4932 34822 5006 4 gnd
rlabel metal3 s 37530 4932 37662 5006 4 gnd
rlabel metal3 s 18606 2506 18738 2580 4 gnd
rlabel metal3 s 9522 4932 9654 5006 4 gnd
rlabel metal3 s 46614 2506 46746 2580 4 gnd
rlabel metal3 s 33388 2506 33520 2580 4 gnd
rlabel metal3 s 3046 2506 3178 2580 4 gnd
rlabel metal3 s 21970 4932 22102 5006 4 gnd
rlabel metal3 s 31824 6100 31890 6232 4 gnd
rlabel metal3 s 458 4932 590 5006 4 gnd
rlabel metal3 s 11604 2506 11736 2580 4 gnd
rlabel metal3 s 34418 4932 34550 5006 4 gnd
rlabel metal3 s 20940 2506 21072 2580 4 gnd
rlabel metal3 s 25608 2506 25740 2580 4 gnd
rlabel metal3 s 39612 2506 39744 2580 4 gnd
rlabel metal3 s 11350 4932 11482 5006 4 gnd
rlabel metal3 s 17574 4932 17706 5006 4 gnd
rlabel metal3 s 704 6100 770 6232 4 gnd
rlabel metal3 s 3298 4932 3430 5006 4 gnd
rlabel metal3 s 38834 2506 38966 2580 4 gnd
rlabel metal3 s 12382 2506 12514 2580 4 gnd
rlabel metal3 s 42470 4932 42602 5006 4 gnd
rlabel metal3 s 40914 4932 41046 5006 4 gnd
rlabel metal3 s 7966 4932 8098 5006 4 gnd
rlabel metal3 s 33380 6100 33446 6232 4 gnd
rlabel metal3 s 14708 6100 14774 6232 4 gnd
rlabel metal3 s 48422 4932 48554 5006 4 gnd
rlabel metal3 s 4854 4932 4986 5006 4 gnd
rlabel metal3 s 26638 4932 26770 5006 4 gnd
rlabel metal3 s 48940 6100 49006 6232 4 gnd
rlabel metal3 s 31578 4932 31710 5006 4 gnd
rlabel metal3 s 22242 4932 22374 5006 4 gnd
rlabel metal3 s 14716 2506 14848 2580 4 gnd
rlabel metal3 s 38056 2506 38188 2580 4 gnd
rlabel metal3 s 19384 2506 19516 2580 4 gnd
rlabel metal3 s 25600 6100 25666 6232 4 gnd
rlabel metal3 s 17050 2506 17182 2580 4 gnd
rlabel metal3 s 35722 2506 35854 2580 4 gnd
rlabel metal3 s 31832 2506 31964 2580 4 gnd
rlabel metal3 s 3824 2506 3956 2580 4 gnd
rlabel metal3 s 7714 2506 7846 2580 4 gnd
rlabel metal3 s 10040 6100 10106 6232 4 gnd
rlabel metal3 s 9794 4932 9926 5006 4 gnd
rlabel metal3 s 19376 6100 19442 6232 4 gnd
rlabel metal3 s 36246 4932 36378 5006 4 gnd
rlabel metal3 s 18858 4932 18990 5006 4 gnd
rlabel metal3 s 39086 4932 39218 5006 4 gnd
rlabel metal3 s 36500 2506 36632 2580 4 gnd
rlabel metal3 s 24044 6100 24110 6232 4 gnd
rlabel metal3 s 44026 4932 44158 5006 4 gnd
rlabel metal3 s 2014 4932 2146 5006 4 gnd
rlabel metal3 s 41946 2506 42078 2580 4 gnd
rlabel metal3 s 1742 4932 1874 5006 4 gnd
rlabel metal3 s 31306 4932 31438 5006 4 gnd
rlabel metal3 s 23274 2506 23406 2580 4 gnd
rlabel metal3 s 12906 4932 13038 5006 4 gnd
rlabel metal3 s 25354 4932 25486 5006 4 gnd
rlabel metal3 s 17820 6100 17886 6232 4 gnd
rlabel metal3 s 24052 2506 24184 2580 4 gnd
rlabel metal3 s 28466 4932 28598 5006 4 gnd
rlabel metal3 s 6410 4932 6542 5006 4 gnd
rlabel metal3 s 14462 4932 14594 5006 4 gnd
rlabel metal3 s 48694 4932 48826 5006 4 gnd
rlabel metal3 s 26386 2506 26518 2580 4 gnd
rlabel metal3 s 13160 2506 13292 2580 4 gnd
rlabel metal3 s 3570 4932 3702 5006 4 gnd
rlabel metal3 s 10048 2506 10180 2580 4 gnd
rlabel metal3 s 19130 4932 19262 5006 4 gnd
<< properties >>
string FIXED_BBOX 0 0 50570 5956
string GDS_FILE sram_0rw2r1w_32_128_sky130A.gds
string GDS_END 2476104
string GDS_START 2331472
<< end >>
