magic
tech sky130A
magscale 1 2
timestamp 1643678851
<< checkpaint >>
rect -1260 -1294 3129 7454
<< locali >>
rect 0 6143 227 6177
rect 261 6143 986 6177
rect 1020 6143 1833 6177
rect 1661 5415 1695 5449
rect 0 4603 227 4637
rect 261 4603 986 4637
rect 1020 4603 1833 4637
rect 1661 3791 1695 3825
rect 0 3063 227 3097
rect 261 3063 986 3097
rect 1020 3063 1833 3097
rect 1661 2335 1695 2369
rect 0 1523 227 1557
rect 261 1523 986 1557
rect 1020 1523 1833 1557
rect 1661 711 1695 745
rect 0 -17 227 17
rect 261 -17 986 17
rect 1020 -17 1833 17
<< viali >>
rect 227 6143 261 6177
rect 986 6143 1020 6177
rect 1143 5853 1177 5887
rect 1243 5605 1277 5639
rect 227 4603 261 4637
rect 986 4603 1020 4637
rect 1243 3601 1277 3635
rect 1143 3353 1177 3387
rect 227 3063 261 3097
rect 986 3063 1020 3097
rect 1143 2773 1177 2807
rect 1243 2525 1277 2559
rect 336 2335 370 2369
rect 468 2335 502 2369
rect 227 1523 261 1557
rect 986 1523 1020 1557
rect 336 711 370 745
rect 468 711 502 745
rect 1243 521 1277 555
rect 1143 273 1177 307
rect 227 -17 261 17
rect 986 -17 1020 17
<< metal1 >>
rect 215 6175 218 6183
rect 189 6145 218 6175
rect 215 6137 218 6145
rect 270 6175 273 6183
rect 974 6175 977 6183
rect 270 6145 300 6175
rect 948 6145 977 6175
rect 270 6137 273 6145
rect 974 6137 977 6145
rect 1029 6175 1032 6183
rect 1029 6145 1059 6175
rect 1029 6137 1032 6145
rect 108 5856 815 5884
rect 1131 5887 1189 5893
rect 1131 5884 1143 5887
rect 867 5856 1143 5884
rect 1131 5853 1143 5856
rect 1177 5853 1189 5887
rect 1131 5847 1189 5853
rect 176 5608 883 5636
rect 1231 5639 1289 5645
rect 1231 5636 1243 5639
rect 935 5608 1243 5636
rect 1231 5605 1243 5608
rect 1277 5605 1289 5639
rect 1231 5599 1289 5605
rect 215 4635 218 4643
rect 189 4605 218 4635
rect 215 4597 218 4605
rect 270 4635 273 4643
rect 974 4635 977 4643
rect 270 4605 300 4635
rect 948 4605 977 4635
rect 270 4597 273 4605
rect 974 4597 977 4605
rect 1029 4635 1032 4643
rect 1029 4605 1059 4635
rect 1029 4597 1032 4605
rect 1231 3635 1289 3641
rect 1231 3632 1243 3635
rect 935 3604 1243 3632
rect 1231 3601 1243 3604
rect 1277 3601 1289 3635
rect 1231 3595 1289 3601
rect 1131 3387 1189 3393
rect 1131 3384 1143 3387
rect 731 3356 1143 3384
rect 1131 3353 1143 3356
rect 1177 3353 1189 3387
rect 1131 3347 1189 3353
rect 215 3095 218 3103
rect 189 3065 218 3095
rect 215 3057 218 3065
rect 270 3095 273 3103
rect 974 3095 977 3103
rect 270 3065 300 3095
rect 948 3065 977 3095
rect 270 3057 273 3065
rect 974 3057 977 3065
rect 1029 3095 1032 3103
rect 1029 3065 1059 3095
rect 1029 3057 1032 3065
rect 609 3008 747 3036
rect 324 2369 382 2375
rect 324 2366 336 2369
rect 176 2338 336 2366
rect 324 2335 336 2338
rect 370 2335 382 2369
rect 324 2329 382 2335
rect 456 2369 514 2375
rect 456 2335 468 2369
rect 502 2366 514 2369
rect 609 2366 637 3008
rect 1131 2807 1189 2813
rect 1131 2804 1143 2807
rect 867 2776 1143 2804
rect 1131 2773 1143 2776
rect 1177 2773 1189 2807
rect 1131 2767 1189 2773
rect 1231 2559 1289 2565
rect 1231 2556 1243 2559
rect 799 2528 1243 2556
rect 1231 2525 1243 2528
rect 1277 2525 1289 2559
rect 1231 2519 1289 2525
rect 502 2338 637 2366
rect 502 2335 514 2338
rect 456 2329 514 2335
rect 215 1555 218 1563
rect 189 1525 218 1555
rect 215 1517 218 1525
rect 270 1555 273 1563
rect 974 1555 977 1563
rect 270 1525 300 1555
rect 948 1525 977 1555
rect 270 1517 273 1525
rect 974 1517 977 1525
rect 1029 1555 1032 1563
rect 1029 1525 1059 1555
rect 1029 1517 1032 1525
rect 609 1468 679 1496
rect 324 745 382 751
rect 324 742 336 745
rect 108 714 336 742
rect 324 711 336 714
rect 370 711 382 745
rect 324 705 382 711
rect 456 745 514 751
rect 456 711 468 745
rect 502 742 514 745
rect 609 742 637 1468
rect 502 714 637 742
rect 502 711 514 714
rect 456 705 514 711
rect 1231 555 1289 561
rect 1231 552 1243 555
rect 799 524 1243 552
rect 1231 521 1243 524
rect 1277 521 1289 555
rect 1231 515 1289 521
rect 1131 307 1189 313
rect 1131 304 1143 307
rect 731 276 1143 304
rect 1131 273 1143 276
rect 1177 273 1189 307
rect 1131 267 1189 273
rect 215 15 218 23
rect 189 -15 218 15
rect 215 -23 218 -15
rect 270 15 273 23
rect 974 15 977 23
rect 270 -15 300 15
rect 948 -15 977 15
rect 270 -23 273 -15
rect 974 -23 977 -15
rect 1029 15 1032 23
rect 1029 -15 1059 15
rect 1029 -23 1032 -15
<< via1 >>
rect 218 6177 270 6186
rect 218 6143 227 6177
rect 227 6143 261 6177
rect 261 6143 270 6177
rect 977 6177 1029 6186
rect 218 6134 270 6143
rect 977 6143 986 6177
rect 986 6143 1020 6177
rect 1020 6143 1029 6177
rect 977 6134 1029 6143
rect 56 5844 108 5896
rect 815 5844 867 5896
rect 124 5596 176 5648
rect 883 5596 935 5648
rect 218 4637 270 4646
rect 218 4603 227 4637
rect 227 4603 261 4637
rect 261 4603 270 4637
rect 977 4637 1029 4646
rect 218 4594 270 4603
rect 977 4603 986 4637
rect 986 4603 1020 4637
rect 1020 4603 1029 4637
rect 977 4594 1029 4603
rect 883 3592 935 3644
rect 679 3344 731 3396
rect 218 3097 270 3106
rect 218 3063 227 3097
rect 227 3063 261 3097
rect 261 3063 270 3097
rect 977 3097 1029 3106
rect 218 3054 270 3063
rect 977 3063 986 3097
rect 986 3063 1020 3097
rect 1020 3063 1029 3097
rect 977 3054 1029 3063
rect 124 2326 176 2378
rect 747 2996 799 3048
rect 815 2764 867 2816
rect 747 2516 799 2568
rect 218 1557 270 1566
rect 218 1523 227 1557
rect 227 1523 261 1557
rect 261 1523 270 1557
rect 977 1557 1029 1566
rect 218 1514 270 1523
rect 977 1523 986 1557
rect 986 1523 1020 1557
rect 1020 1523 1029 1557
rect 977 1514 1029 1523
rect 56 702 108 754
rect 679 1456 731 1508
rect 747 512 799 564
rect 679 264 731 316
rect 218 17 270 26
rect 218 -17 227 17
rect 227 -17 261 17
rect 261 -17 270 17
rect 977 17 1029 26
rect 218 -26 270 -17
rect 977 -17 986 17
rect 986 -17 1020 17
rect 1020 -17 1029 17
rect 977 -26 1029 -17
<< metal2 >>
rect 224 6188 264 6194
rect 983 6188 1023 6194
rect 68 5896 96 6160
rect 68 754 96 5844
rect 136 5648 164 6160
rect 224 6126 264 6132
rect 136 2378 164 5596
rect 224 4648 264 4654
rect 224 4586 264 4592
rect 691 3396 719 6160
rect 224 3108 264 3114
rect 224 3046 264 3052
rect 68 68 96 702
rect 136 68 164 2326
rect 224 1568 264 1574
rect 224 1506 264 1512
rect 691 1508 719 3344
rect 759 3048 787 6160
rect 827 5896 855 6160
rect 759 2568 787 2996
rect 827 2816 855 5844
rect 895 5648 923 6160
rect 983 6126 1023 6132
rect 895 3644 923 5596
rect 983 4648 1023 4654
rect 983 4586 1023 4592
rect 691 316 719 1456
rect 759 564 787 2516
rect 691 68 719 264
rect 759 68 787 512
rect 827 68 855 2764
rect 895 68 923 3592
rect 983 3108 1023 3114
rect 983 3046 1023 3052
rect 983 1568 1023 1574
rect 983 1506 1023 1512
rect 224 28 264 34
rect 983 28 1023 34
rect 224 -34 264 -28
rect 983 -34 1023 -28
<< via2 >>
rect 216 6186 272 6188
rect 216 6134 218 6186
rect 218 6134 270 6186
rect 270 6134 272 6186
rect 975 6186 1031 6188
rect 216 6132 272 6134
rect 216 4646 272 4648
rect 216 4594 218 4646
rect 218 4594 270 4646
rect 270 4594 272 4646
rect 216 4592 272 4594
rect 216 3106 272 3108
rect 216 3054 218 3106
rect 218 3054 270 3106
rect 270 3054 272 3106
rect 216 3052 272 3054
rect 216 1566 272 1568
rect 216 1514 218 1566
rect 218 1514 270 1566
rect 270 1514 272 1566
rect 216 1512 272 1514
rect 975 6134 977 6186
rect 977 6134 1029 6186
rect 1029 6134 1031 6186
rect 975 6132 1031 6134
rect 975 4646 1031 4648
rect 975 4594 977 4646
rect 977 4594 1029 4646
rect 1029 4594 1031 4646
rect 975 4592 1031 4594
rect 975 3106 1031 3108
rect 975 3054 977 3106
rect 977 3054 1029 3106
rect 1029 3054 1031 3106
rect 975 3052 1031 3054
rect 975 1566 1031 1568
rect 975 1514 977 1566
rect 977 1514 1029 1566
rect 1029 1514 1031 1566
rect 975 1512 1031 1514
rect 216 26 272 28
rect 216 -26 218 26
rect 218 -26 270 26
rect 270 -26 272 26
rect 216 -28 272 -26
rect 975 26 1031 28
rect 975 -26 977 26
rect 977 -26 1029 26
rect 1029 -26 1031 26
rect 975 -28 1031 -26
<< metal3 >>
rect 178 6188 310 6193
rect 178 6132 216 6188
rect 272 6132 310 6188
rect 178 6127 310 6132
rect 937 6188 1069 6193
rect 937 6132 975 6188
rect 1031 6132 1069 6188
rect 937 6127 1069 6132
rect 178 4648 310 4653
rect 178 4592 216 4648
rect 272 4592 310 4648
rect 178 4587 310 4592
rect 937 4648 1069 4653
rect 937 4592 975 4648
rect 1031 4592 1069 4648
rect 937 4587 1069 4592
rect 178 3108 310 3113
rect 178 3052 216 3108
rect 272 3052 310 3108
rect 178 3047 310 3052
rect 937 3108 1069 3113
rect 937 3052 975 3108
rect 1031 3052 1069 3108
rect 937 3047 1069 3052
rect 178 1568 310 1573
rect 178 1512 216 1568
rect 272 1512 310 1568
rect 178 1507 310 1512
rect 937 1568 1069 1573
rect 937 1512 975 1568
rect 1031 1512 1069 1568
rect 937 1507 1069 1512
rect 178 28 310 33
rect 178 -28 216 28
rect 272 -28 310 28
rect 178 -33 310 -28
rect 937 28 1069 33
rect 937 -28 975 28
rect 1031 -28 1069 28
rect 937 -33 1069 -28
use contact_18  contact_18_0
timestamp 1643678851
transform 1 0 937 0 1 6127
box 0 0 1 1
use contact_17  contact_17_0
timestamp 1643678851
transform 1 0 988 0 1 6145
box 0 0 1 1
use contact_13  contact_13_0
timestamp 1643678851
transform 1 0 974 0 1 6137
box 0 0 1 1
use contact_18  contact_18_1
timestamp 1643678851
transform 1 0 178 0 1 6127
box 0 0 1 1
use contact_17  contact_17_1
timestamp 1643678851
transform 1 0 229 0 1 6145
box 0 0 1 1
use contact_13  contact_13_1
timestamp 1643678851
transform 1 0 215 0 1 6137
box 0 0 1 1
use contact_18  contact_18_2
timestamp 1643678851
transform 1 0 937 0 1 4587
box 0 0 1 1
use contact_17  contact_17_2
timestamp 1643678851
transform 1 0 988 0 1 4605
box 0 0 1 1
use contact_13  contact_13_2
timestamp 1643678851
transform 1 0 974 0 1 4597
box 0 0 1 1
use contact_18  contact_18_3
timestamp 1643678851
transform 1 0 178 0 1 4587
box 0 0 1 1
use contact_17  contact_17_3
timestamp 1643678851
transform 1 0 229 0 1 4605
box 0 0 1 1
use contact_13  contact_13_3
timestamp 1643678851
transform 1 0 215 0 1 4597
box 0 0 1 1
use contact_18  contact_18_4
timestamp 1643678851
transform 1 0 937 0 1 3047
box 0 0 1 1
use contact_17  contact_17_4
timestamp 1643678851
transform 1 0 988 0 1 3065
box 0 0 1 1
use contact_13  contact_13_4
timestamp 1643678851
transform 1 0 974 0 1 3057
box 0 0 1 1
use contact_18  contact_18_5
timestamp 1643678851
transform 1 0 178 0 1 3047
box 0 0 1 1
use contact_17  contact_17_5
timestamp 1643678851
transform 1 0 229 0 1 3065
box 0 0 1 1
use contact_13  contact_13_5
timestamp 1643678851
transform 1 0 215 0 1 3057
box 0 0 1 1
use contact_18  contact_18_6
timestamp 1643678851
transform 1 0 937 0 1 4587
box 0 0 1 1
use contact_17  contact_17_6
timestamp 1643678851
transform 1 0 988 0 1 4605
box 0 0 1 1
use contact_13  contact_13_6
timestamp 1643678851
transform 1 0 974 0 1 4597
box 0 0 1 1
use contact_18  contact_18_7
timestamp 1643678851
transform 1 0 178 0 1 4587
box 0 0 1 1
use contact_17  contact_17_7
timestamp 1643678851
transform 1 0 229 0 1 4605
box 0 0 1 1
use contact_13  contact_13_7
timestamp 1643678851
transform 1 0 215 0 1 4597
box 0 0 1 1
use contact_18  contact_18_8
timestamp 1643678851
transform 1 0 937 0 1 3047
box 0 0 1 1
use contact_17  contact_17_8
timestamp 1643678851
transform 1 0 988 0 1 3065
box 0 0 1 1
use contact_13  contact_13_8
timestamp 1643678851
transform 1 0 974 0 1 3057
box 0 0 1 1
use contact_18  contact_18_9
timestamp 1643678851
transform 1 0 178 0 1 3047
box 0 0 1 1
use contact_17  contact_17_9
timestamp 1643678851
transform 1 0 229 0 1 3065
box 0 0 1 1
use contact_13  contact_13_9
timestamp 1643678851
transform 1 0 215 0 1 3057
box 0 0 1 1
use contact_18  contact_18_10
timestamp 1643678851
transform 1 0 937 0 1 1507
box 0 0 1 1
use contact_17  contact_17_10
timestamp 1643678851
transform 1 0 988 0 1 1525
box 0 0 1 1
use contact_13  contact_13_10
timestamp 1643678851
transform 1 0 974 0 1 1517
box 0 0 1 1
use contact_18  contact_18_11
timestamp 1643678851
transform 1 0 178 0 1 1507
box 0 0 1 1
use contact_17  contact_17_11
timestamp 1643678851
transform 1 0 229 0 1 1525
box 0 0 1 1
use contact_13  contact_13_11
timestamp 1643678851
transform 1 0 215 0 1 1517
box 0 0 1 1
use contact_18  contact_18_12
timestamp 1643678851
transform 1 0 937 0 1 -33
box 0 0 1 1
use contact_17  contact_17_12
timestamp 1643678851
transform 1 0 988 0 1 -15
box 0 0 1 1
use contact_13  contact_13_12
timestamp 1643678851
transform 1 0 974 0 1 -23
box 0 0 1 1
use contact_18  contact_18_13
timestamp 1643678851
transform 1 0 178 0 1 -33
box 0 0 1 1
use contact_17  contact_17_13
timestamp 1643678851
transform 1 0 229 0 1 -15
box 0 0 1 1
use contact_13  contact_13_13
timestamp 1643678851
transform 1 0 215 0 1 -23
box 0 0 1 1
use contact_18  contact_18_14
timestamp 1643678851
transform 1 0 937 0 1 1507
box 0 0 1 1
use contact_17  contact_17_14
timestamp 1643678851
transform 1 0 988 0 1 1525
box 0 0 1 1
use contact_13  contact_13_14
timestamp 1643678851
transform 1 0 974 0 1 1517
box 0 0 1 1
use contact_18  contact_18_15
timestamp 1643678851
transform 1 0 178 0 1 1507
box 0 0 1 1
use contact_17  contact_17_15
timestamp 1643678851
transform 1 0 229 0 1 1525
box 0 0 1 1
use contact_13  contact_13_15
timestamp 1643678851
transform 1 0 215 0 1 1517
box 0 0 1 1
use contact_17  contact_17_16
timestamp 1643678851
transform 1 0 894 0 1 5607
box 0 0 1 1
use contact_17  contact_17_17
timestamp 1643678851
transform 1 0 135 0 1 5607
box 0 0 1 1
use contact_17  contact_17_18
timestamp 1643678851
transform 1 0 826 0 1 5855
box 0 0 1 1
use contact_17  contact_17_19
timestamp 1643678851
transform 1 0 67 0 1 5855
box 0 0 1 1
use contact_14  contact_14_0
timestamp 1643678851
transform 1 0 758 0 1 3007
box 0 0 1 1
use contact_13  contact_13_16
timestamp 1643678851
transform 1 0 456 0 1 2329
box 0 0 1 1
use contact_14  contact_14_1
timestamp 1643678851
transform 1 0 690 0 1 1467
box 0 0 1 1
use contact_13  contact_13_17
timestamp 1643678851
transform 1 0 456 0 1 705
box 0 0 1 1
use contact_15  contact_15_0
timestamp 1643678851
transform 1 0 1231 0 1 5599
box 0 0 1 1
use contact_14  contact_14_2
timestamp 1643678851
transform 1 0 894 0 1 5607
box 0 0 1 1
use contact_13  contact_13_18
timestamp 1643678851
transform 1 0 1131 0 1 5847
box 0 0 1 1
use contact_14  contact_14_3
timestamp 1643678851
transform 1 0 826 0 1 5855
box 0 0 1 1
use contact_15  contact_15_1
timestamp 1643678851
transform 1 0 1231 0 1 3595
box 0 0 1 1
use contact_14  contact_14_4
timestamp 1643678851
transform 1 0 894 0 1 3603
box 0 0 1 1
use contact_13  contact_13_19
timestamp 1643678851
transform 1 0 1131 0 1 3347
box 0 0 1 1
use contact_14  contact_14_5
timestamp 1643678851
transform 1 0 690 0 1 3355
box 0 0 1 1
use contact_15  contact_15_2
timestamp 1643678851
transform 1 0 1231 0 1 2519
box 0 0 1 1
use contact_14  contact_14_6
timestamp 1643678851
transform 1 0 758 0 1 2527
box 0 0 1 1
use contact_13  contact_13_20
timestamp 1643678851
transform 1 0 1131 0 1 2767
box 0 0 1 1
use contact_14  contact_14_7
timestamp 1643678851
transform 1 0 826 0 1 2775
box 0 0 1 1
use contact_15  contact_15_3
timestamp 1643678851
transform 1 0 1231 0 1 515
box 0 0 1 1
use contact_14  contact_14_8
timestamp 1643678851
transform 1 0 758 0 1 523
box 0 0 1 1
use contact_13  contact_13_21
timestamp 1643678851
transform 1 0 1131 0 1 267
box 0 0 1 1
use contact_14  contact_14_9
timestamp 1643678851
transform 1 0 690 0 1 275
box 0 0 1 1
use contact_14  contact_14_10
timestamp 1643678851
transform 1 0 135 0 1 2337
box 0 0 1 1
use contact_13  contact_13_22
timestamp 1643678851
transform 1 0 324 0 1 2329
box 0 0 1 1
use contact_14  contact_14_11
timestamp 1643678851
transform 1 0 67 0 1 713
box 0 0 1 1
use contact_13  contact_13_23
timestamp 1643678851
transform 1 0 324 0 1 705
box 0 0 1 1
use and2_dec  and2_dec_0
timestamp 1643678851
transform 1 0 1031 0 -1 6160
box -36 -17 838 1597
use and2_dec  and2_dec_1
timestamp 1643678851
transform 1 0 1031 0 1 3080
box -36 -17 838 1597
use and2_dec  and2_dec_2
timestamp 1643678851
transform 1 0 1031 0 -1 3080
box -36 -17 838 1597
use and2_dec  and2_dec_3
timestamp 1643678851
transform 1 0 1031 0 1 0
box -36 -17 838 1597
use pinv  pinv_0
timestamp 1643678851
transform 1 0 272 0 -1 3080
box -36 -17 387 1597
use pinv  pinv_1
timestamp 1643678851
transform 1 0 272 0 1 0
box -36 -17 387 1597
<< labels >>
rlabel metal2 s 67 713 97 743 4 in_0
rlabel metal2 s 135 2337 165 2367 4 in_1
rlabel locali s 1678 728 1678 728 4 out_0
rlabel locali s 1678 2352 1678 2352 4 out_1
rlabel locali s 1678 3808 1678 3808 4 out_2
rlabel locali s 1678 5432 1678 5432 4 out_3
rlabel metal3 s 178 4587 310 4653 4 vdd
rlabel metal3 s 937 4587 1069 4653 4 vdd
rlabel metal3 s 937 1507 1069 1573 4 vdd
rlabel metal3 s 178 1507 310 1573 4 vdd
rlabel metal3 s 178 3047 310 3113 4 gnd
rlabel metal3 s 178 -33 310 33 4 gnd
rlabel metal3 s 937 6127 1069 6193 4 gnd
rlabel metal3 s 937 -33 1069 33 4 gnd
rlabel metal3 s 937 3047 1069 3113 4 gnd
rlabel metal3 s 178 6127 310 6193 4 gnd
<< properties >>
string FIXED_BBOX 937 -33 1069 0
string GDS_FILE sram_0rw2r1w_16_128_sky130A.gds
string GDS_END 1847720
string GDS_START 1837248
<< end >>
