magic
tech sky130A
magscale 1 2
timestamp 1644969367
<< checkpaint >>
rect -1260 -1260 60126 106280
<< locali >>
rect 5124 4029 5158 4063
<< viali >>
rect 5865 5328 5899 5362
rect 6178 4951 6212 4985
rect 5865 4490 5899 4524
rect 6178 4029 6212 4063
rect 5865 3652 5899 3686
<< metal1 >>
rect 8155 104264 8296 104292
rect 8155 104166 8183 104264
rect 8155 104156 8296 104166
rect 8006 104138 8296 104156
rect 8006 104128 8183 104138
rect 8155 104030 8183 104128
rect 8006 104002 8183 104030
rect 8155 103912 8296 103940
rect 8155 103804 8183 103912
rect 8006 103776 8183 103804
rect 8155 102852 8296 102880
rect 8155 102764 8183 102852
rect 8006 102736 8183 102764
rect 8155 102626 8296 102654
rect 8155 102538 8183 102626
rect 8006 102528 8183 102538
rect 8006 102510 8296 102528
rect 8155 102500 8296 102510
rect 8155 102412 8183 102500
rect 8006 102384 8183 102412
rect 8155 101184 8296 101212
rect 8155 101086 8183 101184
rect 8155 101080 8296 101086
rect 8006 101058 8296 101080
rect 8006 101052 8183 101058
rect 8155 100954 8183 101052
rect 8006 100926 8183 100954
rect 8155 100832 8296 100860
rect 8155 100728 8183 100832
rect 8006 100700 8183 100728
rect 8155 99772 8296 99800
rect 8155 99688 8183 99772
rect 8006 99660 8183 99688
rect 8155 99546 8296 99574
rect 8155 99462 8183 99546
rect 8006 99448 8183 99462
rect 8006 99434 8296 99448
rect 8155 99420 8296 99434
rect 8155 99336 8183 99420
rect 8006 99308 8183 99336
rect 8155 98104 8296 98132
rect 8155 98006 8183 98104
rect 8155 98004 8296 98006
rect 8006 97978 8296 98004
rect 8006 97976 8183 97978
rect 8155 97878 8183 97976
rect 8006 97850 8183 97878
rect 8155 97752 8296 97780
rect 8155 97652 8183 97752
rect 8006 97624 8183 97652
rect 8155 96692 8296 96720
rect 8155 96612 8183 96692
rect 8006 96584 8183 96612
rect 8155 96466 8296 96494
rect 8155 96386 8183 96466
rect 8006 96368 8183 96386
rect 8006 96358 8296 96368
rect 8155 96340 8296 96358
rect 8155 96260 8183 96340
rect 8006 96232 8183 96260
rect 8155 95024 8296 95052
rect 8155 94928 8183 95024
rect 8006 94926 8183 94928
rect 8006 94900 8296 94926
rect 8155 94898 8296 94900
rect 8155 94802 8183 94898
rect 8006 94774 8183 94802
rect 8155 94672 8296 94700
rect 8155 94576 8183 94672
rect 8006 94548 8183 94576
rect 8155 93612 8296 93640
rect 8155 93536 8183 93612
rect 8006 93508 8183 93536
rect 8155 93386 8296 93414
rect 8155 93310 8183 93386
rect 8006 93288 8183 93310
rect 8006 93282 8296 93288
rect 8155 93260 8296 93282
rect 8155 93184 8183 93260
rect 8006 93156 8183 93184
rect 8155 91944 8296 91972
rect 8155 91852 8183 91944
rect 8006 91846 8183 91852
rect 8006 91824 8296 91846
rect 8155 91818 8296 91824
rect 8155 91726 8183 91818
rect 8006 91698 8183 91726
rect 8155 91592 8296 91620
rect 8155 91500 8183 91592
rect 8006 91472 8183 91500
rect 8155 90532 8296 90560
rect 8155 90460 8183 90532
rect 8006 90432 8183 90460
rect 8155 90306 8296 90334
rect 8155 90234 8183 90306
rect 8006 90208 8183 90234
rect 8006 90206 8296 90208
rect 8155 90180 8296 90206
rect 8155 90108 8183 90180
rect 8006 90080 8183 90108
rect 8155 88864 8296 88892
rect 8155 88776 8183 88864
rect 8006 88766 8183 88776
rect 8006 88748 8296 88766
rect 8155 88738 8296 88748
rect 8155 88650 8183 88738
rect 8006 88622 8183 88650
rect 8155 88512 8296 88540
rect 8155 88424 8183 88512
rect 8006 88396 8183 88424
rect 8155 87452 8296 87480
rect 8155 87384 8183 87452
rect 8006 87356 8183 87384
rect 8155 87226 8296 87254
rect 8155 87158 8183 87226
rect 8006 87130 8183 87158
rect 8155 87100 8296 87128
rect 8155 87032 8183 87100
rect 8006 87004 8183 87032
rect 8155 85784 8296 85812
rect 8155 85700 8183 85784
rect 8006 85686 8183 85700
rect 8006 85672 8296 85686
rect 8155 85658 8296 85672
rect 8155 85574 8183 85658
rect 8006 85546 8183 85574
rect 8155 85432 8296 85460
rect 8155 85348 8183 85432
rect 8006 85320 8183 85348
rect 8155 84372 8296 84400
rect 8155 84308 8183 84372
rect 8006 84280 8183 84308
rect 8155 84146 8296 84174
rect 8155 84082 8183 84146
rect 8006 84054 8183 84082
rect 8155 84020 8296 84048
rect 8155 83956 8183 84020
rect 8006 83928 8183 83956
rect 8155 82704 8296 82732
rect 8155 82624 8183 82704
rect 8006 82606 8183 82624
rect 8006 82596 8296 82606
rect 8155 82578 8296 82596
rect 8155 82498 8183 82578
rect 8006 82470 8183 82498
rect 8155 82352 8296 82380
rect 8155 82272 8183 82352
rect 8006 82244 8183 82272
rect 8155 81292 8296 81320
rect 8155 81232 8183 81292
rect 8006 81204 8183 81232
rect 8155 81066 8296 81094
rect 8155 81006 8183 81066
rect 8006 80978 8183 81006
rect 8155 80940 8296 80968
rect 8155 80880 8183 80940
rect 8006 80852 8183 80880
rect 8155 79624 8296 79652
rect 8155 79548 8183 79624
rect 8006 79526 8183 79548
rect 8006 79520 8296 79526
rect 8155 79498 8296 79520
rect 8155 79422 8183 79498
rect 8006 79394 8183 79422
rect 8155 79272 8296 79300
rect 8155 79196 8183 79272
rect 8006 79168 8183 79196
rect 8155 78212 8296 78240
rect 8155 78156 8183 78212
rect 8006 78128 8183 78156
rect 8155 77986 8296 78014
rect 8155 77930 8183 77986
rect 8006 77902 8183 77930
rect 8155 77860 8296 77888
rect 8155 77804 8183 77860
rect 8006 77776 8183 77804
rect 8155 76544 8296 76572
rect 8155 76472 8183 76544
rect 8006 76446 8183 76472
rect 8006 76444 8296 76446
rect 8155 76418 8296 76444
rect 8155 76346 8183 76418
rect 8006 76318 8183 76346
rect 8155 76192 8296 76220
rect 8155 76120 8183 76192
rect 8006 76092 8183 76120
rect 8155 75132 8296 75160
rect 8155 75080 8183 75132
rect 8006 75052 8183 75080
rect 8155 74906 8296 74934
rect 8155 74854 8183 74906
rect 8006 74826 8183 74854
rect 8155 74780 8296 74808
rect 8155 74728 8183 74780
rect 8006 74700 8183 74728
rect 8155 73464 8296 73492
rect 8155 73396 8183 73464
rect 8006 73368 8183 73396
rect 8155 73338 8296 73366
rect 8155 73270 8183 73338
rect 8006 73242 8183 73270
rect 8155 73112 8296 73140
rect 8155 73044 8183 73112
rect 8006 73016 8183 73044
rect 8155 72052 8296 72080
rect 8155 72004 8183 72052
rect 8006 71976 8183 72004
rect 8155 71826 8296 71854
rect 8155 71778 8183 71826
rect 8006 71750 8183 71778
rect 8155 71700 8296 71728
rect 8155 71652 8183 71700
rect 8006 71624 8183 71652
rect 8155 70384 8296 70412
rect 8155 70320 8183 70384
rect 8006 70292 8183 70320
rect 8155 70258 8296 70286
rect 8155 70194 8183 70258
rect 8006 70166 8183 70194
rect 8155 70032 8296 70060
rect 8155 69968 8183 70032
rect 8006 69940 8183 69968
rect 8155 68972 8296 69000
rect 8155 68928 8183 68972
rect 8006 68900 8183 68928
rect 8155 68746 8296 68774
rect 8155 68702 8183 68746
rect 8006 68674 8183 68702
rect 8155 68620 8296 68648
rect 8155 68576 8183 68620
rect 8006 68548 8183 68576
rect 8155 67304 8296 67332
rect 8155 67244 8183 67304
rect 8006 67216 8183 67244
rect 8155 67178 8296 67206
rect 8155 67118 8183 67178
rect 8006 67090 8183 67118
rect 8155 66952 8296 66980
rect 8155 66892 8183 66952
rect 8006 66864 8183 66892
rect 8155 65892 8296 65920
rect 8155 65852 8183 65892
rect 8006 65824 8183 65852
rect 8155 65666 8296 65694
rect 8155 65626 8183 65666
rect 8006 65598 8183 65626
rect 8155 65540 8296 65568
rect 8155 65500 8183 65540
rect 8006 65472 8183 65500
rect 8155 64224 8296 64252
rect 8155 64168 8183 64224
rect 8006 64140 8183 64168
rect 8155 64098 8296 64126
rect 8155 64042 8183 64098
rect 8006 64014 8183 64042
rect 8155 63872 8296 63900
rect 8155 63816 8183 63872
rect 8006 63788 8183 63816
rect 8155 62812 8296 62840
rect 8155 62776 8183 62812
rect 8006 62748 8183 62776
rect 8155 62586 8296 62614
rect 8155 62550 8183 62586
rect 8006 62522 8183 62550
rect 8155 62460 8296 62488
rect 8155 62424 8183 62460
rect 8006 62396 8183 62424
rect 8155 61144 8296 61172
rect 8155 61092 8183 61144
rect 8006 61064 8183 61092
rect 8155 61018 8296 61046
rect 8155 60966 8183 61018
rect 8006 60938 8183 60966
rect 8155 60792 8296 60820
rect 8155 60740 8183 60792
rect 8006 60712 8183 60740
rect 8155 59732 8296 59760
rect 8155 59700 8183 59732
rect 8006 59672 8183 59700
rect 8155 59506 8296 59534
rect 8155 59474 8183 59506
rect 8006 59446 8183 59474
rect 8155 59380 8296 59408
rect 8155 59348 8183 59380
rect 8006 59320 8183 59348
rect 8155 58064 8296 58092
rect 8155 58016 8183 58064
rect 8006 57988 8183 58016
rect 8155 57938 8296 57966
rect 8155 57890 8183 57938
rect 8006 57862 8183 57890
rect 8155 57712 8296 57740
rect 8155 57664 8183 57712
rect 8006 57636 8183 57664
rect 8155 56652 8296 56680
rect 8155 56624 8183 56652
rect 8006 56596 8183 56624
rect 8155 56426 8296 56454
rect 8155 56398 8183 56426
rect 8006 56370 8183 56398
rect 8155 56300 8296 56328
rect 8155 56272 8183 56300
rect 8006 56244 8183 56272
rect 8155 54984 8296 55012
rect 8155 54940 8183 54984
rect 8006 54912 8183 54940
rect 8155 54858 8296 54886
rect 8155 54814 8183 54858
rect 8006 54786 8183 54814
rect 8155 54632 8296 54660
rect 8155 54588 8183 54632
rect 8006 54560 8183 54588
rect 8155 53572 8296 53600
rect 8155 53548 8183 53572
rect 8006 53520 8183 53548
rect 8155 53346 8296 53374
rect 8155 53322 8183 53346
rect 8006 53294 8183 53322
rect 8155 53220 8296 53248
rect 8155 53196 8183 53220
rect 8006 53168 8183 53196
rect 8155 51904 8296 51932
rect 8155 51864 8183 51904
rect 8006 51836 8183 51864
rect 8155 51778 8296 51806
rect 8155 51738 8183 51778
rect 8006 51710 8183 51738
rect 8155 51552 8296 51580
rect 8155 51512 8183 51552
rect 8006 51484 8183 51512
rect 8155 50492 8296 50520
rect 8155 50472 8183 50492
rect 8006 50444 8183 50472
rect 8155 50266 8296 50294
rect 8155 50246 8183 50266
rect 8006 50218 8183 50246
rect 8155 50140 8296 50168
rect 8155 50120 8183 50140
rect 8006 50092 8183 50120
rect 8155 48824 8296 48852
rect 8155 48788 8183 48824
rect 8006 48760 8183 48788
rect 8155 48698 8296 48726
rect 8155 48662 8183 48698
rect 8006 48634 8183 48662
rect 8155 48472 8296 48500
rect 8155 48436 8183 48472
rect 8006 48408 8183 48436
rect 8155 47412 8296 47440
rect 8155 47396 8183 47412
rect 8006 47368 8183 47396
rect 8155 47186 8296 47214
rect 8155 47170 8183 47186
rect 8006 47142 8183 47170
rect 8155 47060 8296 47088
rect 8155 47044 8183 47060
rect 8006 47016 8183 47044
rect 8155 45744 8296 45772
rect 8155 45712 8183 45744
rect 8006 45684 8183 45712
rect 8155 45618 8296 45646
rect 8155 45586 8183 45618
rect 8006 45558 8183 45586
rect 8155 45392 8296 45420
rect 8155 45360 8183 45392
rect 8006 45332 8183 45360
rect 8155 44332 8296 44360
rect 8155 44320 8183 44332
rect 8006 44292 8183 44320
rect 8155 44106 8296 44134
rect 8155 44094 8183 44106
rect 8006 44066 8183 44094
rect 8155 43980 8296 44008
rect 8155 43968 8183 43980
rect 8006 43940 8183 43968
rect 8155 42664 8296 42692
rect 8155 42636 8183 42664
rect 8006 42608 8183 42636
rect 8155 42538 8296 42566
rect 8155 42510 8183 42538
rect 8006 42482 8183 42510
rect 8155 42312 8296 42340
rect 8155 42284 8183 42312
rect 8006 42256 8183 42284
rect 8155 41252 8296 41280
rect 8155 41244 8183 41252
rect 8006 41216 8183 41244
rect 8155 41026 8296 41054
rect 8155 41018 8183 41026
rect 8006 40990 8183 41018
rect 8155 40900 8296 40928
rect 8155 40892 8183 40900
rect 8006 40864 8183 40892
rect 8155 39584 8296 39612
rect 8155 39560 8183 39584
rect 8006 39532 8183 39560
rect 8155 39458 8296 39486
rect 8155 39434 8183 39458
rect 8006 39406 8183 39434
rect 8155 39232 8296 39260
rect 8155 39208 8183 39232
rect 8006 39180 8183 39208
rect 8155 38172 8296 38200
rect 8155 38168 8183 38172
rect 8006 38140 8183 38168
rect 8155 37946 8296 37974
rect 8155 37942 8183 37946
rect 8006 37914 8183 37942
rect 8155 37820 8296 37848
rect 8155 37816 8183 37820
rect 8006 37788 8183 37816
rect 8155 36504 8296 36532
rect 8155 36484 8183 36504
rect 8006 36456 8183 36484
rect 8155 36378 8296 36406
rect 8155 36358 8183 36378
rect 8006 36330 8183 36358
rect 8155 36152 8296 36180
rect 8155 36132 8183 36152
rect 8006 36104 8183 36132
rect 8155 35092 8296 35120
rect 8006 35064 8183 35092
rect 8155 34866 8296 34894
rect 8006 34838 8183 34866
rect 8155 34740 8296 34768
rect 8006 34712 8183 34740
rect 8155 33424 8296 33452
rect 8155 33408 8183 33424
rect 8006 33380 8183 33408
rect 8155 33298 8296 33326
rect 8155 33282 8183 33298
rect 8006 33254 8183 33282
rect 8155 33072 8296 33100
rect 8155 33056 8183 33072
rect 8006 33028 8183 33056
rect 8155 32016 8296 32040
rect 8006 32012 8296 32016
rect 8006 31988 8183 32012
rect 8155 31790 8296 31814
rect 8006 31786 8296 31790
rect 8006 31762 8183 31786
rect 8155 31664 8296 31688
rect 8006 31660 8296 31664
rect 8006 31636 8183 31660
rect 8155 30344 8296 30372
rect 8155 30332 8183 30344
rect 8006 30304 8183 30332
rect 8155 30218 8296 30246
rect 8155 30206 8183 30218
rect 8006 30178 8183 30206
rect 8155 29992 8296 30020
rect 8155 29980 8183 29992
rect 8006 29952 8183 29980
rect 8155 28940 8296 28960
rect 8006 28932 8296 28940
rect 8006 28912 8183 28932
rect 8155 28714 8296 28734
rect 8006 28706 8296 28714
rect 8006 28686 8183 28706
rect 8155 28588 8296 28608
rect 8006 28580 8296 28588
rect 8006 28560 8183 28580
rect 8155 27264 8296 27292
rect 8155 27256 8183 27264
rect 8006 27228 8183 27256
rect 8155 27138 8296 27166
rect 8155 27130 8183 27138
rect 8006 27102 8183 27130
rect 8155 26912 8296 26940
rect 8155 26904 8183 26912
rect 8006 26876 8183 26904
rect 8155 25864 8296 25880
rect 8006 25852 8296 25864
rect 8006 25836 8183 25852
rect 8155 25638 8296 25654
rect 8006 25626 8296 25638
rect 8006 25610 8183 25626
rect 8155 25512 8296 25528
rect 8006 25500 8296 25512
rect 8006 25484 8183 25500
rect 8155 24184 8296 24212
rect 8155 24180 8183 24184
rect 8006 24152 8183 24180
rect 8155 24058 8296 24086
rect 8155 24054 8183 24058
rect 8006 24026 8183 24054
rect 8155 23832 8296 23860
rect 8155 23828 8183 23832
rect 8006 23800 8183 23828
rect 8155 22788 8296 22800
rect 8006 22772 8296 22788
rect 8006 22760 8183 22772
rect 8155 22562 8296 22574
rect 8006 22546 8296 22562
rect 8006 22534 8183 22546
rect 8155 22436 8296 22448
rect 8006 22420 8296 22436
rect 8006 22408 8183 22420
rect 8155 21104 8296 21132
rect 8006 21076 8183 21104
rect 8155 20978 8296 21006
rect 8006 20950 8183 20978
rect 8155 20752 8296 20780
rect 8006 20724 8183 20752
rect 8155 19712 8296 19720
rect 8006 19692 8296 19712
rect 8006 19684 8183 19692
rect 8155 19486 8296 19494
rect 8006 19466 8296 19486
rect 8006 19458 8183 19466
rect 8155 19360 8296 19368
rect 8006 19340 8296 19360
rect 8006 19332 8183 19340
rect 8155 18028 8296 18052
rect 8006 18024 8296 18028
rect 8006 18000 8183 18024
rect 8155 17902 8296 17926
rect 8006 17898 8296 17902
rect 8006 17874 8183 17898
rect 8155 17676 8296 17700
rect 8006 17672 8296 17676
rect 8006 17648 8183 17672
rect 8155 16636 8296 16640
rect 8006 16612 8296 16636
rect 8006 16608 8183 16612
rect 8155 16410 8296 16414
rect 8006 16386 8296 16410
rect 8006 16382 8183 16386
rect 8155 16284 8296 16288
rect 8006 16260 8296 16284
rect 8006 16256 8183 16260
rect 8155 14952 8296 14972
rect 8006 14944 8296 14952
rect 8006 14924 8183 14944
rect 8155 14826 8296 14846
rect 8006 14818 8296 14826
rect 8006 14798 8183 14818
rect 8155 14600 8296 14620
rect 8006 14592 8296 14600
rect 8006 14572 8183 14592
rect 8006 13532 8296 13560
rect 8006 13306 8296 13334
rect 8006 13180 8296 13208
rect 8155 11876 8296 11892
rect 8006 11864 8296 11876
rect 8006 11848 8183 11864
rect 8155 11750 8296 11766
rect 8006 11738 8296 11750
rect 8006 11722 8183 11738
rect 8155 11524 8296 11540
rect 8006 11512 8296 11524
rect 8006 11496 8183 11512
rect 8006 10480 8183 10484
rect 8006 10456 8296 10480
rect 8155 10452 8296 10456
rect 8006 10254 8183 10258
rect 8006 10230 8296 10254
rect 8155 10226 8296 10230
rect 8006 10128 8183 10132
rect 8006 10104 8296 10128
rect 8155 10100 8296 10104
rect 8155 8800 8296 8812
rect 8006 8784 8296 8800
rect 8006 8772 8183 8784
rect 8155 8674 8296 8686
rect 8006 8658 8296 8674
rect 8006 8646 8183 8658
rect 8155 8448 8296 8460
rect 8006 8432 8296 8448
rect 8006 8420 8183 8432
rect 8006 7400 8183 7408
rect 8006 7380 8296 7400
rect 8155 7372 8296 7380
rect 8006 7174 8183 7182
rect 8006 7154 8296 7174
rect 8155 7146 8296 7154
rect 8006 7048 8183 7056
rect 8006 7028 8296 7048
rect 8155 7020 8296 7028
rect 7906 5812 7912 5864
rect 7964 5852 7970 5864
rect 7964 5824 32958 5852
rect 7964 5812 7970 5824
rect 5850 5319 5856 5371
rect 5908 5319 5914 5371
rect 4776 4942 4782 4994
rect 4834 4982 4840 4994
rect 6166 4985 6224 4991
rect 6166 4982 6178 4985
rect 4834 4954 6178 4982
rect 4834 4942 4840 4954
rect 6166 4951 6178 4954
rect 6212 4951 6224 4985
rect 6166 4945 6224 4951
rect 5850 4481 5856 4533
rect 5908 4481 5914 4533
rect 4868 4020 4874 4072
rect 4926 4060 4932 4072
rect 6166 4063 6224 4069
rect 6166 4060 6178 4063
rect 4926 4032 6178 4060
rect 4926 4020 4932 4032
rect 6166 4029 6178 4032
rect 6212 4029 6224 4063
rect 6166 4023 6224 4029
rect 5850 3643 5856 3695
rect 5908 3643 5914 3695
rect 4868 3422 4874 3474
rect 4926 3462 4932 3474
rect 4926 3434 8310 3462
rect 4926 3422 4932 3434
rect 4776 3342 4782 3394
rect 4834 3382 4840 3394
rect 4834 3354 8310 3382
rect 4834 3342 4840 3354
rect 58380 1531 58386 1543
rect 33581 1503 58386 1531
rect 58380 1491 58386 1503
rect 58438 1491 58444 1543
<< via1 >>
rect 7912 5812 7964 5864
rect 5856 5362 5908 5371
rect 5856 5328 5865 5362
rect 5865 5328 5899 5362
rect 5899 5328 5908 5362
rect 5856 5319 5908 5328
rect 4782 4942 4834 4994
rect 5856 4524 5908 4533
rect 5856 4490 5865 4524
rect 5865 4490 5899 4524
rect 5899 4490 5908 4524
rect 5856 4481 5908 4490
rect 4874 4020 4926 4072
rect 5856 3686 5908 3695
rect 5856 3652 5865 3686
rect 5865 3652 5899 3686
rect 5899 3652 5908 3686
rect 5856 3643 5908 3652
rect 4874 3422 4926 3474
rect 4782 3342 4834 3394
rect 58386 1491 58438 1543
<< metal2 >>
rect 6802 104794 6830 104822
rect 18 6376 46 43328
rect 102 6376 130 43328
rect 186 6376 214 43328
rect 270 6376 298 43328
rect 354 6376 382 43328
rect 438 6376 466 43328
rect 522 6376 550 43328
rect 606 6376 634 43328
rect 7924 5870 7952 5956
rect 8881 5908 8935 5936
rect 10437 5908 10491 5936
rect 11993 5908 12047 5936
rect 13549 5908 13603 5936
rect 15105 5908 15159 5936
rect 16661 5908 16715 5936
rect 18217 5908 18271 5936
rect 19773 5908 19827 5936
rect 21329 5908 21383 5936
rect 22885 5908 22939 5936
rect 24441 5908 24495 5936
rect 25997 5908 26051 5936
rect 27553 5908 27607 5936
rect 29109 5908 29163 5936
rect 30665 5908 30719 5936
rect 32221 5908 32275 5936
rect 33777 5908 33831 5936
rect 35333 5908 35387 5936
rect 36889 5908 36943 5936
rect 38445 5908 38499 5936
rect 40001 5908 40055 5936
rect 41557 5908 41611 5936
rect 43113 5908 43167 5936
rect 44669 5908 44723 5936
rect 46225 5908 46279 5936
rect 47781 5908 47835 5936
rect 49337 5908 49391 5936
rect 50893 5908 50947 5936
rect 52449 5908 52503 5936
rect 54005 5908 54059 5936
rect 55561 5908 55615 5936
rect 57117 5908 57171 5936
rect 7912 5864 7964 5870
rect 7912 5806 7964 5812
rect 5854 5373 5910 5382
rect 5854 5308 5910 5317
rect 4782 4994 4834 5000
rect 4782 4936 4834 4942
rect 4794 3400 4822 4936
rect 5854 4535 5910 4544
rect 5854 4470 5910 4479
rect 4874 4072 4926 4078
rect 4874 4014 4926 4020
rect 4886 3480 4914 4014
rect 5854 3697 5910 3706
rect 5854 3632 5910 3641
rect 4874 3474 4926 3480
rect 4874 3416 4926 3422
rect 4782 3394 4834 3400
rect 4782 3336 4834 3342
rect 7924 0 7952 5806
rect 8615 4764 8643 5004
rect 8887 4764 8915 5004
rect 10171 4764 10199 5004
rect 10443 4764 10471 5004
rect 11727 4764 11755 5004
rect 11999 4764 12027 5004
rect 13283 4764 13311 5004
rect 13555 4764 13583 5004
rect 14839 4764 14867 5004
rect 15111 4764 15139 5004
rect 16395 4764 16423 5004
rect 16667 4764 16695 5004
rect 17951 4764 17979 5004
rect 18223 4764 18251 5004
rect 19507 4764 19535 5004
rect 19779 4764 19807 5004
rect 21063 4764 21091 5004
rect 21335 4764 21363 5004
rect 22619 4764 22647 5004
rect 22891 4764 22919 5004
rect 24175 4764 24203 5004
rect 24447 4764 24475 5004
rect 25731 4764 25759 5004
rect 26003 4764 26031 5004
rect 27287 4764 27315 5004
rect 27559 4764 27587 5004
rect 28843 4764 28871 5004
rect 29115 4764 29143 5004
rect 30399 4764 30427 5004
rect 30671 4764 30699 5004
rect 31955 4764 31983 5004
rect 32227 4764 32255 5004
rect 58398 1549 58426 105020
rect 58386 1543 58438 1549
rect 58386 1485 58438 1491
rect 58398 0 58426 1485
<< via2 >>
rect 5854 5371 5910 5373
rect 5854 5319 5856 5371
rect 5856 5319 5908 5371
rect 5908 5319 5910 5371
rect 5854 5317 5910 5319
rect 5854 4533 5910 4535
rect 5854 4481 5856 4533
rect 5856 4481 5908 4533
rect 5908 4481 5910 4533
rect 5854 4479 5910 4481
rect 5854 3695 5910 3697
rect 5854 3643 5856 3695
rect 5856 3643 5908 3695
rect 5908 3643 5910 3695
rect 5854 3641 5910 3643
<< metal3 >>
rect 6400 104771 6532 104845
rect 7940 104771 8072 104845
rect 6400 103233 6532 103307
rect 7940 103233 8072 103307
rect 6400 101695 6532 101769
rect 7940 101695 8072 101769
rect 6400 100157 6532 100231
rect 7940 100157 8072 100231
rect 6400 98619 6532 98693
rect 7940 98619 8072 98693
rect 6400 97081 6532 97155
rect 7940 97081 8072 97155
rect 6400 95543 6532 95617
rect 7940 95543 8072 95617
rect 6400 94005 6532 94079
rect 7940 94005 8072 94079
rect 6400 92467 6532 92541
rect 7940 92467 8072 92541
rect 6400 90929 6532 91003
rect 7940 90929 8072 91003
rect 6400 89391 6532 89465
rect 7940 89391 8072 89465
rect 6400 87853 6532 87927
rect 7940 87853 8072 87927
rect 6400 86315 6532 86389
rect 7940 86315 8072 86389
rect 6400 84777 6532 84851
rect 7940 84777 8072 84851
rect 6400 83239 6532 83313
rect 7940 83239 8072 83313
rect 6400 81701 6532 81775
rect 7940 81701 8072 81775
rect 6400 80163 6532 80237
rect 7940 80163 8072 80237
rect 6400 78625 6532 78699
rect 7940 78625 8072 78699
rect 6400 77087 6532 77161
rect 7940 77087 8072 77161
rect 6400 75549 6532 75623
rect 7940 75549 8072 75623
rect 6400 74011 6532 74085
rect 7940 74011 8072 74085
rect 6400 72473 6532 72547
rect 7940 72473 8072 72547
rect 6400 70935 6532 71009
rect 7940 70935 8072 71009
rect 6400 69397 6532 69471
rect 7940 69397 8072 69471
rect 6400 67859 6532 67933
rect 7940 67859 8072 67933
rect 6400 66321 6532 66395
rect 7940 66321 8072 66395
rect 6400 64783 6532 64857
rect 7940 64783 8072 64857
rect 6400 63245 6532 63319
rect 7940 63245 8072 63319
rect 6400 61707 6532 61781
rect 7940 61707 8072 61781
rect 6400 60169 6532 60243
rect 7940 60169 8072 60243
rect 6400 58631 6532 58705
rect 7940 58631 8072 58705
rect 6400 57093 6532 57167
rect 7940 57093 8072 57167
rect 6400 55555 6532 55629
rect 7940 55555 8072 55629
rect 6400 54017 6532 54091
rect 7940 54017 8072 54091
rect 6400 52479 6532 52553
rect 7940 52479 8072 52553
rect 6400 50941 6532 51015
rect 7940 50941 8072 51015
rect 6400 49403 6532 49477
rect 7940 49403 8072 49477
rect 6400 47865 6532 47939
rect 7940 47865 8072 47939
rect 6400 46327 6532 46401
rect 7940 46327 8072 46401
rect 6400 44789 6532 44863
rect 7940 44789 8072 44863
rect 1044 43291 1176 43365
rect 2084 43291 2216 43365
rect 6400 43251 6532 43325
rect 7940 43251 8072 43325
rect 1044 41751 1176 41825
rect 2084 41751 2216 41825
rect 6400 41713 6532 41787
rect 7940 41713 8072 41787
rect 1044 40211 1176 40285
rect 2084 40211 2216 40285
rect 6400 40175 6532 40249
rect 7940 40175 8072 40249
rect 1044 38671 1176 38745
rect 2084 38671 2216 38745
rect 6400 38637 6532 38711
rect 7940 38637 8072 38711
rect 1044 37131 1176 37205
rect 2084 37131 2216 37205
rect 6400 37099 6532 37173
rect 7940 37099 8072 37173
rect 1044 35591 1176 35665
rect 2084 35591 2216 35665
rect 6400 35561 6532 35635
rect 7940 35561 8072 35635
rect 1044 34051 1176 34125
rect 2084 34051 2216 34125
rect 6400 34023 6532 34097
rect 7940 34023 8072 34097
rect 1044 32511 1176 32585
rect 2084 32511 2216 32585
rect 6400 32485 6532 32559
rect 7940 32485 8072 32559
rect 1044 30971 1176 31045
rect 2084 30971 2216 31045
rect 6400 30947 6532 31021
rect 7940 30947 8072 31021
rect 6400 29409 6532 29483
rect 7940 29409 8072 29483
rect 1044 27895 1176 27969
rect 2084 27895 2216 27969
rect 6400 27871 6532 27945
rect 7940 27871 8072 27945
rect 1044 26355 1176 26429
rect 2084 26355 2216 26429
rect 6400 26333 6532 26407
rect 7940 26333 8072 26407
rect 1044 24815 1176 24889
rect 2084 24815 2216 24889
rect 6400 24795 6532 24869
rect 7940 24795 8072 24869
rect 1044 23275 1176 23349
rect 2084 23275 2216 23349
rect 6400 23257 6532 23331
rect 7940 23257 8072 23331
rect 1044 21735 1176 21809
rect 2084 21735 2216 21809
rect 6400 21719 6532 21793
rect 7940 21719 8072 21793
rect 1044 20195 1176 20269
rect 2084 20195 2216 20269
rect 6400 20181 6532 20255
rect 7940 20181 8072 20255
rect 1044 18655 1176 18729
rect 2084 18655 2216 18729
rect 6400 18643 6532 18717
rect 7940 18643 8072 18717
rect 1044 17115 1176 17189
rect 2084 17115 2216 17189
rect 6400 17105 6532 17179
rect 7940 17105 8072 17179
rect 1044 15575 1176 15649
rect 2084 15575 2216 15649
rect 6400 15567 6532 15641
rect 7940 15567 8072 15641
rect 6400 14029 6532 14103
rect 7940 14029 8072 14103
rect 1392 12499 1524 12573
rect 2264 12499 2396 12573
rect 6400 12491 6532 12565
rect 7940 12491 8072 12565
rect 1392 10959 1524 11033
rect 2264 10959 2396 11033
rect 6400 10953 6532 11027
rect 7940 10953 8072 11027
rect 1392 9419 1524 9493
rect 2264 9419 2396 9493
rect 6400 9415 6532 9489
rect 7940 9415 8072 9489
rect 1392 7879 1524 7953
rect 2264 7879 2396 7953
rect 6400 7877 6532 7951
rect 7940 7877 8072 7951
rect 1392 6339 1524 6413
rect 2264 6339 2396 6413
rect 6400 6339 6532 6413
rect 7940 6339 8072 6413
rect 9001 6100 9067 6232
rect 10557 6100 10623 6232
rect 12113 6100 12179 6232
rect 13669 6100 13735 6232
rect 15225 6100 15291 6232
rect 16781 6100 16847 6232
rect 18337 6100 18403 6232
rect 19893 6100 19959 6232
rect 21449 6100 21515 6232
rect 23005 6100 23071 6232
rect 24561 6100 24627 6232
rect 26117 6100 26183 6232
rect 27673 6100 27739 6232
rect 29229 6100 29295 6232
rect 30785 6100 30851 6232
rect 32341 6100 32407 6232
rect 33897 6100 33963 6232
rect 35453 6100 35519 6232
rect 37009 6100 37075 6232
rect 38565 6100 38631 6232
rect 40121 6100 40187 6232
rect 41677 6100 41743 6232
rect 43233 6100 43299 6232
rect 44789 6100 44855 6232
rect 46345 6100 46411 6232
rect 47901 6100 47967 6232
rect 49457 6100 49523 6232
rect 51013 6100 51079 6232
rect 52569 6100 52635 6232
rect 54125 6100 54191 6232
rect 55681 6100 55747 6232
rect 57237 6100 57303 6232
rect 5816 5373 5948 5382
rect 5816 5317 5854 5373
rect 5910 5317 5948 5373
rect 5816 5308 5948 5317
rect 9001 5268 9067 5400
rect 10557 5268 10623 5400
rect 12113 5268 12179 5400
rect 13669 5268 13735 5400
rect 15225 5268 15291 5400
rect 16781 5268 16847 5400
rect 18337 5268 18403 5400
rect 19893 5268 19959 5400
rect 21449 5268 21515 5400
rect 23005 5268 23071 5400
rect 24561 5268 24627 5400
rect 26117 5268 26183 5400
rect 27673 5268 27739 5400
rect 29229 5268 29295 5400
rect 30785 5268 30851 5400
rect 32341 5268 32407 5400
rect 33897 5268 33963 5400
rect 35453 5268 35519 5400
rect 37009 5268 37075 5400
rect 38565 5268 38631 5400
rect 40121 5268 40187 5400
rect 41677 5268 41743 5400
rect 43233 5268 43299 5400
rect 44789 5268 44855 5400
rect 46345 5268 46411 5400
rect 47901 5268 47967 5400
rect 49457 5268 49523 5400
rect 51013 5268 51079 5400
rect 52569 5268 52635 5400
rect 54125 5268 54191 5400
rect 55681 5268 55747 5400
rect 57237 5268 57303 5400
rect 8483 4933 8615 5007
rect 8755 4933 8887 5007
rect 10039 4933 10171 5007
rect 10311 4933 10443 5007
rect 11595 4933 11727 5007
rect 11867 4933 11999 5007
rect 13151 4933 13283 5007
rect 13423 4933 13555 5007
rect 14707 4933 14839 5007
rect 14979 4933 15111 5007
rect 16263 4933 16395 5007
rect 16535 4933 16667 5007
rect 17819 4933 17951 5007
rect 18091 4933 18223 5007
rect 19375 4933 19507 5007
rect 19647 4933 19779 5007
rect 20931 4933 21063 5007
rect 21203 4933 21335 5007
rect 22487 4933 22619 5007
rect 22759 4933 22891 5007
rect 24043 4933 24175 5007
rect 24315 4933 24447 5007
rect 25599 4933 25731 5007
rect 25871 4933 26003 5007
rect 27155 4933 27287 5007
rect 27427 4933 27559 5007
rect 28711 4933 28843 5007
rect 28983 4933 29115 5007
rect 30267 4933 30399 5007
rect 30539 4933 30671 5007
rect 31823 4933 31955 5007
rect 32095 4933 32227 5007
rect 33379 4933 33511 5007
rect 33651 4933 33783 5007
rect 34935 4933 35067 5007
rect 35207 4933 35339 5007
rect 36491 4933 36623 5007
rect 36763 4933 36895 5007
rect 38047 4933 38179 5007
rect 38319 4933 38451 5007
rect 39603 4933 39735 5007
rect 39875 4933 40007 5007
rect 41159 4933 41291 5007
rect 41431 4933 41563 5007
rect 42715 4933 42847 5007
rect 42987 4933 43119 5007
rect 44271 4933 44403 5007
rect 44543 4933 44675 5007
rect 45827 4933 45959 5007
rect 46099 4933 46231 5007
rect 47383 4933 47515 5007
rect 47655 4933 47787 5007
rect 48939 4933 49071 5007
rect 49211 4933 49343 5007
rect 50495 4933 50627 5007
rect 50767 4933 50899 5007
rect 52051 4933 52183 5007
rect 52323 4933 52455 5007
rect 53607 4933 53739 5007
rect 53879 4933 54011 5007
rect 55163 4933 55295 5007
rect 55435 4933 55567 5007
rect 56719 4933 56851 5007
rect 56991 4933 57123 5007
rect 5816 4535 5948 4544
rect 5816 4479 5854 4535
rect 5910 4479 5948 4535
rect 5816 4470 5948 4479
rect 8483 3987 8615 4061
rect 8755 3987 8887 4061
rect 10039 3987 10171 4061
rect 10311 3987 10443 4061
rect 11595 3987 11727 4061
rect 11867 3987 11999 4061
rect 13151 3987 13283 4061
rect 13423 3987 13555 4061
rect 14707 3987 14839 4061
rect 14979 3987 15111 4061
rect 16263 3987 16395 4061
rect 16535 3987 16667 4061
rect 17819 3987 17951 4061
rect 18091 3987 18223 4061
rect 19375 3987 19507 4061
rect 19647 3987 19779 4061
rect 20931 3987 21063 4061
rect 21203 3987 21335 4061
rect 22487 3987 22619 4061
rect 22759 3987 22891 4061
rect 24043 3987 24175 4061
rect 24315 3987 24447 4061
rect 25599 3987 25731 4061
rect 25871 3987 26003 4061
rect 27155 3987 27287 4061
rect 27427 3987 27559 4061
rect 28711 3987 28843 4061
rect 28983 3987 29115 4061
rect 30267 3987 30399 4061
rect 30539 3987 30671 4061
rect 31823 3987 31955 4061
rect 32095 3987 32227 4061
rect 33379 3987 33511 4061
rect 33651 3987 33783 4061
rect 34935 3987 35067 4061
rect 35207 3987 35339 4061
rect 36491 3987 36623 4061
rect 36763 3987 36895 4061
rect 38047 3987 38179 4061
rect 38319 3987 38451 4061
rect 39603 3987 39735 4061
rect 39875 3987 40007 4061
rect 41159 3987 41291 4061
rect 41431 3987 41563 4061
rect 42715 3987 42847 4061
rect 42987 3987 43119 4061
rect 44271 3987 44403 4061
rect 44543 3987 44675 4061
rect 45827 3987 45959 4061
rect 46099 3987 46231 4061
rect 47383 3987 47515 4061
rect 47655 3987 47787 4061
rect 48939 3987 49071 4061
rect 49211 3987 49343 4061
rect 50495 3987 50627 4061
rect 50767 3987 50899 4061
rect 52051 3987 52183 4061
rect 52323 3987 52455 4061
rect 53607 3987 53739 4061
rect 53879 3987 54011 4061
rect 55163 3987 55295 4061
rect 55435 3987 55567 4061
rect 56719 3987 56851 4061
rect 56991 3987 57123 4061
rect 5816 3697 5948 3706
rect 5816 3641 5854 3697
rect 5910 3641 5948 3697
rect 5816 3632 5948 3641
rect 9008 2506 9140 2580
rect 9786 2506 9918 2580
rect 10564 2506 10696 2580
rect 11342 2506 11474 2580
rect 12120 2506 12252 2580
rect 12898 2506 13030 2580
rect 13676 2506 13808 2580
rect 14454 2506 14586 2580
rect 15232 2506 15364 2580
rect 16010 2506 16142 2580
rect 16788 2506 16920 2580
rect 17566 2506 17698 2580
rect 18344 2506 18476 2580
rect 19122 2506 19254 2580
rect 19900 2506 20032 2580
rect 20678 2506 20810 2580
rect 21456 2506 21588 2580
rect 22234 2506 22366 2580
rect 23012 2506 23144 2580
rect 23790 2506 23922 2580
rect 24568 2506 24700 2580
rect 25346 2506 25478 2580
rect 26124 2506 26256 2580
rect 26902 2506 27034 2580
rect 27680 2506 27812 2580
rect 28458 2506 28590 2580
rect 29236 2506 29368 2580
rect 30014 2506 30146 2580
rect 30792 2506 30924 2580
rect 31570 2506 31702 2580
rect 32348 2506 32480 2580
rect 33126 2506 33258 2580
rect 33904 2506 34036 2580
rect 34682 2506 34814 2580
rect 35460 2506 35592 2580
rect 36238 2506 36370 2580
rect 37016 2506 37148 2580
rect 37794 2506 37926 2580
rect 38572 2506 38704 2580
rect 39350 2506 39482 2580
rect 40128 2506 40260 2580
rect 40906 2506 41038 2580
rect 41684 2506 41816 2580
rect 42462 2506 42594 2580
rect 43240 2506 43372 2580
rect 44018 2506 44150 2580
rect 44796 2506 44928 2580
rect 45574 2506 45706 2580
rect 46352 2506 46484 2580
rect 47130 2506 47262 2580
rect 47908 2506 48040 2580
rect 48686 2506 48818 2580
rect 49464 2506 49596 2580
rect 50242 2506 50374 2580
rect 51020 2506 51152 2580
rect 51798 2506 51930 2580
rect 52576 2506 52708 2580
rect 53354 2506 53486 2580
rect 54132 2506 54264 2580
rect 54910 2506 55042 2580
rect 55688 2506 55820 2580
rect 56466 2506 56598 2580
rect 57244 2506 57376 2580
rect 58022 2506 58154 2580
rect 8456 548 8522 680
rect 9234 548 9300 680
rect 10012 548 10078 680
rect 10790 548 10856 680
rect 11568 548 11634 680
rect 12346 548 12412 680
rect 13124 548 13190 680
rect 13902 548 13968 680
rect 14680 548 14746 680
rect 15458 548 15524 680
rect 16236 548 16302 680
rect 17014 548 17080 680
rect 17792 548 17858 680
rect 18570 548 18636 680
rect 19348 548 19414 680
rect 20126 548 20192 680
rect 20904 548 20970 680
rect 21682 548 21748 680
rect 22460 548 22526 680
rect 23238 548 23304 680
rect 24016 548 24082 680
rect 24794 548 24860 680
rect 25572 548 25638 680
rect 26350 548 26416 680
rect 27128 548 27194 680
rect 27906 548 27972 680
rect 28684 548 28750 680
rect 29462 548 29528 680
rect 30240 548 30306 680
rect 31018 548 31084 680
rect 31796 548 31862 680
rect 32574 548 32640 680
rect 33352 548 33418 680
rect 34130 548 34196 680
rect 34908 548 34974 680
rect 35686 548 35752 680
rect 36464 548 36530 680
rect 37242 548 37308 680
rect 38020 548 38086 680
rect 38798 548 38864 680
rect 39576 548 39642 680
rect 40354 548 40420 680
rect 41132 548 41198 680
rect 41910 548 41976 680
rect 42688 548 42754 680
rect 43466 548 43532 680
rect 44244 548 44310 680
rect 45022 548 45088 680
rect 45800 548 45866 680
rect 46578 548 46644 680
rect 47356 548 47422 680
rect 48134 548 48200 680
rect 48912 548 48978 680
rect 49690 548 49756 680
rect 50468 548 50534 680
rect 51246 548 51312 680
rect 52024 548 52090 680
rect 52802 548 52868 680
rect 53580 548 53646 680
rect 54358 548 54424 680
rect 55136 548 55202 680
rect 55914 548 55980 680
rect 56692 548 56758 680
rect 57470 548 57536 680
rect 58248 548 58314 680
use contact_18  contact_18_0
timestamp 1644969367
transform 1 0 5816 0 1 5308
box 0 0 1 1
use contact_17  contact_17_0
timestamp 1644969367
transform 1 0 5850 0 1 5313
box 0 0 1 1
use contact_13  contact_13_0
timestamp 1644969367
transform 1 0 5853 0 1 5322
box 0 0 1 1
use contact_18  contact_18_1
timestamp 1644969367
transform 1 0 5816 0 1 3632
box 0 0 1 1
use contact_17  contact_17_1
timestamp 1644969367
transform 1 0 5850 0 1 3637
box 0 0 1 1
use contact_13  contact_13_1
timestamp 1644969367
transform 1 0 5853 0 1 3646
box 0 0 1 1
use contact_18  contact_18_2
timestamp 1644969367
transform 1 0 5816 0 1 4470
box 0 0 1 1
use contact_17  contact_17_2
timestamp 1644969367
transform 1 0 5850 0 1 4475
box 0 0 1 1
use contact_13  contact_13_2
timestamp 1644969367
transform 1 0 5853 0 1 4484
box 0 0 1 1
use contact_17  contact_17_3
timestamp 1644969367
transform 1 0 58380 0 1 1485
box 0 0 1 1
use contact_17  contact_17_4
timestamp 1644969367
transform 1 0 7906 0 1 5806
box 0 0 1 1
use contact_17  contact_17_5
timestamp 1644969367
transform 1 0 4868 0 1 3416
box 0 0 1 1
use contact_13  contact_13_3
timestamp 1644969367
transform 1 0 6166 0 1 4023
box 0 0 1 1
use contact_17  contact_17_6
timestamp 1644969367
transform 1 0 4868 0 1 4014
box 0 0 1 1
use contact_17  contact_17_7
timestamp 1644969367
transform 1 0 4776 0 1 3336
box 0 0 1 1
use contact_13  contact_13_4
timestamp 1644969367
transform 1 0 6166 0 1 4945
box 0 0 1 1
use contact_17  contact_17_8
timestamp 1644969367
transform 1 0 4776 0 1 4936
box 0 0 1 1
use pinvbuf  pinvbuf_0
timestamp 1644969367
transform 1 0 5060 0 1 3652
box -36 0 1644 1710
use port_address  port_address_0
timestamp 1644969367
transform 1 0 0 0 1 6376
box 0 -42 8072 98474
use port_data  port_data_0
timestamp 1644969367
transform 1 0 8296 0 1 0
box 0 490 50570 6232
use replica_bitcell_array  replica_bitcell_array_0
timestamp 1644969367
transform 1 0 8296 0 1 6376
box 0 -42 49792 98602
<< labels >>
rlabel metal2 s 7924 0 7952 5956 4 w_en
rlabel metal2 s 6802 104794 6830 104822 4 wl_en
rlabel metal2 s 58398 0 58426 105020 4 p_en_bar
rlabel metal2 s 8880 5908 8934 5936 4 din0_0
rlabel metal2 s 10436 5908 10490 5936 4 din0_1
rlabel metal2 s 11992 5908 12046 5936 4 din0_2
rlabel metal2 s 13548 5908 13602 5936 4 din0_3
rlabel metal2 s 15104 5908 15158 5936 4 din0_4
rlabel metal2 s 16660 5908 16714 5936 4 din0_5
rlabel metal2 s 18216 5908 18270 5936 4 din0_6
rlabel metal2 s 19772 5908 19826 5936 4 din0_7
rlabel metal2 s 21328 5908 21382 5936 4 din0_8
rlabel metal2 s 22884 5908 22938 5936 4 din0_9
rlabel metal2 s 24440 5908 24494 5936 4 din0_10
rlabel metal2 s 25996 5908 26050 5936 4 din0_11
rlabel metal2 s 27552 5908 27606 5936 4 din0_12
rlabel metal2 s 29108 5908 29162 5936 4 din0_13
rlabel metal2 s 30664 5908 30718 5936 4 din0_14
rlabel metal2 s 32220 5908 32274 5936 4 din0_15
rlabel metal2 s 33776 5908 33830 5936 4 din0_16
rlabel metal2 s 35332 5908 35386 5936 4 din0_17
rlabel metal2 s 36888 5908 36942 5936 4 din0_18
rlabel metal2 s 38444 5908 38498 5936 4 din0_19
rlabel metal2 s 40000 5908 40054 5936 4 din0_20
rlabel metal2 s 41556 5908 41610 5936 4 din0_21
rlabel metal2 s 43112 5908 43166 5936 4 din0_22
rlabel metal2 s 44668 5908 44722 5936 4 din0_23
rlabel metal2 s 46224 5908 46278 5936 4 din0_24
rlabel metal2 s 47780 5908 47834 5936 4 din0_25
rlabel metal2 s 49336 5908 49390 5936 4 din0_26
rlabel metal2 s 50892 5908 50946 5936 4 din0_27
rlabel metal2 s 52448 5908 52502 5936 4 din0_28
rlabel metal2 s 54004 5908 54058 5936 4 din0_29
rlabel metal2 s 55560 5908 55614 5936 4 din0_30
rlabel metal2 s 57116 5908 57170 5936 4 din0_31
rlabel metal2 s 8614 4764 8642 5004 4 dout0_0
rlabel metal2 s 8629 4884 8629 4884 4 dout1_0
rlabel metal2 s 8886 4764 8914 5004 4 dout0_1
rlabel metal2 s 8901 4884 8901 4884 4 dout1_1
rlabel metal2 s 10170 4764 10198 5004 4 dout0_2
rlabel metal2 s 10185 4884 10185 4884 4 dout1_2
rlabel metal2 s 10442 4764 10470 5004 4 dout0_3
rlabel metal2 s 10457 4884 10457 4884 4 dout1_3
rlabel metal2 s 11726 4764 11754 5004 4 dout0_4
rlabel metal2 s 11741 4884 11741 4884 4 dout1_4
rlabel metal2 s 11998 4764 12026 5004 4 dout0_5
rlabel metal2 s 12013 4884 12013 4884 4 dout1_5
rlabel metal2 s 13282 4764 13310 5004 4 dout0_6
rlabel metal2 s 13297 4884 13297 4884 4 dout1_6
rlabel metal2 s 13554 4764 13582 5004 4 dout0_7
rlabel metal2 s 13569 4884 13569 4884 4 dout1_7
rlabel metal2 s 14838 4764 14866 5004 4 dout0_8
rlabel metal2 s 14853 4884 14853 4884 4 dout1_8
rlabel metal2 s 15110 4764 15138 5004 4 dout0_9
rlabel metal2 s 15125 4884 15125 4884 4 dout1_9
rlabel metal2 s 16394 4764 16422 5004 4 dout0_10
rlabel metal2 s 16409 4884 16409 4884 4 dout1_10
rlabel metal2 s 16666 4764 16694 5004 4 dout0_11
rlabel metal2 s 16681 4884 16681 4884 4 dout1_11
rlabel metal2 s 17950 4764 17978 5004 4 dout0_12
rlabel metal2 s 17965 4884 17965 4884 4 dout1_12
rlabel metal2 s 18222 4764 18250 5004 4 dout0_13
rlabel metal2 s 18237 4884 18237 4884 4 dout1_13
rlabel metal2 s 19506 4764 19534 5004 4 dout0_14
rlabel metal2 s 19521 4884 19521 4884 4 dout1_14
rlabel metal2 s 19778 4764 19806 5004 4 dout0_15
rlabel metal2 s 19793 4884 19793 4884 4 dout1_15
rlabel metal2 s 21062 4764 21090 5004 4 dout0_16
rlabel metal2 s 21077 4884 21077 4884 4 dout1_16
rlabel metal2 s 21334 4764 21362 5004 4 dout0_17
rlabel metal2 s 21349 4884 21349 4884 4 dout1_17
rlabel metal2 s 22618 4764 22646 5004 4 dout0_18
rlabel metal2 s 22633 4884 22633 4884 4 dout1_18
rlabel metal2 s 22890 4764 22918 5004 4 dout0_19
rlabel metal2 s 22905 4884 22905 4884 4 dout1_19
rlabel metal2 s 24174 4764 24202 5004 4 dout0_20
rlabel metal2 s 24189 4884 24189 4884 4 dout1_20
rlabel metal2 s 24446 4764 24474 5004 4 dout0_21
rlabel metal2 s 24461 4884 24461 4884 4 dout1_21
rlabel metal2 s 25730 4764 25758 5004 4 dout0_22
rlabel metal2 s 25745 4884 25745 4884 4 dout1_22
rlabel metal2 s 26002 4764 26030 5004 4 dout0_23
rlabel metal2 s 26017 4884 26017 4884 4 dout1_23
rlabel metal2 s 27286 4764 27314 5004 4 dout0_24
rlabel metal2 s 27301 4884 27301 4884 4 dout1_24
rlabel metal2 s 27558 4764 27586 5004 4 dout0_25
rlabel metal2 s 27573 4884 27573 4884 4 dout1_25
rlabel metal2 s 28842 4764 28870 5004 4 dout0_26
rlabel metal2 s 28857 4884 28857 4884 4 dout1_26
rlabel metal2 s 29114 4764 29142 5004 4 dout0_27
rlabel metal2 s 29129 4884 29129 4884 4 dout1_27
rlabel metal2 s 30398 4764 30426 5004 4 dout0_28
rlabel metal2 s 30413 4884 30413 4884 4 dout1_28
rlabel metal2 s 30670 4764 30698 5004 4 dout0_29
rlabel metal2 s 30685 4884 30685 4884 4 dout1_29
rlabel metal2 s 31954 4764 31982 5004 4 dout0_30
rlabel metal2 s 31969 4884 31969 4884 4 dout1_30
rlabel metal2 s 32226 4764 32254 5004 4 dout0_31
rlabel metal2 s 32241 4884 32241 4884 4 dout1_31
rlabel metal2 s 18 6376 46 43328 4 addr1
rlabel metal2 s 102 6376 130 43328 4 addr2
rlabel metal2 s 186 6376 214 43328 4 addr3
rlabel metal2 s 270 6376 298 43328 4 addr4
rlabel metal2 s 354 6376 382 43328 4 addr5
rlabel metal2 s 438 6376 466 43328 4 addr6
rlabel metal2 s 522 6376 550 43328 4 addr7
rlabel metal2 s 606 6376 634 43328 4 addr8
rlabel locali s 5141 4046 5141 4046 4 addr0
rlabel metal3 s 27672 5268 27738 5400 4 vdd
rlabel metal3 s 8456 548 8522 680 4 vdd
rlabel metal3 s 42714 3986 42846 4060 4 vdd
rlabel metal3 s 31796 548 31862 680 4 vdd
rlabel metal3 s 1044 32510 1176 32584 4 vdd
rlabel metal3 s 7940 17104 8072 17178 4 vdd
rlabel metal3 s 8482 3986 8614 4060 4 vdd
rlabel metal3 s 55434 3986 55566 4060 4 vdd
rlabel metal3 s 54358 548 54424 680 4 vdd
rlabel metal3 s 1392 10958 1524 11032 4 vdd
rlabel metal3 s 6400 84776 6532 84850 4 vdd
rlabel metal3 s 7940 100156 8072 100230 4 vdd
rlabel metal3 s 13902 548 13968 680 4 vdd
rlabel metal3 s 7940 7876 8072 7950 4 vdd
rlabel metal3 s 24042 3986 24174 4060 4 vdd
rlabel metal3 s 45022 548 45088 680 4 vdd
rlabel metal3 s 6400 50940 6532 51014 4 vdd
rlabel metal3 s 26350 548 26416 680 4 vdd
rlabel metal3 s 7940 20180 8072 20254 4 vdd
rlabel metal3 s 27154 3986 27286 4060 4 vdd
rlabel metal3 s 6400 44788 6532 44862 4 vdd
rlabel metal3 s 7940 54016 8072 54090 4 vdd
rlabel metal3 s 50494 3986 50626 4060 4 vdd
rlabel metal3 s 32094 3986 32226 4060 4 vdd
rlabel metal3 s 32574 548 32640 680 4 vdd
rlabel metal3 s 44788 5268 44854 5400 4 vdd
rlabel metal3 s 31018 548 31084 680 4 vdd
rlabel metal3 s 6400 69396 6532 69470 4 vdd
rlabel metal3 s 18336 5268 18402 5400 4 vdd
rlabel metal3 s 47654 3986 47786 4060 4 vdd
rlabel metal3 s 47356 548 47422 680 4 vdd
rlabel metal3 s 5816 4470 5948 4544 4 vdd
rlabel metal3 s 22758 3986 22890 4060 4 vdd
rlabel metal3 s 16534 3986 16666 4060 4 vdd
rlabel metal3 s 57236 5268 57302 5400 4 vdd
rlabel metal3 s 11866 3986 11998 4060 4 vdd
rlabel metal3 s 43466 548 43532 680 4 vdd
rlabel metal3 s 45800 548 45866 680 4 vdd
rlabel metal3 s 7940 32484 8072 32558 4 vdd
rlabel metal3 s 7940 103232 8072 103306 4 vdd
rlabel metal3 s 29462 548 29528 680 4 vdd
rlabel metal3 s 7940 44788 8072 44862 4 vdd
rlabel metal3 s 28684 548 28750 680 4 vdd
rlabel metal3 s 10556 5268 10622 5400 4 vdd
rlabel metal3 s 35452 5268 35518 5400 4 vdd
rlabel metal3 s 6400 97080 6532 97154 4 vdd
rlabel metal3 s 6400 100156 6532 100230 4 vdd
rlabel metal3 s 2084 26354 2216 26428 4 vdd
rlabel metal3 s 24560 5268 24626 5400 4 vdd
rlabel metal3 s 1044 17114 1176 17188 4 vdd
rlabel metal3 s 2264 10958 2396 11032 4 vdd
rlabel metal3 s 55162 3986 55294 4060 4 vdd
rlabel metal3 s 11594 3986 11726 4060 4 vdd
rlabel metal3 s 35686 548 35752 680 4 vdd
rlabel metal3 s 39576 548 39642 680 4 vdd
rlabel metal3 s 7940 60168 8072 60242 4 vdd
rlabel metal3 s 2084 23274 2216 23348 4 vdd
rlabel metal3 s 47900 5268 47966 5400 4 vdd
rlabel metal3 s 1044 26354 1176 26428 4 vdd
rlabel metal3 s 32340 5268 32406 5400 4 vdd
rlabel metal3 s 1044 41750 1176 41824 4 vdd
rlabel metal3 s 48134 548 48200 680 4 vdd
rlabel metal3 s 36490 3986 36622 4060 4 vdd
rlabel metal3 s 19348 548 19414 680 4 vdd
rlabel metal3 s 6400 17104 6532 17178 4 vdd
rlabel metal3 s 53606 3986 53738 4060 4 vdd
rlabel metal3 s 44244 548 44310 680 4 vdd
rlabel metal3 s 6400 29408 6532 29482 4 vdd
rlabel metal3 s 6400 60168 6532 60242 4 vdd
rlabel metal3 s 16236 548 16302 680 4 vdd
rlabel metal3 s 51246 548 51312 680 4 vdd
rlabel metal3 s 21682 548 21748 680 4 vdd
rlabel metal3 s 6400 78624 6532 78698 4 vdd
rlabel metal3 s 33352 548 33418 680 4 vdd
rlabel metal3 s 7940 38636 8072 38710 4 vdd
rlabel metal3 s 2084 17114 2216 17188 4 vdd
rlabel metal3 s 27426 3986 27558 4060 4 vdd
rlabel metal3 s 7940 81700 8072 81774 4 vdd
rlabel metal3 s 41158 3986 41290 4060 4 vdd
rlabel metal3 s 6400 14028 6532 14102 4 vdd
rlabel metal3 s 6400 103232 6532 103306 4 vdd
rlabel metal3 s 48938 3986 49070 4060 4 vdd
rlabel metal3 s 17792 548 17858 680 4 vdd
rlabel metal3 s 10790 548 10856 680 4 vdd
rlabel metal3 s 34908 548 34974 680 4 vdd
rlabel metal3 s 24314 3986 24446 4060 4 vdd
rlabel metal3 s 9234 548 9300 680 4 vdd
rlabel metal3 s 17818 3986 17950 4060 4 vdd
rlabel metal3 s 37242 548 37308 680 4 vdd
rlabel metal3 s 30266 3986 30398 4060 4 vdd
rlabel metal3 s 1392 7878 1524 7952 4 vdd
rlabel metal3 s 2084 35590 2216 35664 4 vdd
rlabel metal3 s 21448 5268 21514 5400 4 vdd
rlabel metal3 s 7940 57092 8072 57166 4 vdd
rlabel metal3 s 36464 548 36530 680 4 vdd
rlabel metal3 s 46098 3986 46230 4060 4 vdd
rlabel metal3 s 38318 3986 38450 4060 4 vdd
rlabel metal3 s 34130 548 34196 680 4 vdd
rlabel metal3 s 25598 3986 25730 4060 4 vdd
rlabel metal3 s 7940 50940 8072 51014 4 vdd
rlabel metal3 s 6400 38636 6532 38710 4 vdd
rlabel metal3 s 20126 548 20192 680 4 vdd
rlabel metal3 s 38564 5268 38630 5400 4 vdd
rlabel metal3 s 24016 548 24082 680 4 vdd
rlabel metal3 s 40120 5268 40186 5400 4 vdd
rlabel metal3 s 1044 20194 1176 20268 4 vdd
rlabel metal3 s 6400 57092 6532 57166 4 vdd
rlabel metal3 s 10038 3986 10170 4060 4 vdd
rlabel metal3 s 30240 548 30306 680 4 vdd
rlabel metal3 s 6400 7876 6532 7950 4 vdd
rlabel metal3 s 53878 3986 54010 4060 4 vdd
rlabel metal3 s 42688 548 42754 680 4 vdd
rlabel metal3 s 35206 3986 35338 4060 4 vdd
rlabel metal3 s 45826 3986 45958 4060 4 vdd
rlabel metal3 s 6400 35560 6532 35634 4 vdd
rlabel metal3 s 18570 548 18636 680 4 vdd
rlabel metal3 s 12346 548 12412 680 4 vdd
rlabel metal3 s 2264 7878 2396 7952 4 vdd
rlabel metal3 s 19892 5268 19958 5400 4 vdd
rlabel metal3 s 24794 548 24860 680 4 vdd
rlabel metal3 s 47382 3986 47514 4060 4 vdd
rlabel metal3 s 41676 5268 41742 5400 4 vdd
rlabel metal3 s 44270 3986 44402 4060 4 vdd
rlabel metal3 s 2084 20194 2216 20268 4 vdd
rlabel metal3 s 14706 3986 14838 4060 4 vdd
rlabel metal3 s 16780 5268 16846 5400 4 vdd
rlabel metal3 s 6400 63244 6532 63318 4 vdd
rlabel metal3 s 9000 5268 9066 5400 4 vdd
rlabel metal3 s 20904 548 20970 680 4 vdd
rlabel metal3 s 11568 548 11634 680 4 vdd
rlabel metal3 s 6400 32484 6532 32558 4 vdd
rlabel metal3 s 42986 3986 43118 4060 4 vdd
rlabel metal3 s 34934 3986 35066 4060 4 vdd
rlabel metal3 s 27128 548 27194 680 4 vdd
rlabel metal3 s 52568 5268 52634 5400 4 vdd
rlabel metal3 s 57470 548 57536 680 4 vdd
rlabel metal3 s 6400 47864 6532 47938 4 vdd
rlabel metal3 s 30538 3986 30670 4060 4 vdd
rlabel metal3 s 46578 548 46644 680 4 vdd
rlabel metal3 s 7940 87852 8072 87926 4 vdd
rlabel metal3 s 54124 5268 54190 5400 4 vdd
rlabel metal3 s 7940 35560 8072 35634 4 vdd
rlabel metal3 s 48912 548 48978 680 4 vdd
rlabel metal3 s 33378 3986 33510 4060 4 vdd
rlabel metal3 s 52802 548 52868 680 4 vdd
rlabel metal3 s 41132 548 41198 680 4 vdd
rlabel metal3 s 7940 29408 8072 29482 4 vdd
rlabel metal3 s 7940 84776 8072 84850 4 vdd
rlabel metal3 s 25870 3986 26002 4060 4 vdd
rlabel metal3 s 37008 5268 37074 5400 4 vdd
rlabel metal3 s 6400 20180 6532 20254 4 vdd
rlabel metal3 s 13422 3986 13554 4060 4 vdd
rlabel metal3 s 7940 75548 8072 75622 4 vdd
rlabel metal3 s 7940 97080 8072 97154 4 vdd
rlabel metal3 s 7940 47864 8072 47938 4 vdd
rlabel metal3 s 41430 3986 41562 4060 4 vdd
rlabel metal3 s 7940 72472 8072 72546 4 vdd
rlabel metal3 s 53580 548 53646 680 4 vdd
rlabel metal3 s 36762 3986 36894 4060 4 vdd
rlabel metal3 s 28982 3986 29114 4060 4 vdd
rlabel metal3 s 6400 75548 6532 75622 4 vdd
rlabel metal3 s 33896 5268 33962 5400 4 vdd
rlabel metal3 s 6400 41712 6532 41786 4 vdd
rlabel metal3 s 10310 3986 10442 4060 4 vdd
rlabel metal3 s 16262 3986 16394 4060 4 vdd
rlabel metal3 s 39602 3986 39734 4060 4 vdd
rlabel metal3 s 50766 3986 50898 4060 4 vdd
rlabel metal3 s 56718 3986 56850 4060 4 vdd
rlabel metal3 s 13150 3986 13282 4060 4 vdd
rlabel metal3 s 15458 548 15524 680 4 vdd
rlabel metal3 s 7940 41712 8072 41786 4 vdd
rlabel metal3 s 7940 94004 8072 94078 4 vdd
rlabel metal3 s 13668 5268 13734 5400 4 vdd
rlabel metal3 s 13124 548 13190 680 4 vdd
rlabel metal3 s 2084 41750 2216 41824 4 vdd
rlabel metal3 s 6400 90928 6532 91002 4 vdd
rlabel metal3 s 14680 548 14746 680 4 vdd
rlabel metal3 s 21202 3986 21334 4060 4 vdd
rlabel metal3 s 7940 66320 8072 66394 4 vdd
rlabel metal3 s 7940 63244 8072 63318 4 vdd
rlabel metal3 s 55914 548 55980 680 4 vdd
rlabel metal3 s 2084 32510 2216 32584 4 vdd
rlabel metal3 s 1044 38670 1176 38744 4 vdd
rlabel metal3 s 49210 3986 49342 4060 4 vdd
rlabel metal3 s 58248 548 58314 680 4 vdd
rlabel metal3 s 7940 14028 8072 14102 4 vdd
rlabel metal3 s 49690 548 49756 680 4 vdd
rlabel metal3 s 38046 3986 38178 4060 4 vdd
rlabel metal3 s 31822 3986 31954 4060 4 vdd
rlabel metal3 s 6400 54016 6532 54090 4 vdd
rlabel metal3 s 40354 548 40420 680 4 vdd
rlabel metal3 s 8754 3986 8886 4060 4 vdd
rlabel metal3 s 7940 69396 8072 69470 4 vdd
rlabel metal3 s 19374 3986 19506 4060 4 vdd
rlabel metal3 s 39874 3986 40006 4060 4 vdd
rlabel metal3 s 7940 78624 8072 78698 4 vdd
rlabel metal3 s 56990 3986 57122 4060 4 vdd
rlabel metal3 s 23238 548 23304 680 4 vdd
rlabel metal3 s 33650 3986 33782 4060 4 vdd
rlabel metal3 s 23004 5268 23070 5400 4 vdd
rlabel metal3 s 26116 5268 26182 5400 4 vdd
rlabel metal3 s 7940 23256 8072 23330 4 vdd
rlabel metal3 s 55680 5268 55746 5400 4 vdd
rlabel metal3 s 52050 3986 52182 4060 4 vdd
rlabel metal3 s 14978 3986 15110 4060 4 vdd
rlabel metal3 s 44542 3986 44674 4060 4 vdd
rlabel metal3 s 6400 10952 6532 11026 4 vdd
rlabel metal3 s 6400 66320 6532 66394 4 vdd
rlabel metal3 s 29228 5268 29294 5400 4 vdd
rlabel metal3 s 30784 5268 30850 5400 4 vdd
rlabel metal3 s 28710 3986 28842 4060 4 vdd
rlabel metal3 s 43232 5268 43298 5400 4 vdd
rlabel metal3 s 41910 548 41976 680 4 vdd
rlabel metal3 s 6400 81700 6532 81774 4 vdd
rlabel metal3 s 7940 10952 8072 11026 4 vdd
rlabel metal3 s 6400 94004 6532 94078 4 vdd
rlabel metal3 s 49456 5268 49522 5400 4 vdd
rlabel metal3 s 22486 3986 22618 4060 4 vdd
rlabel metal3 s 38020 548 38086 680 4 vdd
rlabel metal3 s 12112 5268 12178 5400 4 vdd
rlabel metal3 s 6400 26332 6532 26406 4 vdd
rlabel metal3 s 7940 90928 8072 91002 4 vdd
rlabel metal3 s 51012 5268 51078 5400 4 vdd
rlabel metal3 s 6400 72472 6532 72546 4 vdd
rlabel metal3 s 1044 23274 1176 23348 4 vdd
rlabel metal3 s 6400 87852 6532 87926 4 vdd
rlabel metal3 s 1044 35590 1176 35664 4 vdd
rlabel metal3 s 19646 3986 19778 4060 4 vdd
rlabel metal3 s 52024 548 52090 680 4 vdd
rlabel metal3 s 20930 3986 21062 4060 4 vdd
rlabel metal3 s 6400 23256 6532 23330 4 vdd
rlabel metal3 s 10012 548 10078 680 4 vdd
rlabel metal3 s 50468 548 50534 680 4 vdd
rlabel metal3 s 38798 548 38864 680 4 vdd
rlabel metal3 s 56692 548 56758 680 4 vdd
rlabel metal3 s 27906 548 27972 680 4 vdd
rlabel metal3 s 22460 548 22526 680 4 vdd
rlabel metal3 s 18090 3986 18222 4060 4 vdd
rlabel metal3 s 17014 548 17080 680 4 vdd
rlabel metal3 s 25572 548 25638 680 4 vdd
rlabel metal3 s 15224 5268 15290 5400 4 vdd
rlabel metal3 s 7940 26332 8072 26406 4 vdd
rlabel metal3 s 46344 5268 46410 5400 4 vdd
rlabel metal3 s 52322 3986 52454 4060 4 vdd
rlabel metal3 s 2084 38670 2216 38744 4 vdd
rlabel metal3 s 55136 548 55202 680 4 vdd
rlabel metal3 s 10564 2506 10696 2580 4 gnd
rlabel metal3 s 1044 27894 1176 27968 4 gnd
rlabel metal3 s 32348 2506 32480 2580 4 gnd
rlabel metal3 s 6400 58630 6532 58704 4 gnd
rlabel metal3 s 33904 2506 34036 2580 4 gnd
rlabel metal3 s 39350 2506 39482 2580 4 gnd
rlabel metal3 s 37008 6100 37074 6232 4 gnd
rlabel metal3 s 19646 4932 19778 5006 4 gnd
rlabel metal3 s 16780 6100 16846 6232 4 gnd
rlabel metal3 s 23004 6100 23070 6232 4 gnd
rlabel metal3 s 21448 6100 21514 6232 4 gnd
rlabel metal3 s 22486 4932 22618 5006 4 gnd
rlabel metal3 s 7940 12490 8072 12564 4 gnd
rlabel metal3 s 40906 2506 41038 2580 4 gnd
rlabel metal3 s 1044 34050 1176 34124 4 gnd
rlabel metal3 s 37794 2506 37926 2580 4 gnd
rlabel metal3 s 44542 4932 44674 5006 4 gnd
rlabel metal3 s 11594 4932 11726 5006 4 gnd
rlabel metal3 s 27426 4932 27558 5006 4 gnd
rlabel metal3 s 28982 4932 29114 5006 4 gnd
rlabel metal3 s 1044 15574 1176 15648 4 gnd
rlabel metal3 s 6400 12490 6532 12564 4 gnd
rlabel metal3 s 7940 64782 8072 64856 4 gnd
rlabel metal3 s 7940 86314 8072 86388 4 gnd
rlabel metal3 s 45826 4932 45958 5006 4 gnd
rlabel metal3 s 6400 6338 6532 6412 4 gnd
rlabel metal3 s 28458 2506 28590 2580 4 gnd
rlabel metal3 s 49464 2506 49596 2580 4 gnd
rlabel metal3 s 52568 6100 52634 6232 4 gnd
rlabel metal3 s 47900 6100 47966 6232 4 gnd
rlabel metal3 s 51798 2506 51930 2580 4 gnd
rlabel metal3 s 28710 4932 28842 5006 4 gnd
rlabel metal3 s 6400 95542 6532 95616 4 gnd
rlabel metal3 s 1392 9418 1524 9492 4 gnd
rlabel metal3 s 29228 6100 29294 6232 4 gnd
rlabel metal3 s 7940 104770 8072 104844 4 gnd
rlabel metal3 s 7940 80162 8072 80236 4 gnd
rlabel metal3 s 23790 2506 23922 2580 4 gnd
rlabel metal3 s 6400 40174 6532 40248 4 gnd
rlabel metal3 s 51020 2506 51152 2580 4 gnd
rlabel metal3 s 33126 2506 33258 2580 4 gnd
rlabel metal3 s 45574 2506 45706 2580 4 gnd
rlabel metal3 s 25346 2506 25478 2580 4 gnd
rlabel metal3 s 7940 18642 8072 18716 4 gnd
rlabel metal3 s 16010 2506 16142 2580 4 gnd
rlabel metal3 s 6400 77086 6532 77160 4 gnd
rlabel metal3 s 19892 6100 19958 6232 4 gnd
rlabel metal3 s 6400 80162 6532 80236 4 gnd
rlabel metal3 s 44270 4932 44402 5006 4 gnd
rlabel metal3 s 46344 6100 46410 6232 4 gnd
rlabel metal3 s 14706 4932 14838 5006 4 gnd
rlabel metal3 s 7940 92466 8072 92540 4 gnd
rlabel metal3 s 56466 2506 56598 2580 4 gnd
rlabel metal3 s 6400 98618 6532 98692 4 gnd
rlabel metal3 s 7940 46326 8072 46400 4 gnd
rlabel metal3 s 46098 4932 46230 5006 4 gnd
rlabel metal3 s 7940 98618 8072 98692 4 gnd
rlabel metal3 s 35206 4932 35338 5006 4 gnd
rlabel metal3 s 7940 43250 8072 43324 4 gnd
rlabel metal3 s 33378 4932 33510 5006 4 gnd
rlabel metal3 s 2084 27894 2216 27968 4 gnd
rlabel metal3 s 9786 2506 9918 2580 4 gnd
rlabel metal3 s 5816 3632 5948 3706 4 gnd
rlabel metal3 s 34934 4932 35066 5006 4 gnd
rlabel metal3 s 46352 2506 46484 2580 4 gnd
rlabel metal3 s 24314 4932 24446 5006 4 gnd
rlabel metal3 s 30014 2506 30146 2580 4 gnd
rlabel metal3 s 1044 18654 1176 18728 4 gnd
rlabel metal3 s 8482 4932 8614 5006 4 gnd
rlabel metal3 s 54132 2506 54264 2580 4 gnd
rlabel metal3 s 24560 6100 24626 6232 4 gnd
rlabel metal3 s 30784 6100 30850 6232 4 gnd
rlabel metal3 s 48938 4932 49070 5006 4 gnd
rlabel metal3 s 20678 2506 20810 2580 4 gnd
rlabel metal3 s 14454 2506 14586 2580 4 gnd
rlabel metal3 s 7940 61706 8072 61780 4 gnd
rlabel metal3 s 6400 21718 6532 21792 4 gnd
rlabel metal3 s 43240 2506 43372 2580 4 gnd
rlabel metal3 s 2084 34050 2216 34124 4 gnd
rlabel metal3 s 12120 2506 12252 2580 4 gnd
rlabel metal3 s 47908 2506 48040 2580 4 gnd
rlabel metal3 s 7940 89390 8072 89464 4 gnd
rlabel metal3 s 1044 30970 1176 31044 4 gnd
rlabel metal3 s 13676 2506 13808 2580 4 gnd
rlabel metal3 s 13422 4932 13554 5006 4 gnd
rlabel metal3 s 17818 4932 17950 5006 4 gnd
rlabel metal3 s 23012 2506 23144 2580 4 gnd
rlabel metal3 s 42986 4932 43118 5006 4 gnd
rlabel metal3 s 44788 6100 44854 6232 4 gnd
rlabel metal3 s 47382 4932 47514 5006 4 gnd
rlabel metal3 s 7940 49402 8072 49476 4 gnd
rlabel metal3 s 7940 27870 8072 27944 4 gnd
rlabel metal3 s 1044 43290 1176 43364 4 gnd
rlabel metal3 s 7940 52478 8072 52552 4 gnd
rlabel metal3 s 6400 104770 6532 104844 4 gnd
rlabel metal3 s 6400 46326 6532 46400 4 gnd
rlabel metal3 s 6400 74010 6532 74084 4 gnd
rlabel metal3 s 55162 4932 55294 5006 4 gnd
rlabel metal3 s 55688 2506 55820 2580 4 gnd
rlabel metal3 s 6400 70934 6532 71008 4 gnd
rlabel metal3 s 57244 2506 57376 2580 4 gnd
rlabel metal3 s 54910 2506 55042 2580 4 gnd
rlabel metal3 s 7940 34022 8072 34096 4 gnd
rlabel metal3 s 41158 4932 41290 5006 4 gnd
rlabel metal3 s 48686 2506 48818 2580 4 gnd
rlabel metal3 s 7940 9414 8072 9488 4 gnd
rlabel metal3 s 7940 74010 8072 74084 4 gnd
rlabel metal3 s 44018 2506 44150 2580 4 gnd
rlabel metal3 s 6400 43250 6532 43324 4 gnd
rlabel metal3 s 35452 6100 35518 6232 4 gnd
rlabel metal3 s 41684 2506 41816 2580 4 gnd
rlabel metal3 s 7940 37098 8072 37172 4 gnd
rlabel metal3 s 58022 2506 58154 2580 4 gnd
rlabel metal3 s 18344 2506 18476 2580 4 gnd
rlabel metal3 s 6400 49402 6532 49476 4 gnd
rlabel metal3 s 27154 4932 27286 5006 4 gnd
rlabel metal3 s 6400 83238 6532 83312 4 gnd
rlabel metal3 s 2084 15574 2216 15648 4 gnd
rlabel metal3 s 47654 4932 47786 5006 4 gnd
rlabel metal3 s 52576 2506 52708 2580 4 gnd
rlabel metal3 s 55680 6100 55746 6232 4 gnd
rlabel metal3 s 33896 6100 33962 6232 4 gnd
rlabel metal3 s 2264 12498 2396 12572 4 gnd
rlabel metal3 s 7940 83238 8072 83312 4 gnd
rlabel metal3 s 47130 2506 47262 2580 4 gnd
rlabel metal3 s 8754 4932 8886 5006 4 gnd
rlabel metal3 s 19122 2506 19254 2580 4 gnd
rlabel metal3 s 41676 6100 41742 6232 4 gnd
rlabel metal3 s 6400 89390 6532 89464 4 gnd
rlabel metal3 s 53878 4932 54010 5006 4 gnd
rlabel metal3 s 2084 18654 2216 18728 4 gnd
rlabel metal3 s 7940 67858 8072 67932 4 gnd
rlabel metal3 s 31822 4932 31954 5006 4 gnd
rlabel metal3 s 12898 2506 13030 2580 4 gnd
rlabel metal3 s 6400 64782 6532 64856 4 gnd
rlabel metal3 s 2084 30970 2216 31044 4 gnd
rlabel metal3 s 11342 2506 11474 2580 4 gnd
rlabel metal3 s 19374 4932 19506 5006 4 gnd
rlabel metal3 s 21202 4932 21334 5006 4 gnd
rlabel metal3 s 36490 4932 36622 5006 4 gnd
rlabel metal3 s 40120 6100 40186 6232 4 gnd
rlabel metal3 s 6400 37098 6532 37172 4 gnd
rlabel metal3 s 5816 5308 5948 5382 4 gnd
rlabel metal3 s 15224 6100 15290 6232 4 gnd
rlabel metal3 s 1392 6338 1524 6412 4 gnd
rlabel metal3 s 33650 4932 33782 5006 4 gnd
rlabel metal3 s 22758 4932 22890 5006 4 gnd
rlabel metal3 s 17566 2506 17698 2580 4 gnd
rlabel metal3 s 12112 6100 12178 6232 4 gnd
rlabel metal3 s 27672 6100 27738 6232 4 gnd
rlabel metal3 s 50242 2506 50374 2580 4 gnd
rlabel metal3 s 2084 21734 2216 21808 4 gnd
rlabel metal3 s 6400 24794 6532 24868 4 gnd
rlabel metal3 s 7940 6338 8072 6412 4 gnd
rlabel metal3 s 38046 4932 38178 5006 4 gnd
rlabel metal3 s 16788 2506 16920 2580 4 gnd
rlabel metal3 s 2084 43290 2216 43364 4 gnd
rlabel metal3 s 49210 4932 49342 5006 4 gnd
rlabel metal3 s 2084 40210 2216 40284 4 gnd
rlabel metal3 s 42714 4932 42846 5006 4 gnd
rlabel metal3 s 39874 4932 40006 5006 4 gnd
rlabel metal3 s 6400 61706 6532 61780 4 gnd
rlabel metal3 s 21456 2506 21588 2580 4 gnd
rlabel metal3 s 20930 4932 21062 5006 4 gnd
rlabel metal3 s 16534 4932 16666 5006 4 gnd
rlabel metal3 s 37016 2506 37148 2580 4 gnd
rlabel metal3 s 40128 2506 40260 2580 4 gnd
rlabel metal3 s 7940 95542 8072 95616 4 gnd
rlabel metal3 s 7940 24794 8072 24868 4 gnd
rlabel metal3 s 32340 6100 32406 6232 4 gnd
rlabel metal3 s 6400 55554 6532 55628 4 gnd
rlabel metal3 s 6400 27870 6532 27944 4 gnd
rlabel metal3 s 13150 4932 13282 5006 4 gnd
rlabel metal3 s 42462 2506 42594 2580 4 gnd
rlabel metal3 s 56990 4932 57122 5006 4 gnd
rlabel metal3 s 7940 70934 8072 71008 4 gnd
rlabel metal3 s 31570 2506 31702 2580 4 gnd
rlabel metal3 s 52050 4932 52182 5006 4 gnd
rlabel metal3 s 10556 6100 10622 6232 4 gnd
rlabel metal3 s 10038 4932 10170 5006 4 gnd
rlabel metal3 s 29236 2506 29368 2580 4 gnd
rlabel metal3 s 7940 77086 8072 77160 4 gnd
rlabel metal3 s 36238 2506 36370 2580 4 gnd
rlabel metal3 s 18336 6100 18402 6232 4 gnd
rlabel metal3 s 18090 4932 18222 5006 4 gnd
rlabel metal3 s 1044 40210 1176 40284 4 gnd
rlabel metal3 s 2084 37130 2216 37204 4 gnd
rlabel metal3 s 39602 4932 39734 5006 4 gnd
rlabel metal3 s 6400 52478 6532 52552 4 gnd
rlabel metal3 s 43232 6100 43298 6232 4 gnd
rlabel metal3 s 1044 21734 1176 21808 4 gnd
rlabel metal3 s 16262 4932 16394 5006 4 gnd
rlabel metal3 s 36762 4932 36894 5006 4 gnd
rlabel metal3 s 1044 24814 1176 24888 4 gnd
rlabel metal3 s 15232 2506 15364 2580 4 gnd
rlabel metal3 s 25598 4932 25730 5006 4 gnd
rlabel metal3 s 34682 2506 34814 2580 4 gnd
rlabel metal3 s 9000 6100 9066 6232 4 gnd
rlabel metal3 s 24042 4932 24174 5006 4 gnd
rlabel metal3 s 25870 4932 26002 5006 4 gnd
rlabel metal3 s 30266 4932 30398 5006 4 gnd
rlabel metal3 s 38564 6100 38630 6232 4 gnd
rlabel metal3 s 38318 4932 38450 5006 4 gnd
rlabel metal3 s 30538 4932 30670 5006 4 gnd
rlabel metal3 s 27680 2506 27812 2580 4 gnd
rlabel metal3 s 7940 40174 8072 40248 4 gnd
rlabel metal3 s 6400 30946 6532 31020 4 gnd
rlabel metal3 s 11866 4932 11998 5006 4 gnd
rlabel metal3 s 54124 6100 54190 6232 4 gnd
rlabel metal3 s 52322 4932 52454 5006 4 gnd
rlabel metal3 s 57236 6100 57302 6232 4 gnd
rlabel metal3 s 30792 2506 30924 2580 4 gnd
rlabel metal3 s 1044 37130 1176 37204 4 gnd
rlabel metal3 s 19900 2506 20032 2580 4 gnd
rlabel metal3 s 55434 4932 55566 5006 4 gnd
rlabel metal3 s 41430 4932 41562 5006 4 gnd
rlabel metal3 s 49456 6100 49522 6232 4 gnd
rlabel metal3 s 6400 34022 6532 34096 4 gnd
rlabel metal3 s 7940 21718 8072 21792 4 gnd
rlabel metal3 s 13668 6100 13734 6232 4 gnd
rlabel metal3 s 24568 2506 24700 2580 4 gnd
rlabel metal3 s 50494 4932 50626 5006 4 gnd
rlabel metal3 s 35460 2506 35592 2580 4 gnd
rlabel metal3 s 53606 4932 53738 5006 4 gnd
rlabel metal3 s 53354 2506 53486 2580 4 gnd
rlabel metal3 s 2084 24814 2216 24888 4 gnd
rlabel metal3 s 7940 30946 8072 31020 4 gnd
rlabel metal3 s 26902 2506 27034 2580 4 gnd
rlabel metal3 s 14978 4932 15110 5006 4 gnd
rlabel metal3 s 32094 4932 32226 5006 4 gnd
rlabel metal3 s 6400 18642 6532 18716 4 gnd
rlabel metal3 s 51012 6100 51078 6232 4 gnd
rlabel metal3 s 26116 6100 26182 6232 4 gnd
rlabel metal3 s 6400 9414 6532 9488 4 gnd
rlabel metal3 s 9008 2506 9140 2580 4 gnd
rlabel metal3 s 6400 101694 6532 101768 4 gnd
rlabel metal3 s 7940 58630 8072 58704 4 gnd
rlabel metal3 s 6400 15566 6532 15640 4 gnd
rlabel metal3 s 7940 101694 8072 101768 4 gnd
rlabel metal3 s 44796 2506 44928 2580 4 gnd
rlabel metal3 s 56718 4932 56850 5006 4 gnd
rlabel metal3 s 7940 55554 8072 55628 4 gnd
rlabel metal3 s 6400 92466 6532 92540 4 gnd
rlabel metal3 s 6400 86314 6532 86388 4 gnd
rlabel metal3 s 7940 15566 8072 15640 4 gnd
rlabel metal3 s 1392 12498 1524 12572 4 gnd
rlabel metal3 s 50766 4932 50898 5006 4 gnd
rlabel metal3 s 38572 2506 38704 2580 4 gnd
rlabel metal3 s 26124 2506 26256 2580 4 gnd
rlabel metal3 s 2264 9418 2396 9492 4 gnd
rlabel metal3 s 22234 2506 22366 2580 4 gnd
rlabel metal3 s 2264 6338 2396 6412 4 gnd
rlabel metal3 s 6400 67858 6532 67932 4 gnd
rlabel metal3 s 10310 4932 10442 5006 4 gnd
<< properties >>
string FIXED_BBOX 0 0 58950 105020
string GDS_FILE sram_0rw2r1w_32_128_sky130A.gds
string GDS_END 474952
string GDS_START 298668
<< end >>
