magic
tech sky130A
magscale 1 2
timestamp 1644951705
<< checkpaint >>
rect -1296 -1277 1764 2857
<< nwell >>
rect -36 739 504 1597
<< pwell >>
rect 358 51 408 133
<< psubdiff >>
rect 358 109 408 133
rect 358 75 366 109
rect 400 75 408 109
rect 358 51 408 75
<< nsubdiff >>
rect 358 1465 408 1489
rect 358 1431 366 1465
rect 400 1431 408 1465
rect 358 1407 408 1431
<< psubdiffcont >>
rect 366 75 400 109
<< nsubdiffcont >>
rect 366 1431 400 1465
<< poly >>
rect 114 323 144 1211
rect 214 447 244 1211
rect 196 431 262 447
rect 196 397 212 431
rect 246 397 262 431
rect 196 381 262 397
rect 96 307 162 323
rect 96 273 112 307
rect 146 273 162 307
rect 96 257 162 273
rect 114 245 144 257
rect 214 245 244 381
<< polycont >>
rect 212 397 246 431
rect 112 273 146 307
<< locali >>
rect 0 1523 468 1557
rect 62 1330 96 1523
rect 262 1330 296 1523
rect 366 1465 400 1523
rect 366 1415 400 1431
rect 162 1280 196 1330
rect 162 1246 364 1280
rect 196 431 262 447
rect 196 397 212 431
rect 246 397 262 431
rect 196 381 262 397
rect 96 307 162 323
rect 96 273 112 307
rect 146 273 162 307
rect 96 257 162 273
rect 330 253 364 1246
rect 262 219 364 253
rect 262 168 296 219
rect 366 109 400 125
rect 62 17 96 102
rect 366 17 400 75
rect 0 -17 468 17
use contact_12  contact_12_0
timestamp 1644951705
transform 1 0 196 0 1 381
box 0 0 1 1
use contact_12  contact_12_1
timestamp 1644951705
transform 1 0 96 0 1 257
box 0 0 1 1
use contact_11  contact_11_0
timestamp 1644951705
transform 1 0 358 0 1 51
box 0 0 1 1
use contact_10  contact_10_0
timestamp 1644951705
transform 1 0 358 0 1 1407
box 0 0 1 1
use nmos_m1_w0_840_sactive_dli  nmos_m1_w0_840_sactive_dli_0
timestamp 1644951705
transform 1 0 154 0 1 51
box 0 -26 150 194
use nmos_m1_w0_840_sli_dactive  nmos_m1_w0_840_sli_dactive_0
timestamp 1644951705
transform 1 0 54 0 1 51
box 0 -26 150 194
use pmos_m1_w1_260_sli_dli  pmos_m1_w1_260_sli_dli_0
timestamp 1644951705
transform 1 0 154 0 1 1237
box -59 -54 209 306
use pmos_m1_w1_260_sli_dli  pmos_m1_w1_260_sli_dli_1
timestamp 1644951705
transform 1 0 54 0 1 1237
box -59 -54 209 306
<< labels >>
rlabel locali s 347 1263 347 1263 4 Z
rlabel locali s 234 0 234 0 4 gnd
rlabel locali s 234 1540 234 1540 4 vdd
rlabel locali s 129 290 129 290 4 A
rlabel locali s 229 414 229 414 4 B
<< properties >>
string FIXED_BBOX 0 0 468 1540
string GDS_FILE sram_0rw2r1w_16_128_sky130A.gds
string GDS_END 1790262
string GDS_START 1787870
<< end >>
