magic
tech sky130A
magscale 1 2
timestamp 1643678851
<< checkpaint >>
rect -712 -1260 98552 2310
<< via1 >>
rect 658 954 710 1006
rect 3770 954 3822 1006
rect 6882 954 6934 1006
rect 9994 954 10046 1006
rect 13106 954 13158 1006
rect 16218 954 16270 1006
rect 19330 954 19382 1006
rect 22442 954 22494 1006
rect 25554 954 25606 1006
rect 28666 954 28718 1006
rect 31778 954 31830 1006
rect 34890 954 34942 1006
rect 38002 954 38054 1006
rect 41114 954 41166 1006
rect 44226 954 44278 1006
rect 47338 954 47390 1006
rect 50450 954 50502 1006
rect 53562 954 53614 1006
rect 56674 954 56726 1006
rect 59786 954 59838 1006
rect 62898 954 62950 1006
rect 66010 954 66062 1006
rect 69122 954 69174 1006
rect 72234 954 72286 1006
rect 75346 954 75398 1006
rect 78458 954 78510 1006
rect 81570 954 81622 1006
rect 84682 954 84734 1006
rect 87794 954 87846 1006
rect 90906 954 90958 1006
rect 94018 954 94070 1006
rect 97130 954 97182 1006
rect 658 8 710 60
rect 3770 8 3822 60
rect 6882 8 6934 60
rect 9994 8 10046 60
rect 13106 8 13158 60
rect 16218 8 16270 60
rect 19330 8 19382 60
rect 22442 8 22494 60
rect 25554 8 25606 60
rect 28666 8 28718 60
rect 31778 8 31830 60
rect 34890 8 34942 60
rect 38002 8 38054 60
rect 41114 8 41166 60
rect 44226 8 44278 60
rect 47338 8 47390 60
rect 50450 8 50502 60
rect 53562 8 53614 60
rect 56674 8 56726 60
rect 59786 8 59838 60
rect 62898 8 62950 60
rect 66010 8 66062 60
rect 69122 8 69174 60
rect 72234 8 72286 60
rect 75346 8 75398 60
rect 78458 8 78510 60
rect 81570 8 81622 60
rect 84682 8 84734 60
rect 87794 8 87846 60
rect 90906 8 90958 60
rect 94018 8 94070 60
rect 97130 8 97182 60
<< metal2 >>
rect 664 1008 704 1014
rect 3776 1008 3816 1014
rect 6888 1008 6928 1014
rect 10000 1008 10040 1014
rect 13112 1008 13152 1014
rect 16224 1008 16264 1014
rect 19336 1008 19376 1014
rect 22448 1008 22488 1014
rect 25560 1008 25600 1014
rect 28672 1008 28712 1014
rect 31784 1008 31824 1014
rect 34896 1008 34936 1014
rect 38008 1008 38048 1014
rect 41120 1008 41160 1014
rect 44232 1008 44272 1014
rect 47344 1008 47384 1014
rect 50456 1008 50496 1014
rect 53568 1008 53608 1014
rect 56680 1008 56720 1014
rect 59792 1008 59832 1014
rect 62904 1008 62944 1014
rect 66016 1008 66056 1014
rect 69128 1008 69168 1014
rect 72240 1008 72280 1014
rect 75352 1008 75392 1014
rect 78464 1008 78504 1014
rect 81576 1008 81616 1014
rect 84688 1008 84728 1014
rect 87800 1008 87840 1014
rect 90912 1008 90952 1014
rect 94024 1008 94064 1014
rect 97136 1008 97176 1014
rect 664 946 704 952
rect 3776 946 3816 952
rect 6888 946 6928 952
rect 10000 946 10040 952
rect 13112 946 13152 952
rect 16224 946 16264 952
rect 19336 946 19376 952
rect 22448 946 22488 952
rect 25560 946 25600 952
rect 28672 946 28712 952
rect 31784 946 31824 952
rect 34896 946 34936 952
rect 38008 946 38048 952
rect 41120 946 41160 952
rect 44232 946 44272 952
rect 47344 946 47384 952
rect 50456 946 50496 952
rect 53568 946 53608 952
rect 56680 946 56720 952
rect 59792 946 59832 952
rect 62904 946 62944 952
rect 66016 946 66056 952
rect 69128 946 69168 952
rect 72240 946 72280 952
rect 75352 946 75392 952
rect 78464 946 78504 952
rect 81576 946 81616 952
rect 84688 946 84728 952
rect 87800 946 87840 952
rect 90912 946 90952 952
rect 94024 946 94064 952
rect 97136 946 97176 952
rect 562 0 590 240
rect 664 62 704 68
rect 664 0 704 6
rect 750 0 778 240
rect 3674 0 3702 240
rect 3776 62 3816 68
rect 3776 0 3816 6
rect 3862 0 3890 240
rect 6786 0 6814 240
rect 6888 62 6928 68
rect 6888 0 6928 6
rect 6974 0 7002 240
rect 9898 0 9926 240
rect 10000 62 10040 68
rect 10000 0 10040 6
rect 10086 0 10114 240
rect 13010 0 13038 240
rect 13112 62 13152 68
rect 13112 0 13152 6
rect 13198 0 13226 240
rect 16122 0 16150 240
rect 16224 62 16264 68
rect 16224 0 16264 6
rect 16310 0 16338 240
rect 19234 0 19262 240
rect 19336 62 19376 68
rect 19336 0 19376 6
rect 19422 0 19450 240
rect 22346 0 22374 240
rect 22448 62 22488 68
rect 22448 0 22488 6
rect 22534 0 22562 240
rect 25458 0 25486 240
rect 25560 62 25600 68
rect 25560 0 25600 6
rect 25646 0 25674 240
rect 28570 0 28598 240
rect 28672 62 28712 68
rect 28672 0 28712 6
rect 28758 0 28786 240
rect 31682 0 31710 240
rect 31784 62 31824 68
rect 31784 0 31824 6
rect 31870 0 31898 240
rect 34794 0 34822 240
rect 34896 62 34936 68
rect 34896 0 34936 6
rect 34982 0 35010 240
rect 37906 0 37934 240
rect 38008 62 38048 68
rect 38008 0 38048 6
rect 38094 0 38122 240
rect 41018 0 41046 240
rect 41120 62 41160 68
rect 41120 0 41160 6
rect 41206 0 41234 240
rect 44130 0 44158 240
rect 44232 62 44272 68
rect 44232 0 44272 6
rect 44318 0 44346 240
rect 47242 0 47270 240
rect 47344 62 47384 68
rect 47344 0 47384 6
rect 47430 0 47458 240
rect 50354 0 50382 240
rect 50456 62 50496 68
rect 50456 0 50496 6
rect 50542 0 50570 240
rect 53466 0 53494 240
rect 53568 62 53608 68
rect 53568 0 53608 6
rect 53654 0 53682 240
rect 56578 0 56606 240
rect 56680 62 56720 68
rect 56680 0 56720 6
rect 56766 0 56794 240
rect 59690 0 59718 240
rect 59792 62 59832 68
rect 59792 0 59832 6
rect 59878 0 59906 240
rect 62802 0 62830 240
rect 62904 62 62944 68
rect 62904 0 62944 6
rect 62990 0 63018 240
rect 65914 0 65942 240
rect 66016 62 66056 68
rect 66016 0 66056 6
rect 66102 0 66130 240
rect 69026 0 69054 240
rect 69128 62 69168 68
rect 69128 0 69168 6
rect 69214 0 69242 240
rect 72138 0 72166 240
rect 72240 62 72280 68
rect 72240 0 72280 6
rect 72326 0 72354 240
rect 75250 0 75278 240
rect 75352 62 75392 68
rect 75352 0 75392 6
rect 75438 0 75466 240
rect 78362 0 78390 240
rect 78464 62 78504 68
rect 78464 0 78504 6
rect 78550 0 78578 240
rect 81474 0 81502 240
rect 81576 62 81616 68
rect 81576 0 81616 6
rect 81662 0 81690 240
rect 84586 0 84614 240
rect 84688 62 84728 68
rect 84688 0 84728 6
rect 84774 0 84802 240
rect 87698 0 87726 240
rect 87800 62 87840 68
rect 87800 0 87840 6
rect 87886 0 87914 240
rect 90810 0 90838 240
rect 90912 62 90952 68
rect 90912 0 90952 6
rect 90998 0 91026 240
rect 93922 0 93950 240
rect 94024 62 94064 68
rect 94024 0 94064 6
rect 94110 0 94138 240
rect 97034 0 97062 240
rect 97136 62 97176 68
rect 97136 0 97176 6
rect 97222 0 97250 240
<< via2 >>
rect 656 1006 712 1008
rect 656 954 658 1006
rect 658 954 710 1006
rect 710 954 712 1006
rect 656 952 712 954
rect 3768 1006 3824 1008
rect 3768 954 3770 1006
rect 3770 954 3822 1006
rect 3822 954 3824 1006
rect 3768 952 3824 954
rect 6880 1006 6936 1008
rect 6880 954 6882 1006
rect 6882 954 6934 1006
rect 6934 954 6936 1006
rect 6880 952 6936 954
rect 9992 1006 10048 1008
rect 9992 954 9994 1006
rect 9994 954 10046 1006
rect 10046 954 10048 1006
rect 9992 952 10048 954
rect 13104 1006 13160 1008
rect 13104 954 13106 1006
rect 13106 954 13158 1006
rect 13158 954 13160 1006
rect 13104 952 13160 954
rect 16216 1006 16272 1008
rect 16216 954 16218 1006
rect 16218 954 16270 1006
rect 16270 954 16272 1006
rect 16216 952 16272 954
rect 19328 1006 19384 1008
rect 19328 954 19330 1006
rect 19330 954 19382 1006
rect 19382 954 19384 1006
rect 19328 952 19384 954
rect 22440 1006 22496 1008
rect 22440 954 22442 1006
rect 22442 954 22494 1006
rect 22494 954 22496 1006
rect 22440 952 22496 954
rect 25552 1006 25608 1008
rect 25552 954 25554 1006
rect 25554 954 25606 1006
rect 25606 954 25608 1006
rect 25552 952 25608 954
rect 28664 1006 28720 1008
rect 28664 954 28666 1006
rect 28666 954 28718 1006
rect 28718 954 28720 1006
rect 28664 952 28720 954
rect 31776 1006 31832 1008
rect 31776 954 31778 1006
rect 31778 954 31830 1006
rect 31830 954 31832 1006
rect 31776 952 31832 954
rect 34888 1006 34944 1008
rect 34888 954 34890 1006
rect 34890 954 34942 1006
rect 34942 954 34944 1006
rect 34888 952 34944 954
rect 38000 1006 38056 1008
rect 38000 954 38002 1006
rect 38002 954 38054 1006
rect 38054 954 38056 1006
rect 38000 952 38056 954
rect 41112 1006 41168 1008
rect 41112 954 41114 1006
rect 41114 954 41166 1006
rect 41166 954 41168 1006
rect 41112 952 41168 954
rect 44224 1006 44280 1008
rect 44224 954 44226 1006
rect 44226 954 44278 1006
rect 44278 954 44280 1006
rect 44224 952 44280 954
rect 47336 1006 47392 1008
rect 47336 954 47338 1006
rect 47338 954 47390 1006
rect 47390 954 47392 1006
rect 47336 952 47392 954
rect 50448 1006 50504 1008
rect 50448 954 50450 1006
rect 50450 954 50502 1006
rect 50502 954 50504 1006
rect 50448 952 50504 954
rect 53560 1006 53616 1008
rect 53560 954 53562 1006
rect 53562 954 53614 1006
rect 53614 954 53616 1006
rect 53560 952 53616 954
rect 56672 1006 56728 1008
rect 56672 954 56674 1006
rect 56674 954 56726 1006
rect 56726 954 56728 1006
rect 56672 952 56728 954
rect 59784 1006 59840 1008
rect 59784 954 59786 1006
rect 59786 954 59838 1006
rect 59838 954 59840 1006
rect 59784 952 59840 954
rect 62896 1006 62952 1008
rect 62896 954 62898 1006
rect 62898 954 62950 1006
rect 62950 954 62952 1006
rect 62896 952 62952 954
rect 66008 1006 66064 1008
rect 66008 954 66010 1006
rect 66010 954 66062 1006
rect 66062 954 66064 1006
rect 66008 952 66064 954
rect 69120 1006 69176 1008
rect 69120 954 69122 1006
rect 69122 954 69174 1006
rect 69174 954 69176 1006
rect 69120 952 69176 954
rect 72232 1006 72288 1008
rect 72232 954 72234 1006
rect 72234 954 72286 1006
rect 72286 954 72288 1006
rect 72232 952 72288 954
rect 75344 1006 75400 1008
rect 75344 954 75346 1006
rect 75346 954 75398 1006
rect 75398 954 75400 1006
rect 75344 952 75400 954
rect 78456 1006 78512 1008
rect 78456 954 78458 1006
rect 78458 954 78510 1006
rect 78510 954 78512 1006
rect 78456 952 78512 954
rect 81568 1006 81624 1008
rect 81568 954 81570 1006
rect 81570 954 81622 1006
rect 81622 954 81624 1006
rect 81568 952 81624 954
rect 84680 1006 84736 1008
rect 84680 954 84682 1006
rect 84682 954 84734 1006
rect 84734 954 84736 1006
rect 84680 952 84736 954
rect 87792 1006 87848 1008
rect 87792 954 87794 1006
rect 87794 954 87846 1006
rect 87846 954 87848 1006
rect 87792 952 87848 954
rect 90904 1006 90960 1008
rect 90904 954 90906 1006
rect 90906 954 90958 1006
rect 90958 954 90960 1006
rect 90904 952 90960 954
rect 94016 1006 94072 1008
rect 94016 954 94018 1006
rect 94018 954 94070 1006
rect 94070 954 94072 1006
rect 94016 952 94072 954
rect 97128 1006 97184 1008
rect 97128 954 97130 1006
rect 97130 954 97182 1006
rect 97182 954 97184 1006
rect 97128 952 97184 954
rect 656 60 712 62
rect 656 8 658 60
rect 658 8 710 60
rect 710 8 712 60
rect 656 6 712 8
rect 3768 60 3824 62
rect 3768 8 3770 60
rect 3770 8 3822 60
rect 3822 8 3824 60
rect 3768 6 3824 8
rect 6880 60 6936 62
rect 6880 8 6882 60
rect 6882 8 6934 60
rect 6934 8 6936 60
rect 6880 6 6936 8
rect 9992 60 10048 62
rect 9992 8 9994 60
rect 9994 8 10046 60
rect 10046 8 10048 60
rect 9992 6 10048 8
rect 13104 60 13160 62
rect 13104 8 13106 60
rect 13106 8 13158 60
rect 13158 8 13160 60
rect 13104 6 13160 8
rect 16216 60 16272 62
rect 16216 8 16218 60
rect 16218 8 16270 60
rect 16270 8 16272 60
rect 16216 6 16272 8
rect 19328 60 19384 62
rect 19328 8 19330 60
rect 19330 8 19382 60
rect 19382 8 19384 60
rect 19328 6 19384 8
rect 22440 60 22496 62
rect 22440 8 22442 60
rect 22442 8 22494 60
rect 22494 8 22496 60
rect 22440 6 22496 8
rect 25552 60 25608 62
rect 25552 8 25554 60
rect 25554 8 25606 60
rect 25606 8 25608 60
rect 25552 6 25608 8
rect 28664 60 28720 62
rect 28664 8 28666 60
rect 28666 8 28718 60
rect 28718 8 28720 60
rect 28664 6 28720 8
rect 31776 60 31832 62
rect 31776 8 31778 60
rect 31778 8 31830 60
rect 31830 8 31832 60
rect 31776 6 31832 8
rect 34888 60 34944 62
rect 34888 8 34890 60
rect 34890 8 34942 60
rect 34942 8 34944 60
rect 34888 6 34944 8
rect 38000 60 38056 62
rect 38000 8 38002 60
rect 38002 8 38054 60
rect 38054 8 38056 60
rect 38000 6 38056 8
rect 41112 60 41168 62
rect 41112 8 41114 60
rect 41114 8 41166 60
rect 41166 8 41168 60
rect 41112 6 41168 8
rect 44224 60 44280 62
rect 44224 8 44226 60
rect 44226 8 44278 60
rect 44278 8 44280 60
rect 44224 6 44280 8
rect 47336 60 47392 62
rect 47336 8 47338 60
rect 47338 8 47390 60
rect 47390 8 47392 60
rect 47336 6 47392 8
rect 50448 60 50504 62
rect 50448 8 50450 60
rect 50450 8 50502 60
rect 50502 8 50504 60
rect 50448 6 50504 8
rect 53560 60 53616 62
rect 53560 8 53562 60
rect 53562 8 53614 60
rect 53614 8 53616 60
rect 53560 6 53616 8
rect 56672 60 56728 62
rect 56672 8 56674 60
rect 56674 8 56726 60
rect 56726 8 56728 60
rect 56672 6 56728 8
rect 59784 60 59840 62
rect 59784 8 59786 60
rect 59786 8 59838 60
rect 59838 8 59840 60
rect 59784 6 59840 8
rect 62896 60 62952 62
rect 62896 8 62898 60
rect 62898 8 62950 60
rect 62950 8 62952 60
rect 62896 6 62952 8
rect 66008 60 66064 62
rect 66008 8 66010 60
rect 66010 8 66062 60
rect 66062 8 66064 60
rect 66008 6 66064 8
rect 69120 60 69176 62
rect 69120 8 69122 60
rect 69122 8 69174 60
rect 69174 8 69176 60
rect 69120 6 69176 8
rect 72232 60 72288 62
rect 72232 8 72234 60
rect 72234 8 72286 60
rect 72286 8 72288 60
rect 72232 6 72288 8
rect 75344 60 75400 62
rect 75344 8 75346 60
rect 75346 8 75398 60
rect 75398 8 75400 60
rect 75344 6 75400 8
rect 78456 60 78512 62
rect 78456 8 78458 60
rect 78458 8 78510 60
rect 78510 8 78512 60
rect 78456 6 78512 8
rect 81568 60 81624 62
rect 81568 8 81570 60
rect 81570 8 81622 60
rect 81622 8 81624 60
rect 81568 6 81624 8
rect 84680 60 84736 62
rect 84680 8 84682 60
rect 84682 8 84734 60
rect 84734 8 84736 60
rect 84680 6 84736 8
rect 87792 60 87848 62
rect 87792 8 87794 60
rect 87794 8 87846 60
rect 87846 8 87848 60
rect 87792 6 87848 8
rect 90904 60 90960 62
rect 90904 8 90906 60
rect 90906 8 90958 60
rect 90958 8 90960 60
rect 90904 6 90960 8
rect 94016 60 94072 62
rect 94016 8 94018 60
rect 94018 8 94070 60
rect 94070 8 94072 60
rect 94016 6 94072 8
rect 97128 60 97184 62
rect 97128 8 97130 60
rect 97130 8 97182 60
rect 97182 8 97184 60
rect 97128 6 97184 8
<< metal3 >>
rect 618 1008 750 1013
rect 618 952 656 1008
rect 712 952 750 1008
rect 618 947 750 952
rect 3730 1008 3862 1013
rect 3730 952 3768 1008
rect 3824 952 3862 1008
rect 3730 947 3862 952
rect 6842 1008 6974 1013
rect 6842 952 6880 1008
rect 6936 952 6974 1008
rect 6842 947 6974 952
rect 9954 1008 10086 1013
rect 9954 952 9992 1008
rect 10048 952 10086 1008
rect 9954 947 10086 952
rect 13066 1008 13198 1013
rect 13066 952 13104 1008
rect 13160 952 13198 1008
rect 13066 947 13198 952
rect 16178 1008 16310 1013
rect 16178 952 16216 1008
rect 16272 952 16310 1008
rect 16178 947 16310 952
rect 19290 1008 19422 1013
rect 19290 952 19328 1008
rect 19384 952 19422 1008
rect 19290 947 19422 952
rect 22402 1008 22534 1013
rect 22402 952 22440 1008
rect 22496 952 22534 1008
rect 22402 947 22534 952
rect 25514 1008 25646 1013
rect 25514 952 25552 1008
rect 25608 952 25646 1008
rect 25514 947 25646 952
rect 28626 1008 28758 1013
rect 28626 952 28664 1008
rect 28720 952 28758 1008
rect 28626 947 28758 952
rect 31738 1008 31870 1013
rect 31738 952 31776 1008
rect 31832 952 31870 1008
rect 31738 947 31870 952
rect 34850 1008 34982 1013
rect 34850 952 34888 1008
rect 34944 952 34982 1008
rect 34850 947 34982 952
rect 37962 1008 38094 1013
rect 37962 952 38000 1008
rect 38056 952 38094 1008
rect 37962 947 38094 952
rect 41074 1008 41206 1013
rect 41074 952 41112 1008
rect 41168 952 41206 1008
rect 41074 947 41206 952
rect 44186 1008 44318 1013
rect 44186 952 44224 1008
rect 44280 952 44318 1008
rect 44186 947 44318 952
rect 47298 1008 47430 1013
rect 47298 952 47336 1008
rect 47392 952 47430 1008
rect 47298 947 47430 952
rect 50410 1008 50542 1013
rect 50410 952 50448 1008
rect 50504 952 50542 1008
rect 50410 947 50542 952
rect 53522 1008 53654 1013
rect 53522 952 53560 1008
rect 53616 952 53654 1008
rect 53522 947 53654 952
rect 56634 1008 56766 1013
rect 56634 952 56672 1008
rect 56728 952 56766 1008
rect 56634 947 56766 952
rect 59746 1008 59878 1013
rect 59746 952 59784 1008
rect 59840 952 59878 1008
rect 59746 947 59878 952
rect 62858 1008 62990 1013
rect 62858 952 62896 1008
rect 62952 952 62990 1008
rect 62858 947 62990 952
rect 65970 1008 66102 1013
rect 65970 952 66008 1008
rect 66064 952 66102 1008
rect 65970 947 66102 952
rect 69082 1008 69214 1013
rect 69082 952 69120 1008
rect 69176 952 69214 1008
rect 69082 947 69214 952
rect 72194 1008 72326 1013
rect 72194 952 72232 1008
rect 72288 952 72326 1008
rect 72194 947 72326 952
rect 75306 1008 75438 1013
rect 75306 952 75344 1008
rect 75400 952 75438 1008
rect 75306 947 75438 952
rect 78418 1008 78550 1013
rect 78418 952 78456 1008
rect 78512 952 78550 1008
rect 78418 947 78550 952
rect 81530 1008 81662 1013
rect 81530 952 81568 1008
rect 81624 952 81662 1008
rect 81530 947 81662 952
rect 84642 1008 84774 1013
rect 84642 952 84680 1008
rect 84736 952 84774 1008
rect 84642 947 84774 952
rect 87754 1008 87886 1013
rect 87754 952 87792 1008
rect 87848 952 87886 1008
rect 87754 947 87886 952
rect 90866 1008 90998 1013
rect 90866 952 90904 1008
rect 90960 952 90998 1008
rect 90866 947 90998 952
rect 93978 1008 94110 1013
rect 93978 952 94016 1008
rect 94072 952 94110 1008
rect 93978 947 94110 952
rect 97090 1008 97222 1013
rect 97090 952 97128 1008
rect 97184 952 97222 1008
rect 97090 947 97222 952
rect 618 62 750 67
rect 618 6 656 62
rect 712 6 750 62
rect 618 1 750 6
rect 3730 62 3862 67
rect 3730 6 3768 62
rect 3824 6 3862 62
rect 3730 1 3862 6
rect 6842 62 6974 67
rect 6842 6 6880 62
rect 6936 6 6974 62
rect 6842 1 6974 6
rect 9954 62 10086 67
rect 9954 6 9992 62
rect 10048 6 10086 62
rect 9954 1 10086 6
rect 13066 62 13198 67
rect 13066 6 13104 62
rect 13160 6 13198 62
rect 13066 1 13198 6
rect 16178 62 16310 67
rect 16178 6 16216 62
rect 16272 6 16310 62
rect 16178 1 16310 6
rect 19290 62 19422 67
rect 19290 6 19328 62
rect 19384 6 19422 62
rect 19290 1 19422 6
rect 22402 62 22534 67
rect 22402 6 22440 62
rect 22496 6 22534 62
rect 22402 1 22534 6
rect 25514 62 25646 67
rect 25514 6 25552 62
rect 25608 6 25646 62
rect 25514 1 25646 6
rect 28626 62 28758 67
rect 28626 6 28664 62
rect 28720 6 28758 62
rect 28626 1 28758 6
rect 31738 62 31870 67
rect 31738 6 31776 62
rect 31832 6 31870 62
rect 31738 1 31870 6
rect 34850 62 34982 67
rect 34850 6 34888 62
rect 34944 6 34982 62
rect 34850 1 34982 6
rect 37962 62 38094 67
rect 37962 6 38000 62
rect 38056 6 38094 62
rect 37962 1 38094 6
rect 41074 62 41206 67
rect 41074 6 41112 62
rect 41168 6 41206 62
rect 41074 1 41206 6
rect 44186 62 44318 67
rect 44186 6 44224 62
rect 44280 6 44318 62
rect 44186 1 44318 6
rect 47298 62 47430 67
rect 47298 6 47336 62
rect 47392 6 47430 62
rect 47298 1 47430 6
rect 50410 62 50542 67
rect 50410 6 50448 62
rect 50504 6 50542 62
rect 50410 1 50542 6
rect 53522 62 53654 67
rect 53522 6 53560 62
rect 53616 6 53654 62
rect 53522 1 53654 6
rect 56634 62 56766 67
rect 56634 6 56672 62
rect 56728 6 56766 62
rect 56634 1 56766 6
rect 59746 62 59878 67
rect 59746 6 59784 62
rect 59840 6 59878 62
rect 59746 1 59878 6
rect 62858 62 62990 67
rect 62858 6 62896 62
rect 62952 6 62990 62
rect 62858 1 62990 6
rect 65970 62 66102 67
rect 65970 6 66008 62
rect 66064 6 66102 62
rect 65970 1 66102 6
rect 69082 62 69214 67
rect 69082 6 69120 62
rect 69176 6 69214 62
rect 69082 1 69214 6
rect 72194 62 72326 67
rect 72194 6 72232 62
rect 72288 6 72326 62
rect 72194 1 72326 6
rect 75306 62 75438 67
rect 75306 6 75344 62
rect 75400 6 75438 62
rect 75306 1 75438 6
rect 78418 62 78550 67
rect 78418 6 78456 62
rect 78512 6 78550 62
rect 78418 1 78550 6
rect 81530 62 81662 67
rect 81530 6 81568 62
rect 81624 6 81662 62
rect 81530 1 81662 6
rect 84642 62 84774 67
rect 84642 6 84680 62
rect 84736 6 84774 62
rect 84642 1 84774 6
rect 87754 62 87886 67
rect 87754 6 87792 62
rect 87848 6 87886 62
rect 87754 1 87886 6
rect 90866 62 90998 67
rect 90866 6 90904 62
rect 90960 6 90998 62
rect 90866 1 90998 6
rect 93978 62 94110 67
rect 93978 6 94016 62
rect 94072 6 94110 62
rect 93978 1 94110 6
rect 97090 62 97222 67
rect 97090 6 97128 62
rect 97184 6 97222 62
rect 97090 1 97222 6
use contact_18  contact_18_0
timestamp 1643678851
transform 1 0 97090 0 1 947
box 0 0 1 1
use contact_17  contact_17_0
timestamp 1643678851
transform 1 0 97141 0 1 965
box 0 0 1 1
use contact_18  contact_18_1
timestamp 1643678851
transform 1 0 97090 0 1 1
box 0 0 1 1
use contact_17  contact_17_1
timestamp 1643678851
transform 1 0 97141 0 1 19
box 0 0 1 1
use contact_18  contact_18_2
timestamp 1643678851
transform 1 0 93978 0 1 947
box 0 0 1 1
use contact_17  contact_17_2
timestamp 1643678851
transform 1 0 94029 0 1 965
box 0 0 1 1
use contact_18  contact_18_3
timestamp 1643678851
transform 1 0 93978 0 1 1
box 0 0 1 1
use contact_17  contact_17_3
timestamp 1643678851
transform 1 0 94029 0 1 19
box 0 0 1 1
use contact_18  contact_18_4
timestamp 1643678851
transform 1 0 90866 0 1 947
box 0 0 1 1
use contact_17  contact_17_4
timestamp 1643678851
transform 1 0 90917 0 1 965
box 0 0 1 1
use contact_18  contact_18_5
timestamp 1643678851
transform 1 0 90866 0 1 1
box 0 0 1 1
use contact_17  contact_17_5
timestamp 1643678851
transform 1 0 90917 0 1 19
box 0 0 1 1
use contact_18  contact_18_6
timestamp 1643678851
transform 1 0 87754 0 1 947
box 0 0 1 1
use contact_17  contact_17_6
timestamp 1643678851
transform 1 0 87805 0 1 965
box 0 0 1 1
use contact_18  contact_18_7
timestamp 1643678851
transform 1 0 87754 0 1 1
box 0 0 1 1
use contact_17  contact_17_7
timestamp 1643678851
transform 1 0 87805 0 1 19
box 0 0 1 1
use contact_18  contact_18_8
timestamp 1643678851
transform 1 0 84642 0 1 947
box 0 0 1 1
use contact_17  contact_17_8
timestamp 1643678851
transform 1 0 84693 0 1 965
box 0 0 1 1
use contact_18  contact_18_9
timestamp 1643678851
transform 1 0 84642 0 1 1
box 0 0 1 1
use contact_17  contact_17_9
timestamp 1643678851
transform 1 0 84693 0 1 19
box 0 0 1 1
use contact_18  contact_18_10
timestamp 1643678851
transform 1 0 81530 0 1 947
box 0 0 1 1
use contact_17  contact_17_10
timestamp 1643678851
transform 1 0 81581 0 1 965
box 0 0 1 1
use contact_18  contact_18_11
timestamp 1643678851
transform 1 0 81530 0 1 1
box 0 0 1 1
use contact_17  contact_17_11
timestamp 1643678851
transform 1 0 81581 0 1 19
box 0 0 1 1
use contact_18  contact_18_12
timestamp 1643678851
transform 1 0 78418 0 1 947
box 0 0 1 1
use contact_17  contact_17_12
timestamp 1643678851
transform 1 0 78469 0 1 965
box 0 0 1 1
use contact_18  contact_18_13
timestamp 1643678851
transform 1 0 78418 0 1 1
box 0 0 1 1
use contact_17  contact_17_13
timestamp 1643678851
transform 1 0 78469 0 1 19
box 0 0 1 1
use contact_18  contact_18_14
timestamp 1643678851
transform 1 0 75306 0 1 947
box 0 0 1 1
use contact_17  contact_17_14
timestamp 1643678851
transform 1 0 75357 0 1 965
box 0 0 1 1
use contact_18  contact_18_15
timestamp 1643678851
transform 1 0 75306 0 1 1
box 0 0 1 1
use contact_17  contact_17_15
timestamp 1643678851
transform 1 0 75357 0 1 19
box 0 0 1 1
use contact_18  contact_18_16
timestamp 1643678851
transform 1 0 72194 0 1 947
box 0 0 1 1
use contact_17  contact_17_16
timestamp 1643678851
transform 1 0 72245 0 1 965
box 0 0 1 1
use contact_18  contact_18_17
timestamp 1643678851
transform 1 0 72194 0 1 1
box 0 0 1 1
use contact_17  contact_17_17
timestamp 1643678851
transform 1 0 72245 0 1 19
box 0 0 1 1
use contact_18  contact_18_18
timestamp 1643678851
transform 1 0 69082 0 1 947
box 0 0 1 1
use contact_17  contact_17_18
timestamp 1643678851
transform 1 0 69133 0 1 965
box 0 0 1 1
use contact_18  contact_18_19
timestamp 1643678851
transform 1 0 69082 0 1 1
box 0 0 1 1
use contact_17  contact_17_19
timestamp 1643678851
transform 1 0 69133 0 1 19
box 0 0 1 1
use contact_18  contact_18_20
timestamp 1643678851
transform 1 0 65970 0 1 947
box 0 0 1 1
use contact_17  contact_17_20
timestamp 1643678851
transform 1 0 66021 0 1 965
box 0 0 1 1
use contact_18  contact_18_21
timestamp 1643678851
transform 1 0 65970 0 1 1
box 0 0 1 1
use contact_17  contact_17_21
timestamp 1643678851
transform 1 0 66021 0 1 19
box 0 0 1 1
use contact_18  contact_18_22
timestamp 1643678851
transform 1 0 62858 0 1 947
box 0 0 1 1
use contact_17  contact_17_22
timestamp 1643678851
transform 1 0 62909 0 1 965
box 0 0 1 1
use contact_18  contact_18_23
timestamp 1643678851
transform 1 0 62858 0 1 1
box 0 0 1 1
use contact_17  contact_17_23
timestamp 1643678851
transform 1 0 62909 0 1 19
box 0 0 1 1
use contact_18  contact_18_24
timestamp 1643678851
transform 1 0 59746 0 1 947
box 0 0 1 1
use contact_17  contact_17_24
timestamp 1643678851
transform 1 0 59797 0 1 965
box 0 0 1 1
use contact_18  contact_18_25
timestamp 1643678851
transform 1 0 59746 0 1 1
box 0 0 1 1
use contact_17  contact_17_25
timestamp 1643678851
transform 1 0 59797 0 1 19
box 0 0 1 1
use contact_18  contact_18_26
timestamp 1643678851
transform 1 0 56634 0 1 947
box 0 0 1 1
use contact_17  contact_17_26
timestamp 1643678851
transform 1 0 56685 0 1 965
box 0 0 1 1
use contact_18  contact_18_27
timestamp 1643678851
transform 1 0 56634 0 1 1
box 0 0 1 1
use contact_17  contact_17_27
timestamp 1643678851
transform 1 0 56685 0 1 19
box 0 0 1 1
use contact_18  contact_18_28
timestamp 1643678851
transform 1 0 53522 0 1 947
box 0 0 1 1
use contact_17  contact_17_28
timestamp 1643678851
transform 1 0 53573 0 1 965
box 0 0 1 1
use contact_18  contact_18_29
timestamp 1643678851
transform 1 0 53522 0 1 1
box 0 0 1 1
use contact_17  contact_17_29
timestamp 1643678851
transform 1 0 53573 0 1 19
box 0 0 1 1
use contact_18  contact_18_30
timestamp 1643678851
transform 1 0 50410 0 1 947
box 0 0 1 1
use contact_17  contact_17_30
timestamp 1643678851
transform 1 0 50461 0 1 965
box 0 0 1 1
use contact_18  contact_18_31
timestamp 1643678851
transform 1 0 50410 0 1 1
box 0 0 1 1
use contact_17  contact_17_31
timestamp 1643678851
transform 1 0 50461 0 1 19
box 0 0 1 1
use contact_18  contact_18_32
timestamp 1643678851
transform 1 0 47298 0 1 947
box 0 0 1 1
use contact_17  contact_17_32
timestamp 1643678851
transform 1 0 47349 0 1 965
box 0 0 1 1
use contact_18  contact_18_33
timestamp 1643678851
transform 1 0 47298 0 1 1
box 0 0 1 1
use contact_17  contact_17_33
timestamp 1643678851
transform 1 0 47349 0 1 19
box 0 0 1 1
use contact_18  contact_18_34
timestamp 1643678851
transform 1 0 44186 0 1 947
box 0 0 1 1
use contact_17  contact_17_34
timestamp 1643678851
transform 1 0 44237 0 1 965
box 0 0 1 1
use contact_18  contact_18_35
timestamp 1643678851
transform 1 0 44186 0 1 1
box 0 0 1 1
use contact_17  contact_17_35
timestamp 1643678851
transform 1 0 44237 0 1 19
box 0 0 1 1
use contact_18  contact_18_36
timestamp 1643678851
transform 1 0 41074 0 1 947
box 0 0 1 1
use contact_17  contact_17_36
timestamp 1643678851
transform 1 0 41125 0 1 965
box 0 0 1 1
use contact_18  contact_18_37
timestamp 1643678851
transform 1 0 41074 0 1 1
box 0 0 1 1
use contact_17  contact_17_37
timestamp 1643678851
transform 1 0 41125 0 1 19
box 0 0 1 1
use contact_18  contact_18_38
timestamp 1643678851
transform 1 0 37962 0 1 947
box 0 0 1 1
use contact_17  contact_17_38
timestamp 1643678851
transform 1 0 38013 0 1 965
box 0 0 1 1
use contact_18  contact_18_39
timestamp 1643678851
transform 1 0 37962 0 1 1
box 0 0 1 1
use contact_17  contact_17_39
timestamp 1643678851
transform 1 0 38013 0 1 19
box 0 0 1 1
use contact_18  contact_18_40
timestamp 1643678851
transform 1 0 34850 0 1 947
box 0 0 1 1
use contact_17  contact_17_40
timestamp 1643678851
transform 1 0 34901 0 1 965
box 0 0 1 1
use contact_18  contact_18_41
timestamp 1643678851
transform 1 0 34850 0 1 1
box 0 0 1 1
use contact_17  contact_17_41
timestamp 1643678851
transform 1 0 34901 0 1 19
box 0 0 1 1
use contact_18  contact_18_42
timestamp 1643678851
transform 1 0 31738 0 1 947
box 0 0 1 1
use contact_17  contact_17_42
timestamp 1643678851
transform 1 0 31789 0 1 965
box 0 0 1 1
use contact_18  contact_18_43
timestamp 1643678851
transform 1 0 31738 0 1 1
box 0 0 1 1
use contact_17  contact_17_43
timestamp 1643678851
transform 1 0 31789 0 1 19
box 0 0 1 1
use contact_18  contact_18_44
timestamp 1643678851
transform 1 0 28626 0 1 947
box 0 0 1 1
use contact_17  contact_17_44
timestamp 1643678851
transform 1 0 28677 0 1 965
box 0 0 1 1
use contact_18  contact_18_45
timestamp 1643678851
transform 1 0 28626 0 1 1
box 0 0 1 1
use contact_17  contact_17_45
timestamp 1643678851
transform 1 0 28677 0 1 19
box 0 0 1 1
use contact_18  contact_18_46
timestamp 1643678851
transform 1 0 25514 0 1 947
box 0 0 1 1
use contact_17  contact_17_46
timestamp 1643678851
transform 1 0 25565 0 1 965
box 0 0 1 1
use contact_18  contact_18_47
timestamp 1643678851
transform 1 0 25514 0 1 1
box 0 0 1 1
use contact_17  contact_17_47
timestamp 1643678851
transform 1 0 25565 0 1 19
box 0 0 1 1
use contact_18  contact_18_48
timestamp 1643678851
transform 1 0 22402 0 1 947
box 0 0 1 1
use contact_17  contact_17_48
timestamp 1643678851
transform 1 0 22453 0 1 965
box 0 0 1 1
use contact_18  contact_18_49
timestamp 1643678851
transform 1 0 22402 0 1 1
box 0 0 1 1
use contact_17  contact_17_49
timestamp 1643678851
transform 1 0 22453 0 1 19
box 0 0 1 1
use contact_18  contact_18_50
timestamp 1643678851
transform 1 0 19290 0 1 947
box 0 0 1 1
use contact_17  contact_17_50
timestamp 1643678851
transform 1 0 19341 0 1 965
box 0 0 1 1
use contact_18  contact_18_51
timestamp 1643678851
transform 1 0 19290 0 1 1
box 0 0 1 1
use contact_17  contact_17_51
timestamp 1643678851
transform 1 0 19341 0 1 19
box 0 0 1 1
use contact_18  contact_18_52
timestamp 1643678851
transform 1 0 16178 0 1 947
box 0 0 1 1
use contact_17  contact_17_52
timestamp 1643678851
transform 1 0 16229 0 1 965
box 0 0 1 1
use contact_18  contact_18_53
timestamp 1643678851
transform 1 0 16178 0 1 1
box 0 0 1 1
use contact_17  contact_17_53
timestamp 1643678851
transform 1 0 16229 0 1 19
box 0 0 1 1
use contact_18  contact_18_54
timestamp 1643678851
transform 1 0 13066 0 1 947
box 0 0 1 1
use contact_17  contact_17_54
timestamp 1643678851
transform 1 0 13117 0 1 965
box 0 0 1 1
use contact_18  contact_18_55
timestamp 1643678851
transform 1 0 13066 0 1 1
box 0 0 1 1
use contact_17  contact_17_55
timestamp 1643678851
transform 1 0 13117 0 1 19
box 0 0 1 1
use contact_18  contact_18_56
timestamp 1643678851
transform 1 0 9954 0 1 947
box 0 0 1 1
use contact_17  contact_17_56
timestamp 1643678851
transform 1 0 10005 0 1 965
box 0 0 1 1
use contact_18  contact_18_57
timestamp 1643678851
transform 1 0 9954 0 1 1
box 0 0 1 1
use contact_17  contact_17_57
timestamp 1643678851
transform 1 0 10005 0 1 19
box 0 0 1 1
use contact_18  contact_18_58
timestamp 1643678851
transform 1 0 6842 0 1 947
box 0 0 1 1
use contact_17  contact_17_58
timestamp 1643678851
transform 1 0 6893 0 1 965
box 0 0 1 1
use contact_18  contact_18_59
timestamp 1643678851
transform 1 0 6842 0 1 1
box 0 0 1 1
use contact_17  contact_17_59
timestamp 1643678851
transform 1 0 6893 0 1 19
box 0 0 1 1
use contact_18  contact_18_60
timestamp 1643678851
transform 1 0 3730 0 1 947
box 0 0 1 1
use contact_17  contact_17_60
timestamp 1643678851
transform 1 0 3781 0 1 965
box 0 0 1 1
use contact_18  contact_18_61
timestamp 1643678851
transform 1 0 3730 0 1 1
box 0 0 1 1
use contact_17  contact_17_61
timestamp 1643678851
transform 1 0 3781 0 1 19
box 0 0 1 1
use contact_18  contact_18_62
timestamp 1643678851
transform 1 0 618 0 1 947
box 0 0 1 1
use contact_17  contact_17_62
timestamp 1643678851
transform 1 0 669 0 1 965
box 0 0 1 1
use contact_18  contact_18_63
timestamp 1643678851
transform 1 0 618 0 1 1
box 0 0 1 1
use contact_17  contact_17_63
timestamp 1643678851
transform 1 0 669 0 1 19
box 0 0 1 1
use sense_amp_multiport  sense_amp_multiport_0
timestamp 1643678851
transform 1 0 97020 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_1
timestamp 1643678851
transform 1 0 93908 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_2
timestamp 1643678851
transform 1 0 90796 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_3
timestamp 1643678851
transform 1 0 87684 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_4
timestamp 1643678851
transform 1 0 84572 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_5
timestamp 1643678851
transform 1 0 81460 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_6
timestamp 1643678851
transform 1 0 78348 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_7
timestamp 1643678851
transform 1 0 75236 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_8
timestamp 1643678851
transform 1 0 72124 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_9
timestamp 1643678851
transform 1 0 69012 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_10
timestamp 1643678851
transform 1 0 65900 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_11
timestamp 1643678851
transform 1 0 62788 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_12
timestamp 1643678851
transform 1 0 59676 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_13
timestamp 1643678851
transform 1 0 56564 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_14
timestamp 1643678851
transform 1 0 53452 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_15
timestamp 1643678851
transform 1 0 50340 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_16
timestamp 1643678851
transform 1 0 47228 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_17
timestamp 1643678851
transform 1 0 44116 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_18
timestamp 1643678851
transform 1 0 41004 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_19
timestamp 1643678851
transform 1 0 37892 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_20
timestamp 1643678851
transform 1 0 34780 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_21
timestamp 1643678851
transform 1 0 31668 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_22
timestamp 1643678851
transform 1 0 28556 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_23
timestamp 1643678851
transform 1 0 25444 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_24
timestamp 1643678851
transform 1 0 22332 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_25
timestamp 1643678851
transform 1 0 19220 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_26
timestamp 1643678851
transform 1 0 16108 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_27
timestamp 1643678851
transform 1 0 12996 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_28
timestamp 1643678851
transform 1 0 9884 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_29
timestamp 1643678851
transform 1 0 6772 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_30
timestamp 1643678851
transform 1 0 3660 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_31
timestamp 1643678851
transform 1 0 548 0 1 0
box 0 0 272 1050
<< labels >>
rlabel metal3 s 34850 1 34982 67 4 gnd
rlabel metal3 s 13066 1 13198 67 4 gnd
rlabel metal3 s 28626 1 28758 67 4 gnd
rlabel metal3 s 37962 1 38094 67 4 gnd
rlabel metal3 s 97090 1 97222 67 4 gnd
rlabel metal3 s 25514 1 25646 67 4 gnd
rlabel metal3 s 62858 1 62990 67 4 gnd
rlabel metal3 s 75306 1 75438 67 4 gnd
rlabel metal3 s 84642 1 84774 67 4 gnd
rlabel metal3 s 90866 1 90998 67 4 gnd
rlabel metal3 s 78418 1 78550 67 4 gnd
rlabel metal3 s 9954 1 10086 67 4 gnd
rlabel metal3 s 81530 1 81662 67 4 gnd
rlabel metal3 s 41074 1 41206 67 4 gnd
rlabel metal3 s 72194 1 72326 67 4 gnd
rlabel metal3 s 93978 1 94110 67 4 gnd
rlabel metal3 s 618 1 750 67 4 gnd
rlabel metal3 s 69082 1 69214 67 4 gnd
rlabel metal3 s 22402 1 22534 67 4 gnd
rlabel metal3 s 31738 1 31870 67 4 gnd
rlabel metal3 s 19290 1 19422 67 4 gnd
rlabel metal3 s 53522 1 53654 67 4 gnd
rlabel metal3 s 59746 1 59878 67 4 gnd
rlabel metal3 s 50410 1 50542 67 4 gnd
rlabel metal3 s 47298 1 47430 67 4 gnd
rlabel metal3 s 16178 1 16310 67 4 gnd
rlabel metal3 s 65970 1 66102 67 4 gnd
rlabel metal3 s 3730 1 3862 67 4 gnd
rlabel metal3 s 6842 1 6974 67 4 gnd
rlabel metal3 s 44186 1 44318 67 4 gnd
rlabel metal3 s 87754 1 87886 67 4 gnd
rlabel metal3 s 56634 1 56766 67 4 gnd
rlabel metal3 s 3730 947 3862 1013 4 vdd
rlabel metal3 s 69082 947 69214 1013 4 vdd
rlabel metal3 s 47298 947 47430 1013 4 vdd
rlabel metal3 s 65970 947 66102 1013 4 vdd
rlabel metal3 s 81530 947 81662 1013 4 vdd
rlabel metal3 s 59746 947 59878 1013 4 vdd
rlabel metal3 s 44186 947 44318 1013 4 vdd
rlabel metal3 s 56634 947 56766 1013 4 vdd
rlabel metal3 s 53522 947 53654 1013 4 vdd
rlabel metal3 s 41074 947 41206 1013 4 vdd
rlabel metal3 s 31738 947 31870 1013 4 vdd
rlabel metal3 s 9954 947 10086 1013 4 vdd
rlabel metal3 s 90866 947 90998 1013 4 vdd
rlabel metal3 s 84642 947 84774 1013 4 vdd
rlabel metal3 s 25514 947 25646 1013 4 vdd
rlabel metal3 s 50410 947 50542 1013 4 vdd
rlabel metal3 s 34850 947 34982 1013 4 vdd
rlabel metal3 s 19290 947 19422 1013 4 vdd
rlabel metal3 s 78418 947 78550 1013 4 vdd
rlabel metal3 s 75306 947 75438 1013 4 vdd
rlabel metal3 s 72194 947 72326 1013 4 vdd
rlabel metal3 s 62858 947 62990 1013 4 vdd
rlabel metal3 s 87754 947 87886 1013 4 vdd
rlabel metal3 s 618 947 750 1013 4 vdd
rlabel metal3 s 28626 947 28758 1013 4 vdd
rlabel metal3 s 6842 947 6974 1013 4 vdd
rlabel metal3 s 97090 947 97222 1013 4 vdd
rlabel metal3 s 93978 947 94110 1013 4 vdd
rlabel metal3 s 22402 947 22534 1013 4 vdd
rlabel metal3 s 13066 947 13198 1013 4 vdd
rlabel metal3 s 16178 947 16310 1013 4 vdd
rlabel metal3 s 37962 947 38094 1013 4 vdd
rlabel metal2 s 562 0 590 240 4 rbl_0
rlabel metal2 s 750 0 778 240 4 data_0
rlabel metal2 s 3674 0 3702 240 4 rbl_1
rlabel metal2 s 3862 0 3890 240 4 data_1
rlabel metal2 s 6786 0 6814 240 4 rbl_2
rlabel metal2 s 6974 0 7002 240 4 data_2
rlabel metal2 s 9898 0 9926 240 4 rbl_3
rlabel metal2 s 10086 0 10114 240 4 data_3
rlabel metal2 s 13010 0 13038 240 4 rbl_4
rlabel metal2 s 13198 0 13226 240 4 data_4
rlabel metal2 s 16122 0 16150 240 4 rbl_5
rlabel metal2 s 16310 0 16338 240 4 data_5
rlabel metal2 s 19234 0 19262 240 4 rbl_6
rlabel metal2 s 19422 0 19450 240 4 data_6
rlabel metal2 s 22346 0 22374 240 4 rbl_7
rlabel metal2 s 22534 0 22562 240 4 data_7
rlabel metal2 s 25458 0 25486 240 4 rbl_8
rlabel metal2 s 25646 0 25674 240 4 data_8
rlabel metal2 s 28570 0 28598 240 4 rbl_9
rlabel metal2 s 28758 0 28786 240 4 data_9
rlabel metal2 s 31682 0 31710 240 4 rbl_10
rlabel metal2 s 31870 0 31898 240 4 data_10
rlabel metal2 s 34794 0 34822 240 4 rbl_11
rlabel metal2 s 34982 0 35010 240 4 data_11
rlabel metal2 s 37906 0 37934 240 4 rbl_12
rlabel metal2 s 38094 0 38122 240 4 data_12
rlabel metal2 s 41018 0 41046 240 4 rbl_13
rlabel metal2 s 41206 0 41234 240 4 data_13
rlabel metal2 s 44130 0 44158 240 4 rbl_14
rlabel metal2 s 44318 0 44346 240 4 data_14
rlabel metal2 s 47242 0 47270 240 4 rbl_15
rlabel metal2 s 47430 0 47458 240 4 data_15
rlabel metal2 s 50354 0 50382 240 4 rbl_16
rlabel metal2 s 50542 0 50570 240 4 data_16
rlabel metal2 s 53466 0 53494 240 4 rbl_17
rlabel metal2 s 53654 0 53682 240 4 data_17
rlabel metal2 s 56578 0 56606 240 4 rbl_18
rlabel metal2 s 56766 0 56794 240 4 data_18
rlabel metal2 s 59690 0 59718 240 4 rbl_19
rlabel metal2 s 59878 0 59906 240 4 data_19
rlabel metal2 s 62802 0 62830 240 4 rbl_20
rlabel metal2 s 62990 0 63018 240 4 data_20
rlabel metal2 s 65914 0 65942 240 4 rbl_21
rlabel metal2 s 66102 0 66130 240 4 data_21
rlabel metal2 s 69026 0 69054 240 4 rbl_22
rlabel metal2 s 69214 0 69242 240 4 data_22
rlabel metal2 s 72138 0 72166 240 4 rbl_23
rlabel metal2 s 72326 0 72354 240 4 data_23
rlabel metal2 s 75250 0 75278 240 4 rbl_24
rlabel metal2 s 75438 0 75466 240 4 data_24
rlabel metal2 s 78362 0 78390 240 4 rbl_25
rlabel metal2 s 78550 0 78578 240 4 data_25
rlabel metal2 s 81474 0 81502 240 4 rbl_26
rlabel metal2 s 81662 0 81690 240 4 data_26
rlabel metal2 s 84586 0 84614 240 4 rbl_27
rlabel metal2 s 84774 0 84802 240 4 data_27
rlabel metal2 s 87698 0 87726 240 4 rbl_28
rlabel metal2 s 87886 0 87914 240 4 data_28
rlabel metal2 s 90810 0 90838 240 4 rbl_29
rlabel metal2 s 90998 0 91026 240 4 data_29
rlabel metal2 s 93922 0 93950 240 4 rbl_30
rlabel metal2 s 94110 0 94138 240 4 data_30
rlabel metal2 s 97034 0 97062 240 4 rbl_31
rlabel metal2 s 97222 0 97250 240 4 data_31
<< properties >>
string FIXED_BBOX 0 0 97292 1050
string GDS_FILE sram_0rw2r1w_16_128_sky130A.gds
string GDS_END 1520782
string GDS_START 1485854
<< end >>
