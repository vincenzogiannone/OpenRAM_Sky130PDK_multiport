magic
tech sky130A
magscale 1 2
timestamp 1643678851
<< checkpaint >>
rect -1260 -1294 3616 4646
<< locali >>
rect 0 3335 419 3369
rect 453 3335 1514 3369
rect 1548 3335 2320 3369
rect 2148 2958 2182 2992
rect 0 2497 419 2531
rect 453 2497 1514 2531
rect 1548 2497 2320 2531
rect 2148 2036 2182 2070
rect 0 1659 419 1693
rect 453 1659 1514 1693
rect 1548 1659 2320 1693
rect 2148 1282 2182 1316
rect 0 821 419 855
rect 453 821 1514 855
rect 1548 821 2320 855
rect 2148 360 2182 394
rect 0 -17 419 17
rect 453 -17 1514 17
rect 1548 -17 2320 17
<< viali >>
rect 419 3335 453 3369
rect 1514 3335 1548 3369
rect 1703 3045 1737 3079
rect 1803 2797 1837 2831
rect 419 2497 453 2531
rect 1514 2497 1548 2531
rect 1803 2197 1837 2231
rect 1703 1949 1737 1983
rect 419 1659 453 1693
rect 1514 1659 1548 1693
rect 1703 1369 1737 1403
rect 560 1282 594 1316
rect 692 1282 726 1316
rect 1803 1121 1837 1155
rect 419 821 453 855
rect 1514 821 1548 855
rect 1803 521 1837 555
rect 560 360 594 394
rect 692 360 726 394
rect 1703 273 1737 307
rect 419 -17 453 17
rect 1514 -17 1548 17
<< metal1 >>
rect 407 3367 410 3375
rect 381 3337 410 3367
rect 407 3329 410 3337
rect 462 3367 465 3375
rect 1502 3367 1505 3375
rect 462 3337 492 3367
rect 1476 3337 1505 3367
rect 462 3329 465 3337
rect 1502 3329 1505 3337
rect 1557 3367 1560 3375
rect 1557 3337 1587 3367
rect 1557 3329 1560 3337
rect 164 3048 1207 3076
rect 1691 3079 1749 3085
rect 1691 3076 1703 3079
rect 1259 3048 1703 3076
rect 1691 3045 1703 3048
rect 1737 3045 1749 3079
rect 1691 3039 1749 3045
rect 288 2800 1331 2828
rect 1791 2831 1849 2837
rect 1791 2828 1803 2831
rect 1383 2800 1803 2828
rect 1791 2797 1803 2800
rect 1837 2797 1849 2831
rect 1791 2791 1849 2797
rect 407 2529 410 2537
rect 381 2499 410 2529
rect 407 2491 410 2499
rect 462 2529 465 2537
rect 1502 2529 1505 2537
rect 462 2499 492 2529
rect 1476 2499 1505 2529
rect 462 2491 465 2499
rect 1502 2491 1505 2499
rect 1557 2529 1560 2537
rect 1557 2499 1587 2529
rect 1557 2491 1560 2499
rect 1791 2231 1849 2237
rect 1791 2228 1803 2231
rect 1383 2200 1803 2228
rect 1791 2197 1803 2200
rect 1837 2197 1849 2231
rect 1791 2191 1849 2197
rect 1691 1983 1749 1989
rect 1691 1980 1703 1983
rect 1011 1952 1703 1980
rect 1691 1949 1703 1952
rect 1737 1949 1749 1983
rect 1691 1943 1749 1949
rect 407 1691 410 1699
rect 381 1661 410 1691
rect 407 1653 410 1661
rect 462 1691 465 1699
rect 1502 1691 1505 1699
rect 462 1661 492 1691
rect 1476 1661 1505 1691
rect 462 1653 465 1661
rect 1502 1653 1505 1661
rect 1557 1691 1560 1699
rect 1557 1661 1587 1691
rect 1557 1653 1560 1661
rect 833 1604 1083 1632
rect 548 1316 606 1322
rect 548 1313 560 1316
rect 288 1285 560 1313
rect 548 1282 560 1285
rect 594 1282 606 1316
rect 548 1276 606 1282
rect 680 1316 738 1322
rect 680 1282 692 1316
rect 726 1313 738 1316
rect 833 1313 861 1604
rect 1691 1403 1749 1409
rect 1691 1400 1703 1403
rect 1259 1372 1703 1400
rect 1691 1369 1703 1372
rect 1737 1369 1749 1403
rect 1691 1363 1749 1369
rect 726 1285 861 1313
rect 726 1282 738 1285
rect 680 1276 738 1282
rect 1791 1155 1849 1161
rect 1791 1152 1803 1155
rect 1135 1124 1803 1152
rect 1791 1121 1803 1124
rect 1837 1121 1849 1155
rect 1791 1115 1849 1121
rect 407 853 410 861
rect 381 823 410 853
rect 407 815 410 823
rect 462 853 465 861
rect 1502 853 1505 861
rect 462 823 492 853
rect 1476 823 1505 853
rect 462 815 465 823
rect 1502 815 1505 823
rect 1557 853 1560 861
rect 1557 823 1587 853
rect 1557 815 1560 823
rect 833 766 959 794
rect 548 394 606 400
rect 548 391 560 394
rect 164 363 560 391
rect 548 360 560 363
rect 594 360 606 394
rect 548 354 606 360
rect 680 394 738 400
rect 680 360 692 394
rect 726 391 738 394
rect 833 391 861 766
rect 1791 555 1849 561
rect 1791 552 1803 555
rect 1135 524 1803 552
rect 1791 521 1803 524
rect 1837 521 1849 555
rect 1791 515 1849 521
rect 726 363 861 391
rect 726 360 738 363
rect 680 354 738 360
rect 1691 307 1749 313
rect 1691 304 1703 307
rect 1011 276 1703 304
rect 1691 273 1703 276
rect 1737 273 1749 307
rect 1691 267 1749 273
rect 407 15 410 23
rect 381 -15 410 15
rect 407 -23 410 -15
rect 462 15 465 23
rect 1502 15 1505 23
rect 462 -15 492 15
rect 1476 -15 1505 15
rect 462 -23 465 -15
rect 1502 -23 1505 -15
rect 1557 15 1560 23
rect 1557 -15 1587 15
rect 1557 -23 1560 -15
<< via1 >>
rect 410 3369 462 3378
rect 410 3335 419 3369
rect 419 3335 453 3369
rect 453 3335 462 3369
rect 1505 3369 1557 3378
rect 410 3326 462 3335
rect 1505 3335 1514 3369
rect 1514 3335 1548 3369
rect 1548 3335 1557 3369
rect 1505 3326 1557 3335
rect 112 3036 164 3088
rect 1207 3036 1259 3088
rect 236 2788 288 2840
rect 1331 2788 1383 2840
rect 410 2531 462 2540
rect 410 2497 419 2531
rect 419 2497 453 2531
rect 453 2497 462 2531
rect 1505 2531 1557 2540
rect 410 2488 462 2497
rect 1505 2497 1514 2531
rect 1514 2497 1548 2531
rect 1548 2497 1557 2531
rect 1505 2488 1557 2497
rect 1331 2188 1383 2240
rect 959 1940 1011 1992
rect 410 1693 462 1702
rect 410 1659 419 1693
rect 419 1659 453 1693
rect 453 1659 462 1693
rect 1505 1693 1557 1702
rect 410 1650 462 1659
rect 1505 1659 1514 1693
rect 1514 1659 1548 1693
rect 1548 1659 1557 1693
rect 1505 1650 1557 1659
rect 236 1273 288 1325
rect 1083 1592 1135 1644
rect 1207 1360 1259 1412
rect 1083 1112 1135 1164
rect 410 855 462 864
rect 410 821 419 855
rect 419 821 453 855
rect 453 821 462 855
rect 1505 855 1557 864
rect 410 812 462 821
rect 1505 821 1514 855
rect 1514 821 1548 855
rect 1548 821 1557 855
rect 1505 812 1557 821
rect 112 351 164 403
rect 959 754 1011 806
rect 1083 512 1135 564
rect 959 264 1011 316
rect 410 17 462 26
rect 410 -17 419 17
rect 419 -17 453 17
rect 453 -17 462 17
rect 1505 17 1557 26
rect 410 -26 462 -17
rect 1505 -17 1514 17
rect 1514 -17 1548 17
rect 1548 -17 1557 17
rect 1505 -26 1557 -17
<< metal2 >>
rect 416 3380 456 3386
rect 1511 3380 1551 3386
rect 124 3088 152 3352
rect 124 403 152 3036
rect 248 2840 276 3352
rect 416 3318 456 3324
rect 248 1325 276 2788
rect 416 2542 456 2548
rect 416 2480 456 2486
rect 971 1992 999 3352
rect 416 1704 456 1710
rect 416 1642 456 1648
rect 124 124 152 351
rect 248 124 276 1273
rect 416 866 456 872
rect 416 804 456 810
rect 971 806 999 1940
rect 1095 1644 1123 3352
rect 1219 3088 1247 3352
rect 1095 1164 1123 1592
rect 1219 1412 1247 3036
rect 1343 2840 1371 3352
rect 1511 3318 1551 3324
rect 1343 2240 1371 2788
rect 1511 2542 1551 2548
rect 1511 2480 1551 2486
rect 971 316 999 754
rect 1095 564 1123 1112
rect 971 124 999 264
rect 1095 124 1123 512
rect 1219 124 1247 1360
rect 1343 124 1371 2188
rect 1511 1704 1551 1710
rect 1511 1642 1551 1648
rect 1511 866 1551 872
rect 1511 804 1551 810
rect 416 28 456 34
rect 1511 28 1551 34
rect 416 -34 456 -28
rect 1511 -34 1551 -28
<< via2 >>
rect 408 3378 464 3380
rect 408 3326 410 3378
rect 410 3326 462 3378
rect 462 3326 464 3378
rect 1503 3378 1559 3380
rect 408 3324 464 3326
rect 408 2540 464 2542
rect 408 2488 410 2540
rect 410 2488 462 2540
rect 462 2488 464 2540
rect 408 2486 464 2488
rect 408 1702 464 1704
rect 408 1650 410 1702
rect 410 1650 462 1702
rect 462 1650 464 1702
rect 408 1648 464 1650
rect 408 864 464 866
rect 408 812 410 864
rect 410 812 462 864
rect 462 812 464 864
rect 408 810 464 812
rect 1503 3326 1505 3378
rect 1505 3326 1557 3378
rect 1557 3326 1559 3378
rect 1503 3324 1559 3326
rect 1503 2540 1559 2542
rect 1503 2488 1505 2540
rect 1505 2488 1557 2540
rect 1557 2488 1559 2540
rect 1503 2486 1559 2488
rect 1503 1702 1559 1704
rect 1503 1650 1505 1702
rect 1505 1650 1557 1702
rect 1557 1650 1559 1702
rect 1503 1648 1559 1650
rect 1503 864 1559 866
rect 1503 812 1505 864
rect 1505 812 1557 864
rect 1557 812 1559 864
rect 1503 810 1559 812
rect 408 26 464 28
rect 408 -26 410 26
rect 410 -26 462 26
rect 462 -26 464 26
rect 408 -28 464 -26
rect 1503 26 1559 28
rect 1503 -26 1505 26
rect 1505 -26 1557 26
rect 1557 -26 1559 26
rect 1503 -28 1559 -26
<< metal3 >>
rect 370 3380 502 3385
rect 370 3324 408 3380
rect 464 3324 502 3380
rect 370 3319 502 3324
rect 1465 3380 1597 3385
rect 1465 3324 1503 3380
rect 1559 3324 1597 3380
rect 1465 3319 1597 3324
rect 370 2542 502 2547
rect 370 2486 408 2542
rect 464 2486 502 2542
rect 370 2481 502 2486
rect 1465 2542 1597 2547
rect 1465 2486 1503 2542
rect 1559 2486 1597 2542
rect 1465 2481 1597 2486
rect 370 1704 502 1709
rect 370 1648 408 1704
rect 464 1648 502 1704
rect 370 1643 502 1648
rect 1465 1704 1597 1709
rect 1465 1648 1503 1704
rect 1559 1648 1597 1704
rect 1465 1643 1597 1648
rect 370 866 502 871
rect 370 810 408 866
rect 464 810 502 866
rect 370 805 502 810
rect 1465 866 1597 871
rect 1465 810 1503 866
rect 1559 810 1597 866
rect 1465 805 1597 810
rect 370 28 502 33
rect 370 -28 408 28
rect 464 -28 502 28
rect 370 -33 502 -28
rect 1465 28 1597 33
rect 1465 -28 1503 28
rect 1559 -28 1597 28
rect 1465 -33 1597 -28
use contact_18  contact_18_0
timestamp 1643678851
transform 1 0 1465 0 1 3319
box 0 0 1 1
use contact_17  contact_17_0
timestamp 1643678851
transform 1 0 1516 0 1 3337
box 0 0 1 1
use contact_13  contact_13_0
timestamp 1643678851
transform 1 0 1502 0 1 3329
box 0 0 1 1
use contact_18  contact_18_1
timestamp 1643678851
transform 1 0 370 0 1 3319
box 0 0 1 1
use contact_17  contact_17_1
timestamp 1643678851
transform 1 0 421 0 1 3337
box 0 0 1 1
use contact_13  contact_13_1
timestamp 1643678851
transform 1 0 407 0 1 3329
box 0 0 1 1
use contact_18  contact_18_2
timestamp 1643678851
transform 1 0 1465 0 1 2481
box 0 0 1 1
use contact_17  contact_17_2
timestamp 1643678851
transform 1 0 1516 0 1 2499
box 0 0 1 1
use contact_13  contact_13_2
timestamp 1643678851
transform 1 0 1502 0 1 2491
box 0 0 1 1
use contact_18  contact_18_3
timestamp 1643678851
transform 1 0 370 0 1 2481
box 0 0 1 1
use contact_17  contact_17_3
timestamp 1643678851
transform 1 0 421 0 1 2499
box 0 0 1 1
use contact_13  contact_13_3
timestamp 1643678851
transform 1 0 407 0 1 2491
box 0 0 1 1
use contact_18  contact_18_4
timestamp 1643678851
transform 1 0 1465 0 1 1643
box 0 0 1 1
use contact_17  contact_17_4
timestamp 1643678851
transform 1 0 1516 0 1 1661
box 0 0 1 1
use contact_13  contact_13_4
timestamp 1643678851
transform 1 0 1502 0 1 1653
box 0 0 1 1
use contact_18  contact_18_5
timestamp 1643678851
transform 1 0 370 0 1 1643
box 0 0 1 1
use contact_17  contact_17_5
timestamp 1643678851
transform 1 0 421 0 1 1661
box 0 0 1 1
use contact_13  contact_13_5
timestamp 1643678851
transform 1 0 407 0 1 1653
box 0 0 1 1
use contact_18  contact_18_6
timestamp 1643678851
transform 1 0 1465 0 1 2481
box 0 0 1 1
use contact_17  contact_17_6
timestamp 1643678851
transform 1 0 1516 0 1 2499
box 0 0 1 1
use contact_13  contact_13_6
timestamp 1643678851
transform 1 0 1502 0 1 2491
box 0 0 1 1
use contact_18  contact_18_7
timestamp 1643678851
transform 1 0 370 0 1 2481
box 0 0 1 1
use contact_17  contact_17_7
timestamp 1643678851
transform 1 0 421 0 1 2499
box 0 0 1 1
use contact_13  contact_13_7
timestamp 1643678851
transform 1 0 407 0 1 2491
box 0 0 1 1
use contact_18  contact_18_8
timestamp 1643678851
transform 1 0 1465 0 1 1643
box 0 0 1 1
use contact_17  contact_17_8
timestamp 1643678851
transform 1 0 1516 0 1 1661
box 0 0 1 1
use contact_13  contact_13_8
timestamp 1643678851
transform 1 0 1502 0 1 1653
box 0 0 1 1
use contact_18  contact_18_9
timestamp 1643678851
transform 1 0 370 0 1 1643
box 0 0 1 1
use contact_17  contact_17_9
timestamp 1643678851
transform 1 0 421 0 1 1661
box 0 0 1 1
use contact_13  contact_13_9
timestamp 1643678851
transform 1 0 407 0 1 1653
box 0 0 1 1
use contact_18  contact_18_10
timestamp 1643678851
transform 1 0 1465 0 1 805
box 0 0 1 1
use contact_17  contact_17_10
timestamp 1643678851
transform 1 0 1516 0 1 823
box 0 0 1 1
use contact_13  contact_13_10
timestamp 1643678851
transform 1 0 1502 0 1 815
box 0 0 1 1
use contact_18  contact_18_11
timestamp 1643678851
transform 1 0 370 0 1 805
box 0 0 1 1
use contact_17  contact_17_11
timestamp 1643678851
transform 1 0 421 0 1 823
box 0 0 1 1
use contact_13  contact_13_11
timestamp 1643678851
transform 1 0 407 0 1 815
box 0 0 1 1
use contact_18  contact_18_12
timestamp 1643678851
transform 1 0 1465 0 1 -33
box 0 0 1 1
use contact_17  contact_17_12
timestamp 1643678851
transform 1 0 1516 0 1 -15
box 0 0 1 1
use contact_13  contact_13_12
timestamp 1643678851
transform 1 0 1502 0 1 -23
box 0 0 1 1
use contact_18  contact_18_13
timestamp 1643678851
transform 1 0 370 0 1 -33
box 0 0 1 1
use contact_17  contact_17_13
timestamp 1643678851
transform 1 0 421 0 1 -15
box 0 0 1 1
use contact_13  contact_13_13
timestamp 1643678851
transform 1 0 407 0 1 -23
box 0 0 1 1
use contact_18  contact_18_14
timestamp 1643678851
transform 1 0 1465 0 1 805
box 0 0 1 1
use contact_17  contact_17_14
timestamp 1643678851
transform 1 0 1516 0 1 823
box 0 0 1 1
use contact_13  contact_13_14
timestamp 1643678851
transform 1 0 1502 0 1 815
box 0 0 1 1
use contact_18  contact_18_15
timestamp 1643678851
transform 1 0 370 0 1 805
box 0 0 1 1
use contact_17  contact_17_15
timestamp 1643678851
transform 1 0 421 0 1 823
box 0 0 1 1
use contact_13  contact_13_15
timestamp 1643678851
transform 1 0 407 0 1 815
box 0 0 1 1
use contact_17  contact_17_16
timestamp 1643678851
transform 1 0 1342 0 1 2799
box 0 0 1 1
use contact_17  contact_17_17
timestamp 1643678851
transform 1 0 247 0 1 2799
box 0 0 1 1
use contact_17  contact_17_18
timestamp 1643678851
transform 1 0 1218 0 1 3047
box 0 0 1 1
use contact_17  contact_17_19
timestamp 1643678851
transform 1 0 123 0 1 3047
box 0 0 1 1
use contact_14  contact_14_0
timestamp 1643678851
transform 1 0 1094 0 1 1603
box 0 0 1 1
use contact_13  contact_13_16
timestamp 1643678851
transform 1 0 680 0 1 1276
box 0 0 1 1
use contact_14  contact_14_1
timestamp 1643678851
transform 1 0 970 0 1 765
box 0 0 1 1
use contact_13  contact_13_17
timestamp 1643678851
transform 1 0 680 0 1 354
box 0 0 1 1
use contact_15  contact_15_0
timestamp 1643678851
transform 1 0 1791 0 1 2791
box 0 0 1 1
use contact_14  contact_14_2
timestamp 1643678851
transform 1 0 1342 0 1 2799
box 0 0 1 1
use contact_13  contact_13_18
timestamp 1643678851
transform 1 0 1691 0 1 3039
box 0 0 1 1
use contact_14  contact_14_3
timestamp 1643678851
transform 1 0 1218 0 1 3047
box 0 0 1 1
use contact_15  contact_15_1
timestamp 1643678851
transform 1 0 1791 0 1 2191
box 0 0 1 1
use contact_14  contact_14_4
timestamp 1643678851
transform 1 0 1342 0 1 2199
box 0 0 1 1
use contact_13  contact_13_19
timestamp 1643678851
transform 1 0 1691 0 1 1943
box 0 0 1 1
use contact_14  contact_14_5
timestamp 1643678851
transform 1 0 970 0 1 1951
box 0 0 1 1
use contact_15  contact_15_2
timestamp 1643678851
transform 1 0 1791 0 1 1115
box 0 0 1 1
use contact_14  contact_14_6
timestamp 1643678851
transform 1 0 1094 0 1 1123
box 0 0 1 1
use contact_13  contact_13_20
timestamp 1643678851
transform 1 0 1691 0 1 1363
box 0 0 1 1
use contact_14  contact_14_7
timestamp 1643678851
transform 1 0 1218 0 1 1371
box 0 0 1 1
use contact_15  contact_15_3
timestamp 1643678851
transform 1 0 1791 0 1 515
box 0 0 1 1
use contact_14  contact_14_8
timestamp 1643678851
transform 1 0 1094 0 1 523
box 0 0 1 1
use contact_13  contact_13_21
timestamp 1643678851
transform 1 0 1691 0 1 267
box 0 0 1 1
use contact_14  contact_14_9
timestamp 1643678851
transform 1 0 970 0 1 275
box 0 0 1 1
use contact_14  contact_14_10
timestamp 1643678851
transform 1 0 247 0 1 1284
box 0 0 1 1
use contact_13  contact_13_22
timestamp 1643678851
transform 1 0 548 0 1 1276
box 0 0 1 1
use contact_14  contact_14_11
timestamp 1643678851
transform 1 0 123 0 1 362
box 0 0 1 1
use contact_13  contact_13_23
timestamp 1643678851
transform 1 0 548 0 1 354
box 0 0 1 1
use pand2  pand2_0
timestamp 1643678851
transform 1 0 1591 0 -1 3352
box -36 -17 765 895
use pand2  pand2_1
timestamp 1643678851
transform 1 0 1591 0 1 1676
box -36 -17 765 895
use pand2  pand2_2
timestamp 1643678851
transform 1 0 1591 0 -1 1676
box -36 -17 765 895
use pand2  pand2_3
timestamp 1643678851
transform 1 0 1591 0 1 0
box -36 -17 765 895
use pinv_1  pinv_1_0
timestamp 1643678851
transform 1 0 496 0 -1 1676
box -36 -17 387 895
use pinv_1  pinv_1_1
timestamp 1643678851
transform 1 0 496 0 1 0
box -36 -17 387 895
<< labels >>
rlabel metal2 s 123 362 153 392 4 in_0
rlabel metal2 s 247 1284 277 1314 4 in_1
rlabel locali s 2165 377 2165 377 4 out_0
rlabel locali s 2165 1299 2165 1299 4 out_1
rlabel locali s 2165 2053 2165 2053 4 out_2
rlabel locali s 2165 2975 2165 2975 4 out_3
rlabel metal3 s 370 805 502 871 4 vdd
rlabel metal3 s 1465 2481 1597 2547 4 vdd
rlabel metal3 s 370 2481 502 2547 4 vdd
rlabel metal3 s 1465 805 1597 871 4 vdd
rlabel metal3 s 1465 -33 1597 33 4 gnd
rlabel metal3 s 1465 1643 1597 1709 4 gnd
rlabel metal3 s 370 3319 502 3385 4 gnd
rlabel metal3 s 370 1643 502 1709 4 gnd
rlabel metal3 s 1465 3319 1597 3385 4 gnd
rlabel metal3 s 370 -33 502 33 4 gnd
<< properties >>
string FIXED_BBOX 1465 -33 1597 0
string GDS_FILE sram_0rw2r1w_16_128_sky130A.gds
string GDS_END 1993850
string GDS_START 1983382
<< end >>
