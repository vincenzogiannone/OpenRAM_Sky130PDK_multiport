magic
tech sky130A
magscale 1 2
timestamp 1644969367
<< checkpaint >>
rect -1296 -1277 5252 2155
<< nwell >>
rect -36 402 3992 895
<< locali >>
rect 0 821 3956 855
rect 48 344 114 410
rect 196 360 449 394
rect 551 353 925 387
rect 1260 353 1833 387
rect 2799 353 2833 387
rect 0 -17 3956 17
use pinv_13  pinv_13_0
timestamp 1644969367
transform 1 0 1752 0 1 0
box -36 -17 2240 895
use pinv_12  pinv_12_0
timestamp 1644969367
transform 1 0 844 0 1 0
box -36 -17 944 895
use pinv_11  pinv_11_0
timestamp 1644969367
transform 1 0 368 0 1 0
box -36 -17 512 895
use pinv_6  pinv_6_0
timestamp 1644969367
transform 1 0 0 0 1 0
box -36 -17 404 895
<< labels >>
rlabel locali s 2816 370 2816 370 4 Z
rlabel locali s 81 377 81 377 4 A
rlabel locali s 1978 0 1978 0 4 gnd
rlabel locali s 1978 838 1978 838 4 vdd
<< properties >>
string FIXED_BBOX 0 0 3956 838
string GDS_FILE sram_0rw2r1w_32_128_sky130A.gds
string GDS_END 3373908
string GDS_START 3372630
<< end >>
