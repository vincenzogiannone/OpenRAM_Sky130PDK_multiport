magic
tech sky130A
magscale 1 2
timestamp 1643678851
<< checkpaint >>
rect -1296 -1277 3996 2155
<< nwell >>
rect -36 402 2736 895
<< locali >>
rect 0 821 2700 855
rect 48 344 114 410
rect 196 360 432 394
rect 547 360 783 394
rect 993 356 1458 390
rect 1992 356 2026 390
rect 0 -17 2700 17
use pinv_12  pinv_12_0
timestamp 1643678851
transform 1 0 1377 0 1 0
box -36 -17 1359 895
use pinv_11  pinv_11_0
timestamp 1643678851
transform 1 0 702 0 1 0
box -36 -17 711 895
use pinv_0  pinv_0_0
timestamp 1643678851
transform 1 0 351 0 1 0
box -36 -17 387 895
use pinv_0  pinv_0_1
timestamp 1643678851
transform 1 0 0 0 1 0
box -36 -17 387 895
<< labels >>
rlabel locali s 2009 373 2009 373 4 Z
rlabel locali s 81 377 81 377 4 A
rlabel locali s 1350 0 1350 0 4 gnd
rlabel locali s 1350 838 1350 838 4 vdd
<< properties >>
string FIXED_BBOX 0 0 2700 838
string GDS_FILE sram_0rw2r1w_16_128_sky130A.gds
string GDS_END 2096102
string GDS_START 2094826
<< end >>
