magic
tech sky130A
magscale 1 2
timestamp 1643678851
<< checkpaint >>
rect -1296 -1277 4185 2155
<< locali >>
rect 0 821 2889 855
rect 196 505 262 571
rect 330 388 364 561
rect 330 354 459 388
rect 1639 354 1673 388
rect 96 257 162 323
rect 0 -17 2889 17
use pdriver_3  pdriver_3_0
timestamp 1643678851
transform 1 0 378 0 1 0
box -36 -17 2547 895
use pnand2_0  pnand2_0_0
timestamp 1643678851
transform 1 0 0 0 1 0
box -36 -17 414 895
<< labels >>
rlabel locali s 1656 371 1656 371 4 Z
rlabel locali s 129 290 129 290 4 A
rlabel locali s 229 538 229 538 4 B
rlabel locali s 1444 0 1444 0 4 gnd
rlabel locali s 1444 838 1444 838 4 vdd
<< properties >>
string FIXED_BBOX 0 0 2889 838
string GDS_FILE sram_0rw2r1w_16_128_sky130A.gds
string GDS_END 2106660
string GDS_START 2105526
<< end >>
