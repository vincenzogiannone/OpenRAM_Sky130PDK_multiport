magic
tech sky130A
magscale 1 2
timestamp 1644949024
<< checkpaint >>
rect -1260 -854 5150 5248
<< metal1 >>
rect 0 3580 3092 3608
rect 0 1419 3890 1447
<< metal2 >>
rect 196 3664 250 3692
rect 994 3664 1048 3692
rect 1792 3664 1846 3692
rect 2590 3664 2644 3692
rect 630 3012 658 3642
rect 202 2520 230 2760
rect 474 2520 502 2760
rect 980 2520 1008 2760
rect 1252 2520 1280 2760
rect 70 420 98 1458
rect 532 420 560 1458
rect 848 420 876 1458
rect 1310 420 1338 1458
rect 1626 420 1654 1458
rect 2088 420 2116 1458
rect 2404 420 2432 1458
rect 2866 420 2894 1458
<< metal3 >>
rect 316 3856 382 3988
rect 1114 3856 1180 3988
rect 1912 3856 1978 3988
rect 2710 3856 2776 3988
rect 316 3024 382 3156
rect 1114 3024 1180 3156
rect 1912 3024 1978 3156
rect 2710 3024 2776 3156
rect 70 2689 202 2763
rect 342 2689 474 2763
rect 848 2689 980 2763
rect 1120 2689 1252 2763
rect 1626 2689 1758 2763
rect 1898 2689 2030 2763
rect 2404 2689 2536 2763
rect 2676 2689 2808 2763
rect 70 1743 202 1817
rect 342 1743 474 1817
rect 848 1743 980 1817
rect 1120 1743 1252 1817
rect 1626 1743 1758 1817
rect 1898 1743 2030 1817
rect 2404 1743 2536 1817
rect 2676 1743 2808 1817
rect 160 464 226 596
rect 938 464 1004 596
rect 1716 464 1782 596
rect 2494 464 2560 596
rect 3272 464 3338 596
use write_driver_array  write_driver_array_0
timestamp 1644949024
transform 1 0 0 0 -1 3964
box 0 -24 3092 952
use sense_amp_array  sense_amp_array_0
timestamp 1644949024
transform 1 0 0 0 -1 2760
box 0 -3 2878 1050
use precharge_array_multiport  precharge_array_multiport_0
timestamp 1644949024
transform 1 0 0 0 -1 1458
box 0 -8 3890 1052
<< labels >>
rlabel metal2 s 196 3664 250 3692 4 din0_0
rlabel metal2 s 994 3664 1048 3692 4 din0_1
rlabel metal2 s 1792 3664 1846 3692 4 din0_2
rlabel metal2 s 2590 3664 2644 3692 4 din0_3
rlabel metal2 s 202 2520 230 2760 4 dout0_0
rlabel metal2 s 216 2640 216 2640 4 dout1_0
rlabel metal2 s 474 2520 502 2760 4 dout0_1
rlabel metal2 s 488 2640 488 2640 4 dout1_1
rlabel metal2 s 980 2520 1008 2760 4 dout0_2
rlabel metal2 s 994 2640 994 2640 4 dout1_2
rlabel metal2 s 1252 2520 1280 2760 4 dout0_3
rlabel metal2 s 1266 2640 1266 2640 4 dout1_3
rlabel metal2 s 70 420 98 1458 4 rbl0_0
rlabel metal2 s 532 420 560 1458 4 rbl1_0
rlabel metal2 s 848 420 876 1458 4 rbl0_1
rlabel metal2 s 1310 420 1338 1458 4 rbl1_1
rlabel metal2 s 1626 420 1654 1458 4 rbl0_2
rlabel metal2 s 2088 420 2116 1458 4 rbl1_2
rlabel metal2 s 2404 420 2432 1458 4 rbl0_3
rlabel metal2 s 2866 420 2894 1458 4 rbl1_3
rlabel metal2 s 630 3012 658 3642 4 wbl0_0
rlabel metal1 s 0 1418 3890 1446 4 p_en_bar
rlabel metal1 s 0 3580 3092 3608 4 w_en
rlabel metal3 s 2676 1742 2808 1816 4 vdd
rlabel metal3 s 316 3024 382 3156 4 vdd
rlabel metal3 s 1716 464 1782 596 4 vdd
rlabel metal3 s 1912 3024 1978 3156 4 vdd
rlabel metal3 s 2404 1742 2536 1816 4 vdd
rlabel metal3 s 2710 3024 2776 3156 4 vdd
rlabel metal3 s 3272 464 3338 596 4 vdd
rlabel metal3 s 938 464 1004 596 4 vdd
rlabel metal3 s 1626 1742 1758 1816 4 vdd
rlabel metal3 s 1898 1742 2030 1816 4 vdd
rlabel metal3 s 342 1742 474 1816 4 vdd
rlabel metal3 s 848 1742 980 1816 4 vdd
rlabel metal3 s 1114 3024 1180 3156 4 vdd
rlabel metal3 s 70 1742 202 1816 4 vdd
rlabel metal3 s 160 464 226 596 4 vdd
rlabel metal3 s 1120 1742 1252 1816 4 vdd
rlabel metal3 s 2494 464 2560 596 4 vdd
rlabel metal3 s 1626 2688 1758 2762 4 gnd
rlabel metal3 s 1120 2688 1252 2762 4 gnd
rlabel metal3 s 2676 2688 2808 2762 4 gnd
rlabel metal3 s 848 2688 980 2762 4 gnd
rlabel metal3 s 1898 2688 2030 2762 4 gnd
rlabel metal3 s 316 3856 382 3988 4 gnd
rlabel metal3 s 342 2688 474 2762 4 gnd
rlabel metal3 s 2710 3856 2776 3988 4 gnd
rlabel metal3 s 1114 3856 1180 3988 4 gnd
rlabel metal3 s 2404 2688 2536 2762 4 gnd
rlabel metal3 s 70 2688 202 2762 4 gnd
rlabel metal3 s 1912 3856 1978 3988 4 gnd
<< properties >>
string FIXED_BBOX 0 0 3890 3796
string GDS_FILE sram_0rw2r1w_4_16_sky130A.gds
string GDS_END 190312
string GDS_START 180296
<< end >>
