magic
tech sky130A
magscale 1 2
timestamp 1643593061
<< checkpaint >>
rect -1260 -1290 3340 7450
<< locali >>
rect 0 6143 291 6177
rect 325 6143 1163 6177
rect 1197 6143 2044 6177
rect 1855 5415 1889 5449
rect 0 4603 291 4637
rect 325 4603 1163 4637
rect 1197 4603 2044 4637
rect 1855 3791 1889 3825
rect 0 3063 291 3097
rect 325 3063 1163 3097
rect 1197 3063 2044 3097
rect 1855 2335 1889 2369
rect 0 1523 291 1557
rect 325 1523 1163 1557
rect 1197 1523 2044 1557
rect 1855 711 1889 745
rect 0 -17 291 17
rect 325 -17 1163 17
rect 1197 -17 2044 17
<< viali >>
rect 291 6143 325 6177
rect 1163 6143 1197 6177
rect 1320 5853 1354 5887
rect 1420 5613 1454 5647
rect 291 4603 325 4637
rect 1163 4603 1197 4637
rect 1420 3593 1454 3627
rect 1320 3353 1354 3387
rect 291 3063 325 3097
rect 1163 3063 1197 3097
rect 1320 2773 1354 2807
rect 1420 2533 1454 2567
rect 400 2335 434 2369
rect 532 2335 566 2369
rect 291 1523 325 1557
rect 1163 1523 1197 1557
rect 400 711 434 745
rect 532 711 566 745
rect 1420 513 1454 547
rect 1320 273 1354 307
rect 291 -17 325 17
rect 1163 -17 1197 17
<< metal1 >>
rect 276 6134 282 6186
rect 334 6134 340 6186
rect 1148 6134 1154 6186
rect 1206 6134 1212 6186
rect 66 5844 72 5896
rect 124 5884 130 5896
rect 938 5884 944 5896
rect 124 5856 944 5884
rect 124 5844 130 5856
rect 938 5844 944 5856
rect 996 5884 1002 5896
rect 1308 5887 1366 5893
rect 1308 5884 1320 5887
rect 996 5856 1320 5884
rect 996 5844 1002 5856
rect 1308 5853 1320 5856
rect 1354 5853 1366 5887
rect 1308 5847 1366 5853
rect 150 5604 156 5656
rect 208 5644 214 5656
rect 1022 5644 1028 5656
rect 208 5616 1028 5644
rect 208 5604 214 5616
rect 1022 5604 1028 5616
rect 1080 5644 1086 5656
rect 1408 5647 1466 5653
rect 1408 5644 1420 5647
rect 1080 5616 1420 5644
rect 1080 5604 1086 5616
rect 1408 5613 1420 5616
rect 1454 5613 1466 5647
rect 1408 5607 1466 5613
rect 276 4594 282 4646
rect 334 4594 340 4646
rect 1148 4594 1154 4646
rect 1206 4594 1212 4646
rect 1022 3584 1028 3636
rect 1080 3624 1086 3636
rect 1408 3627 1466 3633
rect 1408 3624 1420 3627
rect 1080 3596 1420 3624
rect 1080 3584 1086 3596
rect 1408 3593 1420 3596
rect 1454 3593 1466 3627
rect 1408 3587 1466 3593
rect 770 3344 776 3396
rect 828 3384 834 3396
rect 1308 3387 1366 3393
rect 1308 3384 1320 3387
rect 828 3356 1320 3384
rect 828 3344 834 3356
rect 1308 3353 1320 3356
rect 1354 3353 1366 3387
rect 1308 3347 1366 3353
rect 276 3054 282 3106
rect 334 3054 340 3106
rect 1148 3054 1154 3106
rect 1206 3054 1212 3106
rect 854 3014 860 3026
rect 690 2986 860 3014
rect 150 2326 156 2378
rect 208 2366 214 2378
rect 388 2369 446 2375
rect 388 2366 400 2369
rect 208 2338 400 2366
rect 208 2326 214 2338
rect 388 2335 400 2338
rect 434 2335 446 2369
rect 388 2329 446 2335
rect 520 2369 578 2375
rect 520 2335 532 2369
rect 566 2366 578 2369
rect 690 2366 718 2986
rect 854 2974 860 2986
rect 912 2974 918 3026
rect 938 2764 944 2816
rect 996 2804 1002 2816
rect 1308 2807 1366 2813
rect 1308 2804 1320 2807
rect 996 2776 1320 2804
rect 996 2764 1002 2776
rect 1308 2773 1320 2776
rect 1354 2773 1366 2807
rect 1308 2767 1366 2773
rect 854 2524 860 2576
rect 912 2564 918 2576
rect 1408 2567 1466 2573
rect 1408 2564 1420 2567
rect 912 2536 1420 2564
rect 912 2524 918 2536
rect 1408 2533 1420 2536
rect 1454 2533 1466 2567
rect 1408 2527 1466 2533
rect 566 2338 718 2366
rect 566 2335 578 2338
rect 520 2329 578 2335
rect 276 1514 282 1566
rect 334 1514 340 1566
rect 1148 1514 1154 1566
rect 1206 1514 1212 1566
rect 770 1474 776 1486
rect 690 1446 776 1474
rect 66 702 72 754
rect 124 742 130 754
rect 388 745 446 751
rect 388 742 400 745
rect 124 714 400 742
rect 124 702 130 714
rect 388 711 400 714
rect 434 711 446 745
rect 388 705 446 711
rect 520 745 578 751
rect 520 711 532 745
rect 566 742 578 745
rect 690 742 718 1446
rect 770 1434 776 1446
rect 828 1434 834 1486
rect 566 714 718 742
rect 566 711 578 714
rect 520 705 578 711
rect 854 504 860 556
rect 912 544 918 556
rect 1408 547 1466 553
rect 1408 544 1420 547
rect 912 516 1420 544
rect 912 504 918 516
rect 1408 513 1420 516
rect 1454 513 1466 547
rect 1408 507 1466 513
rect 770 264 776 316
rect 828 304 834 316
rect 1308 307 1366 313
rect 1308 304 1320 307
rect 828 276 1320 304
rect 828 264 834 276
rect 1308 273 1320 276
rect 1354 273 1366 307
rect 1308 267 1366 273
rect 276 -26 282 26
rect 334 -26 340 26
rect 1148 -26 1154 26
rect 1206 -26 1212 26
<< via1 >>
rect 282 6177 334 6186
rect 282 6143 291 6177
rect 291 6143 325 6177
rect 325 6143 334 6177
rect 282 6134 334 6143
rect 1154 6177 1206 6186
rect 1154 6143 1163 6177
rect 1163 6143 1197 6177
rect 1197 6143 1206 6177
rect 1154 6134 1206 6143
rect 72 5844 124 5896
rect 944 5844 996 5896
rect 156 5604 208 5656
rect 1028 5604 1080 5656
rect 282 4637 334 4646
rect 282 4603 291 4637
rect 291 4603 325 4637
rect 325 4603 334 4637
rect 282 4594 334 4603
rect 1154 4637 1206 4646
rect 1154 4603 1163 4637
rect 1163 4603 1197 4637
rect 1197 4603 1206 4637
rect 1154 4594 1206 4603
rect 1028 3584 1080 3636
rect 776 3344 828 3396
rect 282 3097 334 3106
rect 282 3063 291 3097
rect 291 3063 325 3097
rect 325 3063 334 3097
rect 282 3054 334 3063
rect 1154 3097 1206 3106
rect 1154 3063 1163 3097
rect 1163 3063 1197 3097
rect 1197 3063 1206 3097
rect 1154 3054 1206 3063
rect 156 2326 208 2378
rect 860 2974 912 3026
rect 944 2764 996 2816
rect 860 2524 912 2576
rect 282 1557 334 1566
rect 282 1523 291 1557
rect 291 1523 325 1557
rect 325 1523 334 1557
rect 282 1514 334 1523
rect 1154 1557 1206 1566
rect 1154 1523 1163 1557
rect 1163 1523 1197 1557
rect 1197 1523 1206 1557
rect 1154 1514 1206 1523
rect 72 702 124 754
rect 776 1434 828 1486
rect 860 504 912 556
rect 776 264 828 316
rect 282 17 334 26
rect 282 -17 291 17
rect 291 -17 325 17
rect 325 -17 334 17
rect 282 -26 334 -17
rect 1154 17 1206 26
rect 1154 -17 1163 17
rect 1163 -17 1197 17
rect 1197 -17 1206 17
rect 1154 -26 1206 -17
<< metal2 >>
rect 84 5896 112 6160
rect 84 754 112 5844
rect 168 5656 196 6160
rect 168 2378 196 5604
rect 788 3396 816 6160
rect 84 84 112 702
rect 168 84 196 2326
rect 788 1486 816 3344
rect 872 3026 900 6160
rect 956 5896 984 6160
rect 872 2576 900 2974
rect 956 2816 984 5844
rect 1040 5656 1068 6160
rect 1040 3636 1068 5604
rect 788 316 816 1434
rect 872 556 900 2524
rect 788 84 816 264
rect 872 84 900 504
rect 956 84 984 2764
rect 1040 84 1068 3584
<< via2 >>
rect 280 6186 336 6188
rect 280 6134 282 6186
rect 282 6134 334 6186
rect 334 6134 336 6186
rect 1152 6186 1208 6188
rect 280 6132 336 6134
rect 280 4646 336 4648
rect 280 4594 282 4646
rect 282 4594 334 4646
rect 334 4594 336 4646
rect 280 4592 336 4594
rect 280 3106 336 3108
rect 280 3054 282 3106
rect 282 3054 334 3106
rect 334 3054 336 3106
rect 280 3052 336 3054
rect 280 1566 336 1568
rect 280 1514 282 1566
rect 282 1514 334 1566
rect 334 1514 336 1566
rect 280 1512 336 1514
rect 1152 6134 1154 6186
rect 1154 6134 1206 6186
rect 1206 6134 1208 6186
rect 1152 6132 1208 6134
rect 1152 4646 1208 4648
rect 1152 4594 1154 4646
rect 1154 4594 1206 4646
rect 1206 4594 1208 4646
rect 1152 4592 1208 4594
rect 1152 3106 1208 3108
rect 1152 3054 1154 3106
rect 1154 3054 1206 3106
rect 1206 3054 1208 3106
rect 1152 3052 1208 3054
rect 1152 1566 1208 1568
rect 1152 1514 1154 1566
rect 1154 1514 1206 1566
rect 1206 1514 1208 1566
rect 1152 1512 1208 1514
rect 280 26 336 28
rect 280 -26 282 26
rect 282 -26 334 26
rect 334 -26 336 26
rect 280 -28 336 -26
rect 1152 26 1208 28
rect 1152 -26 1154 26
rect 1154 -26 1206 26
rect 1206 -26 1208 26
rect 1152 -28 1208 -26
<< metal3 >>
rect 278 6188 338 6190
rect 278 6132 280 6188
rect 336 6132 338 6188
rect 278 6130 338 6132
rect 1150 6188 1210 6190
rect 1150 6132 1152 6188
rect 1208 6132 1210 6188
rect 1150 6130 1210 6132
rect 278 4648 338 4650
rect 278 4592 280 4648
rect 336 4592 338 4648
rect 278 4590 338 4592
rect 1150 4648 1210 4650
rect 1150 4592 1152 4648
rect 1208 4592 1210 4648
rect 1150 4590 1210 4592
rect 278 3108 338 3110
rect 278 3052 280 3108
rect 336 3052 338 3108
rect 278 3050 338 3052
rect 1150 3108 1210 3110
rect 1150 3052 1152 3108
rect 1208 3052 1210 3108
rect 1150 3050 1210 3052
rect 278 1568 338 1570
rect 278 1512 280 1568
rect 336 1512 338 1568
rect 278 1510 338 1512
rect 1150 1568 1210 1570
rect 1150 1512 1152 1568
rect 1208 1512 1210 1568
rect 1150 1510 1210 1512
rect 278 28 338 30
rect 278 -28 280 28
rect 336 -28 338 28
rect 278 -30 338 -28
rect 1150 28 1210 30
rect 1150 -28 1152 28
rect 1208 -28 1210 28
rect 1150 -30 1210 -28
use contact_18  contact_18_0
timestamp 1643593061
transform 1 0 1150 0 1 6130
box 0 0 1 1
use contact_17  contact_17_0
timestamp 1643593061
transform 1 0 1148 0 1 6134
box 0 0 1 1
use contact_13  contact_13_0
timestamp 1643593061
transform 1 0 1151 0 1 6137
box 0 0 1 1
use contact_18  contact_18_1
timestamp 1643593061
transform 1 0 278 0 1 6130
box 0 0 1 1
use contact_17  contact_17_1
timestamp 1643593061
transform 1 0 276 0 1 6134
box 0 0 1 1
use contact_13  contact_13_1
timestamp 1643593061
transform 1 0 279 0 1 6137
box 0 0 1 1
use contact_18  contact_18_2
timestamp 1643593061
transform 1 0 1150 0 1 4590
box 0 0 1 1
use contact_17  contact_17_2
timestamp 1643593061
transform 1 0 1148 0 1 4594
box 0 0 1 1
use contact_13  contact_13_2
timestamp 1643593061
transform 1 0 1151 0 1 4597
box 0 0 1 1
use contact_18  contact_18_3
timestamp 1643593061
transform 1 0 278 0 1 4590
box 0 0 1 1
use contact_17  contact_17_3
timestamp 1643593061
transform 1 0 276 0 1 4594
box 0 0 1 1
use contact_13  contact_13_3
timestamp 1643593061
transform 1 0 279 0 1 4597
box 0 0 1 1
use contact_18  contact_18_4
timestamp 1643593061
transform 1 0 1150 0 1 3050
box 0 0 1 1
use contact_17  contact_17_4
timestamp 1643593061
transform 1 0 1148 0 1 3054
box 0 0 1 1
use contact_13  contact_13_4
timestamp 1643593061
transform 1 0 1151 0 1 3057
box 0 0 1 1
use contact_18  contact_18_5
timestamp 1643593061
transform 1 0 278 0 1 3050
box 0 0 1 1
use contact_17  contact_17_5
timestamp 1643593061
transform 1 0 276 0 1 3054
box 0 0 1 1
use contact_13  contact_13_5
timestamp 1643593061
transform 1 0 279 0 1 3057
box 0 0 1 1
use contact_18  contact_18_6
timestamp 1643593061
transform 1 0 1150 0 1 4590
box 0 0 1 1
use contact_17  contact_17_6
timestamp 1643593061
transform 1 0 1148 0 1 4594
box 0 0 1 1
use contact_13  contact_13_6
timestamp 1643593061
transform 1 0 1151 0 1 4597
box 0 0 1 1
use contact_18  contact_18_7
timestamp 1643593061
transform 1 0 278 0 1 4590
box 0 0 1 1
use contact_17  contact_17_7
timestamp 1643593061
transform 1 0 276 0 1 4594
box 0 0 1 1
use contact_13  contact_13_7
timestamp 1643593061
transform 1 0 279 0 1 4597
box 0 0 1 1
use contact_18  contact_18_8
timestamp 1643593061
transform 1 0 1150 0 1 3050
box 0 0 1 1
use contact_17  contact_17_8
timestamp 1643593061
transform 1 0 1148 0 1 3054
box 0 0 1 1
use contact_13  contact_13_8
timestamp 1643593061
transform 1 0 1151 0 1 3057
box 0 0 1 1
use contact_18  contact_18_9
timestamp 1643593061
transform 1 0 278 0 1 3050
box 0 0 1 1
use contact_17  contact_17_9
timestamp 1643593061
transform 1 0 276 0 1 3054
box 0 0 1 1
use contact_13  contact_13_9
timestamp 1643593061
transform 1 0 279 0 1 3057
box 0 0 1 1
use contact_18  contact_18_10
timestamp 1643593061
transform 1 0 1150 0 1 1510
box 0 0 1 1
use contact_17  contact_17_10
timestamp 1643593061
transform 1 0 1148 0 1 1514
box 0 0 1 1
use contact_13  contact_13_10
timestamp 1643593061
transform 1 0 1151 0 1 1517
box 0 0 1 1
use contact_18  contact_18_11
timestamp 1643593061
transform 1 0 278 0 1 1510
box 0 0 1 1
use contact_17  contact_17_11
timestamp 1643593061
transform 1 0 276 0 1 1514
box 0 0 1 1
use contact_13  contact_13_11
timestamp 1643593061
transform 1 0 279 0 1 1517
box 0 0 1 1
use contact_18  contact_18_12
timestamp 1643593061
transform 1 0 1150 0 1 -30
box 0 0 1 1
use contact_17  contact_17_12
timestamp 1643593061
transform 1 0 1148 0 1 -26
box 0 0 1 1
use contact_13  contact_13_12
timestamp 1643593061
transform 1 0 1151 0 1 -23
box 0 0 1 1
use contact_18  contact_18_13
timestamp 1643593061
transform 1 0 278 0 1 -30
box 0 0 1 1
use contact_17  contact_17_13
timestamp 1643593061
transform 1 0 276 0 1 -26
box 0 0 1 1
use contact_13  contact_13_13
timestamp 1643593061
transform 1 0 279 0 1 -23
box 0 0 1 1
use contact_18  contact_18_14
timestamp 1643593061
transform 1 0 1150 0 1 1510
box 0 0 1 1
use contact_17  contact_17_14
timestamp 1643593061
transform 1 0 1148 0 1 1514
box 0 0 1 1
use contact_13  contact_13_14
timestamp 1643593061
transform 1 0 1151 0 1 1517
box 0 0 1 1
use contact_18  contact_18_15
timestamp 1643593061
transform 1 0 278 0 1 1510
box 0 0 1 1
use contact_17  contact_17_15
timestamp 1643593061
transform 1 0 276 0 1 1514
box 0 0 1 1
use contact_13  contact_13_15
timestamp 1643593061
transform 1 0 279 0 1 1517
box 0 0 1 1
use contact_17  contact_17_16
timestamp 1643593061
transform 1 0 1022 0 1 5604
box 0 0 1 1
use contact_17  contact_17_17
timestamp 1643593061
transform 1 0 150 0 1 5604
box 0 0 1 1
use contact_17  contact_17_18
timestamp 1643593061
transform 1 0 938 0 1 5844
box 0 0 1 1
use contact_17  contact_17_19
timestamp 1643593061
transform 1 0 66 0 1 5844
box 0 0 1 1
use contact_14  contact_14_0
timestamp 1643593061
transform 1 0 854 0 1 2974
box 0 0 1 1
use contact_13  contact_13_16
timestamp 1643593061
transform 1 0 520 0 1 2329
box 0 0 1 1
use contact_14  contact_14_1
timestamp 1643593061
transform 1 0 770 0 1 1434
box 0 0 1 1
use contact_13  contact_13_17
timestamp 1643593061
transform 1 0 520 0 1 705
box 0 0 1 1
use contact_15  contact_15_0
timestamp 1643593061
transform 1 0 1408 0 1 5607
box 0 0 1 1
use contact_14  contact_14_2
timestamp 1643593061
transform 1 0 1022 0 1 5604
box 0 0 1 1
use contact_13  contact_13_18
timestamp 1643593061
transform 1 0 1308 0 1 5847
box 0 0 1 1
use contact_14  contact_14_3
timestamp 1643593061
transform 1 0 938 0 1 5844
box 0 0 1 1
use contact_15  contact_15_1
timestamp 1643593061
transform 1 0 1408 0 1 3587
box 0 0 1 1
use contact_14  contact_14_4
timestamp 1643593061
transform 1 0 1022 0 1 3584
box 0 0 1 1
use contact_13  contact_13_19
timestamp 1643593061
transform 1 0 1308 0 1 3347
box 0 0 1 1
use contact_14  contact_14_5
timestamp 1643593061
transform 1 0 770 0 1 3344
box 0 0 1 1
use contact_15  contact_15_2
timestamp 1643593061
transform 1 0 1408 0 1 2527
box 0 0 1 1
use contact_14  contact_14_6
timestamp 1643593061
transform 1 0 854 0 1 2524
box 0 0 1 1
use contact_13  contact_13_20
timestamp 1643593061
transform 1 0 1308 0 1 2767
box 0 0 1 1
use contact_14  contact_14_7
timestamp 1643593061
transform 1 0 938 0 1 2764
box 0 0 1 1
use contact_15  contact_15_3
timestamp 1643593061
transform 1 0 1408 0 1 507
box 0 0 1 1
use contact_14  contact_14_8
timestamp 1643593061
transform 1 0 854 0 1 504
box 0 0 1 1
use contact_13  contact_13_21
timestamp 1643593061
transform 1 0 1308 0 1 267
box 0 0 1 1
use contact_14  contact_14_9
timestamp 1643593061
transform 1 0 770 0 1 264
box 0 0 1 1
use contact_14  contact_14_10
timestamp 1643593061
transform 1 0 150 0 1 2326
box 0 0 1 1
use contact_13  contact_13_22
timestamp 1643593061
transform 1 0 388 0 1 2329
box 0 0 1 1
use contact_14  contact_14_11
timestamp 1643593061
transform 1 0 66 0 1 702
box 0 0 1 1
use contact_13  contact_13_23
timestamp 1643593061
transform 1 0 388 0 1 705
box 0 0 1 1
use and2_dec  and2_dec_0
timestamp 1643593061
transform 1 0 1208 0 -1 6160
box -36 -17 872 1597
use and2_dec  and2_dec_1
timestamp 1643593061
transform 1 0 1208 0 1 3080
box -36 -17 872 1597
use and2_dec  and2_dec_2
timestamp 1643593061
transform 1 0 1208 0 -1 3080
box -36 -17 872 1597
use and2_dec  and2_dec_3
timestamp 1643593061
transform 1 0 1208 0 1 0
box -36 -17 872 1597
use pinv  pinv_0
timestamp 1643593061
transform 1 0 336 0 -1 3080
box -36 -17 404 1597
use pinv  pinv_1
timestamp 1643593061
transform 1 0 336 0 1 0
box -36 -17 404 1597
<< labels >>
rlabel metal2 s 72 702 124 754 4 in_0
rlabel metal2 s 156 2326 208 2378 4 in_1
rlabel locali s 1872 728 1872 728 4 out_0
rlabel locali s 1872 2352 1872 2352 4 out_1
rlabel locali s 1872 3808 1872 3808 4 out_2
rlabel locali s 1872 5432 1872 5432 4 out_3
rlabel metal3 s 1150 4590 1210 4650 4 vdd
rlabel metal3 s 278 1510 338 1570 4 vdd
rlabel metal3 s 1150 1510 1210 1570 4 vdd
rlabel metal3 s 278 4590 338 4650 4 vdd
rlabel metal3 s 278 6130 338 6190 4 gnd
rlabel metal3 s 278 3050 338 3110 4 gnd
rlabel metal3 s 1150 3050 1210 3110 4 gnd
rlabel metal3 s 278 -30 338 30 4 gnd
rlabel metal3 s 1150 -30 1210 30 4 gnd
rlabel metal3 s 1150 6130 1210 6190 4 gnd
<< properties >>
string FIXED_BBOX 1150 -30 1210 -26
string GDS_FILE sram_0rw2r1w_2_16_sky130A.gds
string GDS_END 397146
string GDS_START 386674
<< end >>
