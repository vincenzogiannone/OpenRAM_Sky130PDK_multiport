magic
tech sky130A
magscale 1 2
timestamp 1643671299
<< checkpaint >>
rect -1296 -1260 2853 2970
<< locali >>
rect 0 1676 1593 1710
rect 213 1299 891 1333
rect 1101 1299 1135 1333
rect 0 838 1593 872
rect 64 377 98 411
rect 213 377 449 411
rect 551 377 908 411
rect 1101 377 1135 411
rect 0 0 1593 34
<< viali >>
rect 179 1299 213 1333
rect 179 377 213 411
<< metal1 >>
rect 167 1333 225 1339
rect 167 1299 179 1333
rect 213 1299 225 1333
rect 167 1293 225 1299
rect 182 417 210 1293
rect 167 411 225 417
rect 167 377 179 411
rect 213 377 225 411
rect 167 371 225 377
use contact_13  contact_13_0
timestamp 1643671299
transform 1 0 167 0 1 371
box 0 0 1 1
use contact_13  contact_13_1
timestamp 1643671299
transform 1 0 167 0 1 1293
box 0 0 1 1
use pinv_2  pinv_2_0
timestamp 1643671299
transform 1 0 810 0 -1 1693
box -36 -17 711 895
use pinv_2  pinv_2_1
timestamp 1643671299
transform 1 0 810 0 1 17
box -36 -17 711 895
use pinv_1  pinv_1_0
timestamp 1643671299
transform 1 0 351 0 1 17
box -36 -17 495 895
use pinv_0  pinv_0_0
timestamp 1643671299
transform 1 0 0 0 1 17
box -36 -17 387 895
<< labels >>
rlabel locali s 796 855 796 855 4 vdd
rlabel locali s 796 17 796 17 4 gnd
rlabel locali s 796 1693 796 1693 4 gnd
rlabel locali s 1118 1316 1118 1316 4 Z
rlabel locali s 1118 394 1118 394 4 Zb
rlabel locali s 81 394 81 394 4 A
<< properties >>
string FIXED_BBOX 0 0 1593 1693
string GDS_FILE sram_0rw2r1w_16_32_sky130A.gds
string GDS_END 1098508
string GDS_START 1096914
<< end >>
