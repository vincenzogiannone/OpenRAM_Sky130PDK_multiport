magic
tech sky130A
magscale 1 2
timestamp 1643678851
<< checkpaint >>
rect -1271 -1302 7894 50518
<< metal1 >>
rect 5501 48606 5914 48634
rect 5501 48514 5529 48606
rect 6540 48536 6568 48564
rect 5410 48486 5612 48514
rect 5410 48368 5438 48486
rect 5357 48340 5438 48368
rect 5357 47868 5385 48340
rect 5410 47868 5438 48340
rect 5501 47868 5529 48486
rect 6540 48410 6568 48438
rect 6540 48184 6568 48212
rect 5336 47840 5529 47868
rect 5357 47746 5385 47840
rect 5336 47718 5385 47746
rect 5410 47600 5438 47840
rect 5336 47572 5438 47600
rect 6540 47144 6568 47172
rect 5357 46988 5434 47016
rect 5357 46296 5385 46988
rect 6540 46918 6568 46946
rect 5410 46842 5612 46870
rect 5410 46296 5438 46842
rect 6540 46792 6568 46820
rect 5336 46268 5438 46296
rect 5501 46722 5914 46750
rect 5357 46150 5385 46268
rect 5336 46122 5385 46150
rect 5501 46028 5529 46722
rect 5336 46000 5529 46028
rect 5501 45530 5914 45558
rect 5501 45438 5529 45530
rect 6540 45460 6568 45488
rect 5410 45410 5612 45438
rect 5410 45292 5438 45410
rect 5357 45264 5438 45292
rect 5357 44840 5385 45264
rect 5410 44840 5438 45264
rect 5501 44840 5529 45410
rect 6540 45334 6568 45362
rect 6540 45108 6568 45136
rect 5336 44812 5529 44840
rect 5357 44718 5385 44812
rect 5336 44690 5385 44718
rect 5410 44572 5438 44812
rect 5336 44544 5438 44572
rect 6540 44068 6568 44096
rect 5357 43912 5434 43940
rect 5357 43268 5385 43912
rect 6540 43842 6568 43870
rect 5410 43766 5612 43794
rect 5410 43268 5438 43766
rect 6540 43716 6568 43744
rect 5336 43240 5438 43268
rect 5501 43646 5914 43674
rect 5357 43122 5385 43240
rect 5336 43094 5385 43122
rect 5501 43000 5529 43646
rect 5336 42972 5529 43000
rect 5501 42454 5914 42482
rect 5501 42362 5529 42454
rect 6540 42384 6568 42412
rect 5410 42334 5612 42362
rect 5410 42216 5438 42334
rect 5357 42188 5438 42216
rect 5357 41812 5385 42188
rect 5410 41812 5438 42188
rect 5501 41812 5529 42334
rect 6540 42258 6568 42286
rect 6540 42032 6568 42060
rect 5336 41784 5529 41812
rect 5357 41690 5385 41784
rect 5336 41662 5385 41690
rect 5410 41544 5438 41784
rect 5336 41516 5438 41544
rect 6540 40992 6568 41020
rect 5357 40836 5434 40864
rect 5357 40240 5385 40836
rect 6540 40766 6568 40794
rect 5410 40690 5612 40718
rect 5410 40240 5438 40690
rect 6540 40640 6568 40668
rect 5336 40212 5438 40240
rect 5501 40570 5914 40598
rect 5357 40094 5385 40212
rect 5336 40066 5385 40094
rect 5501 39972 5529 40570
rect 5336 39944 5529 39972
rect 5501 39378 5914 39406
rect 5501 39286 5529 39378
rect 6540 39308 6568 39336
rect 5410 39258 5612 39286
rect 5410 39140 5438 39258
rect 5357 39112 5438 39140
rect 5357 38784 5385 39112
rect 5410 38784 5438 39112
rect 5501 38784 5529 39258
rect 6540 39182 6568 39210
rect 6540 38956 6568 38984
rect 5336 38756 5529 38784
rect 5357 38662 5385 38756
rect 5336 38634 5385 38662
rect 5410 38516 5438 38756
rect 5336 38488 5438 38516
rect 6540 37916 6568 37944
rect 5357 37760 5434 37788
rect 5357 37212 5385 37760
rect 6540 37690 6568 37718
rect 5410 37614 5612 37642
rect 5410 37212 5438 37614
rect 6540 37564 6568 37592
rect 5336 37184 5438 37212
rect 5501 37494 5914 37522
rect 5357 37066 5385 37184
rect 5336 37038 5385 37066
rect 5501 36944 5529 37494
rect 5336 36916 5529 36944
rect 5501 36302 5914 36330
rect 5501 36210 5529 36302
rect 6540 36232 6568 36260
rect 5410 36182 5612 36210
rect 5410 36064 5438 36182
rect 5357 36036 5438 36064
rect 5357 35756 5385 36036
rect 5410 35756 5438 36036
rect 5501 35756 5529 36182
rect 6540 36106 6568 36134
rect 6540 35880 6568 35908
rect 5336 35728 5529 35756
rect 5357 35634 5385 35728
rect 5336 35606 5385 35634
rect 5410 35488 5438 35728
rect 5336 35460 5438 35488
rect 6540 34840 6568 34868
rect 5357 34684 5434 34712
rect 5357 34184 5385 34684
rect 6540 34614 6568 34642
rect 5410 34538 5612 34566
rect 5410 34184 5438 34538
rect 6540 34488 6568 34516
rect 5336 34156 5438 34184
rect 5501 34418 5914 34446
rect 5357 34038 5385 34156
rect 5336 34010 5385 34038
rect 5501 33916 5529 34418
rect 5336 33888 5529 33916
rect 5501 33226 5914 33254
rect 5501 33134 5529 33226
rect 6540 33156 6568 33184
rect 5410 33106 5612 33134
rect 5410 32988 5438 33106
rect 5357 32960 5438 32988
rect 5357 32728 5385 32960
rect 5410 32728 5438 32960
rect 5501 32728 5529 33106
rect 6540 33030 6568 33058
rect 6540 32804 6568 32832
rect 5336 32700 5529 32728
rect 5357 32606 5385 32700
rect 5336 32578 5385 32606
rect 5410 32460 5438 32700
rect 5336 32432 5438 32460
rect 6540 31764 6568 31792
rect 5357 31608 5434 31636
rect 5357 31156 5385 31608
rect 6540 31538 6568 31566
rect 5410 31462 5612 31490
rect 5410 31156 5438 31462
rect 6540 31412 6568 31440
rect 5336 31128 5438 31156
rect 5501 31342 5914 31370
rect 5357 31010 5385 31128
rect 5336 30982 5385 31010
rect 5501 30888 5529 31342
rect 5336 30860 5529 30888
rect 5501 30150 5914 30178
rect 5501 30058 5529 30150
rect 6540 30080 6568 30108
rect 5410 30030 5612 30058
rect 5410 29912 5438 30030
rect 5357 29884 5438 29912
rect 5357 29700 5385 29884
rect 5410 29700 5438 29884
rect 5501 29700 5529 30030
rect 6540 29954 6568 29982
rect 6540 29728 6568 29756
rect 5336 29672 5529 29700
rect 5357 29578 5385 29672
rect 5336 29550 5385 29578
rect 5410 29432 5438 29672
rect 5336 29404 5438 29432
rect 6540 28688 6568 28716
rect 5357 28532 5434 28560
rect 5357 28128 5385 28532
rect 6540 28462 6568 28490
rect 5410 28386 5612 28414
rect 5410 28128 5438 28386
rect 6540 28336 6568 28364
rect 5336 28100 5438 28128
rect 5501 28266 5914 28294
rect 5357 27982 5385 28100
rect 5336 27954 5385 27982
rect 5501 27860 5529 28266
rect 5336 27832 5529 27860
rect 5501 27074 5914 27102
rect 5501 26982 5529 27074
rect 6540 27004 6568 27032
rect 5410 26954 5612 26982
rect 5410 26836 5438 26954
rect 5357 26808 5438 26836
rect 5357 26672 5385 26808
rect 5410 26672 5438 26808
rect 5501 26672 5529 26954
rect 6540 26878 6568 26906
rect 5336 26644 5529 26672
rect 6540 26652 6568 26680
rect 5357 26550 5385 26644
rect 5336 26522 5385 26550
rect 5410 26404 5438 26644
rect 5336 26376 5438 26404
rect 6540 25612 6568 25640
rect 5357 25456 5434 25484
rect 5357 25100 5385 25456
rect 6540 25386 6568 25414
rect 5410 25310 5612 25338
rect 5410 25100 5438 25310
rect 6540 25260 6568 25288
rect 5336 25072 5438 25100
rect 5501 25190 5914 25218
rect 5357 24954 5385 25072
rect 5336 24926 5385 24954
rect 5501 24832 5529 25190
rect 5336 24804 5529 24832
rect 5501 23998 5914 24026
rect 5501 23906 5529 23998
rect 6540 23928 6568 23956
rect 5410 23878 5612 23906
rect 5410 23760 5438 23878
rect 5357 23732 5438 23760
rect 5357 23644 5385 23732
rect 5410 23644 5438 23732
rect 5501 23644 5529 23878
rect 6540 23802 6568 23830
rect 5336 23616 5529 23644
rect 5357 23522 5385 23616
rect 5336 23494 5385 23522
rect 5410 23376 5438 23616
rect 6540 23576 6568 23604
rect 5336 23348 5438 23376
rect 6540 22536 6568 22564
rect 5357 22380 5434 22408
rect 5357 22072 5385 22380
rect 6540 22310 6568 22338
rect 5410 22234 5612 22262
rect 5410 22072 5438 22234
rect 6540 22184 6568 22212
rect 5336 22044 5438 22072
rect 5501 22114 5914 22142
rect 5357 21926 5385 22044
rect 5336 21898 5385 21926
rect 5501 21804 5529 22114
rect 5336 21776 5529 21804
rect 5501 20922 5914 20950
rect 5501 20830 5529 20922
rect 6540 20852 6568 20880
rect 5410 20802 5612 20830
rect 5410 20684 5438 20802
rect 5357 20656 5438 20684
rect 5357 20616 5385 20656
rect 5410 20616 5438 20656
rect 5501 20616 5529 20802
rect 6540 20726 6568 20754
rect 5336 20588 5529 20616
rect 5357 20494 5385 20588
rect 5336 20466 5385 20494
rect 5410 20348 5438 20588
rect 6540 20500 6568 20528
rect 5336 20320 5438 20348
rect 6540 19460 6568 19488
rect 5357 19304 5434 19332
rect 5357 19044 5385 19304
rect 6540 19234 6568 19262
rect 5410 19158 5612 19186
rect 5410 19044 5438 19158
rect 6540 19108 6568 19136
rect 5336 19016 5438 19044
rect 5501 19038 5914 19066
rect 5357 18898 5385 19016
rect 5336 18870 5385 18898
rect 5501 18776 5529 19038
rect 5336 18748 5529 18776
rect 5501 17846 5914 17874
rect 5501 17754 5529 17846
rect 6540 17776 6568 17804
rect 5410 17726 5612 17754
rect 5410 17608 5438 17726
rect 5357 17588 5438 17608
rect 5501 17588 5529 17726
rect 6540 17650 6568 17678
rect 5336 17560 5529 17588
rect 5357 17466 5385 17560
rect 5336 17438 5385 17466
rect 5410 17320 5438 17560
rect 6540 17424 6568 17452
rect 5336 17292 5438 17320
rect 6540 16384 6568 16412
rect 5357 16228 5434 16256
rect 5357 16016 5385 16228
rect 6540 16158 6568 16186
rect 5410 16082 5612 16110
rect 5410 16016 5438 16082
rect 6540 16032 6568 16060
rect 5336 15988 5438 16016
rect 5357 15870 5385 15988
rect 5336 15842 5385 15870
rect 5501 15962 5914 15990
rect 5501 15748 5529 15962
rect 5336 15720 5529 15748
rect 5501 14770 5914 14798
rect 5501 14678 5529 14770
rect 6540 14700 6568 14728
rect 5410 14650 5612 14678
rect 5410 14560 5438 14650
rect 5501 14560 5529 14650
rect 6540 14574 6568 14602
rect 5336 14532 5529 14560
rect 5357 14504 5438 14532
rect 5357 14438 5385 14504
rect 5336 14410 5385 14438
rect 5410 14292 5438 14504
rect 6540 14348 6568 14376
rect 5336 14264 5438 14292
rect 6540 13308 6568 13336
rect 5357 13152 5434 13180
rect 5357 12988 5385 13152
rect 6540 13082 6568 13110
rect 5410 13006 5612 13034
rect 5410 12988 5438 13006
rect 5336 12960 5438 12988
rect 5357 12842 5385 12960
rect 6540 12956 6568 12984
rect 5336 12814 5385 12842
rect 5501 12886 5914 12914
rect 5501 12720 5529 12886
rect 5336 12692 5529 12720
rect 5501 11694 5914 11722
rect 5501 11602 5529 11694
rect 6540 11624 6568 11652
rect 5410 11574 5612 11602
rect 5410 11532 5438 11574
rect 5501 11532 5529 11574
rect 5336 11504 5529 11532
rect 5410 11456 5438 11504
rect 6540 11498 6568 11526
rect 5357 11428 5438 11456
rect 5357 11410 5385 11428
rect 5336 11382 5385 11410
rect 5410 11264 5438 11428
rect 6540 11272 6568 11300
rect 5336 11236 5438 11264
rect 6540 10232 6568 10260
rect 5357 10076 5434 10104
rect 5357 9960 5385 10076
rect 6540 10006 6568 10034
rect 5336 9958 5438 9960
rect 5336 9932 5612 9958
rect 5357 9814 5385 9932
rect 5410 9930 5612 9932
rect 6540 9880 6568 9908
rect 5336 9786 5385 9814
rect 5501 9810 5914 9838
rect 5501 9692 5529 9810
rect 5336 9664 5529 9692
rect 5501 8618 5914 8646
rect 5501 8526 5529 8618
rect 6540 8548 6568 8576
rect 5410 8504 5612 8526
rect 5336 8498 5612 8504
rect 5336 8476 5529 8498
rect 5336 8380 5385 8382
rect 5410 8380 5438 8476
rect 6540 8422 6568 8450
rect 5336 8354 5438 8380
rect 5357 8352 5438 8354
rect 5410 8236 5438 8352
rect 5336 8208 5438 8236
rect 6540 8196 6568 8224
rect 6540 7156 6568 7184
rect 5357 7000 5434 7028
rect 5357 6932 5385 7000
rect 5336 6904 5438 6932
rect 6540 6930 6568 6958
rect 5357 6786 5385 6904
rect 5410 6882 5438 6904
rect 5410 6854 5612 6882
rect 6540 6804 6568 6832
rect 5336 6758 5385 6786
rect 5501 6734 5914 6762
rect 5501 6664 5529 6734
rect 5336 6636 5529 6664
rect 5501 5542 5914 5570
rect 5501 5476 5529 5542
rect 5336 5450 5529 5476
rect 6540 5472 6568 5500
rect 5336 5448 5612 5450
rect 5410 5422 5612 5448
rect 5336 5326 5385 5354
rect 5357 5304 5385 5326
rect 5410 5304 5438 5422
rect 6540 5346 6568 5374
rect 5357 5276 5438 5304
rect 5410 5208 5438 5276
rect 5336 5180 5438 5208
rect 6540 5120 6568 5148
rect 6540 4080 6568 4108
rect 5357 3924 5434 3952
rect 5357 3904 5385 3924
rect 5336 3876 5438 3904
rect 5357 3758 5385 3876
rect 5410 3806 5438 3876
rect 6540 3854 6568 3882
rect 5410 3778 5612 3806
rect 5336 3730 5385 3758
rect 6540 3728 6568 3756
rect 5501 3658 5914 3686
rect 5501 3636 5529 3658
rect 5336 3608 5529 3636
rect 5501 2466 5914 2494
rect 5501 2448 5529 2466
rect 5336 2420 5529 2448
rect 6540 2396 6568 2424
rect 5410 2346 5612 2374
rect 5336 2298 5385 2326
rect 5357 2228 5385 2298
rect 5410 2228 5438 2346
rect 6540 2270 6568 2298
rect 5357 2200 5438 2228
rect 5410 2180 5438 2200
rect 5336 2152 5438 2180
rect 6540 2044 6568 2072
rect 6540 1004 6568 1032
rect 5336 848 5438 876
rect 5357 730 5385 848
rect 5336 702 5385 730
rect 5410 730 5438 848
rect 6540 778 6568 806
rect 5410 702 5612 730
rect 6540 652 6568 680
rect 5501 608 5914 610
rect 5336 582 5914 608
rect 5336 580 5529 582
<< metal2 >>
rect 5178 49202 5392 49230
rect 1 0 29 30792
rect 69 0 97 30792
rect 137 0 165 30792
rect 205 0 233 30792
rect 273 0 301 30792
rect 341 0 369 30792
rect 409 0 437 30792
<< metal3 >>
rect 6502 49183 6634 49249
rect 5298 48415 5430 48481
rect 6502 47645 6634 47711
rect 5298 46901 5430 46967
rect 6502 46107 6634 46173
rect 5298 45387 5430 45453
rect 6502 44569 6634 44635
rect 5298 43873 5430 43939
rect 6502 43031 6634 43097
rect 5298 42359 5430 42425
rect 6502 41493 6634 41559
rect 5298 40845 5430 40911
rect 6502 39955 6634 40021
rect 5298 39331 5430 39397
rect 6502 38417 6634 38483
rect 5298 37817 5430 37883
rect 6502 36879 6634 36945
rect 5298 36303 5430 36369
rect 6502 35341 6634 35407
rect 5298 34789 5430 34855
rect 6502 33803 6634 33869
rect 5298 33275 5430 33341
rect 6502 32265 6634 32331
rect 5298 31761 5430 31827
rect 751 30759 883 30825
rect 1646 30759 1778 30825
rect 6502 30727 6634 30793
rect 5298 30247 5430 30313
rect 751 29219 883 29285
rect 1646 29219 1778 29285
rect 6502 29189 6634 29255
rect 5298 28733 5430 28799
rect 751 27679 883 27745
rect 1646 27679 1778 27745
rect 6502 27651 6634 27717
rect 5298 27219 5430 27285
rect 751 26139 883 26205
rect 1646 26139 1778 26205
rect 6502 26113 6634 26179
rect 5298 25705 5430 25771
rect 751 24599 883 24665
rect 1646 24599 1778 24665
rect 6502 24575 6634 24641
rect 5298 24191 5430 24257
rect 751 23059 883 23125
rect 1646 23059 1778 23125
rect 6502 23037 6634 23103
rect 5298 22677 5430 22743
rect 751 21519 883 21585
rect 1646 21519 1778 21585
rect 6502 21499 6634 21565
rect 5298 21163 5430 21229
rect 751 19979 883 20045
rect 1646 19979 1778 20045
rect 6502 19961 6634 20027
rect 5298 19649 5430 19715
rect 751 18439 883 18505
rect 1646 18439 1778 18505
rect 6502 18423 6634 18489
rect 5298 18135 5430 18201
rect 6502 16885 6634 16951
rect 5298 16621 5430 16687
rect 1045 15363 1177 15429
rect 1804 15363 1936 15429
rect 6502 15347 6634 15413
rect 5298 15107 5430 15173
rect 1045 13823 1177 13889
rect 1804 13823 1936 13889
rect 6502 13809 6634 13875
rect 5298 13593 5430 13659
rect 1045 12283 1177 12349
rect 1804 12283 1936 12349
rect 6502 12271 6634 12337
rect 5298 12079 5430 12145
rect 1045 10743 1177 10809
rect 1804 10743 1936 10809
rect 6502 10733 6634 10799
rect 5298 10565 5430 10631
rect 1045 9203 1177 9269
rect 1804 9203 1936 9269
rect 6502 9195 6634 9261
rect 5298 9051 5430 9117
rect 6502 7657 6634 7723
rect 5298 7537 5430 7603
rect 1045 6127 1177 6193
rect 1804 6127 1936 6193
rect 6502 6119 6634 6185
rect 5298 6023 5430 6089
rect 1045 4587 1177 4653
rect 1804 4587 1936 4653
rect 6502 4581 6634 4647
rect 5298 4509 5430 4575
rect 1045 3047 1177 3113
rect 1804 3047 1936 3113
rect 5298 2995 5430 3061
rect 6502 3043 6634 3109
rect 1045 1507 1177 1573
rect 1804 1507 1936 1573
rect 5298 1481 5430 1547
rect 6502 1505 6634 1571
rect 1045 -33 1177 33
rect 1804 -33 1936 33
rect 5298 -33 5430 33
rect 6502 -33 6634 33
use wordline_driver_array  wordline_driver_array_0
timestamp 1643678851
transform 1 0 5364 0 1 0
box 0 -42 1270 49258
use hierarchical_decoder  hierarchical_decoder_0
timestamp 1643678851
transform 1 0 0 0 1 0
box -11 -42 5430 49244
<< labels >>
rlabel metal2 s 1 0 29 30792 4 addr0
rlabel metal2 s 69 0 97 30792 4 addr1
rlabel metal2 s 137 0 165 30792 4 addr2
rlabel metal2 s 205 0 233 30792 4 addr3
rlabel metal2 s 273 0 301 30792 4 addr4
rlabel metal2 s 341 0 369 30792 4 addr5
rlabel metal2 s 409 0 437 30792 4 addr6
rlabel metal1 s 6540 778 6568 806 4 rwl0_0
rlabel metal1 s 6540 1004 6568 1032 4 rwl1_0
rlabel metal1 s 6540 652 6568 680 4 wwl0_0
rlabel metal1 s 6540 2270 6568 2298 4 rwl0_1
rlabel metal1 s 6540 2044 6568 2072 4 rwl1_1
rlabel metal1 s 6540 2396 6568 2424 4 wwl0_1
rlabel metal1 s 6540 3854 6568 3882 4 rwl0_2
rlabel metal1 s 6540 4080 6568 4108 4 rwl1_2
rlabel metal1 s 6540 3728 6568 3756 4 wwl0_2
rlabel metal1 s 6540 5346 6568 5374 4 rwl0_3
rlabel metal1 s 6540 5120 6568 5148 4 rwl1_3
rlabel metal1 s 6540 5472 6568 5500 4 wwl0_3
rlabel metal1 s 6540 6930 6568 6958 4 rwl0_4
rlabel metal1 s 6540 7156 6568 7184 4 rwl1_4
rlabel metal1 s 6540 6804 6568 6832 4 wwl0_4
rlabel metal1 s 6540 8422 6568 8450 4 rwl0_5
rlabel metal1 s 6540 8196 6568 8224 4 rwl1_5
rlabel metal1 s 6540 8548 6568 8576 4 wwl0_5
rlabel metal1 s 6540 10006 6568 10034 4 rwl0_6
rlabel metal1 s 6540 10232 6568 10260 4 rwl1_6
rlabel metal1 s 6540 9880 6568 9908 4 wwl0_6
rlabel metal1 s 6540 11498 6568 11526 4 rwl0_7
rlabel metal1 s 6540 11272 6568 11300 4 rwl1_7
rlabel metal1 s 6540 11624 6568 11652 4 wwl0_7
rlabel metal1 s 6540 13082 6568 13110 4 rwl0_8
rlabel metal1 s 6540 13308 6568 13336 4 rwl1_8
rlabel metal1 s 6540 12956 6568 12984 4 wwl0_8
rlabel metal1 s 6540 14574 6568 14602 4 rwl0_9
rlabel metal1 s 6540 14348 6568 14376 4 rwl1_9
rlabel metal1 s 6540 14700 6568 14728 4 wwl0_9
rlabel metal1 s 6540 16158 6568 16186 4 rwl0_10
rlabel metal1 s 6540 16384 6568 16412 4 rwl1_10
rlabel metal1 s 6540 16032 6568 16060 4 wwl0_10
rlabel metal1 s 6540 17650 6568 17678 4 rwl0_11
rlabel metal1 s 6540 17424 6568 17452 4 rwl1_11
rlabel metal1 s 6540 17776 6568 17804 4 wwl0_11
rlabel metal1 s 6540 19234 6568 19262 4 rwl0_12
rlabel metal1 s 6540 19460 6568 19488 4 rwl1_12
rlabel metal1 s 6540 19108 6568 19136 4 wwl0_12
rlabel metal1 s 6540 20726 6568 20754 4 rwl0_13
rlabel metal1 s 6540 20500 6568 20528 4 rwl1_13
rlabel metal1 s 6540 20852 6568 20880 4 wwl0_13
rlabel metal1 s 6540 22310 6568 22338 4 rwl0_14
rlabel metal1 s 6540 22536 6568 22564 4 rwl1_14
rlabel metal1 s 6540 22184 6568 22212 4 wwl0_14
rlabel metal1 s 6540 23802 6568 23830 4 rwl0_15
rlabel metal1 s 6540 23576 6568 23604 4 rwl1_15
rlabel metal1 s 6540 23928 6568 23956 4 wwl0_15
rlabel metal1 s 6540 25386 6568 25414 4 rwl0_16
rlabel metal1 s 6540 25612 6568 25640 4 rwl1_16
rlabel metal1 s 6540 25260 6568 25288 4 wwl0_16
rlabel metal1 s 6540 26878 6568 26906 4 rwl0_17
rlabel metal1 s 6540 26652 6568 26680 4 rwl1_17
rlabel metal1 s 6540 27004 6568 27032 4 wwl0_17
rlabel metal1 s 6540 28462 6568 28490 4 rwl0_18
rlabel metal1 s 6540 28688 6568 28716 4 rwl1_18
rlabel metal1 s 6540 28336 6568 28364 4 wwl0_18
rlabel metal1 s 6540 29954 6568 29982 4 rwl0_19
rlabel metal1 s 6540 29728 6568 29756 4 rwl1_19
rlabel metal1 s 6540 30080 6568 30108 4 wwl0_19
rlabel metal1 s 6540 31538 6568 31566 4 rwl0_20
rlabel metal1 s 6540 31764 6568 31792 4 rwl1_20
rlabel metal1 s 6540 31412 6568 31440 4 wwl0_20
rlabel metal1 s 6540 33030 6568 33058 4 rwl0_21
rlabel metal1 s 6540 32804 6568 32832 4 rwl1_21
rlabel metal1 s 6540 33156 6568 33184 4 wwl0_21
rlabel metal1 s 6540 34614 6568 34642 4 rwl0_22
rlabel metal1 s 6540 34840 6568 34868 4 rwl1_22
rlabel metal1 s 6540 34488 6568 34516 4 wwl0_22
rlabel metal1 s 6540 36106 6568 36134 4 rwl0_23
rlabel metal1 s 6540 35880 6568 35908 4 rwl1_23
rlabel metal1 s 6540 36232 6568 36260 4 wwl0_23
rlabel metal1 s 6540 37690 6568 37718 4 rwl0_24
rlabel metal1 s 6540 37916 6568 37944 4 rwl1_24
rlabel metal1 s 6540 37564 6568 37592 4 wwl0_24
rlabel metal1 s 6540 39182 6568 39210 4 rwl0_25
rlabel metal1 s 6540 38956 6568 38984 4 rwl1_25
rlabel metal1 s 6540 39308 6568 39336 4 wwl0_25
rlabel metal1 s 6540 40766 6568 40794 4 rwl0_26
rlabel metal1 s 6540 40992 6568 41020 4 rwl1_26
rlabel metal1 s 6540 40640 6568 40668 4 wwl0_26
rlabel metal1 s 6540 42258 6568 42286 4 rwl0_27
rlabel metal1 s 6540 42032 6568 42060 4 rwl1_27
rlabel metal1 s 6540 42384 6568 42412 4 wwl0_27
rlabel metal1 s 6540 43842 6568 43870 4 rwl0_28
rlabel metal1 s 6540 44068 6568 44096 4 rwl1_28
rlabel metal1 s 6540 43716 6568 43744 4 wwl0_28
rlabel metal1 s 6540 45334 6568 45362 4 rwl0_29
rlabel metal1 s 6540 45108 6568 45136 4 rwl1_29
rlabel metal1 s 6540 45460 6568 45488 4 wwl0_29
rlabel metal1 s 6540 46918 6568 46946 4 rwl0_30
rlabel metal1 s 6540 47144 6568 47172 4 rwl1_30
rlabel metal1 s 6540 46792 6568 46820 4 wwl0_30
rlabel metal1 s 6540 48410 6568 48438 4 rwl0_31
rlabel metal1 s 6540 48184 6568 48212 4 rwl1_31
rlabel metal1 s 6540 48536 6568 48564 4 wwl0_31
rlabel metal2 s 5364 49202 5392 49230 4 wl_en
rlabel metal3 s 5298 1481 5430 1547 4 vdd
rlabel metal3 s 6502 1505 6634 1571 4 vdd
rlabel metal3 s 6502 41493 6634 41559 4 vdd
rlabel metal3 s 6502 32265 6634 32331 4 vdd
rlabel metal3 s 6502 7657 6634 7723 4 vdd
rlabel metal3 s 5298 16621 5430 16687 4 vdd
rlabel metal3 s 1804 4587 1936 4653 4 vdd
rlabel metal3 s 751 29219 883 29285 4 vdd
rlabel metal3 s 5298 40845 5430 40911 4 vdd
rlabel metal3 s 6502 4581 6634 4647 4 vdd
rlabel metal3 s 1646 19979 1778 20045 4 vdd
rlabel metal3 s 6502 38417 6634 38483 4 vdd
rlabel metal3 s 6502 35341 6634 35407 4 vdd
rlabel metal3 s 5298 43873 5430 43939 4 vdd
rlabel metal3 s 5298 4509 5430 4575 4 vdd
rlabel metal3 s 5298 28733 5430 28799 4 vdd
rlabel metal3 s 6502 10733 6634 10799 4 vdd
rlabel metal3 s 5298 31761 5430 31827 4 vdd
rlabel metal3 s 1045 13823 1177 13889 4 vdd
rlabel metal3 s 6502 13809 6634 13875 4 vdd
rlabel metal3 s 751 26139 883 26205 4 vdd
rlabel metal3 s 5298 25705 5430 25771 4 vdd
rlabel metal3 s 6502 23037 6634 23103 4 vdd
rlabel metal3 s 1045 10743 1177 10809 4 vdd
rlabel metal3 s 5298 37817 5430 37883 4 vdd
rlabel metal3 s 1646 26139 1778 26205 4 vdd
rlabel metal3 s 6502 19961 6634 20027 4 vdd
rlabel metal3 s 751 19979 883 20045 4 vdd
rlabel metal3 s 5298 46901 5430 46967 4 vdd
rlabel metal3 s 1646 23059 1778 23125 4 vdd
rlabel metal3 s 1804 13823 1936 13889 4 vdd
rlabel metal3 s 5298 10565 5430 10631 4 vdd
rlabel metal3 s 5298 19649 5430 19715 4 vdd
rlabel metal3 s 6502 47645 6634 47711 4 vdd
rlabel metal3 s 6502 44569 6634 44635 4 vdd
rlabel metal3 s 6502 16885 6634 16951 4 vdd
rlabel metal3 s 1045 4587 1177 4653 4 vdd
rlabel metal3 s 5298 22677 5430 22743 4 vdd
rlabel metal3 s 1804 10743 1936 10809 4 vdd
rlabel metal3 s 1646 29219 1778 29285 4 vdd
rlabel metal3 s 5298 7537 5430 7603 4 vdd
rlabel metal3 s 6502 29189 6634 29255 4 vdd
rlabel metal3 s 5298 13593 5430 13659 4 vdd
rlabel metal3 s 1045 1507 1177 1573 4 vdd
rlabel metal3 s 1804 1507 1936 1573 4 vdd
rlabel metal3 s 6502 26113 6634 26179 4 vdd
rlabel metal3 s 5298 34789 5430 34855 4 vdd
rlabel metal3 s 751 23059 883 23125 4 vdd
rlabel metal3 s 6502 6119 6634 6185 4 gnd
rlabel metal3 s 6502 3043 6634 3109 4 gnd
rlabel metal3 s 5298 48415 5430 48481 4 gnd
rlabel metal3 s 5298 -33 5430 33 4 gnd
rlabel metal3 s 1646 27679 1778 27745 4 gnd
rlabel metal3 s 6502 24575 6634 24641 4 gnd
rlabel metal3 s 1045 3047 1177 3113 4 gnd
rlabel metal3 s 1804 15363 1936 15429 4 gnd
rlabel metal3 s 5298 24191 5430 24257 4 gnd
rlabel metal3 s 1646 21519 1778 21585 4 gnd
rlabel metal3 s 751 24599 883 24665 4 gnd
rlabel metal3 s 5298 6023 5430 6089 4 gnd
rlabel metal3 s 5298 12079 5430 12145 4 gnd
rlabel metal3 s 6502 21499 6634 21565 4 gnd
rlabel metal3 s 1646 24599 1778 24665 4 gnd
rlabel metal3 s 5298 9051 5430 9117 4 gnd
rlabel metal3 s 5298 18135 5430 18201 4 gnd
rlabel metal3 s 5298 27219 5430 27285 4 gnd
rlabel metal3 s 751 27679 883 27745 4 gnd
rlabel metal3 s 5298 33275 5430 33341 4 gnd
rlabel metal3 s 751 18439 883 18505 4 gnd
rlabel metal3 s 5298 2995 5430 3061 4 gnd
rlabel metal3 s 6502 46107 6634 46173 4 gnd
rlabel metal3 s 6502 39955 6634 40021 4 gnd
rlabel metal3 s 6502 27651 6634 27717 4 gnd
rlabel metal3 s 1045 -33 1177 33 4 gnd
rlabel metal3 s 1045 6127 1177 6193 4 gnd
rlabel metal3 s 5298 21163 5430 21229 4 gnd
rlabel metal3 s 6502 12271 6634 12337 4 gnd
rlabel metal3 s 5298 36303 5430 36369 4 gnd
rlabel metal3 s 1045 9203 1177 9269 4 gnd
rlabel metal3 s 1804 3047 1936 3113 4 gnd
rlabel metal3 s 6502 33803 6634 33869 4 gnd
rlabel metal3 s 1045 12283 1177 12349 4 gnd
rlabel metal3 s 6502 9195 6634 9261 4 gnd
rlabel metal3 s 5298 42359 5430 42425 4 gnd
rlabel metal3 s 1646 18439 1778 18505 4 gnd
rlabel metal3 s 5298 30247 5430 30313 4 gnd
rlabel metal3 s 6502 36879 6634 36945 4 gnd
rlabel metal3 s 751 21519 883 21585 4 gnd
rlabel metal3 s 6502 30727 6634 30793 4 gnd
rlabel metal3 s 5298 45387 5430 45453 4 gnd
rlabel metal3 s 5298 39331 5430 39397 4 gnd
rlabel metal3 s 1045 15363 1177 15429 4 gnd
rlabel metal3 s 1646 30759 1778 30825 4 gnd
rlabel metal3 s 1804 12283 1936 12349 4 gnd
rlabel metal3 s 1804 9203 1936 9269 4 gnd
rlabel metal3 s 1804 -33 1936 33 4 gnd
rlabel metal3 s 6502 15347 6634 15413 4 gnd
rlabel metal3 s 5298 15107 5430 15173 4 gnd
rlabel metal3 s 6502 18423 6634 18489 4 gnd
rlabel metal3 s 6502 -33 6634 33 4 gnd
rlabel metal3 s 6502 43031 6634 43097 4 gnd
rlabel metal3 s 6502 49183 6634 49249 4 gnd
rlabel metal3 s 1804 6127 1936 6193 4 gnd
rlabel metal3 s 751 30759 883 30825 4 gnd
<< properties >>
string FIXED_BBOX 0 0 6604 49244
string GDS_FILE sram_0rw2r1w_16_128_sky130A.gds
string GDS_END 1711092
string GDS_START 1628758
<< end >>
