magic
tech sky130A
timestamp 1642355658
<< nwell >>
rect 0 218 741 458
<< nmos >>
rect 54 48 69 90
rect 110 48 125 90
rect 166 48 181 90
rect 222 48 237 90
rect 278 48 293 90
rect 334 48 349 90
rect 390 48 405 90
rect 446 48 461 90
rect 502 48 517 90
rect 558 48 573 90
rect 672 48 687 90
<< pmos >>
rect 54 236 69 371
rect 110 236 125 371
rect 166 236 181 371
rect 222 236 237 371
rect 278 236 293 371
rect 334 236 349 371
rect 390 236 405 371
rect 446 236 461 371
rect 502 236 517 371
rect 558 236 573 371
rect 672 236 687 371
<< ndiff >>
rect 18 77 54 90
rect 18 60 25 77
rect 42 60 54 77
rect 18 48 54 60
rect 69 77 110 90
rect 69 60 81 77
rect 98 60 110 77
rect 69 48 110 60
rect 125 77 166 90
rect 125 60 137 77
rect 154 60 166 77
rect 125 48 166 60
rect 181 77 222 90
rect 181 60 193 77
rect 210 60 222 77
rect 181 48 222 60
rect 237 48 278 90
rect 293 77 334 90
rect 293 60 305 77
rect 322 60 334 77
rect 293 48 334 60
rect 349 77 390 90
rect 349 60 361 77
rect 378 60 390 77
rect 349 48 390 60
rect 405 77 446 90
rect 405 60 417 77
rect 434 60 446 77
rect 405 48 446 60
rect 461 48 502 90
rect 517 77 558 90
rect 517 60 529 77
rect 546 60 558 77
rect 517 48 558 60
rect 573 77 609 90
rect 573 60 585 77
rect 602 60 609 77
rect 573 48 609 60
rect 636 77 672 90
rect 636 60 643 77
rect 660 60 672 77
rect 636 48 672 60
rect 687 77 723 90
rect 687 60 699 77
rect 716 60 723 77
rect 687 48 723 60
<< pdiff >>
rect 18 350 54 371
rect 18 333 25 350
rect 42 333 54 350
rect 18 312 54 333
rect 18 295 25 312
rect 42 295 54 312
rect 18 274 54 295
rect 18 257 25 274
rect 42 257 54 274
rect 18 236 54 257
rect 69 350 110 371
rect 69 333 81 350
rect 98 333 110 350
rect 69 312 110 333
rect 69 295 81 312
rect 98 295 110 312
rect 69 274 110 295
rect 69 257 81 274
rect 98 257 110 274
rect 69 236 110 257
rect 125 350 166 371
rect 125 333 137 350
rect 154 333 166 350
rect 125 312 166 333
rect 125 295 137 312
rect 154 295 166 312
rect 125 274 166 295
rect 125 257 137 274
rect 154 257 166 274
rect 125 236 166 257
rect 181 350 222 371
rect 181 333 193 350
rect 210 333 222 350
rect 181 312 222 333
rect 181 295 193 312
rect 210 295 222 312
rect 181 274 222 295
rect 181 257 193 274
rect 210 257 222 274
rect 181 236 222 257
rect 237 236 278 371
rect 293 350 334 371
rect 293 333 305 350
rect 322 333 334 350
rect 293 312 334 333
rect 293 295 305 312
rect 322 295 334 312
rect 293 274 334 295
rect 293 257 305 274
rect 322 257 334 274
rect 293 236 334 257
rect 349 350 390 371
rect 349 333 361 350
rect 378 333 390 350
rect 349 312 390 333
rect 349 295 361 312
rect 378 295 390 312
rect 349 274 390 295
rect 349 257 361 274
rect 378 257 390 274
rect 349 236 390 257
rect 405 350 446 371
rect 405 333 417 350
rect 434 333 446 350
rect 405 312 446 333
rect 405 295 417 312
rect 434 295 446 312
rect 405 274 446 295
rect 405 257 417 274
rect 434 257 446 274
rect 405 236 446 257
rect 461 236 502 371
rect 517 350 558 371
rect 517 333 529 350
rect 546 333 558 350
rect 517 312 558 333
rect 517 295 529 312
rect 546 295 558 312
rect 517 274 558 295
rect 517 257 529 274
rect 546 257 558 274
rect 517 236 558 257
rect 573 350 609 371
rect 573 333 585 350
rect 602 333 609 350
rect 573 312 609 333
rect 573 295 585 312
rect 602 295 609 312
rect 573 274 609 295
rect 573 257 585 274
rect 602 257 609 274
rect 573 236 609 257
rect 636 350 672 371
rect 636 333 643 350
rect 660 333 672 350
rect 636 312 672 333
rect 636 295 643 312
rect 660 295 672 312
rect 636 274 672 295
rect 636 257 643 274
rect 660 257 672 274
rect 636 236 672 257
rect 687 350 723 371
rect 687 333 699 350
rect 716 333 723 350
rect 687 312 723 333
rect 687 295 699 312
rect 716 295 723 312
rect 687 274 723 295
rect 687 257 699 274
rect 716 257 723 274
rect 687 236 723 257
<< ndiffc >>
rect 25 60 42 77
rect 81 60 98 77
rect 137 60 154 77
rect 193 60 210 77
rect 305 60 322 77
rect 361 60 378 77
rect 417 60 434 77
rect 529 60 546 77
rect 585 60 602 77
rect 643 60 660 77
rect 699 60 716 77
<< pdiffc >>
rect 25 333 42 350
rect 25 295 42 312
rect 25 257 42 274
rect 81 333 98 350
rect 81 295 98 312
rect 81 257 98 274
rect 137 333 154 350
rect 137 295 154 312
rect 137 257 154 274
rect 193 333 210 350
rect 193 295 210 312
rect 193 257 210 274
rect 305 333 322 350
rect 305 295 322 312
rect 305 257 322 274
rect 361 333 378 350
rect 361 295 378 312
rect 361 257 378 274
rect 417 333 434 350
rect 417 295 434 312
rect 417 257 434 274
rect 529 333 546 350
rect 529 295 546 312
rect 529 257 546 274
rect 585 333 602 350
rect 585 295 602 312
rect 585 257 602 274
rect 643 333 660 350
rect 643 295 660 312
rect 643 257 660 274
rect 699 333 716 350
rect 699 295 716 312
rect 699 257 716 274
<< psubdiff >>
rect 70 9 106 21
rect 70 -9 79 9
rect 97 -9 106 9
rect 70 -21 106 -9
rect 211 9 247 21
rect 211 -9 220 9
rect 238 -9 247 9
rect 211 -21 247 -9
rect 352 9 388 21
rect 352 -9 361 9
rect 379 -9 388 9
rect 352 -21 388 -9
rect 493 9 529 21
rect 493 -9 502 9
rect 520 -9 529 9
rect 493 -21 529 -9
rect 634 9 670 21
rect 634 -9 643 9
rect 661 -9 670 9
rect 634 -21 670 -9
<< nsubdiff >>
rect 70 428 106 440
rect 70 410 79 428
rect 97 410 106 428
rect 70 398 106 410
rect 211 428 247 440
rect 211 410 220 428
rect 238 410 247 428
rect 211 398 247 410
rect 352 428 388 440
rect 352 410 361 428
rect 379 410 388 428
rect 352 398 388 410
rect 493 428 529 440
rect 493 410 502 428
rect 520 410 529 428
rect 493 398 529 410
rect 634 428 670 440
rect 634 410 643 428
rect 661 410 670 428
rect 634 398 670 410
<< psubdiffcont >>
rect 79 -9 97 9
rect 220 -9 238 9
rect 361 -9 379 9
rect 502 -9 520 9
rect 643 -9 661 9
<< nsubdiffcont >>
rect 79 410 97 428
rect 220 410 238 428
rect 361 410 379 428
rect 502 410 520 428
rect 643 410 661 428
<< poly >>
rect 54 371 69 384
rect 110 371 125 384
rect 166 371 181 384
rect 222 371 237 384
rect 278 371 293 384
rect 334 371 349 384
rect 390 371 405 384
rect 446 371 461 384
rect 502 371 517 384
rect 558 371 573 384
rect 672 371 687 384
rect 54 185 69 236
rect 0 177 69 185
rect 0 160 5 177
rect 22 170 69 177
rect 22 160 27 170
rect 0 152 27 160
rect 54 90 69 170
rect 110 140 125 236
rect 166 219 181 236
rect 222 219 237 236
rect 278 219 293 236
rect 160 211 187 219
rect 160 194 165 211
rect 182 194 187 211
rect 160 186 187 194
rect 222 211 256 219
rect 222 194 234 211
rect 251 194 256 211
rect 222 186 256 194
rect 278 211 305 219
rect 278 194 283 211
rect 300 194 305 211
rect 278 186 305 194
rect 90 132 125 140
rect 90 115 95 132
rect 112 115 125 132
rect 90 107 125 115
rect 160 132 187 140
rect 160 115 165 132
rect 182 115 187 132
rect 160 107 187 115
rect 222 127 256 135
rect 222 110 234 127
rect 251 110 256 127
rect 110 90 125 107
rect 166 90 181 107
rect 222 102 256 110
rect 222 90 237 102
rect 278 90 293 186
rect 334 165 349 236
rect 390 219 405 236
rect 446 219 461 236
rect 502 219 517 236
rect 384 211 411 219
rect 384 194 389 211
rect 406 194 411 211
rect 384 186 411 194
rect 446 211 480 219
rect 446 194 458 211
rect 475 194 480 211
rect 446 186 480 194
rect 502 211 529 219
rect 502 194 507 211
rect 524 194 529 211
rect 502 186 529 194
rect 314 157 349 165
rect 314 140 319 157
rect 336 140 349 157
rect 314 132 349 140
rect 334 90 349 132
rect 384 132 411 140
rect 384 115 389 132
rect 406 115 411 132
rect 384 107 411 115
rect 446 127 480 135
rect 446 110 458 127
rect 475 110 480 127
rect 390 90 405 107
rect 446 102 480 110
rect 446 90 461 102
rect 502 90 517 186
rect 558 165 573 236
rect 672 219 687 236
rect 660 211 687 219
rect 660 194 665 211
rect 682 194 687 211
rect 660 186 687 194
rect 538 157 573 165
rect 538 140 543 157
rect 560 140 573 157
rect 538 132 573 140
rect 558 90 573 132
rect 672 90 687 186
rect 54 35 69 48
rect 110 35 125 48
rect 166 35 181 48
rect 222 35 237 48
rect 278 35 293 48
rect 334 35 349 48
rect 390 35 405 48
rect 446 35 461 48
rect 502 35 517 48
rect 558 35 573 48
rect 672 35 687 48
<< polycont >>
rect 5 160 22 177
rect 165 194 182 211
rect 234 194 251 211
rect 283 194 300 211
rect 95 115 112 132
rect 165 115 182 132
rect 234 110 251 127
rect 389 194 406 211
rect 458 194 475 211
rect 507 194 524 211
rect 319 140 336 157
rect 389 115 406 132
rect 458 110 475 127
rect 665 194 682 211
rect 543 140 560 157
<< locali >>
rect 79 428 97 436
rect 79 371 97 410
rect 220 428 238 436
rect 220 402 238 410
rect 361 428 379 436
rect 361 405 379 410
rect 312 388 379 405
rect 502 428 520 436
rect 502 402 520 410
rect 643 428 661 436
rect 312 371 329 388
rect 502 385 539 402
rect 522 371 539 385
rect 643 371 661 410
rect 18 350 49 371
rect 18 333 25 350
rect 42 333 49 350
rect 18 312 49 333
rect 18 295 25 312
rect 42 295 49 312
rect 18 274 49 295
rect 18 257 25 274
rect 42 257 49 274
rect 18 236 49 257
rect 74 350 105 371
rect 74 333 81 350
rect 98 333 105 350
rect 74 312 105 333
rect 74 295 81 312
rect 98 295 105 312
rect 74 274 105 295
rect 74 257 81 274
rect 98 257 105 274
rect 74 236 105 257
rect 130 350 161 371
rect 130 333 137 350
rect 154 333 161 350
rect 130 312 161 333
rect 130 295 137 312
rect 154 295 161 312
rect 130 274 161 295
rect 130 257 137 274
rect 154 257 161 274
rect 130 236 161 257
rect 186 350 217 371
rect 186 333 193 350
rect 210 333 217 350
rect 186 312 217 333
rect 186 295 193 312
rect 210 295 217 312
rect 186 274 217 295
rect 186 257 193 274
rect 210 257 217 274
rect 186 236 217 257
rect 298 350 329 371
rect 298 333 305 350
rect 322 333 329 350
rect 298 312 329 333
rect 298 295 305 312
rect 322 295 329 312
rect 298 274 329 295
rect 298 257 305 274
rect 322 257 329 274
rect 298 236 329 257
rect 354 350 385 371
rect 354 333 361 350
rect 378 333 385 350
rect 354 312 385 333
rect 354 295 361 312
rect 378 295 385 312
rect 354 274 385 295
rect 354 257 361 274
rect 378 257 385 274
rect 354 236 385 257
rect 410 350 441 371
rect 410 333 417 350
rect 434 333 441 350
rect 410 312 441 333
rect 410 295 417 312
rect 434 295 441 312
rect 410 274 441 295
rect 410 257 417 274
rect 434 257 441 274
rect 410 236 441 257
rect 522 350 553 371
rect 522 333 529 350
rect 546 333 553 350
rect 522 312 553 333
rect 522 295 529 312
rect 546 295 553 312
rect 522 274 553 295
rect 522 257 529 274
rect 546 257 553 274
rect 522 236 553 257
rect 578 350 609 371
rect 578 333 585 350
rect 602 333 609 350
rect 578 312 609 333
rect 578 295 585 312
rect 602 295 609 312
rect 578 274 609 295
rect 578 257 585 274
rect 602 257 609 274
rect 578 236 609 257
rect 636 350 667 371
rect 636 333 643 350
rect 660 333 667 350
rect 636 312 667 333
rect 636 295 643 312
rect 660 295 667 312
rect 636 274 667 295
rect 636 257 643 274
rect 660 257 667 274
rect 636 236 667 257
rect 692 350 723 371
rect 692 333 699 350
rect 716 333 723 350
rect 692 312 723 333
rect 692 295 699 312
rect 716 295 723 312
rect 692 274 723 295
rect 692 257 699 274
rect 716 257 723 274
rect 692 236 723 257
rect 32 219 49 236
rect 32 202 69 219
rect 5 177 22 185
rect 5 152 22 160
rect 52 135 69 202
rect 32 118 69 135
rect 95 132 112 140
rect 32 90 49 118
rect 95 107 112 115
rect 130 90 147 236
rect 165 211 182 219
rect 165 186 182 194
rect 200 169 217 236
rect 354 219 371 236
rect 234 211 251 219
rect 234 186 251 194
rect 283 211 371 219
rect 300 202 371 211
rect 283 186 300 194
rect 200 157 336 169
rect 200 152 319 157
rect 165 132 182 140
rect 165 107 182 115
rect 200 90 217 152
rect 234 127 251 135
rect 319 132 336 140
rect 234 102 251 110
rect 354 90 371 202
rect 389 211 406 219
rect 389 186 406 194
rect 424 169 441 236
rect 458 211 475 219
rect 458 186 475 194
rect 507 211 524 219
rect 578 211 595 236
rect 665 211 682 219
rect 524 194 665 211
rect 507 186 524 194
rect 424 157 560 169
rect 424 152 543 157
rect 389 132 406 140
rect 389 107 406 115
rect 424 90 441 152
rect 458 127 475 135
rect 543 132 560 140
rect 458 102 475 110
rect 578 90 595 194
rect 665 186 682 194
rect 706 129 723 236
rect 652 112 723 129
rect 706 90 723 112
rect 18 77 49 90
rect 18 60 25 77
rect 42 60 49 77
rect 18 48 49 60
rect 74 77 105 90
rect 74 60 81 77
rect 98 60 105 77
rect 74 48 105 60
rect 130 77 161 90
rect 130 60 137 77
rect 154 60 161 77
rect 130 48 161 60
rect 186 77 217 90
rect 186 60 193 77
rect 210 60 217 77
rect 186 48 217 60
rect 298 77 329 90
rect 298 60 305 77
rect 322 60 329 77
rect 298 48 329 60
rect 354 77 385 90
rect 354 60 361 77
rect 378 60 385 77
rect 354 48 385 60
rect 410 77 441 90
rect 410 60 417 77
rect 434 60 441 77
rect 410 48 441 60
rect 522 77 553 90
rect 522 60 529 77
rect 546 60 553 77
rect 522 48 553 60
rect 578 77 609 90
rect 578 60 585 77
rect 602 60 609 77
rect 578 48 609 60
rect 636 77 667 90
rect 636 60 643 77
rect 660 60 667 77
rect 636 48 667 60
rect 692 77 723 90
rect 692 60 699 77
rect 716 60 723 77
rect 692 48 723 60
rect 79 9 97 48
rect 312 31 329 48
rect 522 34 539 48
rect 79 -17 97 -9
rect 220 9 238 17
rect 312 14 379 31
rect 220 -17 238 -9
rect 361 9 379 14
rect 361 -17 379 -9
rect 502 17 539 34
rect 502 9 520 17
rect 502 -17 520 -9
rect 643 9 661 48
rect 643 -17 661 -9
<< viali >>
rect 79 410 97 428
rect 220 410 238 428
rect 361 410 379 428
rect 502 410 520 428
rect 643 410 661 428
rect 5 160 22 177
rect 95 115 112 132
rect 165 194 182 211
rect 234 194 251 211
rect 165 115 182 132
rect 234 110 251 127
rect 389 194 406 211
rect 458 194 475 211
rect 389 115 406 132
rect 458 110 475 127
rect 635 112 652 129
rect 25 60 42 77
rect 79 -9 97 9
rect 220 -9 238 9
rect 361 -9 379 9
rect 502 -9 520 9
rect 643 -9 661 9
<< metal1 >>
rect 0 428 741 434
rect 0 410 79 428
rect 97 410 220 428
rect 238 410 361 428
rect 379 410 502 428
rect 520 410 643 428
rect 661 410 741 428
rect 0 404 741 410
rect 162 213 185 219
rect 453 217 479 220
rect 13 211 185 213
rect 13 199 165 211
rect 13 185 27 199
rect 162 194 165 199
rect 182 194 185 211
rect 162 186 185 194
rect 229 211 409 217
rect 229 194 234 211
rect 251 203 389 211
rect 251 194 254 203
rect 229 186 254 194
rect 386 194 389 203
rect 406 194 409 211
rect 386 188 409 194
rect 453 188 479 191
rect 0 182 27 185
rect 0 156 1 182
rect 229 169 243 186
rect 0 152 27 156
rect 171 155 243 169
rect 390 174 404 188
rect 390 160 473 174
rect 90 137 117 140
rect 171 138 185 155
rect 90 111 91 137
rect 90 107 117 111
rect 162 132 185 138
rect 162 115 165 132
rect 182 115 185 132
rect 162 109 185 115
rect 230 133 256 136
rect 386 132 409 138
rect 459 133 473 160
rect 631 133 657 136
rect 386 123 389 132
rect 256 115 389 123
rect 406 115 409 132
rect 166 83 180 109
rect 256 109 409 115
rect 455 127 478 133
rect 455 110 458 127
rect 475 110 478 127
rect 230 103 256 107
rect 455 104 478 110
rect 631 104 657 107
rect 19 77 180 83
rect 19 60 25 77
rect 42 69 180 77
rect 42 60 48 69
rect 19 54 48 60
rect 0 9 741 15
rect 0 -9 79 9
rect 97 -9 220 9
rect 238 -9 361 9
rect 379 -9 502 9
rect 520 -9 643 9
rect 661 -9 741 9
rect 0 -15 741 -9
<< via1 >>
rect 453 211 479 217
rect 453 194 458 211
rect 458 194 475 211
rect 475 194 479 211
rect 453 191 479 194
rect 1 177 27 182
rect 1 160 5 177
rect 5 160 22 177
rect 22 160 27 177
rect 1 156 27 160
rect 91 132 117 137
rect 91 115 95 132
rect 95 115 112 132
rect 112 115 117 132
rect 91 111 117 115
rect 230 127 256 133
rect 230 110 234 127
rect 234 110 251 127
rect 251 110 256 127
rect 230 107 256 110
rect 631 129 657 133
rect 631 112 635 129
rect 635 112 652 129
rect 652 112 657 129
rect 631 107 657 112
<< metal2 >>
rect 453 217 479 220
rect 424 197 453 211
rect 1 182 27 185
rect 0 161 1 175
rect 1 152 27 156
rect 13 90 27 152
rect 91 137 117 140
rect 90 116 91 130
rect 91 108 117 111
rect 230 133 256 136
rect 230 104 256 107
rect 242 90 256 104
rect 424 90 438 197
rect 453 188 479 191
rect 631 133 657 136
rect 630 114 631 128
rect 631 104 657 107
rect 13 76 438 90
<< labels >>
flabel metal2 0 167 0 167 0 FreeSans 80 0 0 0 clk
port 2 nsew
flabel metal1 39 423 39 423 0 FreeSans 80 0 0 0 vdd
port 3 nsew
flabel metal1 31 1 31 1 0 FreeSans 80 0 0 0 gnd
port 4 nsew
flabel metal1 34 56 34 56 0 FreeSans 80 0 0 0 clkb
flabel locali 138 166 138 166 0 FreeSans 80 0 0 0 net1
flabel locali 211 177 211 177 0 FreeSans 80 0 0 0 net2
flabel pdiff 258 282 258 282 0 FreeSans 80 0 0 0 net4
flabel ndiff 249 62 249 62 0 FreeSans 80 0 0 0 net5
flabel locali 362 176 362 176 0 FreeSans 80 0 0 0 net3
flabel locali 434 215 434 215 0 FreeSans 80 0 0 0 net6
flabel locali 589 143 589 143 0 FreeSans 80 0 0 0 net7
flabel pdiff 478 276 478 276 0 FreeSans 80 0 0 0 net8
flabel ndiff 480 68 480 68 0 FreeSans 80 0 0 0 net9
flabel metal2 90 121 90 121 0 FreeSans 80 0 0 0 D
port 7 nsew
flabel metal2 630 120 630 120 0 FreeSans 80 0 0 0 Q
port 8 nsew
<< properties >>
string FIXED_BBOX 0 0 741 419
<< end >>
