magic
tech sky130A
magscale 1 2
timestamp 1644949024
<< checkpaint >>
rect -1260 -1302 8060 25929
<< metal1 >>
rect 5166 24026 5460 24028
rect 5166 24000 6080 24026
rect 5432 23998 6080 24000
rect 6706 23928 6734 23956
rect 5166 23878 5778 23906
rect 6706 23802 6734 23830
rect 5166 23732 5600 23760
rect 6706 23576 6734 23604
rect 6706 22536 6734 22564
rect 5166 22380 5600 22408
rect 6706 22310 6734 22338
rect 5166 22234 5778 22262
rect 6706 22184 6734 22212
rect 5432 22140 6080 22142
rect 5166 22114 6080 22140
rect 5166 22112 5460 22114
rect 5166 20950 5460 20952
rect 5166 20924 6080 20950
rect 5432 20922 6080 20924
rect 6706 20852 6734 20880
rect 5166 20802 5778 20830
rect 6706 20726 6734 20754
rect 5166 20656 5600 20684
rect 6706 20500 6734 20528
rect 6706 19460 6734 19488
rect 5166 19304 5600 19332
rect 6706 19234 6734 19262
rect 5166 19158 5778 19186
rect 6706 19108 6734 19136
rect 5432 19064 6080 19066
rect 5166 19038 6080 19064
rect 5166 19036 5460 19038
rect 5166 17874 5460 17876
rect 5166 17848 6080 17874
rect 5432 17846 6080 17848
rect 6706 17776 6734 17804
rect 5166 17726 5778 17754
rect 6706 17650 6734 17678
rect 5166 17580 5600 17608
rect 6706 17424 6734 17452
rect 6706 16384 6734 16412
rect 5166 16228 5600 16256
rect 6706 16158 6734 16186
rect 5166 16082 5778 16110
rect 6706 16032 6734 16060
rect 5432 15988 6080 15990
rect 5166 15962 6080 15988
rect 5166 15960 5460 15962
rect 5166 14798 5460 14800
rect 5166 14772 6080 14798
rect 5432 14770 6080 14772
rect 6706 14700 6734 14728
rect 5166 14650 5778 14678
rect 6706 14574 6734 14602
rect 5166 14504 5600 14532
rect 6706 14348 6734 14376
rect 6706 13308 6734 13336
rect 5166 13152 5600 13180
rect 6706 13082 6734 13110
rect 5166 13006 5778 13034
rect 6706 12956 6734 12984
rect 5432 12912 6080 12914
rect 5166 12886 6080 12912
rect 5166 12884 5460 12886
rect 5166 11722 5460 11724
rect 5166 11696 6080 11722
rect 5432 11694 6080 11696
rect 6706 11624 6734 11652
rect 5166 11574 5778 11602
rect 6706 11498 6734 11526
rect 5166 11428 5600 11456
rect 6706 11272 6734 11300
rect 6706 10232 6734 10260
rect 5166 10076 5600 10104
rect 6706 10006 6734 10034
rect 5166 9930 5778 9958
rect 6706 9880 6734 9908
rect 5432 9836 6080 9838
rect 5166 9810 6080 9836
rect 5166 9808 5460 9810
rect 5166 8646 5460 8648
rect 5166 8620 6080 8646
rect 5432 8618 6080 8620
rect 6706 8548 6734 8576
rect 5166 8498 5778 8526
rect 6706 8422 6734 8450
rect 5166 8352 5600 8380
rect 6706 8196 6734 8224
rect 6706 7156 6734 7184
rect 5166 7000 5600 7028
rect 6706 6930 6734 6958
rect 5166 6854 5778 6882
rect 6706 6804 6734 6832
rect 5432 6760 6080 6762
rect 5166 6734 6080 6760
rect 5166 6732 5460 6734
rect 5166 5570 5460 5572
rect 5166 5544 6080 5570
rect 5432 5542 6080 5544
rect 6706 5472 6734 5500
rect 5166 5422 5778 5450
rect 6706 5346 6734 5374
rect 5166 5276 5600 5304
rect 6706 5120 6734 5148
rect 6706 4080 6734 4108
rect 5166 3924 5600 3952
rect 6706 3854 6734 3882
rect 5166 3778 5778 3806
rect 6706 3728 6734 3756
rect 5432 3684 6080 3686
rect 5166 3658 6080 3684
rect 5166 3656 5460 3658
rect 5166 2494 5460 2496
rect 5166 2468 6080 2494
rect 5432 2466 6080 2468
rect 6706 2396 6734 2424
rect 5166 2346 5778 2374
rect 6706 2270 6734 2298
rect 5166 2200 5600 2228
rect 6706 2044 6734 2072
rect 6706 1004 6734 1032
rect 5166 848 5600 876
rect 6706 778 6734 806
rect 5166 702 5778 730
rect 6706 652 6734 680
rect 5432 608 6080 610
rect 5166 582 6080 608
rect 5166 580 5460 582
<< metal2 >>
rect 18 0 46 24632
rect 102 0 130 24632
rect 186 0 214 24632
rect 270 0 298 24632
rect 354 0 382 24632
rect 438 0 466 24632
rect 5344 24594 5558 24622
<< metal3 >>
rect 792 24595 924 24669
rect 1664 24595 1796 24669
rect 5128 24571 5260 24645
rect 6668 24571 6800 24645
rect 792 23055 924 23129
rect 1664 23055 1796 23129
rect 5128 23033 5260 23107
rect 6668 23033 6800 23107
rect 792 21515 924 21589
rect 1664 21515 1796 21589
rect 5128 21495 5260 21569
rect 6668 21495 6800 21569
rect 792 19975 924 20049
rect 1664 19975 1796 20049
rect 5128 19957 5260 20031
rect 6668 19957 6800 20031
rect 792 18435 924 18509
rect 1664 18435 1796 18509
rect 5128 18419 5260 18493
rect 6668 18419 6800 18493
rect 5128 16881 5260 16955
rect 6668 16881 6800 16955
rect 792 15359 924 15433
rect 1664 15359 1796 15433
rect 5128 15343 5260 15417
rect 6668 15343 6800 15417
rect 792 13819 924 13893
rect 1664 13819 1796 13893
rect 5128 13805 5260 13879
rect 6668 13805 6800 13879
rect 792 12279 924 12353
rect 1664 12279 1796 12353
rect 5128 12267 5260 12341
rect 6668 12267 6800 12341
rect 792 10739 924 10813
rect 1664 10739 1796 10813
rect 5128 10729 5260 10803
rect 6668 10729 6800 10803
rect 792 9199 924 9273
rect 1664 9199 1796 9273
rect 5128 9191 5260 9265
rect 6668 9191 6800 9265
rect 5128 7653 5260 7727
rect 6668 7653 6800 7727
rect 792 6123 924 6197
rect 1664 6123 1796 6197
rect 5128 6115 5260 6189
rect 6668 6115 6800 6189
rect 792 4583 924 4657
rect 1664 4583 1796 4657
rect 5128 4577 5260 4651
rect 6668 4577 6800 4651
rect 792 3043 924 3117
rect 1664 3043 1796 3117
rect 5128 3039 5260 3113
rect 6668 3039 6800 3113
rect 792 1503 924 1577
rect 1664 1503 1796 1577
rect 5128 1501 5260 1575
rect 6668 1501 6800 1575
rect 792 -37 924 37
rect 1664 -37 1796 37
rect 5128 -37 5260 37
rect 6668 -37 6800 37
use wordline_driver_array  wordline_driver_array_0
timestamp 1644949024
transform 1 0 5530 0 1 0
box 0 -42 1270 24650
use hierarchical_decoder  hierarchical_decoder_0
timestamp 1644949024
transform 1 0 0 0 1 0
box 0 -42 5260 24669
<< labels >>
rlabel metal2 s 18 0 46 24632 4 addr0
rlabel metal2 s 102 0 130 24632 4 addr1
rlabel metal2 s 186 0 214 24632 4 addr2
rlabel metal2 s 270 0 298 24632 4 addr3
rlabel metal2 s 354 0 382 24632 4 addr4
rlabel metal2 s 438 0 466 24632 4 addr5
rlabel metal1 s 6706 778 6734 806 4 rwl0_0
rlabel metal1 s 6706 1004 6734 1032 4 rwl1_0
rlabel metal1 s 6706 652 6734 680 4 wwl0_0
rlabel metal1 s 6706 2270 6734 2298 4 rwl0_1
rlabel metal1 s 6706 2044 6734 2072 4 rwl1_1
rlabel metal1 s 6706 2396 6734 2424 4 wwl0_1
rlabel metal1 s 6706 3854 6734 3882 4 rwl0_2
rlabel metal1 s 6706 4080 6734 4108 4 rwl1_2
rlabel metal1 s 6706 3728 6734 3756 4 wwl0_2
rlabel metal1 s 6706 5346 6734 5374 4 rwl0_3
rlabel metal1 s 6706 5120 6734 5148 4 rwl1_3
rlabel metal1 s 6706 5472 6734 5500 4 wwl0_3
rlabel metal1 s 6706 6930 6734 6958 4 rwl0_4
rlabel metal1 s 6706 7156 6734 7184 4 rwl1_4
rlabel metal1 s 6706 6804 6734 6832 4 wwl0_4
rlabel metal1 s 6706 8422 6734 8450 4 rwl0_5
rlabel metal1 s 6706 8196 6734 8224 4 rwl1_5
rlabel metal1 s 6706 8548 6734 8576 4 wwl0_5
rlabel metal1 s 6706 10006 6734 10034 4 rwl0_6
rlabel metal1 s 6706 10232 6734 10260 4 rwl1_6
rlabel metal1 s 6706 9880 6734 9908 4 wwl0_6
rlabel metal1 s 6706 11498 6734 11526 4 rwl0_7
rlabel metal1 s 6706 11272 6734 11300 4 rwl1_7
rlabel metal1 s 6706 11624 6734 11652 4 wwl0_7
rlabel metal1 s 6706 13082 6734 13110 4 rwl0_8
rlabel metal1 s 6706 13308 6734 13336 4 rwl1_8
rlabel metal1 s 6706 12956 6734 12984 4 wwl0_8
rlabel metal1 s 6706 14574 6734 14602 4 rwl0_9
rlabel metal1 s 6706 14348 6734 14376 4 rwl1_9
rlabel metal1 s 6706 14700 6734 14728 4 wwl0_9
rlabel metal1 s 6706 16158 6734 16186 4 rwl0_10
rlabel metal1 s 6706 16384 6734 16412 4 rwl1_10
rlabel metal1 s 6706 16032 6734 16060 4 wwl0_10
rlabel metal1 s 6706 17650 6734 17678 4 rwl0_11
rlabel metal1 s 6706 17424 6734 17452 4 rwl1_11
rlabel metal1 s 6706 17776 6734 17804 4 wwl0_11
rlabel metal1 s 6706 19234 6734 19262 4 rwl0_12
rlabel metal1 s 6706 19460 6734 19488 4 rwl1_12
rlabel metal1 s 6706 19108 6734 19136 4 wwl0_12
rlabel metal1 s 6706 20726 6734 20754 4 rwl0_13
rlabel metal1 s 6706 20500 6734 20528 4 rwl1_13
rlabel metal1 s 6706 20852 6734 20880 4 wwl0_13
rlabel metal1 s 6706 22310 6734 22338 4 rwl0_14
rlabel metal1 s 6706 22536 6734 22564 4 rwl1_14
rlabel metal1 s 6706 22184 6734 22212 4 wwl0_14
rlabel metal1 s 6706 23802 6734 23830 4 rwl0_15
rlabel metal1 s 6706 23576 6734 23604 4 rwl1_15
rlabel metal1 s 6706 23928 6734 23956 4 wwl0_15
rlabel metal2 s 5530 24594 5558 24622 4 wl_en
rlabel metal3 s 1664 19975 1796 20049 4 vdd
rlabel metal3 s 792 19975 924 20049 4 vdd
rlabel metal3 s 5128 10729 5260 10803 4 vdd
rlabel metal3 s 6668 19957 6800 20031 4 vdd
rlabel metal3 s 1664 13819 1796 13893 4 vdd
rlabel metal3 s 792 13819 924 13893 4 vdd
rlabel metal3 s 792 10739 924 10813 4 vdd
rlabel metal3 s 6668 16881 6800 16955 4 vdd
rlabel metal3 s 6668 13805 6800 13879 4 vdd
rlabel metal3 s 5128 23033 5260 23107 4 vdd
rlabel metal3 s 5128 13805 5260 13879 4 vdd
rlabel metal3 s 6668 23033 6800 23107 4 vdd
rlabel metal3 s 5128 7653 5260 7727 4 vdd
rlabel metal3 s 792 23055 924 23129 4 vdd
rlabel metal3 s 1664 23055 1796 23129 4 vdd
rlabel metal3 s 5128 4577 5260 4651 4 vdd
rlabel metal3 s 5128 1501 5260 1575 4 vdd
rlabel metal3 s 1664 1503 1796 1577 4 vdd
rlabel metal3 s 5128 19957 5260 20031 4 vdd
rlabel metal3 s 792 1503 924 1577 4 vdd
rlabel metal3 s 1664 4583 1796 4657 4 vdd
rlabel metal3 s 5128 16881 5260 16955 4 vdd
rlabel metal3 s 6668 4577 6800 4651 4 vdd
rlabel metal3 s 6668 7653 6800 7727 4 vdd
rlabel metal3 s 6668 10729 6800 10803 4 vdd
rlabel metal3 s 792 4583 924 4657 4 vdd
rlabel metal3 s 1664 10739 1796 10813 4 vdd
rlabel metal3 s 6668 1501 6800 1575 4 vdd
rlabel metal3 s 6668 12267 6800 12341 4 gnd
rlabel metal3 s 1664 6123 1796 6197 4 gnd
rlabel metal3 s 5128 24571 5260 24645 4 gnd
rlabel metal3 s 5128 18419 5260 18493 4 gnd
rlabel metal3 s 792 -37 924 37 4 gnd
rlabel metal3 s 5128 12267 5260 12341 4 gnd
rlabel metal3 s 792 21515 924 21589 4 gnd
rlabel metal3 s 6668 6115 6800 6189 4 gnd
rlabel metal3 s 1664 12279 1796 12353 4 gnd
rlabel metal3 s 792 15359 924 15433 4 gnd
rlabel metal3 s 792 12279 924 12353 4 gnd
rlabel metal3 s 5128 21495 5260 21569 4 gnd
rlabel metal3 s 6668 9191 6800 9265 4 gnd
rlabel metal3 s 792 3043 924 3117 4 gnd
rlabel metal3 s 1664 9199 1796 9273 4 gnd
rlabel metal3 s 1664 24595 1796 24669 4 gnd
rlabel metal3 s 792 24595 924 24669 4 gnd
rlabel metal3 s 1664 -37 1796 37 4 gnd
rlabel metal3 s 6668 15343 6800 15417 4 gnd
rlabel metal3 s 792 18435 924 18509 4 gnd
rlabel metal3 s 6668 24571 6800 24645 4 gnd
rlabel metal3 s 1664 15359 1796 15433 4 gnd
rlabel metal3 s 5128 9191 5260 9265 4 gnd
rlabel metal3 s 1664 3043 1796 3117 4 gnd
rlabel metal3 s 5128 6115 5260 6189 4 gnd
rlabel metal3 s 792 6123 924 6197 4 gnd
rlabel metal3 s 792 9199 924 9273 4 gnd
rlabel metal3 s 5128 -37 5260 37 4 gnd
rlabel metal3 s 6668 18419 6800 18493 4 gnd
rlabel metal3 s 1664 18435 1796 18509 4 gnd
rlabel metal3 s 6668 -37 6800 37 4 gnd
rlabel metal3 s 5128 15343 5260 15417 4 gnd
rlabel metal3 s 5128 3039 5260 3113 4 gnd
rlabel metal3 s 6668 3039 6800 3113 4 gnd
rlabel metal3 s 6668 21495 6800 21569 4 gnd
rlabel metal3 s 1664 21515 1796 21589 4 gnd
<< properties >>
string FIXED_BBOX 0 0 6770 24660
string GDS_FILE sram_0rw2r1w_4_16_sky130A.gds
string GDS_END 268042
string GDS_START 230104
<< end >>
