magic
tech sky130A
magscale 1 2
timestamp 1644951705
<< checkpaint >>
rect -1211 -1260 2104 2768
<< pwell >>
rect 753 718 803 800
<< psubdiff >>
rect 753 776 803 800
rect 753 742 761 776
rect 795 742 803 776
rect 753 718 803 742
<< psubdiffcont >>
rect 761 742 795 776
<< poly >>
rect 374 726 404 780
rect 374 28 404 54
<< locali >>
rect 115 1435 456 1469
rect 422 1116 456 1435
rect 761 776 795 792
rect 761 726 795 742
rect 322 73 356 390
rect 322 39 691 73
<< viali >>
rect 81 1435 115 1469
rect 322 1099 356 1133
rect 761 742 795 776
rect 422 373 456 407
rect 691 39 725 73
<< metal1 >>
rect 66 1469 72 1478
rect 124 1469 130 1478
rect 49 1435 72 1469
rect 124 1435 147 1469
rect 66 1426 72 1435
rect 124 1426 130 1435
rect 310 1133 368 1139
rect 310 1099 322 1133
rect 356 1099 368 1133
rect 310 1093 368 1099
rect 325 470 353 1093
rect 694 952 722 1452
rect 84 442 353 470
rect 425 924 722 952
rect 84 56 112 442
rect 425 413 453 924
rect 746 733 752 785
rect 804 733 810 785
rect 410 407 468 413
rect 410 373 422 407
rect 456 373 468 407
rect 410 367 468 373
rect 676 73 682 82
rect 734 73 740 82
rect 659 39 682 73
rect 734 39 757 73
rect 676 30 682 39
rect 734 30 740 39
<< via1 >>
rect 72 1469 124 1478
rect 72 1435 81 1469
rect 81 1435 115 1469
rect 115 1435 124 1469
rect 72 1426 124 1435
rect 752 776 804 785
rect 752 742 761 776
rect 761 742 795 776
rect 795 742 804 776
rect 752 733 804 742
rect 682 73 734 82
rect 682 39 691 73
rect 691 39 725 73
rect 725 39 734 73
rect 682 30 734 39
<< metal2 >>
rect 84 1484 112 1508
rect 72 1478 124 1484
rect 694 1452 722 1508
rect 72 1420 124 1426
rect 750 787 806 796
rect 750 722 806 731
rect 682 82 734 88
rect 84 0 112 56
rect 682 24 734 30
rect 694 0 722 24
<< via2 >>
rect 750 785 806 787
rect 750 733 752 785
rect 752 733 804 785
rect 804 733 806 785
rect 750 731 806 733
<< metal3 >>
rect 712 787 844 796
rect 712 731 750 787
rect 806 731 844 787
rect 712 722 844 731
use contact_18  contact_18_0
timestamp 1644951705
transform 1 0 712 0 1 722
box 0 0 1 1
use contact_17  contact_17_0
timestamp 1644951705
transform 1 0 746 0 1 727
box 0 0 1 1
use contact_13  contact_13_0
timestamp 1644951705
transform 1 0 749 0 1 736
box 0 0 1 1
use contact_25  contact_25_0
timestamp 1644951705
transform 1 0 753 0 1 718
box 0 0 1 1
use contact_13  contact_13_1
timestamp 1644951705
transform 1 0 410 0 1 367
box 0 0 1 1
use contact_13  contact_13_2
timestamp 1644951705
transform 1 0 310 0 1 1093
box 0 0 1 1
use contact_13  contact_13_3
timestamp 1644951705
transform 1 0 679 0 1 33
box 0 0 1 1
use contact_17  contact_17_1
timestamp 1644951705
transform 1 0 676 0 1 24
box 0 0 1 1
use contact_13  contact_13_4
timestamp 1644951705
transform 1 0 69 0 1 1429
box 0 0 1 1
use contact_17  contact_17_2
timestamp 1644951705
transform 1 0 66 0 1 1420
box 0 0 1 1
use nmos_m1_w3_360_sli_dli  nmos_m1_w3_360_sli_dli_0
timestamp 1644951705
transform 1 0 314 0 1 780
box 0 -26 150 698
use nmos_m1_w3_360_sli_dli  nmos_m1_w3_360_sli_dli_1
timestamp 1644951705
transform 1 0 314 0 1 54
box 0 -26 150 698
<< labels >>
rlabel mvvaractor s 389 41 389 41 4 sel
rlabel metal2 s 84 1452 112 1508 4 rbl0
rlabel metal2 s 694 1452 722 1508 4 rbl1
rlabel metal2 s 84 0 112 56 4 rbl0_out
rlabel metal2 s 694 0 722 56 4 rbl1_out
rlabel metal3 s 712 722 844 796 4 gnd
<< properties >>
string FIXED_BBOX 0 0 778 693
string GDS_FILE sram_0rw2r1w_16_128_sky130A.gds
string GDS_END 1595010
string GDS_START 1592034
<< end >>
