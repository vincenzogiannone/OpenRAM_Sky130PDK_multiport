magic
tech sky130A
magscale 1 2
timestamp 1644969367
<< checkpaint >>
rect -1260 -1286 1626 1403
<< scnmos >>
rect 60 0 90 84
rect 168 0 198 84
rect 276 0 306 84
<< ndiff >>
rect 0 59 60 84
rect 0 25 8 59
rect 42 25 60 59
rect 0 0 60 25
rect 90 59 168 84
rect 90 25 112 59
rect 146 25 168 59
rect 90 0 168 25
rect 198 59 276 84
rect 198 25 220 59
rect 254 25 276 59
rect 198 0 276 25
rect 306 59 366 84
rect 306 25 324 59
rect 358 25 366 59
rect 306 0 366 25
<< ndiffc >>
rect 8 25 42 59
rect 112 25 146 59
rect 220 25 254 59
rect 324 25 358 59
<< poly >>
rect 60 110 306 140
rect 60 84 90 110
rect 168 84 198 110
rect 276 84 306 110
rect 60 -26 90 0
rect 168 -26 198 0
rect 276 -26 306 0
<< locali >>
rect 112 109 358 143
rect 8 59 42 75
rect 8 9 42 25
rect 112 59 146 109
rect 112 9 146 25
rect 220 59 254 75
rect 220 9 254 25
rect 324 59 358 109
rect 324 9 358 25
use contact_8  contact_8_0
timestamp 1644969367
transform 1 0 316 0 1 1
box 0 0 1 1
use contact_8  contact_8_1
timestamp 1644969367
transform 1 0 212 0 1 1
box 0 0 1 1
use contact_8  contact_8_2
timestamp 1644969367
transform 1 0 104 0 1 1
box 0 0 1 1
use contact_8  contact_8_3
timestamp 1644969367
transform 1 0 0 0 1 1
box 0 0 1 1
<< labels >>
rlabel mvvaractor s 183 125 183 125 4 G
rlabel locali s 237 42 237 42 4 S
rlabel locali s 25 42 25 42 4 S
rlabel locali s 235 126 235 126 4 D
<< properties >>
string FIXED_BBOX -25 -26 391 143
string GDS_FILE sram_0rw2r1w_32_128_sky130A.gds
string GDS_END 3311052
string GDS_START 3309832
<< end >>
