magic
tech sky130A
magscale 1 2
timestamp 1643678851
<< checkpaint >>
rect -1260 -1260 122464 64800
<< metal2 >>
rect 13004 7245 13032 12430
rect 14705 12420 14733 27410
rect 14773 13612 14801 27410
rect 14841 14096 14869 27410
rect 14909 15288 14937 27410
rect 14977 15772 15005 27410
rect 15045 16964 15073 27410
rect 15113 17448 15141 27410
rect 20068 11545 20096 61230
rect 21190 9871 21218 11960
rect 12121 7231 13032 7245
rect 12121 7217 13084 7231
rect 12952 3038 13084 7217
rect 71664 6210 71692 10556
rect 12952 3010 12990 3038
rect 13046 3010 13084 3038
<< via2 >>
rect 13265 17396 13321 17452
rect 14345 17392 14401 17448
rect 13265 16904 13321 16960
rect 14345 16908 14401 16964
rect 13265 15720 13321 15776
rect 14345 15716 14401 15772
rect 13265 15228 13321 15284
rect 14345 15232 14401 15288
rect 13265 14044 13321 14100
rect 14345 14040 14401 14096
rect 13265 13552 13321 13608
rect 14345 13556 14401 13612
rect 12990 12430 13046 12486
rect 2863 7426 2919 7482
rect 6223 7211 6279 7267
rect 13265 12368 13321 12424
rect 15099 17392 15155 17448
rect 15031 16908 15087 16964
rect 14963 15716 15019 15772
rect 14895 15232 14951 15288
rect 14827 14040 14883 14096
rect 14759 13556 14815 13612
rect 14345 12364 14401 12420
rect 14691 12364 14747 12420
rect 14540 11489 14596 11545
rect 20054 11489 20110 11545
rect 14540 10556 14596 10612
rect 22298 10642 22354 10698
rect 25410 10642 25466 10698
rect 28522 10642 28578 10698
rect 31634 10642 31690 10698
rect 34746 10642 34802 10698
rect 37858 10642 37914 10698
rect 40970 10642 41026 10698
rect 44082 10642 44138 10698
rect 47194 10642 47250 10698
rect 50306 10642 50362 10698
rect 53418 10642 53474 10698
rect 56530 10642 56586 10698
rect 59642 10642 59698 10698
rect 62754 10642 62810 10698
rect 65866 10642 65922 10698
rect 68978 10642 69034 10698
rect 71650 10556 71706 10612
rect 14540 9815 14596 9871
rect 21176 9815 21232 9871
rect 2863 6242 2919 6298
rect 12990 2982 13046 3038
rect 16229 2920 16285 2976
rect 17711 2920 17767 2976
rect 19193 2920 19249 2976
rect 20675 2920 20731 2976
rect 22157 2920 22213 2976
rect 23639 2920 23695 2976
rect 25121 2920 25177 2976
rect 26603 2920 26659 2976
rect 28085 2920 28141 2976
rect 29567 2920 29623 2976
rect 31049 2920 31105 2976
rect 32531 2920 32587 2976
rect 34013 2920 34069 2976
rect 35495 2920 35551 2976
rect 36977 2920 37033 2976
rect 38459 2920 38515 2976
rect 39941 2920 39997 2976
rect 41423 2920 41479 2976
<< metal3 >>
rect 424 63496 121204 63540
rect 424 63432 468 63496
rect 532 63432 680 63496
rect 744 63432 892 63496
rect 956 63432 120672 63496
rect 120736 63432 120884 63496
rect 120948 63432 121096 63496
rect 121160 63432 121204 63496
rect 424 63284 121204 63432
rect 424 63220 468 63284
rect 532 63220 680 63284
rect 744 63220 892 63284
rect 956 63220 120672 63284
rect 120736 63220 120884 63284
rect 120948 63220 121096 63284
rect 121160 63220 121204 63284
rect 424 63072 121204 63220
rect 424 63008 468 63072
rect 532 63008 680 63072
rect 744 63008 892 63072
rect 956 63008 21456 63072
rect 21520 63008 120672 63072
rect 120736 63008 120884 63072
rect 120948 63008 121096 63072
rect 121160 63008 121204 63072
rect 424 62964 121204 63008
rect 1484 62436 120144 62480
rect 1484 62372 1528 62436
rect 1592 62372 1740 62436
rect 1804 62372 1952 62436
rect 2016 62372 119612 62436
rect 119676 62372 119824 62436
rect 119888 62372 120036 62436
rect 120100 62372 120144 62436
rect 1484 62224 120144 62372
rect 1484 62160 1528 62224
rect 1592 62160 1740 62224
rect 1804 62160 1952 62224
rect 2016 62160 119612 62224
rect 119676 62160 119824 62224
rect 119888 62160 120036 62224
rect 120100 62160 120144 62224
rect 1484 62012 120144 62160
rect 1484 61948 1528 62012
rect 1592 61948 1740 62012
rect 1804 61948 1952 62012
rect 2016 61948 21244 62012
rect 21308 61948 119612 62012
rect 119676 61948 119824 62012
rect 119888 61948 120036 62012
rect 120100 61948 120144 62012
rect 1484 61904 120144 61948
rect 21200 61376 21564 61420
rect 21200 61312 21456 61376
rect 21520 61312 21564 61376
rect 21200 61268 21564 61312
rect 21200 61208 21352 61268
rect 20216 61164 21352 61208
rect 20140 61100 20184 61164
rect 20248 61100 21352 61164
rect 20216 61056 21352 61100
rect 19928 60528 21140 60572
rect 19928 60464 20184 60528
rect 20248 60464 21032 60528
rect 21096 60464 21140 60528
rect 19928 60420 21140 60464
rect 21200 59892 21352 59936
rect 21200 59828 21244 59892
rect 21308 59828 21352 59892
rect 21200 59680 21352 59828
rect 21200 59616 21244 59680
rect 21308 59616 21352 59680
rect 21200 59572 21352 59616
rect 19928 59044 21352 59088
rect 19928 58980 21244 59044
rect 21308 58980 21352 59044
rect 19928 58936 21352 58980
rect 19928 58876 20292 58936
rect 19928 58832 21352 58876
rect 19928 58768 21244 58832
rect 21308 58768 21352 58832
rect 19928 58724 21352 58768
rect 21064 58196 21352 58240
rect 20988 58132 21032 58196
rect 21096 58132 21352 58196
rect 21064 58088 21352 58132
rect 21200 57604 21352 58088
rect 19928 57452 21352 57604
rect 19928 57392 20292 57452
rect 19928 57348 21140 57392
rect 19928 57284 21032 57348
rect 21096 57284 21140 57348
rect 19928 57240 21140 57284
rect 21200 56712 21352 56756
rect 21200 56648 21244 56712
rect 21308 56648 21352 56712
rect 21200 56500 21352 56648
rect 21200 56436 21244 56500
rect 21308 56436 21352 56500
rect 21200 56392 21352 56436
rect 19928 56076 21352 56120
rect 19928 56012 21244 56076
rect 21308 56012 21352 56076
rect 19928 55968 21352 56012
rect 19928 55908 20292 55968
rect 19928 55864 21352 55908
rect 19928 55800 21244 55864
rect 21308 55800 21352 55864
rect 19928 55756 21352 55800
rect 21064 55228 21352 55272
rect 20988 55164 21032 55228
rect 21096 55164 21352 55228
rect 21064 55120 21352 55164
rect 21200 54636 21352 55120
rect 19928 54484 21352 54636
rect 19928 54424 20292 54484
rect 19928 54380 21140 54424
rect 19928 54316 21032 54380
rect 21096 54316 21140 54380
rect 19928 54272 21140 54316
rect 20216 53532 21352 53576
rect 20140 53468 20184 53532
rect 20248 53468 21244 53532
rect 21308 53468 21352 53532
rect 20216 53424 21352 53468
rect 19928 52896 21352 52940
rect 19928 52832 20184 52896
rect 20248 52832 21244 52896
rect 21308 52832 21352 52896
rect 19928 52788 21352 52832
rect 21064 52048 21352 52092
rect 20988 51984 21032 52048
rect 21096 51984 21352 52048
rect 21064 51940 21352 51984
rect 21200 51456 21352 51940
rect 19928 51412 21352 51456
rect 19928 51348 19972 51412
rect 20036 51348 21352 51412
rect 19928 51304 21352 51348
rect 21200 50564 21352 50608
rect 21200 50500 21244 50564
rect 21308 50500 21352 50564
rect 21200 50352 21352 50500
rect 21200 50288 21244 50352
rect 21308 50288 21352 50352
rect 21200 50244 21352 50288
rect 19928 49928 21352 49972
rect 19928 49864 20184 49928
rect 20248 49864 21244 49928
rect 21308 49864 21352 49928
rect 19928 49820 21352 49864
rect 20004 49080 21352 49124
rect 19928 49016 19972 49080
rect 20036 49016 21352 49080
rect 20004 48972 21352 49016
rect 21200 48868 21352 48972
rect 21200 48804 21244 48868
rect 21308 48804 21352 48868
rect 21200 48760 21352 48804
rect 19928 48444 21352 48488
rect 19928 48380 21244 48444
rect 21308 48380 21352 48444
rect 19928 48336 21352 48380
rect 19928 48276 20292 48336
rect 19928 48232 21140 48276
rect 19928 48168 21032 48232
rect 21096 48168 21140 48232
rect 19928 48124 21140 48168
rect 20216 47384 21352 47428
rect 20140 47320 20184 47384
rect 20248 47320 21244 47384
rect 21308 47320 21352 47384
rect 20216 47276 21352 47320
rect 19928 46960 21352 47004
rect 19928 46896 21244 46960
rect 21308 46896 21352 46960
rect 19928 46852 21352 46896
rect 19928 46792 20292 46852
rect 19928 46748 21352 46792
rect 19928 46684 21244 46748
rect 21308 46684 21352 46748
rect 19928 46640 21352 46684
rect 21064 45900 21352 45944
rect 20988 45836 21032 45900
rect 21096 45836 21352 45900
rect 21064 45792 21352 45836
rect 21200 45520 21352 45792
rect 19928 45368 21352 45520
rect 19928 45308 20292 45368
rect 19928 45264 21140 45308
rect 19928 45200 21032 45264
rect 21096 45200 21140 45264
rect 19928 45156 21140 45200
rect 21200 44416 21352 44460
rect 21200 44352 21244 44416
rect 21308 44352 21352 44416
rect 21200 44036 21352 44352
rect 19928 43884 21352 44036
rect 19928 43824 20292 43884
rect 19928 43780 21352 43824
rect 19928 43716 21244 43780
rect 21308 43716 21352 43780
rect 19928 43672 21352 43716
rect 15264 42824 16688 42976
rect 21064 42932 21352 42976
rect 20988 42868 21032 42932
rect 21096 42868 21352 42932
rect 21064 42824 21352 42868
rect 15264 42612 15628 42824
rect 16324 42764 16688 42824
rect 16188 42720 16688 42764
rect 16112 42656 16156 42720
rect 16220 42656 16688 42720
rect 16188 42612 16688 42656
rect 21200 42340 21352 42824
rect 19928 42296 21352 42340
rect 19928 42232 19972 42296
rect 20036 42232 21352 42296
rect 19928 42188 21352 42232
rect 15264 41280 15628 41492
rect 16324 41280 16688 41492
rect 15264 41236 16688 41280
rect 20216 41236 21352 41280
rect 15264 41172 15308 41236
rect 15372 41172 16688 41236
rect 20140 41172 20184 41236
rect 20248 41172 21244 41236
rect 21308 41172 21352 41236
rect 15264 41128 16688 41172
rect 20216 41128 21352 41172
rect 19928 40812 21352 40856
rect 19928 40748 20184 40812
rect 20248 40748 21244 40812
rect 21308 40748 21352 40812
rect 19928 40704 21352 40748
rect 15476 39856 16476 40008
rect 15476 39796 15628 39856
rect 16324 39796 16476 39856
rect 15264 39752 16264 39796
rect 15264 39688 16156 39752
rect 16220 39688 16264 39752
rect 15264 39644 16264 39688
rect 16324 39752 16688 39796
rect 20004 39752 21352 39796
rect 16324 39688 16368 39752
rect 16432 39688 16688 39752
rect 19928 39688 19972 39752
rect 20036 39688 21352 39752
rect 16324 39644 16688 39688
rect 20004 39644 21352 39688
rect 21200 39372 21352 39644
rect 19928 39328 21352 39372
rect 19928 39264 20184 39328
rect 20248 39264 21352 39328
rect 19928 39220 21352 39264
rect 15264 38268 15628 38312
rect 15264 38204 15308 38268
rect 15372 38204 15628 38268
rect 15264 38100 15628 38204
rect 16324 38100 16688 38312
rect 15264 38056 16688 38100
rect 15264 37992 15520 38056
rect 15584 37992 16688 38056
rect 15264 37948 16688 37992
rect 21200 38268 21352 38312
rect 21200 38204 21244 38268
rect 21308 38204 21352 38268
rect 21200 37888 21352 38204
rect 19928 37736 21352 37888
rect 19928 37676 20292 37736
rect 19928 37632 21352 37676
rect 19928 37568 21244 37632
rect 21308 37568 21352 37632
rect 19928 37524 21352 37568
rect 15264 36784 16264 36828
rect 15264 36720 16156 36784
rect 16220 36720 16264 36784
rect 15264 36676 16264 36720
rect 15264 36616 15628 36676
rect 16324 36616 16688 36828
rect 20216 36784 21352 36828
rect 20140 36720 20184 36784
rect 20248 36720 21352 36784
rect 20216 36676 21352 36720
rect 15264 36572 16688 36616
rect 15264 36508 16368 36572
rect 16432 36508 16688 36572
rect 15264 36464 16688 36508
rect 21200 36404 21352 36676
rect 19928 36252 21352 36404
rect 19928 36192 20292 36252
rect 19928 36148 21140 36192
rect 19928 36084 21032 36148
rect 21096 36084 21140 36148
rect 19928 36040 21140 36084
rect 15264 35300 15628 35344
rect 15264 35236 15520 35300
rect 15584 35236 15628 35300
rect 15264 35132 15628 35236
rect 16324 35132 16688 35344
rect 15264 35088 16688 35132
rect 15264 35024 15308 35088
rect 15372 35024 16688 35088
rect 15264 34980 16688 35024
rect 21200 35088 21352 35132
rect 21200 35024 21244 35088
rect 21308 35024 21352 35088
rect 21200 34920 21352 35024
rect 15552 34876 16476 34920
rect 15476 34812 15520 34876
rect 15584 34812 16368 34876
rect 16432 34812 16476 34876
rect 15552 34768 16476 34812
rect 19928 34768 21352 34920
rect 19928 34708 20292 34768
rect 19928 34664 21352 34708
rect 19928 34600 21244 34664
rect 21308 34600 21352 34664
rect 19928 34556 21352 34600
rect 15476 33708 16476 33860
rect 15476 33648 15628 33708
rect 16324 33648 16476 33708
rect 15264 33604 16264 33648
rect 15264 33540 15520 33604
rect 15584 33540 16156 33604
rect 16220 33540 16264 33604
rect 15264 33496 16264 33540
rect 16324 33496 16688 33648
rect 21064 33604 21352 33648
rect 20988 33540 21032 33604
rect 21096 33540 21352 33604
rect 21064 33496 21352 33540
rect 21200 33436 21352 33496
rect 19928 33284 21352 33436
rect 19928 33224 20292 33284
rect 19928 33180 21140 33224
rect 19928 33116 21032 33180
rect 21096 33116 21140 33180
rect 19928 33072 21140 33116
rect 15264 32120 15628 32164
rect 15264 32056 15308 32120
rect 15372 32056 15628 32120
rect 15264 31952 15628 32056
rect 16324 31952 16688 32164
rect 21200 32120 21352 32164
rect 21200 32056 21244 32120
rect 21308 32056 21352 32120
rect 21200 31952 21352 32056
rect 15264 31800 17112 31952
rect 16960 31740 17112 31800
rect 20140 31800 21352 31952
rect 20140 31740 20292 31800
rect 16960 31696 21352 31740
rect 16960 31632 21244 31696
rect 21308 31632 21352 31696
rect 16960 31588 21352 31632
rect 15264 30636 16688 30680
rect 21064 30636 21352 30680
rect 15264 30572 16368 30636
rect 16432 30572 16688 30636
rect 20988 30572 21032 30636
rect 21096 30572 21352 30636
rect 15264 30528 16688 30572
rect 21064 30528 21352 30572
rect 15264 30468 15628 30528
rect 15264 30424 16264 30468
rect 15264 30360 16156 30424
rect 16220 30360 16264 30424
rect 15264 30316 16264 30360
rect 16324 30316 16688 30528
rect 21200 30468 21352 30528
rect 20140 30316 21352 30468
rect 20140 30256 20292 30316
rect 19928 30212 21140 30256
rect 19928 30148 21032 30212
rect 21096 30148 21140 30212
rect 19928 30104 21140 30148
rect 21200 28940 21352 28984
rect 21200 28876 21244 28940
rect 21308 28876 21352 28940
rect 21200 28772 21352 28876
rect 19928 28728 21352 28772
rect 19928 28664 20184 28728
rect 20248 28664 21352 28728
rect 19928 28620 21352 28664
rect 15900 27560 16476 27712
rect 15900 27500 16052 27560
rect 16324 27500 16476 27560
rect 15688 27348 16052 27500
rect 16188 27456 16688 27500
rect 21064 27456 21352 27500
rect 16112 27392 16156 27456
rect 16220 27392 16688 27456
rect 20988 27392 21032 27456
rect 21096 27392 21352 27456
rect 16188 27348 16688 27392
rect 21064 27348 21352 27392
rect 15900 27288 16052 27348
rect 21200 27288 21352 27348
rect 15900 27244 16476 27288
rect 15900 27180 16368 27244
rect 16432 27180 16476 27244
rect 15900 27136 16476 27180
rect 19928 27136 21352 27288
rect 19928 27076 20292 27136
rect 19928 27032 21352 27076
rect 19928 26968 21244 27032
rect 21308 26968 21352 27032
rect 19928 26924 21352 26968
rect 15688 25864 16688 26016
rect 20216 25972 21352 26016
rect 20140 25908 20184 25972
rect 20248 25908 21352 25972
rect 20216 25864 21352 25908
rect 15688 25652 16052 25864
rect 16324 25804 16688 25864
rect 21200 25804 21352 25864
rect 16188 25760 16688 25804
rect 16112 25696 16156 25760
rect 16220 25696 16688 25760
rect 16188 25652 16688 25696
rect 19928 25652 21352 25804
rect 19928 25548 20292 25652
rect 19928 25484 19972 25548
rect 20036 25484 20292 25548
rect 19928 25440 20292 25484
rect 15688 24488 16688 24532
rect 15688 24424 16368 24488
rect 16432 24424 16688 24488
rect 15688 24380 16688 24424
rect 15688 24168 16052 24380
rect 16324 24276 16688 24380
rect 21200 24488 21352 24532
rect 21200 24424 21244 24488
rect 21308 24424 21352 24488
rect 21200 24320 21352 24424
rect 16324 24212 16368 24276
rect 16432 24212 16688 24276
rect 16324 24168 16688 24212
rect 19928 24276 21352 24320
rect 19928 24212 21244 24276
rect 21308 24212 21352 24276
rect 19928 24168 21352 24212
rect 19928 23956 20292 24168
rect 15900 22896 16476 23048
rect 15900 22836 16052 22896
rect 16324 22836 16476 22896
rect 15688 22792 16264 22836
rect 15688 22728 16156 22792
rect 16220 22728 16264 22792
rect 15688 22684 16264 22728
rect 16324 22684 17112 22836
rect 16960 22624 17112 22684
rect 19928 22792 21352 22836
rect 19928 22728 19972 22792
rect 20036 22728 21244 22792
rect 21308 22728 21352 22792
rect 19928 22684 21352 22728
rect 19928 22624 20292 22684
rect 16960 22472 20292 22624
rect 15900 21412 16476 21564
rect 15900 21352 16052 21412
rect 16324 21352 16476 21412
rect 15688 21308 16264 21352
rect 15688 21244 16156 21308
rect 16220 21244 16264 21308
rect 15688 21200 16264 21244
rect 16324 21308 16688 21352
rect 16324 21244 16368 21308
rect 16432 21244 16688 21308
rect 16324 21200 16688 21244
rect 20988 21308 21564 21352
rect 20988 21244 21032 21308
rect 21096 21244 21456 21308
rect 21520 21244 21564 21308
rect 20988 21200 21564 21244
rect 21200 21140 21352 21200
rect 19928 20988 21352 21140
rect 13568 19612 13932 19868
rect 21200 19824 21352 19868
rect 21200 19760 21244 19824
rect 21308 19760 21352 19824
rect 21200 19656 21352 19760
rect 13568 19548 13612 19612
rect 13676 19548 13932 19612
rect 13568 19504 13932 19548
rect 19928 19504 21352 19656
rect 20140 19444 20292 19504
rect 20140 19400 21352 19444
rect 20140 19336 21244 19400
rect 21308 19336 21352 19400
rect 20140 19292 21352 19336
rect 13568 18808 13932 19020
rect 13568 18764 15840 18808
rect 13568 18700 13824 18764
rect 13888 18700 15732 18764
rect 15796 18700 15840 18764
rect 13568 18656 15840 18700
rect 15688 18340 16052 18384
rect 16188 18340 16688 18384
rect 15688 18276 15732 18340
rect 15796 18276 16052 18340
rect 16112 18276 16156 18340
rect 16220 18276 16688 18340
rect 15688 18172 16052 18276
rect 16188 18232 16688 18276
rect 16324 18172 16688 18232
rect 21200 18340 21488 18384
rect 21200 18276 21456 18340
rect 21520 18276 21564 18340
rect 21200 18232 21488 18276
rect 21200 18172 21352 18232
rect 13568 18128 13932 18172
rect 13568 18064 13612 18128
rect 13676 18064 13932 18128
rect 13568 17960 13932 18064
rect 15688 18020 16688 18172
rect 19928 18128 21352 18172
rect 19928 18064 20184 18128
rect 20248 18064 21352 18128
rect 19928 18020 21352 18064
rect 13568 17916 15840 17960
rect 13568 17852 13612 17916
rect 13676 17852 15732 17916
rect 15796 17852 15840 17916
rect 13568 17808 15840 17852
rect 0 17452 13508 17536
rect 0 17396 13265 17452
rect 13321 17396 13508 17452
rect 0 17384 13508 17396
rect 14307 17450 14439 17453
rect 15061 17450 15193 17453
rect 14307 17448 15193 17450
rect 14307 17392 14345 17448
rect 14401 17392 15099 17448
rect 15155 17392 15193 17448
rect 14307 17390 15193 17392
rect 14307 17387 14439 17390
rect 15061 17387 15193 17390
rect 13780 17280 13932 17324
rect 13780 17216 13824 17280
rect 13888 17216 13932 17280
rect 13780 17211 13932 17216
rect 13761 17145 13932 17211
rect 13780 17112 13932 17145
rect 13144 16960 13508 17112
rect 13780 17068 14068 17112
rect 13780 17004 14036 17068
rect 14100 17004 14144 17068
rect 13780 16960 14068 17004
rect 14307 16966 14439 16969
rect 14993 16966 15125 16969
rect 14307 16964 15125 16966
rect 13144 16904 13265 16960
rect 13321 16904 13508 16960
rect 13144 16900 13508 16904
rect 14307 16908 14345 16964
rect 14401 16908 15031 16964
rect 15087 16908 15125 16964
rect 14307 16906 15125 16908
rect 14307 16903 14439 16906
rect 14993 16903 15125 16906
rect 0 16748 13508 16900
rect 15688 16644 16688 16688
rect 15688 16580 15732 16644
rect 15796 16580 16688 16644
rect 15688 16536 16688 16580
rect 19928 16644 21352 16688
rect 19928 16580 21244 16644
rect 21308 16580 21352 16644
rect 19928 16536 21352 16580
rect 13568 16432 13932 16476
rect 13568 16368 13612 16432
rect 13676 16368 13932 16432
rect 13568 16220 13932 16368
rect 19928 16432 20292 16536
rect 19928 16368 19972 16432
rect 20036 16368 20292 16432
rect 19928 16324 20292 16368
rect 13568 16156 13824 16220
rect 13888 16156 13932 16220
rect 13568 16112 13932 16156
rect 0 15776 13508 15840
rect 0 15720 13265 15776
rect 13321 15720 13508 15776
rect 0 15688 13508 15720
rect 14307 15774 14439 15777
rect 14925 15774 15057 15777
rect 14307 15772 15057 15774
rect 14307 15716 14345 15772
rect 14401 15716 14963 15772
rect 15019 15716 15057 15772
rect 14307 15714 15057 15716
rect 14307 15711 14439 15714
rect 14925 15711 15057 15714
rect 13780 15584 14144 15628
rect 13780 15535 14036 15584
rect 13761 15520 14036 15535
rect 14100 15520 14144 15584
rect 13761 15476 14144 15520
rect 13761 15469 13932 15476
rect 13780 15416 13932 15469
rect 0 15284 13508 15416
rect 0 15264 13265 15284
rect 13144 15228 13265 15264
rect 13321 15228 13508 15284
rect 13144 15052 13508 15228
rect 13780 15372 14068 15416
rect 20216 15372 21352 15416
rect 13780 15308 14036 15372
rect 14100 15308 14144 15372
rect 20140 15308 20184 15372
rect 20248 15308 21352 15372
rect 13780 15264 14068 15308
rect 14307 15290 14439 15293
rect 14857 15290 14989 15293
rect 14307 15288 14989 15290
rect 13780 15204 13932 15264
rect 14307 15232 14345 15288
rect 14401 15232 14895 15288
rect 14951 15232 14989 15288
rect 20216 15264 21352 15308
rect 14307 15230 14989 15232
rect 14307 15227 14439 15230
rect 14857 15227 14989 15230
rect 21200 15204 21352 15264
rect 13780 15052 14144 15204
rect 13992 14992 14144 15052
rect 15688 15052 16688 15204
rect 19928 15052 21352 15204
rect 15688 14992 15840 15052
rect 13992 14840 15840 14992
rect 19928 14992 20292 15052
rect 19928 14948 21352 14992
rect 19928 14884 21244 14948
rect 21308 14884 21352 14948
rect 19928 14840 21352 14884
rect 13568 14736 13932 14780
rect 13568 14672 13612 14736
rect 13676 14672 13824 14736
rect 13888 14672 13932 14736
rect 13568 14628 13932 14672
rect 0 14100 13508 14144
rect 0 14044 13265 14100
rect 13321 14044 13508 14100
rect 0 13992 13508 14044
rect 14307 14098 14439 14101
rect 14789 14098 14921 14101
rect 14307 14096 14921 14098
rect 14307 14040 14345 14096
rect 14401 14040 14827 14096
rect 14883 14040 14921 14096
rect 14307 14038 14921 14040
rect 14307 14035 14439 14038
rect 14789 14035 14921 14038
rect 13780 13888 14144 13932
rect 13780 13859 13824 13888
rect 13761 13824 13824 13859
rect 13888 13824 14036 13888
rect 14100 13824 14144 13888
rect 13761 13793 14144 13824
rect 13780 13780 14144 13793
rect 0 13608 13508 13720
rect 0 13568 13265 13608
rect 13144 13552 13265 13568
rect 13321 13552 13508 13608
rect 13144 13356 13508 13552
rect 14307 13614 14439 13617
rect 14721 13614 14853 13617
rect 14307 13612 14853 13614
rect 14307 13556 14345 13612
rect 14401 13556 14759 13612
rect 14815 13556 14853 13612
rect 14307 13554 14853 13556
rect 14307 13551 14439 13554
rect 14721 13551 14853 13554
rect 15688 13508 16052 13720
rect 16324 13508 16688 13720
rect 19928 13676 20292 13720
rect 19928 13612 19972 13676
rect 20036 13612 20292 13676
rect 19928 13508 20292 13612
rect 21200 13508 21352 13720
rect 15688 13464 17112 13508
rect 15688 13400 15732 13464
rect 15796 13400 17112 13464
rect 15688 13356 17112 13400
rect 16960 13296 17112 13356
rect 19928 13464 21988 13508
rect 19928 13400 21880 13464
rect 21944 13400 21988 13464
rect 19928 13356 21988 13400
rect 19928 13296 20080 13356
rect 16960 13144 20080 13296
rect 13568 13040 15840 13084
rect 13568 12976 13612 13040
rect 13676 12976 15732 13040
rect 15796 12976 15840 13040
rect 13568 12932 15840 12976
rect 12952 12486 13086 12491
rect 12952 12430 12990 12486
rect 13046 12430 13086 12486
rect 12952 12425 13086 12430
rect 13144 12429 13296 12448
rect 13356 12429 13508 12448
rect 13144 12424 13508 12429
rect 13144 12404 13265 12424
rect 13144 12340 13188 12404
rect 13252 12368 13265 12404
rect 13321 12368 13508 12424
rect 13252 12363 13508 12368
rect 13252 12340 13296 12363
rect 13144 12296 13296 12340
rect 13356 12296 13508 12363
rect 14307 12422 14439 12425
rect 14653 12422 14785 12425
rect 14307 12420 14785 12422
rect 14307 12364 14345 12420
rect 14401 12364 14691 12420
rect 14747 12364 14785 12420
rect 14307 12362 14785 12364
rect 14307 12359 14439 12362
rect 14653 12359 14785 12362
rect 13780 12192 16688 12236
rect 13780 12183 13824 12192
rect 13761 12128 13824 12183
rect 13888 12128 16688 12192
rect 13761 12117 16688 12128
rect 13780 12084 16688 12117
rect 15688 11872 16052 12084
rect 16324 12024 16688 12084
rect 19928 12192 21352 12236
rect 19928 12128 21244 12192
rect 21308 12128 21352 12192
rect 19928 12084 21352 12128
rect 16324 11980 17112 12024
rect 16324 11916 17004 11980
rect 17068 11916 17112 11980
rect 16324 11872 17112 11916
rect 19928 11980 20292 12084
rect 19928 11916 19972 11980
rect 20036 11916 20292 11980
rect 19928 11872 20292 11916
rect 21200 12024 21352 12084
rect 21200 11872 21988 12024
rect 21836 11812 21988 11872
rect 24804 11812 25168 12024
rect 27984 11812 28348 12024
rect 31164 11812 31316 12024
rect 34132 11812 34496 12024
rect 37312 11812 37676 12024
rect 40492 11812 40644 12024
rect 43460 11812 43824 12024
rect 46640 11812 47004 12024
rect 49820 11812 49972 12024
rect 52788 11812 53152 12024
rect 55968 11812 56332 12024
rect 59148 11812 59300 12024
rect 62328 11812 62480 12024
rect 65296 11812 65660 12024
rect 68476 11812 68628 12024
rect 21836 11768 22412 11812
rect 21836 11704 22304 11768
rect 22368 11704 22412 11768
rect 21836 11660 22412 11704
rect 24804 11768 25380 11812
rect 24804 11704 25272 11768
rect 25336 11704 25380 11768
rect 24804 11660 25380 11704
rect 27984 11768 28560 11812
rect 27984 11704 28452 11768
rect 28516 11704 28560 11768
rect 27984 11660 28560 11704
rect 31164 11768 31528 11812
rect 31164 11704 31420 11768
rect 31484 11704 31528 11768
rect 31164 11660 31528 11704
rect 34132 11768 34708 11812
rect 34132 11704 34600 11768
rect 34664 11704 34708 11768
rect 34132 11660 34708 11704
rect 37312 11768 38100 11812
rect 37312 11704 37992 11768
rect 38056 11704 38100 11768
rect 37312 11660 38100 11704
rect 40492 11768 40856 11812
rect 40492 11704 40748 11768
rect 40812 11704 40856 11768
rect 40492 11660 40856 11704
rect 43460 11768 44036 11812
rect 43460 11704 43928 11768
rect 43992 11704 44036 11768
rect 43460 11660 44036 11704
rect 46640 11768 47216 11812
rect 46640 11704 47108 11768
rect 47172 11704 47216 11768
rect 46640 11660 47216 11704
rect 49820 11768 50608 11812
rect 49820 11704 50500 11768
rect 50564 11704 50608 11768
rect 49820 11660 50608 11704
rect 52788 11768 53364 11812
rect 52788 11704 53256 11768
rect 53320 11704 53364 11768
rect 52788 11660 53364 11704
rect 55968 11768 56968 11812
rect 55968 11704 56860 11768
rect 56924 11704 56968 11768
rect 55968 11660 56968 11704
rect 59148 11768 59724 11812
rect 59148 11704 59616 11768
rect 59680 11704 59724 11768
rect 59148 11660 59724 11704
rect 62328 11768 62692 11812
rect 62328 11704 62584 11768
rect 62648 11704 62692 11768
rect 62328 11660 62692 11704
rect 65296 11768 65872 11812
rect 65296 11704 65764 11768
rect 65828 11704 65872 11768
rect 65296 11660 65872 11704
rect 68476 11768 68840 11812
rect 68476 11704 68732 11768
rect 68796 11704 68840 11768
rect 68476 11660 68840 11704
rect 14502 11547 14634 11550
rect 20016 11547 20148 11550
rect 14502 11545 20148 11547
rect 14502 11489 14540 11545
rect 14596 11489 20054 11545
rect 20110 11489 20148 11545
rect 14502 11487 20148 11489
rect 14502 11484 14634 11487
rect 20016 11484 20148 11487
rect 49684 11344 50396 11388
rect 55832 11344 56544 11388
rect 49608 11280 49652 11344
rect 49716 11280 50288 11344
rect 50352 11280 50396 11344
rect 55756 11280 55800 11344
rect 55864 11280 56436 11344
rect 56500 11280 56544 11344
rect 49684 11236 50396 11280
rect 55832 11236 56544 11280
rect 17036 11132 18172 11176
rect 16960 11068 17004 11132
rect 17068 11068 18172 11132
rect 17036 11024 18172 11068
rect 17808 10964 18172 11024
rect 18868 11132 20080 11176
rect 18868 11068 19972 11132
rect 20036 11068 20080 11132
rect 18868 11024 20080 11068
rect 21836 11132 22200 11176
rect 21836 11068 21880 11132
rect 21944 11068 22092 11132
rect 22156 11068 22200 11132
rect 21836 11024 22200 11068
rect 18868 10964 19232 11024
rect 17808 10920 19232 10964
rect 17808 10856 18064 10920
rect 18128 10856 19232 10920
rect 17808 10812 19232 10856
rect 21836 10920 21988 11024
rect 21836 10856 21880 10920
rect 21944 10856 21988 10920
rect 21836 10812 21988 10856
rect 22048 10920 23048 10964
rect 22048 10856 22304 10920
rect 22368 10856 22940 10920
rect 23004 10856 23048 10920
rect 22048 10812 23048 10856
rect 24804 10920 25168 11176
rect 27984 11132 28348 11176
rect 27984 11068 28240 11132
rect 28304 11068 28348 11132
rect 27984 11024 28348 11068
rect 28408 11068 28452 11132
rect 28516 11068 28560 11132
rect 27984 11006 28168 11024
rect 24804 10856 24848 10920
rect 24912 10856 25060 10920
rect 25124 10856 25168 10920
rect 24804 10812 25168 10856
rect 25228 10920 26016 10964
rect 25228 10856 25272 10920
rect 25336 10856 25908 10920
rect 25972 10856 26016 10920
rect 25228 10812 26016 10856
rect 27984 10920 28136 11006
rect 28408 10964 28560 11068
rect 31164 10964 31316 11176
rect 34132 11132 34920 11176
rect 34132 11068 34812 11132
rect 34876 11068 34920 11132
rect 34132 11024 34920 11068
rect 37312 11132 37888 11176
rect 37312 11068 37780 11132
rect 37844 11068 37888 11132
rect 37312 11024 37888 11068
rect 27984 10856 28028 10920
rect 28092 10856 28136 10920
rect 27984 10812 28136 10856
rect 28196 10920 28560 10964
rect 28196 10856 28452 10920
rect 28516 10856 28560 10920
rect 28196 10812 28560 10856
rect 30952 10920 31316 10964
rect 30952 10856 30996 10920
rect 31060 10856 31208 10920
rect 31272 10856 31316 10920
rect 30952 10812 31316 10856
rect 31376 10920 32376 10964
rect 31376 10856 31420 10920
rect 31484 10856 32268 10920
rect 32332 10856 32376 10920
rect 31376 10812 32376 10856
rect 34132 10920 34496 11024
rect 34132 10856 34176 10920
rect 34240 10856 34496 10920
rect 34132 10812 34496 10856
rect 34556 10920 35056 10964
rect 37312 10920 37676 11024
rect 40492 10964 40644 11176
rect 43460 11132 44248 11176
rect 43460 11068 44140 11132
rect 44204 11068 44248 11132
rect 43460 11024 44248 11068
rect 34556 10856 34600 10920
rect 34664 10856 35024 10920
rect 35088 10856 35132 10920
rect 37312 10856 37356 10920
rect 37420 10856 37676 10920
rect 34556 10812 35056 10856
rect 37312 10812 37676 10856
rect 37736 10920 38736 10964
rect 37736 10856 37992 10920
rect 38056 10856 38628 10920
rect 38692 10856 38736 10920
rect 37736 10812 38736 10856
rect 40280 10920 40644 10964
rect 40280 10856 40324 10920
rect 40388 10856 40536 10920
rect 40600 10856 40644 10920
rect 40280 10812 40644 10856
rect 40704 10920 41280 10964
rect 40704 10856 40748 10920
rect 40812 10856 41172 10920
rect 41236 10856 41280 10920
rect 40704 10812 41280 10856
rect 43460 10920 43824 11024
rect 46640 10964 47004 11176
rect 49820 11132 50184 11176
rect 49820 11068 50076 11132
rect 50140 11068 50184 11132
rect 49820 11024 50184 11068
rect 43460 10856 43504 10920
rect 43568 10856 43824 10920
rect 43460 10812 43824 10856
rect 43884 10920 44884 10964
rect 43884 10856 43928 10920
rect 43992 10856 44776 10920
rect 44840 10856 44884 10920
rect 43884 10812 44884 10856
rect 46428 10920 47004 10964
rect 46428 10856 46472 10920
rect 46536 10856 46684 10920
rect 46748 10856 47004 10920
rect 46428 10812 47004 10856
rect 47064 10920 47640 10964
rect 47064 10856 47108 10920
rect 47172 10856 47532 10920
rect 47596 10856 47640 10920
rect 47064 10812 47640 10856
rect 49820 10920 49972 11024
rect 49820 10856 49864 10920
rect 49928 10856 49972 10920
rect 49820 10812 49972 10856
rect 50032 10920 50532 10964
rect 52788 10920 53152 11176
rect 55968 11132 56756 11176
rect 55968 11068 56648 11132
rect 56712 11068 56756 11132
rect 55968 11024 56756 11068
rect 59148 11132 59512 11176
rect 59148 11068 59404 11132
rect 59468 11068 59512 11132
rect 59148 11024 59512 11068
rect 62328 11132 62904 11176
rect 62328 11068 62796 11132
rect 62860 11068 62904 11132
rect 62328 11024 62904 11068
rect 65296 11132 66084 11176
rect 65296 11068 65976 11132
rect 66040 11068 66084 11132
rect 65296 11024 66084 11068
rect 50032 10856 50288 10920
rect 50352 10856 50500 10920
rect 50564 10856 50608 10920
rect 52788 10856 52832 10920
rect 52896 10856 53044 10920
rect 53108 10856 53152 10920
rect 50032 10812 50532 10856
rect 52788 10812 53152 10856
rect 53212 10920 53576 10964
rect 53212 10856 53256 10920
rect 53320 10856 53468 10920
rect 53532 10856 53576 10920
rect 53212 10812 53576 10856
rect 55968 10920 56332 11024
rect 55968 10856 56012 10920
rect 56076 10856 56332 10920
rect 55968 10812 56332 10856
rect 56392 10920 56892 10964
rect 56392 10856 56436 10920
rect 56500 10856 56860 10920
rect 56924 10856 56968 10920
rect 56392 10812 56892 10856
rect 59148 10812 59300 11024
rect 62328 10964 62480 11024
rect 59360 10920 60148 10964
rect 62192 10920 62480 10964
rect 59360 10856 59616 10920
rect 59680 10856 60040 10920
rect 60104 10856 60148 10920
rect 62116 10856 62160 10920
rect 62224 10856 62480 10920
rect 59360 10812 60148 10856
rect 62192 10812 62480 10856
rect 62540 10920 63116 10964
rect 62540 10856 62584 10920
rect 62648 10856 63008 10920
rect 63072 10856 63116 10920
rect 62540 10812 63116 10856
rect 65296 10920 65660 11024
rect 68476 10964 68628 11176
rect 65296 10856 65340 10920
rect 65404 10856 65660 10920
rect 65296 10812 65660 10856
rect 65720 10920 66720 10964
rect 65720 10856 65764 10920
rect 65828 10856 66612 10920
rect 66676 10856 66720 10920
rect 65720 10812 66720 10856
rect 68264 10920 68628 10964
rect 68264 10856 68308 10920
rect 68372 10856 68520 10920
rect 68584 10856 68628 10920
rect 68264 10812 68628 10856
rect 68688 10920 69188 10964
rect 68688 10856 68732 10920
rect 68796 10856 69156 10920
rect 69220 10856 69264 10920
rect 68688 10812 69188 10856
rect 22180 10752 22312 10812
rect 25292 10752 25424 10812
rect 28404 10752 28536 10812
rect 31516 10752 31648 10812
rect 34628 10752 34760 10812
rect 37740 10752 37872 10812
rect 40852 10752 40984 10812
rect 43964 10752 44096 10812
rect 47076 10752 47208 10812
rect 50188 10752 50320 10812
rect 53300 10752 53432 10812
rect 56412 10752 56544 10812
rect 59524 10752 59656 10812
rect 62636 10752 62768 10812
rect 65748 10752 65880 10812
rect 68860 10752 68992 10812
rect 71868 10752 72232 10964
rect 75048 10752 75412 10964
rect 78016 10812 84740 10964
rect 78016 10752 78380 10812
rect 22180 10723 22412 10752
rect 22260 10708 22412 10723
rect 22260 10698 22304 10708
rect 22260 10642 22298 10698
rect 22368 10644 22412 10708
rect 22354 10642 22412 10644
rect 14502 10614 14634 10617
rect 22260 10614 22412 10642
rect 25228 10723 25424 10752
rect 25228 10703 25380 10723
rect 25440 10708 25592 10752
rect 28404 10723 28560 10752
rect 25440 10703 25484 10708
rect 25228 10698 25484 10703
rect 25228 10642 25410 10698
rect 25466 10644 25484 10698
rect 25548 10644 25592 10708
rect 25466 10642 25592 10644
rect 25228 10637 25592 10642
rect 25228 10614 25380 10637
rect 25440 10614 25592 10637
rect 28408 10703 28560 10723
rect 28620 10708 28772 10752
rect 31516 10723 31740 10752
rect 28620 10703 28664 10708
rect 28408 10698 28664 10703
rect 28408 10642 28522 10698
rect 28578 10644 28664 10698
rect 28728 10644 28772 10708
rect 28578 10642 28772 10644
rect 28408 10637 28772 10642
rect 28408 10614 28560 10637
rect 28620 10614 28772 10637
rect 31588 10708 31740 10723
rect 31588 10644 31632 10708
rect 31696 10644 31740 10708
rect 31588 10642 31634 10644
rect 31690 10642 31740 10644
rect 31588 10614 31740 10642
rect 34556 10723 34760 10752
rect 34556 10708 34708 10723
rect 34556 10644 34600 10708
rect 34664 10703 34708 10708
rect 34768 10703 34920 10752
rect 34664 10698 34920 10703
rect 34664 10644 34746 10698
rect 34556 10642 34746 10644
rect 34802 10642 34920 10698
rect 34556 10637 34920 10642
rect 34556 10614 34708 10637
rect 34768 10614 34920 10637
rect 37736 10703 37888 10752
rect 37948 10708 38100 10752
rect 40852 10723 41068 10752
rect 37948 10703 37992 10708
rect 37736 10698 37992 10703
rect 37736 10642 37858 10698
rect 37914 10644 37992 10698
rect 38056 10644 38100 10708
rect 37914 10642 38100 10644
rect 37736 10637 38100 10642
rect 37736 10614 37888 10637
rect 37948 10614 38100 10637
rect 40916 10708 41068 10723
rect 40916 10644 40960 10708
rect 41024 10698 41068 10708
rect 40916 10642 40970 10644
rect 41026 10642 41068 10698
rect 40916 10614 41068 10642
rect 43884 10723 44248 10752
rect 43884 10708 44036 10723
rect 43884 10644 43928 10708
rect 43992 10703 44036 10708
rect 44096 10703 44248 10723
rect 43992 10698 44248 10703
rect 43992 10644 44082 10698
rect 43884 10642 44082 10644
rect 44138 10642 44248 10698
rect 43884 10637 44248 10642
rect 43884 10614 44036 10637
rect 44096 10614 44248 10637
rect 47064 10708 47216 10752
rect 47064 10644 47108 10708
rect 47172 10703 47216 10708
rect 47276 10703 47428 10752
rect 50188 10723 50396 10752
rect 47172 10698 47428 10703
rect 47172 10644 47194 10698
rect 47064 10642 47194 10644
rect 47250 10642 47428 10698
rect 47064 10637 47428 10642
rect 47064 10614 47216 10637
rect 47276 10614 47428 10637
rect 50244 10703 50396 10723
rect 50456 10708 50608 10752
rect 50456 10703 50500 10708
rect 50244 10698 50500 10703
rect 50244 10642 50306 10698
rect 50362 10644 50500 10698
rect 50564 10644 50608 10708
rect 50362 10642 50608 10644
rect 50244 10637 50608 10642
rect 50244 10614 50396 10637
rect 50456 10614 50608 10637
rect 53212 10723 53576 10752
rect 53212 10708 53364 10723
rect 53212 10644 53256 10708
rect 53320 10703 53364 10708
rect 53424 10703 53576 10723
rect 53320 10698 53576 10703
rect 53320 10644 53418 10698
rect 53212 10642 53418 10644
rect 53474 10642 53576 10698
rect 53212 10637 53576 10642
rect 53212 10614 53364 10637
rect 53424 10614 53576 10637
rect 56392 10708 56544 10752
rect 56392 10644 56436 10708
rect 56500 10703 56544 10708
rect 56604 10703 56756 10752
rect 59524 10723 59724 10752
rect 56500 10698 56756 10703
rect 56500 10644 56530 10698
rect 56392 10642 56530 10644
rect 56586 10642 56756 10698
rect 56392 10637 56756 10642
rect 56392 10614 56544 10637
rect 56604 10614 56756 10637
rect 59572 10703 59724 10723
rect 59784 10708 59936 10752
rect 59784 10703 59828 10708
rect 59572 10698 59828 10703
rect 59572 10642 59642 10698
rect 59698 10644 59828 10698
rect 59892 10644 59936 10708
rect 59698 10642 59936 10644
rect 59572 10637 59936 10642
rect 59572 10614 59724 10637
rect 59784 10614 59936 10637
rect 62540 10723 62904 10752
rect 62540 10708 62692 10723
rect 62540 10644 62584 10708
rect 62648 10703 62692 10708
rect 62752 10703 62904 10723
rect 62648 10698 62904 10703
rect 62648 10644 62754 10698
rect 62540 10642 62754 10644
rect 62810 10642 62904 10698
rect 62540 10637 62904 10642
rect 62540 10614 62692 10637
rect 62752 10614 62904 10637
rect 65720 10723 65880 10752
rect 65720 10708 65872 10723
rect 65720 10644 65764 10708
rect 65828 10703 65872 10708
rect 65932 10703 66084 10752
rect 68860 10723 69052 10752
rect 65828 10698 66084 10703
rect 65828 10644 65866 10698
rect 65720 10642 65866 10644
rect 65922 10642 66084 10698
rect 65720 10637 66084 10642
rect 65720 10614 65872 10637
rect 65932 10614 66084 10637
rect 68900 10708 69052 10723
rect 68900 10644 68944 10708
rect 69008 10703 69052 10708
rect 69112 10703 69264 10752
rect 69008 10698 69264 10703
rect 68900 10642 68978 10644
rect 69034 10642 69264 10698
rect 68900 10637 69264 10642
rect 68900 10614 69052 10637
rect 69112 10614 69264 10637
rect 71868 10708 78380 10752
rect 71868 10644 71912 10708
rect 71976 10644 78380 10708
rect 71612 10614 71744 10617
rect 14502 10612 71744 10614
rect 14502 10556 14540 10612
rect 14596 10556 71650 10612
rect 71706 10556 71744 10612
rect 71868 10600 78380 10644
rect 81196 10600 81560 10812
rect 84376 10752 84740 10812
rect 87344 10812 94068 10964
rect 87344 10752 87708 10812
rect 84376 10600 87708 10752
rect 90524 10600 90888 10812
rect 93704 10752 94068 10812
rect 96672 10812 115692 10964
rect 96672 10752 97036 10812
rect 93704 10600 97036 10752
rect 99852 10600 100216 10812
rect 103032 10600 103396 10812
rect 106000 10600 106364 10812
rect 109180 10600 109544 10812
rect 112360 10600 112724 10812
rect 115328 10600 115692 10812
rect 118508 10920 120780 10964
rect 118508 10856 120672 10920
rect 120736 10856 120780 10920
rect 118508 10812 120780 10856
rect 118508 10600 118872 10812
rect 14502 10554 71744 10556
rect 14502 10551 14634 10554
rect 71612 10551 71744 10554
rect 17808 10284 21988 10328
rect 17808 10220 21880 10284
rect 21944 10220 21988 10284
rect 17808 10176 21988 10220
rect 17808 9964 18172 10176
rect 18868 10072 19232 10176
rect 31028 10072 31528 10116
rect 40356 10072 40856 10116
rect 46504 10072 47216 10116
rect 68340 10072 68840 10116
rect 18868 10008 18912 10072
rect 18976 10008 19232 10072
rect 30952 10008 30996 10072
rect 31060 10008 31528 10072
rect 40280 10008 40324 10072
rect 40388 10008 40856 10072
rect 46428 10008 46472 10072
rect 46536 10008 47216 10072
rect 68264 10008 68308 10072
rect 68372 10008 68840 10072
rect 18868 9964 19232 10008
rect 31028 9964 31528 10008
rect 40356 9964 40856 10008
rect 46504 9964 47216 10008
rect 68340 9964 68840 10008
rect 31376 9904 31528 9964
rect 40704 9904 40856 9964
rect 47064 9904 47216 9964
rect 68688 9904 68840 9964
rect 14502 9873 14634 9876
rect 21138 9873 21270 9876
rect 14502 9871 21270 9873
rect 14502 9815 14540 9871
rect 14596 9815 21176 9871
rect 21232 9815 21270 9871
rect 14502 9813 21270 9815
rect 14502 9810 14634 9813
rect 21138 9810 21270 9813
rect 22048 9860 24956 9904
rect 25092 9860 28136 9904
rect 22048 9796 22092 9860
rect 22156 9796 24848 9860
rect 24912 9796 24956 9860
rect 25016 9796 25060 9860
rect 25124 9796 28028 9860
rect 28092 9796 28136 9860
rect 22048 9752 24956 9796
rect 25092 9752 28136 9796
rect 28196 9860 31316 9904
rect 28196 9796 28240 9860
rect 28304 9796 31208 9860
rect 31272 9796 31316 9860
rect 28196 9752 31316 9796
rect 31376 9860 34284 9904
rect 31376 9796 34176 9860
rect 34240 9796 34284 9860
rect 31376 9752 34284 9796
rect 34556 9860 37464 9904
rect 34556 9796 34812 9860
rect 34876 9796 37356 9860
rect 37420 9796 37464 9860
rect 34556 9752 37464 9796
rect 37736 9860 40644 9904
rect 37736 9796 37780 9860
rect 37844 9796 40536 9860
rect 40600 9796 40644 9860
rect 37736 9752 40644 9796
rect 40704 9860 43612 9904
rect 40704 9796 43504 9860
rect 43568 9796 43612 9860
rect 40704 9752 43612 9796
rect 43884 9860 46792 9904
rect 43884 9796 44140 9860
rect 44204 9796 46684 9860
rect 46748 9796 46792 9860
rect 43884 9752 46792 9796
rect 47064 9860 49972 9904
rect 47064 9796 49864 9860
rect 49928 9796 49972 9860
rect 47064 9752 49972 9796
rect 50032 9860 52940 9904
rect 53076 9860 56120 9904
rect 50032 9796 50076 9860
rect 50140 9796 52832 9860
rect 52896 9796 52940 9860
rect 53000 9796 53044 9860
rect 53108 9796 56012 9860
rect 56076 9796 56120 9860
rect 50032 9752 52940 9796
rect 53076 9752 56120 9796
rect 56392 9860 62268 9904
rect 56392 9796 56648 9860
rect 56712 9796 59404 9860
rect 59468 9796 62160 9860
rect 62224 9796 62268 9860
rect 56392 9752 62268 9796
rect 62540 9860 65448 9904
rect 62540 9796 62796 9860
rect 62860 9796 65340 9860
rect 65404 9796 65448 9860
rect 62540 9752 65448 9796
rect 65720 9860 68628 9904
rect 65720 9796 65976 9860
rect 66040 9796 68520 9860
rect 68584 9796 68628 9860
rect 65720 9752 68628 9796
rect 68688 9752 100216 9904
rect 103032 9860 119720 9904
rect 103032 9796 119612 9860
rect 119676 9796 119720 9860
rect 103032 9752 119720 9796
rect 17808 9436 18172 9480
rect 17808 9372 18064 9436
rect 18128 9372 18172 9436
rect 17808 9268 18172 9372
rect 18868 9268 19232 9480
rect 17808 9224 19232 9268
rect 17808 9160 19124 9224
rect 19188 9160 19232 9224
rect 17808 9116 19232 9160
rect 17808 8588 19232 8632
rect 17808 8524 18912 8588
rect 18976 8524 19232 8588
rect 17808 8480 19232 8524
rect 17808 8268 18172 8480
rect 18868 8268 19232 8480
rect 25440 8480 26228 8632
rect 25440 8420 25592 8480
rect 26076 8420 26228 8480
rect 27772 8480 28560 8632
rect 27772 8420 27924 8480
rect 28408 8420 28560 8480
rect 34344 8588 35132 8632
rect 34344 8524 35024 8588
rect 35088 8524 35132 8588
rect 34344 8480 35132 8524
rect 47276 8480 48064 8632
rect 34344 8420 34496 8480
rect 47276 8420 47428 8480
rect 47912 8420 48064 8480
rect 53000 8588 53576 8632
rect 53000 8524 53468 8588
rect 53532 8524 53576 8588
rect 53000 8480 53576 8524
rect 59784 8480 60360 8632
rect 53000 8420 53152 8480
rect 59784 8420 59936 8480
rect 60208 8420 60360 8480
rect 62752 8480 63540 8632
rect 62752 8420 62904 8480
rect 63388 8420 63540 8480
rect 68688 8588 69264 8632
rect 68688 8524 69156 8588
rect 69220 8524 69264 8588
rect 68688 8480 69264 8524
rect 68688 8420 68840 8480
rect 22260 8376 25940 8420
rect 26076 8376 28348 8420
rect 22260 8312 22940 8376
rect 23004 8312 25908 8376
rect 25972 8312 26016 8376
rect 26076 8312 28240 8376
rect 28304 8312 28348 8376
rect 22260 8268 25940 8312
rect 26076 8268 28348 8312
rect 28408 8376 34496 8420
rect 28408 8312 32268 8376
rect 32332 8312 34496 8376
rect 28408 8268 34496 8312
rect 34556 8376 47564 8420
rect 47912 8376 53152 8420
rect 34556 8312 38628 8376
rect 38692 8312 41172 8376
rect 41236 8312 44776 8376
rect 44840 8312 47532 8376
rect 47596 8312 47640 8376
rect 47912 8312 49652 8376
rect 49716 8312 53152 8376
rect 34556 8268 47564 8312
rect 47912 8268 53152 8312
rect 53212 8376 60072 8420
rect 60208 8376 63040 8420
rect 63388 8376 68840 8420
rect 53212 8312 55800 8376
rect 55864 8312 60040 8376
rect 60104 8312 60148 8376
rect 60208 8312 63008 8376
rect 63072 8312 63116 8376
rect 63388 8312 66612 8376
rect 66676 8312 68840 8376
rect 53212 8268 60072 8312
rect 60208 8268 63040 8312
rect 63388 8268 68840 8312
rect 68900 8376 72020 8420
rect 68900 8312 71912 8376
rect 71976 8312 72020 8376
rect 68900 8268 72020 8312
rect 34132 8208 34284 8268
rect 34556 8208 34708 8268
rect 34132 8056 34708 8208
rect 52788 8208 52940 8268
rect 53212 8208 53364 8268
rect 52788 8056 53364 8208
rect 68264 8208 68416 8268
rect 68900 8208 69052 8268
rect 68264 8056 69052 8208
rect 848 7740 2908 7784
rect 848 7676 892 7740
rect 956 7676 2588 7740
rect 2652 7676 2908 7740
rect 848 7632 2908 7676
rect 17808 7572 18172 7784
rect 18868 7740 19232 7784
rect 18868 7676 19124 7740
rect 19188 7676 19232 7740
rect 18868 7572 19232 7676
rect 2825 7482 2957 7487
rect 2825 7426 2863 7482
rect 2919 7426 2957 7482
rect 2825 7421 2957 7426
rect 17808 7420 19232 7572
rect 6148 7267 6512 7360
rect 6148 7211 6223 7267
rect 6279 7211 6512 7267
rect 6148 7104 6512 7211
rect 6148 7040 6192 7104
rect 6256 7040 6512 7104
rect 6148 6996 6512 7040
rect 1908 6892 2908 6936
rect 1908 6828 1952 6892
rect 2016 6828 2908 6892
rect 1908 6784 2908 6828
rect 21624 6572 24320 6724
rect 21624 6360 21988 6572
rect 22472 6360 22624 6572
rect 23108 6360 23472 6572
rect 23956 6512 24320 6572
rect 24804 6512 24956 6724
rect 25440 6572 26652 6724
rect 25440 6512 25804 6572
rect 23956 6360 25804 6512
rect 26288 6512 26652 6572
rect 27136 6512 27288 6724
rect 27772 6512 28136 6724
rect 28620 6512 28984 6724
rect 29468 6512 29620 6724
rect 30104 6512 30468 6724
rect 30952 6512 31316 6724
rect 31800 6572 32800 6724
rect 31800 6512 31952 6572
rect 26288 6468 31952 6512
rect 26288 6404 28876 6468
rect 28940 6404 31952 6468
rect 26288 6360 31952 6404
rect 32436 6512 32800 6572
rect 33284 6572 34284 6724
rect 33284 6512 33648 6572
rect 32436 6360 33648 6512
rect 34132 6512 34284 6572
rect 34768 6512 35132 6724
rect 35616 6572 36616 6724
rect 35616 6512 35980 6572
rect 34132 6360 35980 6512
rect 36464 6512 36616 6572
rect 37100 6512 37464 6724
rect 37948 6572 38948 6724
rect 37948 6512 38312 6572
rect 36464 6360 38312 6512
rect 38796 6512 38948 6572
rect 39432 6572 40644 6724
rect 39432 6512 39796 6572
rect 38796 6360 39796 6512
rect 40280 6512 40644 6572
rect 41128 6572 42976 6724
rect 41128 6512 41280 6572
rect 40280 6360 41280 6512
rect 41764 6360 42128 6572
rect 42612 6512 42976 6572
rect 43460 6512 43612 6724
rect 44096 6572 45308 6724
rect 44096 6512 44460 6572
rect 42612 6360 44460 6512
rect 44944 6512 45308 6572
rect 45792 6512 45944 6724
rect 46428 6512 46792 6724
rect 47276 6512 47640 6724
rect 48124 6512 48276 6724
rect 48760 6512 49124 6724
rect 49608 6572 51456 6724
rect 49608 6512 49972 6572
rect 44944 6360 49972 6512
rect 50456 6360 50608 6572
rect 51092 6512 51456 6572
rect 51940 6572 52940 6724
rect 51940 6512 52304 6572
rect 51092 6360 52304 6512
rect 52788 6512 52940 6572
rect 53424 6572 55272 6724
rect 53424 6512 53788 6572
rect 52788 6360 53788 6512
rect 54272 6360 54636 6572
rect 55120 6512 55272 6572
rect 55756 6512 56120 6724
rect 56604 6512 56968 6724
rect 57452 6512 57604 6724
rect 58088 6512 58452 6724
rect 58936 6512 59300 6724
rect 59784 6572 60784 6724
rect 59784 6512 59936 6572
rect 55120 6360 59936 6512
rect 60420 6512 60784 6572
rect 61268 6512 61632 6724
rect 62116 6572 63964 6724
rect 62116 6512 62268 6572
rect 60420 6360 62268 6512
rect 62752 6360 63116 6572
rect 63600 6512 63964 6572
rect 64448 6512 64600 6724
rect 65084 6512 65448 6724
rect 65932 6512 66296 6724
rect 66780 6512 66932 6724
rect 67416 6572 68628 6724
rect 67416 6512 67780 6572
rect 63600 6360 67780 6512
rect 68264 6512 68628 6572
rect 69112 6572 70112 6724
rect 69112 6512 69264 6572
rect 68264 6360 69264 6512
rect 69748 6512 70112 6572
rect 70596 6572 71596 6724
rect 70596 6512 70960 6572
rect 69748 6360 70960 6512
rect 71444 6360 71596 6572
rect 2825 6298 2957 6303
rect 2825 6242 2863 6298
rect 2919 6242 2957 6298
rect 2825 6237 2957 6242
rect 2544 6044 2908 6088
rect 2544 5980 2588 6044
rect 2652 5980 2908 6044
rect 2544 5936 2908 5980
rect 16536 3544 16900 3756
rect 18020 3544 18384 3756
rect 16536 3500 18384 3544
rect 16536 3436 18064 3500
rect 18128 3436 18384 3500
rect 16536 3392 18384 3436
rect 19504 3544 19868 3756
rect 20988 3544 21352 3756
rect 22472 3604 24320 3756
rect 22472 3544 22836 3604
rect 19504 3392 22836 3544
rect 23956 3544 24320 3604
rect 25440 3544 25804 3756
rect 26924 3544 27288 3756
rect 23956 3500 27288 3544
rect 23956 3436 24212 3500
rect 24276 3436 27288 3500
rect 23956 3392 27288 3436
rect 28408 3712 28984 3756
rect 28408 3648 28876 3712
rect 28940 3648 28984 3712
rect 28408 3604 28984 3648
rect 28408 3544 28772 3604
rect 29892 3544 30256 3756
rect 31376 3544 31740 3756
rect 32860 3544 33224 3756
rect 34344 3544 34708 3756
rect 28408 3500 34708 3544
rect 28408 3436 30148 3500
rect 30212 3436 34708 3500
rect 28408 3392 34708 3436
rect 35828 3604 37676 3756
rect 35828 3392 36192 3604
rect 37312 3500 37676 3604
rect 37312 3436 37356 3500
rect 37420 3436 37676 3500
rect 37312 3392 37676 3436
rect 38796 3544 39160 3756
rect 40280 3604 42128 3756
rect 40280 3544 40644 3604
rect 38796 3500 40644 3544
rect 38796 3436 40324 3500
rect 40388 3436 40644 3500
rect 38796 3392 40644 3436
rect 41764 3392 42128 3604
rect 12952 3040 13084 3043
rect 12952 3038 30870 3040
rect 12952 2982 12990 3038
rect 13046 2982 30870 3038
rect 12952 2980 30870 2982
rect 12952 2977 13084 2980
rect 16191 2976 16323 2980
rect 16191 2920 16229 2976
rect 16285 2920 16323 2976
rect 16191 2908 16323 2920
rect 17673 2976 17805 2980
rect 17673 2920 17711 2976
rect 17767 2920 17805 2976
rect 17673 2908 17805 2920
rect 19155 2976 19287 2980
rect 19155 2920 19193 2976
rect 19249 2920 19287 2976
rect 19155 2908 19287 2920
rect 20637 2976 20769 2980
rect 20637 2920 20675 2976
rect 20731 2920 20769 2976
rect 20637 2908 20769 2920
rect 22119 2976 22251 2980
rect 22119 2920 22157 2976
rect 22213 2920 22251 2976
rect 22119 2908 22251 2920
rect 23601 2976 23733 2980
rect 23601 2920 23639 2976
rect 23695 2920 23733 2976
rect 23601 2908 23733 2920
rect 25083 2976 25215 2980
rect 25083 2920 25121 2976
rect 25177 2920 25215 2976
rect 25083 2908 25215 2920
rect 26565 2976 26697 2980
rect 26565 2920 26603 2976
rect 26659 2920 26697 2976
rect 26565 2908 26697 2920
rect 28047 2976 28179 2980
rect 28047 2920 28085 2976
rect 28141 2920 28179 2976
rect 28047 2908 28179 2920
rect 29529 2976 29661 2980
rect 29529 2920 29567 2976
rect 29623 2920 29661 2976
rect 29529 2908 29661 2920
rect 31011 2976 31143 2981
rect 31011 2920 31049 2976
rect 31105 2920 31143 2976
rect 31011 2908 31143 2920
rect 32493 2976 32625 2981
rect 32493 2920 32531 2976
rect 32587 2920 32625 2976
rect 32493 2908 32625 2920
rect 33975 2976 34107 2981
rect 33975 2920 34013 2976
rect 34069 2920 34107 2976
rect 33975 2908 34107 2920
rect 35457 2976 35589 2981
rect 35457 2920 35495 2976
rect 35551 2920 35589 2976
rect 35457 2908 35589 2920
rect 36939 2976 37071 2981
rect 36939 2920 36977 2976
rect 37033 2920 37071 2976
rect 36939 2908 37071 2920
rect 38421 2976 38553 2981
rect 38421 2920 38459 2976
rect 38515 2920 38553 2976
rect 38421 2908 38553 2920
rect 39903 2976 40035 2981
rect 39903 2920 39941 2976
rect 39997 2920 40035 2976
rect 39903 2908 40035 2920
rect 41385 2976 41517 2981
rect 41385 2920 41423 2976
rect 41479 2920 41517 2976
rect 41385 2908 41517 2920
rect 16112 2864 16476 2908
rect 16112 2800 16156 2864
rect 16220 2800 16476 2864
rect 16112 2756 16476 2800
rect 16536 2696 16900 2908
rect 17596 2864 17960 2908
rect 17596 2800 17640 2864
rect 17704 2800 17960 2864
rect 17596 2756 17960 2800
rect 18020 2696 18384 2908
rect 19080 2864 19444 2908
rect 19080 2800 19336 2864
rect 19400 2800 19444 2864
rect 19080 2756 19444 2800
rect 19504 2696 19868 2908
rect 20564 2864 20928 2908
rect 20564 2800 20608 2864
rect 20672 2800 20928 2864
rect 20564 2756 20928 2800
rect 20988 2696 21352 2908
rect 22048 2864 22412 2908
rect 22048 2800 22092 2864
rect 22156 2800 22412 2864
rect 22048 2756 22412 2800
rect 22472 2696 22836 2908
rect 23532 2864 23896 2908
rect 23532 2800 23788 2864
rect 23852 2800 23896 2864
rect 23532 2756 23896 2800
rect 23956 2696 24320 2908
rect 25016 2864 25380 2908
rect 25016 2800 25272 2864
rect 25336 2800 25380 2864
rect 25016 2756 25380 2800
rect 25440 2696 25804 2908
rect 26500 2864 26864 2908
rect 26500 2800 26756 2864
rect 26820 2800 26864 2864
rect 26500 2756 26864 2800
rect 27136 2735 27288 2908
rect 27984 2864 28348 2908
rect 27984 2800 28240 2864
rect 28304 2800 28348 2864
rect 27984 2756 28348 2800
rect 27099 2696 27288 2735
rect 28408 2696 28772 2908
rect 29468 2864 29832 2908
rect 29468 2800 29512 2864
rect 29576 2800 29832 2864
rect 29468 2756 29832 2800
rect 30104 2735 30256 2908
rect 30952 2864 31316 2908
rect 30952 2800 30996 2864
rect 31060 2800 31316 2864
rect 30952 2756 31316 2800
rect 30063 2696 30256 2735
rect 31376 2696 31740 2908
rect 32436 2864 32800 2908
rect 32436 2800 32480 2864
rect 32544 2800 32800 2864
rect 32436 2756 32800 2800
rect 32860 2696 33224 2908
rect 33920 2864 34284 2908
rect 33920 2800 33964 2864
rect 34028 2800 34284 2864
rect 33920 2756 34284 2800
rect 34344 2696 34708 2908
rect 35404 2864 35768 2908
rect 35404 2800 35660 2864
rect 35724 2800 35768 2864
rect 35404 2756 35768 2800
rect 35828 2696 36192 2908
rect 36888 2864 37252 2908
rect 36888 2800 36932 2864
rect 36996 2800 37252 2864
rect 36888 2756 37252 2800
rect 37312 2696 37676 2908
rect 38372 2864 38736 2908
rect 38372 2800 38628 2864
rect 38692 2800 38736 2864
rect 38372 2756 38736 2800
rect 38796 2696 39160 2908
rect 39856 2864 40220 2908
rect 39856 2800 39900 2864
rect 39964 2800 40220 2864
rect 39856 2756 40220 2800
rect 40280 2696 40644 2908
rect 41340 2864 41704 2908
rect 41340 2800 41596 2864
rect 41660 2800 41704 2864
rect 41340 2756 41704 2800
rect 41764 2696 42128 2908
rect 16536 2652 42128 2696
rect 16536 2588 16792 2652
rect 16856 2588 42128 2652
rect 16536 2544 42128 2588
rect 1484 2016 120144 2060
rect 1484 1952 1528 2016
rect 1592 1952 1740 2016
rect 1804 1952 1952 2016
rect 2016 1952 18064 2016
rect 18128 1952 24212 2016
rect 24276 1952 30148 2016
rect 30212 1952 37356 2016
rect 37420 1952 40324 2016
rect 40388 1952 119612 2016
rect 119676 1952 119824 2016
rect 119888 1952 120036 2016
rect 120100 1952 120144 2016
rect 1484 1804 120144 1952
rect 1484 1740 1528 1804
rect 1592 1740 1740 1804
rect 1804 1740 1952 1804
rect 2016 1740 119612 1804
rect 119676 1740 119824 1804
rect 119888 1740 120036 1804
rect 120100 1740 120144 1804
rect 1484 1592 120144 1740
rect 1484 1528 1528 1592
rect 1592 1528 1740 1592
rect 1804 1528 1952 1592
rect 2016 1528 119612 1592
rect 119676 1528 119824 1592
rect 119888 1528 120036 1592
rect 120100 1528 120144 1592
rect 1484 1484 120144 1528
rect 424 956 121204 1000
rect 424 892 468 956
rect 532 892 680 956
rect 744 892 892 956
rect 956 892 16792 956
rect 16856 892 120672 956
rect 120736 892 120884 956
rect 120948 892 121096 956
rect 121160 892 121204 956
rect 424 744 121204 892
rect 424 680 468 744
rect 532 680 680 744
rect 744 680 892 744
rect 956 680 120672 744
rect 120736 680 120884 744
rect 120948 680 121096 744
rect 121160 680 121204 744
rect 424 532 121204 680
rect 424 468 468 532
rect 532 468 680 532
rect 744 468 892 532
rect 956 468 120672 532
rect 120736 468 120884 532
rect 120948 468 121096 532
rect 121160 468 121204 532
rect 424 424 121204 468
<< via3 >>
rect 468 63432 532 63496
rect 680 63432 744 63496
rect 892 63432 956 63496
rect 120672 63432 120736 63496
rect 120884 63432 120948 63496
rect 121096 63432 121160 63496
rect 468 63220 532 63284
rect 680 63220 744 63284
rect 892 63220 956 63284
rect 120672 63220 120736 63284
rect 120884 63220 120948 63284
rect 121096 63220 121160 63284
rect 468 63008 532 63072
rect 680 63008 744 63072
rect 892 63008 956 63072
rect 21456 63008 21520 63072
rect 120672 63008 120736 63072
rect 120884 63008 120948 63072
rect 121096 63008 121160 63072
rect 1528 62372 1592 62436
rect 1740 62372 1804 62436
rect 1952 62372 2016 62436
rect 119612 62372 119676 62436
rect 119824 62372 119888 62436
rect 120036 62372 120100 62436
rect 1528 62160 1592 62224
rect 1740 62160 1804 62224
rect 1952 62160 2016 62224
rect 119612 62160 119676 62224
rect 119824 62160 119888 62224
rect 120036 62160 120100 62224
rect 1528 61948 1592 62012
rect 1740 61948 1804 62012
rect 1952 61948 2016 62012
rect 21244 61948 21308 62012
rect 119612 61948 119676 62012
rect 119824 61948 119888 62012
rect 120036 61948 120100 62012
rect 21456 61312 21520 61376
rect 20184 61100 20248 61164
rect 20184 60464 20248 60528
rect 21032 60464 21096 60528
rect 21244 59828 21308 59892
rect 21244 59616 21308 59680
rect 21244 58980 21308 59044
rect 21244 58768 21308 58832
rect 21032 58132 21096 58196
rect 21032 57284 21096 57348
rect 21244 56648 21308 56712
rect 21244 56436 21308 56500
rect 21244 56012 21308 56076
rect 21244 55800 21308 55864
rect 21032 55164 21096 55228
rect 21032 54316 21096 54380
rect 20184 53468 20248 53532
rect 21244 53468 21308 53532
rect 20184 52832 20248 52896
rect 21244 52832 21308 52896
rect 21032 51984 21096 52048
rect 19972 51348 20036 51412
rect 21244 50500 21308 50564
rect 21244 50288 21308 50352
rect 20184 49864 20248 49928
rect 21244 49864 21308 49928
rect 19972 49016 20036 49080
rect 21244 48804 21308 48868
rect 21244 48380 21308 48444
rect 21032 48168 21096 48232
rect 20184 47320 20248 47384
rect 21244 47320 21308 47384
rect 21244 46896 21308 46960
rect 21244 46684 21308 46748
rect 21032 45836 21096 45900
rect 21032 45200 21096 45264
rect 21244 44352 21308 44416
rect 21244 43716 21308 43780
rect 21032 42868 21096 42932
rect 16156 42656 16220 42720
rect 19972 42232 20036 42296
rect 15308 41172 15372 41236
rect 20184 41172 20248 41236
rect 21244 41172 21308 41236
rect 20184 40748 20248 40812
rect 21244 40748 21308 40812
rect 16156 39688 16220 39752
rect 16368 39688 16432 39752
rect 19972 39688 20036 39752
rect 20184 39264 20248 39328
rect 15308 38204 15372 38268
rect 15520 37992 15584 38056
rect 21244 38204 21308 38268
rect 21244 37568 21308 37632
rect 16156 36720 16220 36784
rect 20184 36720 20248 36784
rect 16368 36508 16432 36572
rect 21032 36084 21096 36148
rect 15520 35236 15584 35300
rect 15308 35024 15372 35088
rect 21244 35024 21308 35088
rect 15520 34812 15584 34876
rect 16368 34812 16432 34876
rect 21244 34600 21308 34664
rect 15520 33540 15584 33604
rect 16156 33540 16220 33604
rect 21032 33540 21096 33604
rect 21032 33116 21096 33180
rect 15308 32056 15372 32120
rect 21244 32056 21308 32120
rect 21244 31632 21308 31696
rect 16368 30572 16432 30636
rect 21032 30572 21096 30636
rect 16156 30360 16220 30424
rect 21032 30148 21096 30212
rect 21244 28876 21308 28940
rect 20184 28664 20248 28728
rect 16156 27392 16220 27456
rect 21032 27392 21096 27456
rect 16368 27180 16432 27244
rect 21244 26968 21308 27032
rect 20184 25908 20248 25972
rect 16156 25696 16220 25760
rect 19972 25484 20036 25548
rect 16368 24424 16432 24488
rect 21244 24424 21308 24488
rect 16368 24212 16432 24276
rect 21244 24212 21308 24276
rect 16156 22728 16220 22792
rect 19972 22728 20036 22792
rect 21244 22728 21308 22792
rect 16156 21244 16220 21308
rect 16368 21244 16432 21308
rect 21032 21244 21096 21308
rect 21456 21244 21520 21308
rect 21244 19760 21308 19824
rect 13612 19548 13676 19612
rect 21244 19336 21308 19400
rect 13824 18700 13888 18764
rect 15732 18700 15796 18764
rect 15732 18276 15796 18340
rect 16156 18276 16220 18340
rect 21456 18276 21520 18340
rect 13612 18064 13676 18128
rect 20184 18064 20248 18128
rect 13612 17852 13676 17916
rect 15732 17852 15796 17916
rect 13824 17216 13888 17280
rect 14036 17004 14100 17068
rect 15732 16580 15796 16644
rect 21244 16580 21308 16644
rect 13612 16368 13676 16432
rect 19972 16368 20036 16432
rect 13824 16156 13888 16220
rect 14036 15520 14100 15584
rect 14036 15308 14100 15372
rect 20184 15308 20248 15372
rect 21244 14884 21308 14948
rect 13612 14672 13676 14736
rect 13824 14672 13888 14736
rect 13824 13824 13888 13888
rect 14036 13824 14100 13888
rect 19972 13612 20036 13676
rect 15732 13400 15796 13464
rect 21880 13400 21944 13464
rect 13612 12976 13676 13040
rect 15732 12976 15796 13040
rect 13188 12340 13252 12404
rect 13824 12128 13888 12192
rect 21244 12128 21308 12192
rect 17004 11916 17068 11980
rect 19972 11916 20036 11980
rect 22304 11704 22368 11768
rect 25272 11704 25336 11768
rect 28452 11704 28516 11768
rect 31420 11704 31484 11768
rect 34600 11704 34664 11768
rect 37992 11704 38056 11768
rect 40748 11704 40812 11768
rect 43928 11704 43992 11768
rect 47108 11704 47172 11768
rect 50500 11704 50564 11768
rect 53256 11704 53320 11768
rect 56860 11704 56924 11768
rect 59616 11704 59680 11768
rect 62584 11704 62648 11768
rect 65764 11704 65828 11768
rect 68732 11704 68796 11768
rect 49652 11280 49716 11344
rect 50288 11280 50352 11344
rect 55800 11280 55864 11344
rect 56436 11280 56500 11344
rect 17004 11068 17068 11132
rect 19972 11068 20036 11132
rect 21880 11068 21944 11132
rect 22092 11068 22156 11132
rect 18064 10856 18128 10920
rect 21880 10856 21944 10920
rect 22304 10856 22368 10920
rect 22940 10856 23004 10920
rect 28240 11068 28304 11132
rect 28452 11068 28516 11132
rect 24848 10856 24912 10920
rect 25060 10856 25124 10920
rect 25272 10856 25336 10920
rect 25908 10856 25972 10920
rect 34812 11068 34876 11132
rect 37780 11068 37844 11132
rect 28028 10856 28092 10920
rect 28452 10856 28516 10920
rect 30996 10856 31060 10920
rect 31208 10856 31272 10920
rect 31420 10856 31484 10920
rect 32268 10856 32332 10920
rect 34176 10856 34240 10920
rect 44140 11068 44204 11132
rect 34600 10856 34664 10920
rect 35024 10856 35088 10920
rect 37356 10856 37420 10920
rect 37992 10856 38056 10920
rect 38628 10856 38692 10920
rect 40324 10856 40388 10920
rect 40536 10856 40600 10920
rect 40748 10856 40812 10920
rect 41172 10856 41236 10920
rect 50076 11068 50140 11132
rect 43504 10856 43568 10920
rect 43928 10856 43992 10920
rect 44776 10856 44840 10920
rect 46472 10856 46536 10920
rect 46684 10856 46748 10920
rect 47108 10856 47172 10920
rect 47532 10856 47596 10920
rect 49864 10856 49928 10920
rect 56648 11068 56712 11132
rect 59404 11068 59468 11132
rect 62796 11068 62860 11132
rect 65976 11068 66040 11132
rect 50288 10856 50352 10920
rect 50500 10856 50564 10920
rect 52832 10856 52896 10920
rect 53044 10856 53108 10920
rect 53256 10856 53320 10920
rect 53468 10856 53532 10920
rect 56012 10856 56076 10920
rect 56436 10856 56500 10920
rect 56860 10856 56924 10920
rect 59616 10856 59680 10920
rect 60040 10856 60104 10920
rect 62160 10856 62224 10920
rect 62584 10856 62648 10920
rect 63008 10856 63072 10920
rect 65340 10856 65404 10920
rect 65764 10856 65828 10920
rect 66612 10856 66676 10920
rect 68308 10856 68372 10920
rect 68520 10856 68584 10920
rect 68732 10856 68796 10920
rect 69156 10856 69220 10920
rect 22304 10698 22368 10708
rect 22304 10644 22354 10698
rect 22354 10644 22368 10698
rect 25484 10644 25548 10708
rect 28664 10644 28728 10708
rect 31632 10698 31696 10708
rect 31632 10644 31634 10698
rect 31634 10644 31690 10698
rect 31690 10644 31696 10698
rect 34600 10644 34664 10708
rect 37992 10644 38056 10708
rect 40960 10698 41024 10708
rect 40960 10644 40970 10698
rect 40970 10644 41024 10698
rect 43928 10644 43992 10708
rect 47108 10644 47172 10708
rect 50500 10644 50564 10708
rect 53256 10644 53320 10708
rect 56436 10644 56500 10708
rect 59828 10644 59892 10708
rect 62584 10644 62648 10708
rect 65764 10644 65828 10708
rect 68944 10698 69008 10708
rect 68944 10644 68978 10698
rect 68978 10644 69008 10698
rect 71912 10644 71976 10708
rect 120672 10856 120736 10920
rect 21880 10220 21944 10284
rect 18912 10008 18976 10072
rect 30996 10008 31060 10072
rect 40324 10008 40388 10072
rect 46472 10008 46536 10072
rect 68308 10008 68372 10072
rect 22092 9796 22156 9860
rect 24848 9796 24912 9860
rect 25060 9796 25124 9860
rect 28028 9796 28092 9860
rect 28240 9796 28304 9860
rect 31208 9796 31272 9860
rect 34176 9796 34240 9860
rect 34812 9796 34876 9860
rect 37356 9796 37420 9860
rect 37780 9796 37844 9860
rect 40536 9796 40600 9860
rect 43504 9796 43568 9860
rect 44140 9796 44204 9860
rect 46684 9796 46748 9860
rect 49864 9796 49928 9860
rect 50076 9796 50140 9860
rect 52832 9796 52896 9860
rect 53044 9796 53108 9860
rect 56012 9796 56076 9860
rect 56648 9796 56712 9860
rect 59404 9796 59468 9860
rect 62160 9796 62224 9860
rect 62796 9796 62860 9860
rect 65340 9796 65404 9860
rect 65976 9796 66040 9860
rect 68520 9796 68584 9860
rect 119612 9796 119676 9860
rect 18064 9372 18128 9436
rect 19124 9160 19188 9224
rect 18912 8524 18976 8588
rect 35024 8524 35088 8588
rect 53468 8524 53532 8588
rect 69156 8524 69220 8588
rect 22940 8312 23004 8376
rect 25908 8312 25972 8376
rect 28240 8312 28304 8376
rect 32268 8312 32332 8376
rect 38628 8312 38692 8376
rect 41172 8312 41236 8376
rect 44776 8312 44840 8376
rect 47532 8312 47596 8376
rect 49652 8312 49716 8376
rect 55800 8312 55864 8376
rect 60040 8312 60104 8376
rect 63008 8312 63072 8376
rect 66612 8312 66676 8376
rect 71912 8312 71976 8376
rect 892 7676 956 7740
rect 2588 7676 2652 7740
rect 19124 7676 19188 7740
rect 6192 7040 6256 7104
rect 1952 6828 2016 6892
rect 28876 6404 28940 6468
rect 2588 5980 2652 6044
rect 18064 3436 18128 3500
rect 24212 3436 24276 3500
rect 28876 3648 28940 3712
rect 30148 3436 30212 3500
rect 37356 3436 37420 3500
rect 40324 3436 40388 3500
rect 16156 2800 16220 2864
rect 17640 2800 17704 2864
rect 19336 2800 19400 2864
rect 20608 2800 20672 2864
rect 22092 2800 22156 2864
rect 23788 2800 23852 2864
rect 25272 2800 25336 2864
rect 26756 2800 26820 2864
rect 28240 2800 28304 2864
rect 29512 2800 29576 2864
rect 30996 2800 31060 2864
rect 32480 2800 32544 2864
rect 33964 2800 34028 2864
rect 35660 2800 35724 2864
rect 36932 2800 36996 2864
rect 38628 2800 38692 2864
rect 39900 2800 39964 2864
rect 41596 2800 41660 2864
rect 16792 2588 16856 2652
rect 1528 1952 1592 2016
rect 1740 1952 1804 2016
rect 1952 1952 2016 2016
rect 18064 1952 18128 2016
rect 24212 1952 24276 2016
rect 30148 1952 30212 2016
rect 37356 1952 37420 2016
rect 40324 1952 40388 2016
rect 119612 1952 119676 2016
rect 119824 1952 119888 2016
rect 120036 1952 120100 2016
rect 1528 1740 1592 1804
rect 1740 1740 1804 1804
rect 1952 1740 2016 1804
rect 119612 1740 119676 1804
rect 119824 1740 119888 1804
rect 120036 1740 120100 1804
rect 1528 1528 1592 1592
rect 1740 1528 1804 1592
rect 1952 1528 2016 1592
rect 119612 1528 119676 1592
rect 119824 1528 119888 1592
rect 120036 1528 120100 1592
rect 468 892 532 956
rect 680 892 744 956
rect 892 892 956 956
rect 16792 892 16856 956
rect 120672 892 120736 956
rect 120884 892 120948 956
rect 121096 892 121160 956
rect 468 680 532 744
rect 680 680 744 744
rect 892 680 956 744
rect 120672 680 120736 744
rect 120884 680 120948 744
rect 121096 680 121160 744
rect 468 468 532 532
rect 680 468 744 532
rect 892 468 956 532
rect 120672 468 120736 532
rect 120884 468 120948 532
rect 121096 468 121160 532
<< metal4 >>
rect 424 63496 1000 63540
rect 424 63432 468 63496
rect 532 63432 680 63496
rect 744 63432 892 63496
rect 956 63432 1000 63496
rect 424 63284 1000 63432
rect 424 63220 468 63284
rect 532 63220 680 63284
rect 744 63220 892 63284
rect 956 63220 1000 63284
rect 424 63072 1000 63220
rect 120628 63496 121204 63540
rect 120628 63432 120672 63496
rect 120736 63432 120884 63496
rect 120948 63432 121096 63496
rect 121160 63432 121204 63496
rect 120628 63284 121204 63432
rect 120628 63220 120672 63284
rect 120736 63220 120884 63284
rect 120948 63220 121096 63284
rect 121160 63220 121204 63284
rect 424 63008 468 63072
rect 532 63008 680 63072
rect 744 63008 892 63072
rect 956 63008 1000 63072
rect 424 7740 1000 63008
rect 21412 63072 21564 63116
rect 21412 63008 21456 63072
rect 21520 63008 21564 63072
rect 424 7676 892 7740
rect 956 7676 1000 7740
rect 424 956 1000 7676
rect 1484 62436 2060 62480
rect 1484 62372 1528 62436
rect 1592 62372 1740 62436
rect 1804 62372 1952 62436
rect 2016 62372 2060 62436
rect 1484 62224 2060 62372
rect 1484 62160 1528 62224
rect 1592 62160 1740 62224
rect 1804 62160 1952 62224
rect 2016 62160 2060 62224
rect 1484 62012 2060 62160
rect 1484 61948 1528 62012
rect 1592 61948 1740 62012
rect 1804 61948 1952 62012
rect 2016 61948 2060 62012
rect 1484 6892 2060 61948
rect 21200 62012 21352 62056
rect 21200 61948 21244 62012
rect 21308 61948 21352 62012
rect 20140 61164 20292 61208
rect 20140 61100 20184 61164
rect 20248 61100 20292 61164
rect 20140 60528 20292 61100
rect 20140 60496 20184 60528
rect 20170 60464 20184 60496
rect 20248 60496 20292 60528
rect 21018 60528 21110 60542
rect 21018 60496 21032 60528
rect 20248 60464 20262 60496
rect 20170 60450 20262 60464
rect 20988 60464 21032 60496
rect 21096 60496 21110 60528
rect 21096 60464 21140 60496
rect 20988 58196 21140 60464
rect 21200 59892 21352 61948
rect 21412 61376 21564 63008
rect 120628 63072 121204 63220
rect 120628 63008 120672 63072
rect 120736 63008 120884 63072
rect 120948 63008 121096 63072
rect 121160 63008 121204 63072
rect 21412 61344 21456 61376
rect 21442 61312 21456 61344
rect 21520 61344 21564 61376
rect 119568 62436 120144 62480
rect 119568 62372 119612 62436
rect 119676 62372 119824 62436
rect 119888 62372 120036 62436
rect 120100 62372 120144 62436
rect 119568 62224 120144 62372
rect 119568 62160 119612 62224
rect 119676 62160 119824 62224
rect 119888 62160 120036 62224
rect 120100 62160 120144 62224
rect 119568 62012 120144 62160
rect 119568 61948 119612 62012
rect 119676 61948 119824 62012
rect 119888 61948 120036 62012
rect 120100 61948 120144 62012
rect 21520 61312 21534 61344
rect 21442 61298 21534 61312
rect 21200 59860 21244 59892
rect 21230 59828 21244 59860
rect 21308 59860 21352 59892
rect 21308 59828 21322 59860
rect 21230 59814 21322 59828
rect 21200 59680 21352 59724
rect 21200 59616 21244 59680
rect 21308 59616 21352 59680
rect 21200 59044 21352 59616
rect 21200 59012 21244 59044
rect 21230 58980 21244 59012
rect 21308 59012 21352 59044
rect 21308 58980 21322 59012
rect 21230 58966 21322 58980
rect 21230 58832 21322 58846
rect 21230 58800 21244 58832
rect 20988 58132 21032 58196
rect 21096 58132 21140 58196
rect 20988 58088 21140 58132
rect 21200 58768 21244 58800
rect 21308 58800 21322 58832
rect 21308 58768 21352 58800
rect 21018 57348 21110 57362
rect 21018 57316 21032 57348
rect 20988 57284 21032 57316
rect 21096 57316 21110 57348
rect 21096 57284 21140 57316
rect 20988 55228 21140 57284
rect 21200 56712 21352 58768
rect 21200 56648 21244 56712
rect 21308 56648 21352 56712
rect 21200 56604 21352 56648
rect 21200 56500 21352 56544
rect 21200 56436 21244 56500
rect 21308 56436 21352 56500
rect 21200 56076 21352 56436
rect 21200 56044 21244 56076
rect 21230 56012 21244 56044
rect 21308 56044 21352 56076
rect 21308 56012 21322 56044
rect 21230 55998 21322 56012
rect 21230 55864 21322 55878
rect 21230 55832 21244 55864
rect 20988 55164 21032 55228
rect 21096 55164 21140 55228
rect 20988 55120 21140 55164
rect 21200 55800 21244 55832
rect 21308 55832 21322 55864
rect 21308 55800 21352 55832
rect 21018 54380 21110 54394
rect 21018 54348 21032 54380
rect 20988 54316 21032 54348
rect 21096 54348 21110 54380
rect 21096 54316 21140 54348
rect 20140 53532 20292 53576
rect 20140 53468 20184 53532
rect 20248 53468 20292 53532
rect 20140 52896 20292 53468
rect 20140 52864 20184 52896
rect 20170 52832 20184 52864
rect 20248 52864 20292 52896
rect 20248 52832 20262 52864
rect 20170 52818 20262 52832
rect 20988 52048 21140 54316
rect 21200 53532 21352 55800
rect 21200 53468 21244 53532
rect 21308 53468 21352 53532
rect 21200 53424 21352 53468
rect 21230 52896 21322 52910
rect 21230 52864 21244 52896
rect 20988 51984 21032 52048
rect 21096 51984 21140 52048
rect 20988 51940 21140 51984
rect 21200 52832 21244 52864
rect 21308 52864 21322 52896
rect 21308 52832 21352 52864
rect 19958 51412 20050 51426
rect 19958 51380 19972 51412
rect 19928 51348 19972 51380
rect 20036 51380 20050 51412
rect 20036 51348 20080 51380
rect 19928 49080 20080 51348
rect 21200 50564 21352 52832
rect 21200 50500 21244 50564
rect 21308 50500 21352 50564
rect 21200 50456 21352 50500
rect 21200 50352 21352 50396
rect 21200 50288 21244 50352
rect 21308 50288 21352 50352
rect 20170 49928 20262 49942
rect 20170 49896 20184 49928
rect 19928 49016 19972 49080
rect 20036 49016 20080 49080
rect 19928 48972 20080 49016
rect 20140 49864 20184 49896
rect 20248 49896 20262 49928
rect 21200 49928 21352 50288
rect 21200 49896 21244 49928
rect 20248 49864 20292 49896
rect 20140 47384 20292 49864
rect 21230 49864 21244 49896
rect 21308 49896 21352 49928
rect 21308 49864 21322 49896
rect 21230 49850 21322 49864
rect 21200 48868 21352 48912
rect 21200 48804 21244 48868
rect 21308 48804 21352 48868
rect 21200 48444 21352 48804
rect 21200 48412 21244 48444
rect 21230 48380 21244 48412
rect 21308 48412 21352 48444
rect 21308 48380 21322 48412
rect 21230 48366 21322 48380
rect 21018 48232 21110 48246
rect 21018 48200 21032 48232
rect 20140 47320 20184 47384
rect 20248 47320 20292 47384
rect 20140 47276 20292 47320
rect 20988 48168 21032 48200
rect 21096 48200 21110 48232
rect 21096 48168 21140 48200
rect 20988 45900 21140 48168
rect 21200 47384 21352 47428
rect 21200 47320 21244 47384
rect 21308 47320 21352 47384
rect 21200 46960 21352 47320
rect 21200 46928 21244 46960
rect 21230 46896 21244 46928
rect 21308 46928 21352 46960
rect 21308 46896 21322 46928
rect 21230 46882 21322 46896
rect 21230 46748 21322 46762
rect 21230 46716 21244 46748
rect 20988 45836 21032 45900
rect 21096 45836 21140 45900
rect 20988 45792 21140 45836
rect 21200 46684 21244 46716
rect 21308 46716 21322 46748
rect 21308 46684 21352 46716
rect 21018 45264 21110 45278
rect 21018 45232 21032 45264
rect 20988 45200 21032 45232
rect 21096 45232 21110 45264
rect 21096 45200 21140 45232
rect 20988 42932 21140 45200
rect 21200 44416 21352 46684
rect 21200 44352 21244 44416
rect 21308 44352 21352 44416
rect 21200 44308 21352 44352
rect 21230 43780 21322 43794
rect 21230 43748 21244 43780
rect 20988 42868 21032 42932
rect 21096 42868 21140 42932
rect 20988 42824 21140 42868
rect 21200 43716 21244 43748
rect 21308 43748 21322 43780
rect 21308 43716 21352 43748
rect 16112 42720 16264 42764
rect 16112 42656 16156 42720
rect 16220 42656 16264 42720
rect 15294 41236 15386 41250
rect 15294 41204 15308 41236
rect 15264 41172 15308 41204
rect 15372 41204 15386 41236
rect 15372 41172 15416 41204
rect 15264 38268 15416 41172
rect 16112 39752 16264 42656
rect 19958 42296 20050 42310
rect 19958 42264 19972 42296
rect 19928 42232 19972 42264
rect 20036 42264 20050 42296
rect 20036 42232 20080 42264
rect 16112 39720 16156 39752
rect 16142 39688 16156 39720
rect 16220 39720 16264 39752
rect 16324 39752 16476 39796
rect 16220 39688 16234 39720
rect 16142 39674 16234 39688
rect 16324 39688 16368 39752
rect 16432 39688 16476 39752
rect 16324 39584 16476 39688
rect 19928 39752 20080 42232
rect 20140 41236 20292 41280
rect 20140 41172 20184 41236
rect 20248 41172 20292 41236
rect 20140 40812 20292 41172
rect 21200 41236 21352 43716
rect 21200 41172 21244 41236
rect 21308 41172 21352 41236
rect 21200 41128 21352 41172
rect 20140 40780 20184 40812
rect 20170 40748 20184 40780
rect 20248 40780 20292 40812
rect 21230 40812 21322 40826
rect 21230 40780 21244 40812
rect 20248 40748 20262 40780
rect 20170 40734 20262 40748
rect 21200 40748 21244 40780
rect 21308 40780 21322 40812
rect 21308 40748 21352 40780
rect 19928 39688 19972 39752
rect 20036 39688 20080 39752
rect 19928 39644 20080 39688
rect 15264 38204 15308 38268
rect 15372 38204 15416 38268
rect 15264 38160 15416 38204
rect 16112 39432 16476 39584
rect 15506 38056 15598 38070
rect 15506 38024 15520 38056
rect 15476 37992 15520 38024
rect 15584 38024 15598 38056
rect 15584 37992 15628 38024
rect 15476 35300 15628 37992
rect 16112 36784 16264 39432
rect 20170 39328 20262 39342
rect 20170 39296 20184 39328
rect 16112 36752 16156 36784
rect 16142 36720 16156 36752
rect 16220 36752 16264 36784
rect 20140 39264 20184 39296
rect 20248 39296 20262 39328
rect 20248 39264 20292 39296
rect 20140 36784 20292 39264
rect 21200 38268 21352 40748
rect 21200 38204 21244 38268
rect 21308 38204 21352 38268
rect 21200 38160 21352 38204
rect 21230 37632 21322 37646
rect 21230 37600 21244 37632
rect 16220 36720 16234 36752
rect 16142 36706 16234 36720
rect 20140 36720 20184 36784
rect 20248 36720 20292 36784
rect 20140 36676 20292 36720
rect 21200 37568 21244 37600
rect 21308 37600 21322 37632
rect 21308 37568 21352 37600
rect 15476 35236 15520 35300
rect 15584 35236 15628 35300
rect 15476 35192 15628 35236
rect 16324 36572 16476 36616
rect 16324 36508 16368 36572
rect 16432 36508 16476 36572
rect 15264 35088 15416 35132
rect 15264 35024 15308 35088
rect 15372 35024 15416 35088
rect 15264 32120 15416 35024
rect 15476 34876 15628 34920
rect 15476 34812 15520 34876
rect 15584 34812 15628 34876
rect 16324 34876 16476 36508
rect 21018 36148 21110 36162
rect 21018 36116 21032 36148
rect 16324 34844 16368 34876
rect 15476 33604 15628 34812
rect 16354 34812 16368 34844
rect 16432 34844 16476 34876
rect 20988 36084 21032 36116
rect 21096 36116 21110 36148
rect 21096 36084 21140 36116
rect 16432 34812 16446 34844
rect 16354 34798 16446 34812
rect 15476 33572 15520 33604
rect 15506 33540 15520 33572
rect 15584 33572 15628 33604
rect 16142 33604 16234 33618
rect 16142 33572 16156 33604
rect 15584 33540 15598 33572
rect 15506 33526 15598 33540
rect 16112 33540 16156 33572
rect 16220 33572 16234 33604
rect 20988 33604 21140 36084
rect 21200 35088 21352 37568
rect 21200 35024 21244 35088
rect 21308 35024 21352 35088
rect 21200 34980 21352 35024
rect 21230 34664 21322 34678
rect 21230 34632 21244 34664
rect 16220 33540 16264 33572
rect 15264 32088 15308 32120
rect 15294 32056 15308 32088
rect 15372 32088 15416 32120
rect 15372 32056 15386 32088
rect 15294 32042 15386 32056
rect 16112 30680 16264 33540
rect 20988 33540 21032 33604
rect 21096 33540 21140 33604
rect 20988 33496 21140 33540
rect 21200 34600 21244 34632
rect 21308 34632 21322 34664
rect 21308 34600 21352 34632
rect 21018 33180 21110 33194
rect 21018 33148 21032 33180
rect 20988 33116 21032 33148
rect 21096 33148 21110 33180
rect 21096 33116 21140 33148
rect 16112 30636 16476 30680
rect 16112 30572 16368 30636
rect 16432 30572 16476 30636
rect 16112 30528 16476 30572
rect 20988 30636 21140 33116
rect 21200 32120 21352 34600
rect 21200 32056 21244 32120
rect 21308 32056 21352 32120
rect 21200 32012 21352 32056
rect 21230 31696 21322 31710
rect 21230 31664 21244 31696
rect 20988 30572 21032 30636
rect 21096 30572 21140 30636
rect 20988 30528 21140 30572
rect 21200 31632 21244 31664
rect 21308 31664 21322 31696
rect 21308 31632 21352 31664
rect 16142 30424 16234 30438
rect 16142 30392 16156 30424
rect 16112 30360 16156 30392
rect 16220 30392 16234 30424
rect 16220 30360 16264 30392
rect 16112 27456 16264 30360
rect 21018 30212 21110 30226
rect 21018 30180 21032 30212
rect 20988 30148 21032 30180
rect 21096 30180 21110 30212
rect 21096 30148 21140 30180
rect 20170 28728 20262 28742
rect 20170 28696 20184 28728
rect 16112 27392 16156 27456
rect 16220 27392 16264 27456
rect 16112 27348 16264 27392
rect 20140 28664 20184 28696
rect 20248 28696 20262 28728
rect 20248 28664 20292 28696
rect 16354 27244 16446 27258
rect 16354 27212 16368 27244
rect 16324 27180 16368 27212
rect 16432 27212 16446 27244
rect 16432 27180 16476 27212
rect 16112 25760 16264 25804
rect 16112 25696 16156 25760
rect 16220 25696 16264 25760
rect 16112 22792 16264 25696
rect 16324 24488 16476 27180
rect 20140 25972 20292 28664
rect 20988 27456 21140 30148
rect 21200 28940 21352 31632
rect 21200 28876 21244 28940
rect 21308 28876 21352 28940
rect 21200 28832 21352 28876
rect 20988 27392 21032 27456
rect 21096 27392 21140 27456
rect 20988 27348 21140 27392
rect 21230 27032 21322 27046
rect 21230 27000 21244 27032
rect 20140 25908 20184 25972
rect 20248 25908 20292 25972
rect 20140 25864 20292 25908
rect 21200 26968 21244 27000
rect 21308 27000 21322 27032
rect 21308 26968 21352 27000
rect 16324 24424 16368 24488
rect 16432 24424 16476 24488
rect 16324 24380 16476 24424
rect 19928 25548 20080 25592
rect 19928 25484 19972 25548
rect 20036 25484 20080 25548
rect 16112 22760 16156 22792
rect 16142 22728 16156 22760
rect 16220 22760 16264 22792
rect 16324 24276 16476 24320
rect 16324 24212 16368 24276
rect 16432 24212 16476 24276
rect 16220 22728 16234 22760
rect 16142 22714 16234 22728
rect 16142 21308 16234 21322
rect 16142 21276 16156 21308
rect 16112 21244 16156 21276
rect 16220 21276 16234 21308
rect 16324 21308 16476 24212
rect 19928 22792 20080 25484
rect 21200 24488 21352 26968
rect 21200 24424 21244 24488
rect 21308 24424 21352 24488
rect 21200 24380 21352 24424
rect 19928 22760 19972 22792
rect 19958 22728 19972 22760
rect 20036 22760 20080 22792
rect 20988 24276 21352 24320
rect 20988 24212 21244 24276
rect 21308 24212 21352 24276
rect 20988 24168 21352 24212
rect 20036 22728 20050 22760
rect 19958 22714 20050 22728
rect 16324 21276 16368 21308
rect 16220 21244 16264 21276
rect 13598 19612 13690 19626
rect 13598 19580 13612 19612
rect 13568 19548 13612 19580
rect 13676 19580 13690 19612
rect 13676 19548 13720 19580
rect 13568 18128 13720 19548
rect 13810 18764 13902 18778
rect 13810 18732 13824 18764
rect 13568 18064 13612 18128
rect 13676 18064 13720 18128
rect 13568 18020 13720 18064
rect 13780 18700 13824 18732
rect 13888 18732 13902 18764
rect 15718 18764 15810 18778
rect 15718 18732 15732 18764
rect 13888 18700 13932 18732
rect 13568 17916 13720 17960
rect 13568 17852 13612 17916
rect 13676 17852 13720 17916
rect 13568 16432 13720 17852
rect 13780 17280 13932 18700
rect 15688 18700 15732 18732
rect 15796 18732 15810 18764
rect 15796 18700 15840 18732
rect 15688 18340 15840 18700
rect 15688 18276 15732 18340
rect 15796 18276 15840 18340
rect 15688 18232 15840 18276
rect 16112 18340 16264 21244
rect 16354 21244 16368 21276
rect 16432 21276 16476 21308
rect 20988 21308 21140 24168
rect 21230 22792 21322 22806
rect 21230 22760 21244 22792
rect 20988 21276 21032 21308
rect 16432 21244 16446 21276
rect 16354 21230 16446 21244
rect 21018 21244 21032 21276
rect 21096 21276 21140 21308
rect 21200 22728 21244 22760
rect 21308 22760 21322 22792
rect 21308 22728 21352 22760
rect 21096 21244 21110 21276
rect 21018 21230 21110 21244
rect 21200 19824 21352 22728
rect 21442 21308 21534 21322
rect 21442 21276 21456 21308
rect 21200 19760 21244 19824
rect 21308 19760 21352 19824
rect 21200 19716 21352 19760
rect 21412 21244 21456 21276
rect 21520 21276 21534 21308
rect 21520 21244 21564 21276
rect 21230 19400 21322 19414
rect 21230 19368 21244 19400
rect 16112 18276 16156 18340
rect 16220 18276 16264 18340
rect 16112 18232 16264 18276
rect 21200 19336 21244 19368
rect 21308 19368 21322 19400
rect 21308 19336 21352 19368
rect 20170 18128 20262 18142
rect 20170 18096 20184 18128
rect 20140 18064 20184 18096
rect 20248 18096 20262 18128
rect 20248 18064 20292 18096
rect 15718 17916 15810 17930
rect 15718 17884 15732 17916
rect 13780 17216 13824 17280
rect 13888 17216 13932 17280
rect 13780 17172 13932 17216
rect 15688 17852 15732 17884
rect 15796 17884 15810 17916
rect 15796 17852 15840 17884
rect 13568 16400 13612 16432
rect 13598 16368 13612 16400
rect 13676 16400 13720 16432
rect 13992 17068 14144 17112
rect 13992 17004 14036 17068
rect 14100 17004 14144 17068
rect 13676 16368 13690 16400
rect 13598 16354 13690 16368
rect 13810 16220 13902 16234
rect 13810 16188 13824 16220
rect 13780 16156 13824 16188
rect 13888 16188 13902 16220
rect 13888 16156 13932 16188
rect 13598 14736 13690 14750
rect 13598 14704 13612 14736
rect 13568 14672 13612 14704
rect 13676 14704 13690 14736
rect 13780 14736 13932 16156
rect 13992 15584 14144 17004
rect 15688 16644 15840 17852
rect 15688 16580 15732 16644
rect 15796 16580 15840 16644
rect 15688 16536 15840 16580
rect 19958 16432 20050 16446
rect 19958 16400 19972 16432
rect 13992 15552 14036 15584
rect 14022 15520 14036 15552
rect 14100 15552 14144 15584
rect 19928 16368 19972 16400
rect 20036 16400 20050 16432
rect 20036 16368 20080 16400
rect 14100 15520 14114 15552
rect 14022 15506 14114 15520
rect 13676 14672 13720 14704
rect 13568 13040 13720 14672
rect 13780 14672 13824 14736
rect 13888 14672 13932 14736
rect 13780 14628 13932 14672
rect 13992 15372 14144 15416
rect 13992 15308 14036 15372
rect 14100 15308 14144 15372
rect 13810 13888 13902 13902
rect 13810 13856 13824 13888
rect 13568 12976 13612 13040
rect 13676 12976 13720 13040
rect 13568 12932 13720 12976
rect 13780 13824 13824 13856
rect 13888 13856 13902 13888
rect 13992 13888 14144 15308
rect 13992 13856 14036 13888
rect 13888 13824 13932 13856
rect 13174 12404 13266 12418
rect 13174 12372 13188 12404
rect 13144 12340 13188 12372
rect 13252 12372 13266 12404
rect 13252 12340 13296 12372
rect 2574 7740 2666 7754
rect 2574 7708 2588 7740
rect 1484 6828 1952 6892
rect 2016 6828 2060 6892
rect 1484 2016 2060 6828
rect 2544 7676 2588 7708
rect 2652 7708 2666 7740
rect 2652 7676 2696 7708
rect 2544 6044 2696 7676
rect 6178 7104 6270 7118
rect 6178 7072 6192 7104
rect 2544 5980 2588 6044
rect 2652 5980 2696 6044
rect 2544 5936 2696 5980
rect 6148 7040 6192 7072
rect 6256 7072 6270 7104
rect 6256 7040 6300 7072
rect 1484 1952 1528 2016
rect 1592 1952 1740 2016
rect 1804 1952 1952 2016
rect 2016 1952 2060 2016
rect 1484 1804 2060 1952
rect 1484 1740 1528 1804
rect 1592 1740 1740 1804
rect 1804 1740 1952 1804
rect 2016 1740 2060 1804
rect 1484 1592 2060 1740
rect 1484 1528 1528 1592
rect 1592 1528 1740 1592
rect 1804 1528 1952 1592
rect 2016 1528 2060 1592
rect 1484 1484 2060 1528
rect 424 892 468 956
rect 532 892 680 956
rect 744 892 892 956
rect 956 892 1000 956
rect 424 744 1000 892
rect 424 680 468 744
rect 532 680 680 744
rect 744 680 892 744
rect 956 680 1000 744
rect 424 532 1000 680
rect 424 468 468 532
rect 532 468 680 532
rect 744 468 892 532
rect 956 468 1000 532
rect 424 424 1000 468
rect 6148 0 6300 7040
rect 13144 0 13296 12340
rect 13780 12192 13932 13824
rect 14022 13824 14036 13856
rect 14100 13856 14144 13888
rect 14100 13824 14114 13856
rect 14022 13810 14114 13824
rect 19928 13676 20080 16368
rect 20140 15372 20292 18064
rect 21200 16644 21352 19336
rect 21412 18340 21564 21244
rect 21412 18276 21456 18340
rect 21520 18276 21564 18340
rect 21412 18232 21564 18276
rect 21200 16580 21244 16644
rect 21308 16580 21352 16644
rect 21200 16536 21352 16580
rect 20140 15308 20184 15372
rect 20248 15308 20292 15372
rect 20140 15264 20292 15308
rect 21230 14948 21322 14962
rect 21230 14916 21244 14948
rect 19928 13612 19972 13676
rect 20036 13612 20080 13676
rect 19928 13568 20080 13612
rect 21200 14884 21244 14916
rect 21308 14916 21322 14948
rect 21308 14884 21352 14916
rect 15688 13464 15840 13508
rect 15688 13400 15732 13464
rect 15796 13400 15840 13464
rect 15688 13040 15840 13400
rect 15688 13008 15732 13040
rect 15718 12976 15732 13008
rect 15796 13008 15840 13040
rect 15796 12976 15810 13008
rect 15718 12962 15810 12976
rect 13780 12128 13824 12192
rect 13888 12128 13932 12192
rect 13780 12084 13932 12128
rect 21200 12192 21352 14884
rect 21866 13464 21958 13478
rect 21866 13432 21880 13464
rect 21200 12128 21244 12192
rect 21308 12128 21352 12192
rect 21200 12084 21352 12128
rect 21836 13400 21880 13432
rect 21944 13432 21958 13464
rect 21944 13400 21988 13432
rect 16990 11980 17082 11994
rect 16990 11948 17004 11980
rect 16960 11916 17004 11948
rect 17068 11948 17082 11980
rect 19928 11980 20080 12024
rect 17068 11916 17112 11948
rect 16960 11132 17112 11916
rect 16960 11068 17004 11132
rect 17068 11068 17112 11132
rect 19928 11916 19972 11980
rect 20036 11916 20080 11980
rect 19928 11132 20080 11916
rect 19928 11100 19972 11132
rect 16960 11024 17112 11068
rect 19958 11068 19972 11100
rect 20036 11100 20080 11132
rect 21836 11132 21988 13400
rect 22290 11768 22382 11782
rect 22290 11736 22304 11768
rect 22260 11704 22304 11736
rect 22368 11736 22382 11768
rect 25258 11768 25350 11782
rect 25258 11736 25272 11768
rect 22368 11704 22412 11736
rect 20036 11068 20050 11100
rect 19958 11054 20050 11068
rect 21836 11068 21880 11132
rect 21944 11068 21988 11132
rect 22078 11132 22170 11146
rect 22078 11100 22092 11132
rect 21836 11024 21988 11068
rect 22048 11068 22092 11100
rect 22156 11100 22170 11132
rect 22156 11068 22200 11100
rect 18050 10920 18142 10934
rect 18050 10888 18064 10920
rect 18020 10856 18064 10888
rect 18128 10888 18142 10920
rect 21836 10920 21988 10964
rect 18128 10856 18172 10888
rect 18020 9436 18172 10856
rect 21836 10856 21880 10920
rect 21944 10856 21988 10920
rect 21836 10284 21988 10856
rect 21836 10252 21880 10284
rect 21866 10220 21880 10252
rect 21944 10252 21988 10284
rect 21944 10220 21958 10252
rect 21866 10206 21958 10220
rect 18020 9372 18064 9436
rect 18128 9372 18172 9436
rect 18020 9328 18172 9372
rect 18868 10072 19020 10116
rect 18868 10008 18912 10072
rect 18976 10008 19020 10072
rect 18868 8588 19020 10008
rect 22048 9860 22200 11068
rect 22260 10920 22412 11704
rect 25228 11704 25272 11736
rect 25336 11736 25350 11768
rect 28438 11768 28530 11782
rect 28438 11736 28452 11768
rect 25336 11704 25380 11736
rect 22260 10856 22304 10920
rect 22368 10856 22412 10920
rect 22926 10920 23018 10934
rect 22926 10888 22940 10920
rect 22260 10812 22412 10856
rect 22896 10856 22940 10888
rect 23004 10888 23018 10920
rect 24804 10920 24956 10964
rect 23004 10856 23048 10888
rect 22290 10708 22382 10722
rect 22290 10676 22304 10708
rect 22048 9796 22092 9860
rect 22156 9796 22200 9860
rect 22048 9752 22200 9796
rect 22260 10644 22304 10676
rect 22368 10676 22382 10708
rect 22368 10644 22412 10676
rect 18868 8556 18912 8588
rect 18898 8524 18912 8556
rect 18976 8556 19020 8588
rect 19080 9224 19232 9268
rect 19080 9160 19124 9224
rect 19188 9160 19232 9224
rect 18976 8524 18990 8556
rect 18898 8510 18990 8524
rect 19080 7740 19232 9160
rect 19080 7708 19124 7740
rect 19110 7676 19124 7708
rect 19188 7708 19232 7740
rect 19188 7676 19202 7708
rect 19110 7662 19202 7676
rect 18050 3500 18142 3514
rect 18050 3468 18064 3500
rect 18020 3436 18064 3468
rect 18128 3468 18142 3500
rect 18128 3436 18172 3468
rect 16142 2864 16234 2878
rect 16142 2832 16156 2864
rect 16112 2800 16156 2832
rect 16220 2832 16234 2864
rect 17626 2864 17718 2878
rect 17626 2832 17640 2864
rect 16220 2800 16264 2832
rect 16112 0 16264 2800
rect 17596 2800 17640 2832
rect 17704 2832 17718 2864
rect 17704 2800 17748 2832
rect 16778 2652 16870 2666
rect 16778 2620 16792 2652
rect 16748 2588 16792 2620
rect 16856 2620 16870 2652
rect 16856 2588 16900 2620
rect 16748 956 16900 2588
rect 16748 892 16792 956
rect 16856 892 16900 956
rect 16748 848 16900 892
rect 17596 0 17748 2800
rect 18020 2016 18172 3436
rect 19322 2864 19414 2878
rect 19322 2832 19336 2864
rect 18020 1952 18064 2016
rect 18128 1952 18172 2016
rect 18020 1908 18172 1952
rect 19292 2800 19336 2832
rect 19400 2832 19414 2864
rect 20594 2864 20686 2878
rect 20594 2832 20608 2864
rect 19400 2800 19444 2832
rect 19292 0 19444 2800
rect 20564 2800 20608 2832
rect 20672 2832 20686 2864
rect 22078 2864 22170 2878
rect 22078 2832 22092 2864
rect 20672 2800 20716 2832
rect 20564 0 20716 2800
rect 22048 2800 22092 2832
rect 22156 2832 22170 2864
rect 22156 2800 22200 2832
rect 22048 0 22200 2800
rect 22260 0 22412 10644
rect 22896 8376 23048 10856
rect 24804 10856 24848 10920
rect 24912 10856 24956 10920
rect 25046 10920 25138 10934
rect 25046 10888 25060 10920
rect 24804 9860 24956 10856
rect 24804 9828 24848 9860
rect 24834 9796 24848 9828
rect 24912 9828 24956 9860
rect 25016 10856 25060 10888
rect 25124 10888 25138 10920
rect 25228 10920 25380 11704
rect 28408 11704 28452 11736
rect 28516 11736 28530 11768
rect 31406 11768 31498 11782
rect 31406 11736 31420 11768
rect 28516 11704 28560 11736
rect 28226 11132 28318 11146
rect 28226 11100 28240 11132
rect 28196 11068 28240 11100
rect 28304 11100 28318 11132
rect 28408 11132 28560 11704
rect 28304 11068 28348 11100
rect 25124 10856 25168 10888
rect 25016 9860 25168 10856
rect 25228 10856 25272 10920
rect 25336 10856 25380 10920
rect 25894 10920 25986 10934
rect 25894 10888 25908 10920
rect 25228 10812 25380 10856
rect 25864 10856 25908 10888
rect 25972 10888 25986 10920
rect 27984 10920 28136 10964
rect 25972 10856 26016 10888
rect 25470 10708 25562 10722
rect 25470 10676 25484 10708
rect 24912 9796 24926 9828
rect 24834 9782 24926 9796
rect 25016 9796 25060 9860
rect 25124 9796 25168 9860
rect 25016 9752 25168 9796
rect 25440 10644 25484 10676
rect 25548 10676 25562 10708
rect 25548 10644 25592 10676
rect 22896 8312 22940 8376
rect 23004 8312 23048 8376
rect 22896 8268 23048 8312
rect 24198 3500 24290 3514
rect 24198 3468 24212 3500
rect 24168 3436 24212 3468
rect 24276 3468 24290 3500
rect 24276 3436 24320 3468
rect 23774 2864 23866 2878
rect 23774 2832 23788 2864
rect 23744 2800 23788 2832
rect 23852 2832 23866 2864
rect 23852 2800 23896 2832
rect 23744 0 23896 2800
rect 24168 2016 24320 3436
rect 25258 2864 25350 2878
rect 25258 2832 25272 2864
rect 24168 1952 24212 2016
rect 24276 1952 24320 2016
rect 24168 1908 24320 1952
rect 25228 2800 25272 2832
rect 25336 2832 25350 2864
rect 25336 2800 25380 2832
rect 25228 0 25380 2800
rect 25440 0 25592 10644
rect 25864 8376 26016 10856
rect 27984 10856 28028 10920
rect 28092 10856 28136 10920
rect 27984 9860 28136 10856
rect 27984 9828 28028 9860
rect 28014 9796 28028 9828
rect 28092 9828 28136 9860
rect 28196 9860 28348 11068
rect 28408 11068 28452 11132
rect 28516 11068 28560 11132
rect 28408 11024 28560 11068
rect 31376 11704 31420 11736
rect 31484 11736 31498 11768
rect 34586 11768 34678 11782
rect 34586 11736 34600 11768
rect 31484 11704 31528 11736
rect 28092 9796 28106 9828
rect 28014 9782 28106 9796
rect 28196 9796 28240 9860
rect 28304 9796 28348 9860
rect 28196 9752 28348 9796
rect 28408 10920 28560 10964
rect 28408 10856 28452 10920
rect 28516 10856 28560 10920
rect 30982 10920 31074 10934
rect 30982 10888 30996 10920
rect 28408 9692 28560 10856
rect 30952 10856 30996 10888
rect 31060 10888 31074 10920
rect 31164 10920 31316 10964
rect 31060 10856 31104 10888
rect 28650 10708 28742 10722
rect 28650 10676 28664 10708
rect 25864 8312 25908 8376
rect 25972 8312 26016 8376
rect 28196 9540 28560 9692
rect 28620 10644 28664 10676
rect 28728 10676 28742 10708
rect 28728 10644 28772 10676
rect 28196 8376 28348 9540
rect 28196 8344 28240 8376
rect 25864 8268 26016 8312
rect 28226 8312 28240 8344
rect 28304 8344 28348 8376
rect 28304 8312 28318 8344
rect 28226 8298 28318 8312
rect 26742 2864 26834 2878
rect 26742 2832 26756 2864
rect 26712 2800 26756 2832
rect 26820 2832 26834 2864
rect 28226 2864 28318 2878
rect 28226 2832 28240 2864
rect 26820 2800 26864 2832
rect 26712 0 26864 2800
rect 28196 2800 28240 2832
rect 28304 2832 28318 2864
rect 28304 2800 28348 2832
rect 28196 0 28348 2800
rect 28620 0 28772 10644
rect 30952 10072 31104 10856
rect 30952 10008 30996 10072
rect 31060 10008 31104 10072
rect 30952 9964 31104 10008
rect 31164 10856 31208 10920
rect 31272 10856 31316 10920
rect 31164 9860 31316 10856
rect 31376 10920 31528 11704
rect 34556 11704 34600 11736
rect 34664 11736 34678 11768
rect 37978 11768 38070 11782
rect 37978 11736 37992 11768
rect 34664 11704 34708 11736
rect 31376 10856 31420 10920
rect 31484 10856 31528 10920
rect 32254 10920 32346 10934
rect 32254 10888 32268 10920
rect 31376 10812 31528 10856
rect 32224 10856 32268 10888
rect 32332 10888 32346 10920
rect 34132 10920 34284 10964
rect 32332 10856 32376 10888
rect 31618 10708 31710 10722
rect 31618 10676 31632 10708
rect 31164 9828 31208 9860
rect 31194 9796 31208 9828
rect 31272 9828 31316 9860
rect 31588 10644 31632 10676
rect 31696 10676 31710 10708
rect 31696 10644 31740 10676
rect 31272 9796 31286 9828
rect 31194 9782 31286 9796
rect 28832 6468 28984 6512
rect 28832 6404 28876 6468
rect 28940 6404 28984 6468
rect 28832 3712 28984 6404
rect 28832 3680 28876 3712
rect 28862 3648 28876 3680
rect 28940 3680 28984 3712
rect 28940 3648 28954 3680
rect 28862 3634 28954 3648
rect 30134 3500 30226 3514
rect 30134 3468 30148 3500
rect 30104 3436 30148 3468
rect 30212 3468 30226 3500
rect 30212 3436 30256 3468
rect 29498 2864 29590 2878
rect 29498 2832 29512 2864
rect 29468 2800 29512 2832
rect 29576 2832 29590 2864
rect 29576 2800 29620 2832
rect 29468 0 29620 2800
rect 30104 2016 30256 3436
rect 30982 2864 31074 2878
rect 30982 2832 30996 2864
rect 30104 1952 30148 2016
rect 30212 1952 30256 2016
rect 30104 1908 30256 1952
rect 30952 2800 30996 2832
rect 31060 2832 31074 2864
rect 31060 2800 31104 2832
rect 30952 0 31104 2800
rect 31588 0 31740 10644
rect 32224 8376 32376 10856
rect 34132 10856 34176 10920
rect 34240 10856 34284 10920
rect 34132 9860 34284 10856
rect 34556 10920 34708 11704
rect 37948 11704 37992 11736
rect 38056 11736 38070 11768
rect 40734 11768 40826 11782
rect 40734 11736 40748 11768
rect 38056 11704 38100 11736
rect 34798 11132 34890 11146
rect 34798 11100 34812 11132
rect 34556 10856 34600 10920
rect 34664 10856 34708 10920
rect 34556 10812 34708 10856
rect 34768 11068 34812 11100
rect 34876 11100 34890 11132
rect 37766 11132 37858 11146
rect 37766 11100 37780 11132
rect 34876 11068 34920 11100
rect 34586 10708 34678 10722
rect 34586 10676 34600 10708
rect 34132 9828 34176 9860
rect 34162 9796 34176 9828
rect 34240 9828 34284 9860
rect 34556 10644 34600 10676
rect 34664 10676 34678 10708
rect 34664 10644 34708 10676
rect 34240 9796 34254 9828
rect 34162 9782 34254 9796
rect 32224 8312 32268 8376
rect 32332 8312 32376 8376
rect 32224 8268 32376 8312
rect 32466 2864 32558 2878
rect 32466 2832 32480 2864
rect 32436 2800 32480 2832
rect 32544 2832 32558 2864
rect 33950 2864 34042 2878
rect 33950 2832 33964 2864
rect 32544 2800 32588 2832
rect 32436 0 32588 2800
rect 33920 2800 33964 2832
rect 34028 2832 34042 2864
rect 34028 2800 34072 2832
rect 33920 0 34072 2800
rect 34556 0 34708 10644
rect 34768 9860 34920 11068
rect 37736 11068 37780 11100
rect 37844 11100 37858 11132
rect 37844 11068 37888 11100
rect 34768 9796 34812 9860
rect 34876 9796 34920 9860
rect 34768 9752 34920 9796
rect 34980 10920 35132 10964
rect 34980 10856 35024 10920
rect 35088 10856 35132 10920
rect 34980 8588 35132 10856
rect 37312 10920 37464 10964
rect 37312 10856 37356 10920
rect 37420 10856 37464 10920
rect 37312 9860 37464 10856
rect 37312 9828 37356 9860
rect 37342 9796 37356 9828
rect 37420 9828 37464 9860
rect 37736 9860 37888 11068
rect 37948 10920 38100 11704
rect 40704 11704 40748 11736
rect 40812 11736 40826 11768
rect 43914 11768 44006 11782
rect 43914 11736 43928 11768
rect 40812 11704 40856 11736
rect 37948 10856 37992 10920
rect 38056 10856 38100 10920
rect 38614 10920 38706 10934
rect 38614 10888 38628 10920
rect 37948 10812 38100 10856
rect 38584 10856 38628 10888
rect 38692 10888 38706 10920
rect 40310 10920 40402 10934
rect 40310 10888 40324 10920
rect 38692 10856 38736 10888
rect 37978 10708 38070 10722
rect 37978 10676 37992 10708
rect 37420 9796 37434 9828
rect 37342 9782 37434 9796
rect 37736 9796 37780 9860
rect 37844 9796 37888 9860
rect 37736 9752 37888 9796
rect 37948 10644 37992 10676
rect 38056 10676 38070 10708
rect 38056 10644 38100 10676
rect 34980 8556 35024 8588
rect 35010 8524 35024 8556
rect 35088 8556 35132 8588
rect 35088 8524 35102 8556
rect 35010 8510 35102 8524
rect 37342 3500 37434 3514
rect 37342 3468 37356 3500
rect 37312 3436 37356 3468
rect 37420 3468 37434 3500
rect 37420 3436 37464 3468
rect 35646 2864 35738 2878
rect 35646 2832 35660 2864
rect 35616 2800 35660 2832
rect 35724 2832 35738 2864
rect 36918 2864 37010 2878
rect 36918 2832 36932 2864
rect 35724 2800 35768 2832
rect 35616 0 35768 2800
rect 36888 2800 36932 2832
rect 36996 2832 37010 2864
rect 36996 2800 37040 2832
rect 36888 0 37040 2800
rect 37312 2016 37464 3436
rect 37312 1952 37356 2016
rect 37420 1952 37464 2016
rect 37312 1908 37464 1952
rect 37948 0 38100 10644
rect 38584 8376 38736 10856
rect 40280 10856 40324 10888
rect 40388 10888 40402 10920
rect 40492 10920 40644 10964
rect 40388 10856 40432 10888
rect 40280 10072 40432 10856
rect 40280 10008 40324 10072
rect 40388 10008 40432 10072
rect 40280 9964 40432 10008
rect 40492 10856 40536 10920
rect 40600 10856 40644 10920
rect 40492 9860 40644 10856
rect 40704 10920 40856 11704
rect 43884 11704 43928 11736
rect 43992 11736 44006 11768
rect 47094 11768 47186 11782
rect 47094 11736 47108 11768
rect 43992 11704 44036 11736
rect 40704 10856 40748 10920
rect 40812 10856 40856 10920
rect 41158 10920 41250 10934
rect 41158 10888 41172 10920
rect 40704 10812 40856 10856
rect 41128 10856 41172 10888
rect 41236 10888 41250 10920
rect 43460 10920 43612 10964
rect 41236 10856 41280 10888
rect 40946 10708 41038 10722
rect 40946 10676 40960 10708
rect 40492 9828 40536 9860
rect 40522 9796 40536 9828
rect 40600 9828 40644 9860
rect 40916 10644 40960 10676
rect 41024 10676 41038 10708
rect 41024 10644 41068 10676
rect 40600 9796 40614 9828
rect 40522 9782 40614 9796
rect 38584 8312 38628 8376
rect 38692 8312 38736 8376
rect 38584 8268 38736 8312
rect 40310 3500 40402 3514
rect 40310 3468 40324 3500
rect 40280 3436 40324 3468
rect 40388 3468 40402 3500
rect 40388 3436 40432 3468
rect 38614 2864 38706 2878
rect 38614 2832 38628 2864
rect 38584 2800 38628 2832
rect 38692 2832 38706 2864
rect 39886 2864 39978 2878
rect 39886 2832 39900 2864
rect 38692 2800 38736 2832
rect 38584 0 38736 2800
rect 39856 2800 39900 2832
rect 39964 2832 39978 2864
rect 39964 2800 40008 2832
rect 39856 0 40008 2800
rect 40280 2016 40432 3436
rect 40280 1952 40324 2016
rect 40388 1952 40432 2016
rect 40280 1908 40432 1952
rect 40916 0 41068 10644
rect 41128 8376 41280 10856
rect 43460 10856 43504 10920
rect 43568 10856 43612 10920
rect 43460 9860 43612 10856
rect 43884 10920 44036 11704
rect 47064 11704 47108 11736
rect 47172 11736 47186 11768
rect 50486 11768 50578 11782
rect 50486 11736 50500 11768
rect 47172 11704 47216 11736
rect 44126 11132 44218 11146
rect 44126 11100 44140 11132
rect 43884 10856 43928 10920
rect 43992 10856 44036 10920
rect 43884 10812 44036 10856
rect 44096 11068 44140 11100
rect 44204 11100 44218 11132
rect 44204 11068 44248 11100
rect 43914 10708 44006 10722
rect 43914 10676 43928 10708
rect 43460 9828 43504 9860
rect 43490 9796 43504 9828
rect 43568 9828 43612 9860
rect 43884 10644 43928 10676
rect 43992 10676 44006 10708
rect 43992 10644 44036 10676
rect 43568 9796 43582 9828
rect 43490 9782 43582 9796
rect 41128 8312 41172 8376
rect 41236 8312 41280 8376
rect 41128 8268 41280 8312
rect 41582 2864 41674 2878
rect 41582 2832 41596 2864
rect 41552 2800 41596 2832
rect 41660 2832 41674 2864
rect 41660 2800 41704 2832
rect 41552 0 41704 2800
rect 43884 0 44036 10644
rect 44096 9860 44248 11068
rect 44762 10920 44854 10934
rect 44762 10888 44776 10920
rect 44096 9796 44140 9860
rect 44204 9796 44248 9860
rect 44096 9752 44248 9796
rect 44732 10856 44776 10888
rect 44840 10888 44854 10920
rect 46458 10920 46550 10934
rect 46458 10888 46472 10920
rect 44840 10856 44884 10888
rect 44732 8376 44884 10856
rect 46428 10856 46472 10888
rect 46536 10888 46550 10920
rect 46640 10920 46792 10964
rect 46536 10856 46580 10888
rect 46428 10072 46580 10856
rect 46428 10008 46472 10072
rect 46536 10008 46580 10072
rect 46428 9964 46580 10008
rect 46640 10856 46684 10920
rect 46748 10856 46792 10920
rect 46640 9860 46792 10856
rect 47064 10920 47216 11704
rect 50456 11704 50500 11736
rect 50564 11736 50578 11768
rect 53242 11768 53334 11782
rect 53242 11736 53256 11768
rect 50564 11704 50608 11736
rect 49608 11344 49760 11388
rect 49608 11280 49652 11344
rect 49716 11280 49760 11344
rect 50274 11344 50366 11358
rect 50274 11312 50288 11344
rect 47064 10856 47108 10920
rect 47172 10856 47216 10920
rect 47518 10920 47610 10934
rect 47518 10888 47532 10920
rect 47064 10812 47216 10856
rect 47488 10856 47532 10888
rect 47596 10888 47610 10920
rect 47596 10856 47640 10888
rect 47094 10708 47186 10722
rect 47094 10676 47108 10708
rect 46640 9828 46684 9860
rect 46670 9796 46684 9828
rect 46748 9828 46792 9860
rect 47064 10644 47108 10676
rect 47172 10676 47186 10708
rect 47172 10644 47216 10676
rect 46748 9796 46762 9828
rect 46670 9782 46762 9796
rect 44732 8312 44776 8376
rect 44840 8312 44884 8376
rect 44732 8268 44884 8312
rect 47064 0 47216 10644
rect 47488 8376 47640 10856
rect 47488 8312 47532 8376
rect 47596 8312 47640 8376
rect 49608 8376 49760 11280
rect 50244 11280 50288 11312
rect 50352 11312 50366 11344
rect 50352 11280 50396 11312
rect 50062 11132 50154 11146
rect 50062 11100 50076 11132
rect 50032 11068 50076 11100
rect 50140 11100 50154 11132
rect 50140 11068 50184 11100
rect 49820 10920 49972 10964
rect 49820 10856 49864 10920
rect 49928 10856 49972 10920
rect 49820 9860 49972 10856
rect 49820 9828 49864 9860
rect 49850 9796 49864 9828
rect 49928 9828 49972 9860
rect 50032 9860 50184 11068
rect 50244 10920 50396 11280
rect 50244 10856 50288 10920
rect 50352 10856 50396 10920
rect 50244 10812 50396 10856
rect 50456 10920 50608 11704
rect 53212 11704 53256 11736
rect 53320 11736 53334 11768
rect 56846 11768 56938 11782
rect 56846 11736 56860 11768
rect 53320 11704 53364 11736
rect 50456 10856 50500 10920
rect 50564 10856 50608 10920
rect 50456 10812 50608 10856
rect 52788 10920 52940 10964
rect 52788 10856 52832 10920
rect 52896 10856 52940 10920
rect 53030 10920 53122 10934
rect 53030 10888 53044 10920
rect 50486 10708 50578 10722
rect 50486 10676 50500 10708
rect 49928 9796 49942 9828
rect 49850 9782 49942 9796
rect 50032 9796 50076 9860
rect 50140 9796 50184 9860
rect 50032 9752 50184 9796
rect 50456 10644 50500 10676
rect 50564 10676 50578 10708
rect 50564 10644 50608 10676
rect 49608 8344 49652 8376
rect 47488 8268 47640 8312
rect 49638 8312 49652 8344
rect 49716 8344 49760 8376
rect 49716 8312 49730 8344
rect 49638 8298 49730 8312
rect 50456 0 50608 10644
rect 52788 9860 52940 10856
rect 52788 9828 52832 9860
rect 52818 9796 52832 9828
rect 52896 9828 52940 9860
rect 53000 10856 53044 10888
rect 53108 10888 53122 10920
rect 53212 10920 53364 11704
rect 56816 11704 56860 11736
rect 56924 11736 56938 11768
rect 59602 11768 59694 11782
rect 59602 11736 59616 11768
rect 56924 11704 56968 11736
rect 55756 11344 55908 11388
rect 55756 11280 55800 11344
rect 55864 11280 55908 11344
rect 56422 11344 56514 11358
rect 56422 11312 56436 11344
rect 53108 10856 53152 10888
rect 53000 9860 53152 10856
rect 53212 10856 53256 10920
rect 53320 10856 53364 10920
rect 53212 10812 53364 10856
rect 53424 10920 53576 10964
rect 53424 10856 53468 10920
rect 53532 10856 53576 10920
rect 53242 10708 53334 10722
rect 53242 10676 53256 10708
rect 52896 9796 52910 9828
rect 52818 9782 52910 9796
rect 53000 9796 53044 9860
rect 53108 9796 53152 9860
rect 53000 9752 53152 9796
rect 53212 10644 53256 10676
rect 53320 10676 53334 10708
rect 53320 10644 53364 10676
rect 53212 0 53364 10644
rect 53424 8588 53576 10856
rect 53424 8556 53468 8588
rect 53454 8524 53468 8556
rect 53532 8556 53576 8588
rect 53532 8524 53546 8556
rect 53454 8510 53546 8524
rect 55756 8376 55908 11280
rect 56392 11280 56436 11312
rect 56500 11312 56514 11344
rect 56500 11280 56544 11312
rect 55968 10920 56120 10964
rect 55968 10856 56012 10920
rect 56076 10856 56120 10920
rect 55968 9860 56120 10856
rect 56392 10920 56544 11280
rect 56634 11132 56726 11146
rect 56634 11100 56648 11132
rect 56392 10856 56436 10920
rect 56500 10856 56544 10920
rect 56392 10812 56544 10856
rect 56604 11068 56648 11100
rect 56712 11100 56726 11132
rect 56712 11068 56756 11100
rect 56422 10708 56514 10722
rect 56422 10676 56436 10708
rect 55968 9828 56012 9860
rect 55998 9796 56012 9828
rect 56076 9828 56120 9860
rect 56392 10644 56436 10676
rect 56500 10676 56514 10708
rect 56500 10644 56544 10676
rect 56076 9796 56090 9828
rect 55998 9782 56090 9796
rect 55756 8344 55800 8376
rect 55786 8312 55800 8344
rect 55864 8344 55908 8376
rect 55864 8312 55878 8344
rect 55786 8298 55878 8312
rect 56392 0 56544 10644
rect 56604 9860 56756 11068
rect 56816 10920 56968 11704
rect 59572 11704 59616 11736
rect 59680 11736 59694 11768
rect 62570 11768 62662 11782
rect 62570 11736 62584 11768
rect 59680 11704 59724 11736
rect 59390 11132 59482 11146
rect 59390 11100 59404 11132
rect 56816 10856 56860 10920
rect 56924 10856 56968 10920
rect 56816 10812 56968 10856
rect 59360 11068 59404 11100
rect 59468 11100 59482 11132
rect 59468 11068 59512 11100
rect 56604 9796 56648 9860
rect 56712 9796 56756 9860
rect 56604 9752 56756 9796
rect 59360 9860 59512 11068
rect 59572 10920 59724 11704
rect 62540 11704 62584 11736
rect 62648 11736 62662 11768
rect 65750 11768 65842 11782
rect 65750 11736 65764 11768
rect 62648 11704 62692 11736
rect 59572 10856 59616 10920
rect 59680 10856 59724 10920
rect 60026 10920 60118 10934
rect 60026 10888 60040 10920
rect 59572 10812 59724 10856
rect 59996 10856 60040 10888
rect 60104 10888 60118 10920
rect 62116 10920 62268 10964
rect 60104 10856 60148 10888
rect 59814 10708 59906 10722
rect 59814 10676 59828 10708
rect 59360 9796 59404 9860
rect 59468 9796 59512 9860
rect 59360 9752 59512 9796
rect 59784 10644 59828 10676
rect 59892 10676 59906 10708
rect 59892 10644 59936 10676
rect 59784 0 59936 10644
rect 59996 8376 60148 10856
rect 62116 10856 62160 10920
rect 62224 10856 62268 10920
rect 62116 9860 62268 10856
rect 62540 10920 62692 11704
rect 65720 11704 65764 11736
rect 65828 11736 65842 11768
rect 68718 11768 68810 11782
rect 68718 11736 68732 11768
rect 65828 11704 65872 11736
rect 62782 11132 62874 11146
rect 62782 11100 62796 11132
rect 62540 10856 62584 10920
rect 62648 10856 62692 10920
rect 62540 10812 62692 10856
rect 62752 11068 62796 11100
rect 62860 11100 62874 11132
rect 62860 11068 62904 11100
rect 62570 10708 62662 10722
rect 62570 10676 62584 10708
rect 62116 9828 62160 9860
rect 62146 9796 62160 9828
rect 62224 9828 62268 9860
rect 62540 10644 62584 10676
rect 62648 10676 62662 10708
rect 62648 10644 62692 10676
rect 62224 9796 62238 9828
rect 62146 9782 62238 9796
rect 59996 8312 60040 8376
rect 60104 8312 60148 8376
rect 59996 8268 60148 8312
rect 62540 0 62692 10644
rect 62752 9860 62904 11068
rect 62994 10920 63086 10934
rect 62994 10888 63008 10920
rect 62752 9796 62796 9860
rect 62860 9796 62904 9860
rect 62752 9752 62904 9796
rect 62964 10856 63008 10888
rect 63072 10888 63086 10920
rect 65296 10920 65448 10964
rect 63072 10856 63116 10888
rect 62964 8376 63116 10856
rect 65296 10856 65340 10920
rect 65404 10856 65448 10920
rect 65296 9860 65448 10856
rect 65720 10920 65872 11704
rect 68688 11704 68732 11736
rect 68796 11736 68810 11768
rect 68796 11704 68840 11736
rect 65962 11132 66054 11146
rect 65962 11100 65976 11132
rect 65720 10856 65764 10920
rect 65828 10856 65872 10920
rect 65720 10812 65872 10856
rect 65932 11068 65976 11100
rect 66040 11100 66054 11132
rect 66040 11068 66084 11100
rect 65750 10708 65842 10722
rect 65750 10676 65764 10708
rect 65296 9828 65340 9860
rect 65326 9796 65340 9828
rect 65404 9828 65448 9860
rect 65720 10644 65764 10676
rect 65828 10676 65842 10708
rect 65828 10644 65872 10676
rect 65404 9796 65418 9828
rect 65326 9782 65418 9796
rect 62964 8312 63008 8376
rect 63072 8312 63116 8376
rect 62964 8268 63116 8312
rect 65720 0 65872 10644
rect 65932 9860 66084 11068
rect 66598 10920 66690 10934
rect 66598 10888 66612 10920
rect 65932 9796 65976 9860
rect 66040 9796 66084 9860
rect 65932 9752 66084 9796
rect 66568 10856 66612 10888
rect 66676 10888 66690 10920
rect 68294 10920 68386 10934
rect 68294 10888 68308 10920
rect 66676 10856 66720 10888
rect 66568 8376 66720 10856
rect 68264 10856 68308 10888
rect 68372 10888 68386 10920
rect 68476 10920 68628 10964
rect 68372 10856 68416 10888
rect 68264 10072 68416 10856
rect 68264 10008 68308 10072
rect 68372 10008 68416 10072
rect 68264 9964 68416 10008
rect 68476 10856 68520 10920
rect 68584 10856 68628 10920
rect 68476 9860 68628 10856
rect 68688 10920 68840 11704
rect 68688 10856 68732 10920
rect 68796 10856 68840 10920
rect 68688 10812 68840 10856
rect 69112 10920 69264 10964
rect 69112 10856 69156 10920
rect 69220 10856 69264 10920
rect 68930 10708 69022 10722
rect 68930 10676 68944 10708
rect 68476 9828 68520 9860
rect 68506 9796 68520 9828
rect 68584 9828 68628 9860
rect 68900 10644 68944 10676
rect 69008 10676 69022 10708
rect 69008 10644 69052 10676
rect 68584 9796 68598 9828
rect 68506 9782 68598 9796
rect 66568 8312 66612 8376
rect 66676 8312 66720 8376
rect 66568 8268 66720 8312
rect 68900 0 69052 10644
rect 69112 8588 69264 10856
rect 69112 8556 69156 8588
rect 69142 8524 69156 8556
rect 69220 8556 69264 8588
rect 71868 10708 72020 10752
rect 71868 10644 71912 10708
rect 71976 10644 72020 10708
rect 69220 8524 69234 8556
rect 69142 8510 69234 8524
rect 71868 8376 72020 10644
rect 71868 8344 71912 8376
rect 71898 8312 71912 8344
rect 71976 8344 72020 8376
rect 119568 9860 120144 61948
rect 119568 9796 119612 9860
rect 119676 9796 120144 9860
rect 71976 8312 71990 8344
rect 71898 8298 71990 8312
rect 119568 2016 120144 9796
rect 119568 1952 119612 2016
rect 119676 1952 119824 2016
rect 119888 1952 120036 2016
rect 120100 1952 120144 2016
rect 119568 1804 120144 1952
rect 119568 1740 119612 1804
rect 119676 1740 119824 1804
rect 119888 1740 120036 1804
rect 120100 1740 120144 1804
rect 119568 1592 120144 1740
rect 119568 1528 119612 1592
rect 119676 1528 119824 1592
rect 119888 1528 120036 1592
rect 120100 1528 120144 1592
rect 119568 1484 120144 1528
rect 120628 10920 121204 63008
rect 120628 10856 120672 10920
rect 120736 10856 121204 10920
rect 120628 956 121204 10856
rect 120628 892 120672 956
rect 120736 892 120884 956
rect 120948 892 121096 956
rect 121160 892 121204 956
rect 120628 744 121204 892
rect 120628 680 120672 744
rect 120736 680 120884 744
rect 120948 680 121096 744
rect 121160 680 121204 744
rect 120628 532 121204 680
rect 120628 468 120672 532
rect 120736 468 120884 532
rect 120948 468 121096 532
rect 121160 468 121204 532
rect 120628 424 121204 468
use contact_31  contact_31_0
timestamp 1643678851
transform 1 0 120628 0 1 10842
box 0 0 1 1
use contact_31  contact_31_1
timestamp 1643678851
transform 1 0 71868 0 1 10630
box 0 0 1 1
use contact_31  contact_31_2
timestamp 1643678851
transform 1 0 71868 0 1 8298
box 0 0 1 1
use contact_31  contact_31_3
timestamp 1643678851
transform 1 0 68688 0 1 10842
box 0 0 1 1
use contact_31  contact_31_4
timestamp 1643678851
transform 1 0 68688 0 1 11690
box 0 0 1 1
use contact_31  contact_31_5
timestamp 1643678851
transform 1 0 69112 0 1 10842
box 0 0 1 1
use contact_31  contact_31_6
timestamp 1643678851
transform 1 0 69112 0 1 8510
box 0 0 1 1
use contact_31  contact_31_7
timestamp 1643678851
transform 1 0 66568 0 1 8298
box 0 0 1 1
use contact_31  contact_31_8
timestamp 1643678851
transform 1 0 66568 0 1 10842
box 0 0 1 1
use contact_31  contact_31_9
timestamp 1643678851
transform 1 0 65720 0 1 10842
box 0 0 1 1
use contact_31  contact_31_10
timestamp 1643678851
transform 1 0 65720 0 1 11690
box 0 0 1 1
use contact_31  contact_31_11
timestamp 1643678851
transform 1 0 62964 0 1 8298
box 0 0 1 1
use contact_31  contact_31_12
timestamp 1643678851
transform 1 0 62964 0 1 10842
box 0 0 1 1
use contact_31  contact_31_13
timestamp 1643678851
transform 1 0 62540 0 1 10842
box 0 0 1 1
use contact_31  contact_31_14
timestamp 1643678851
transform 1 0 62540 0 1 11690
box 0 0 1 1
use contact_31  contact_31_15
timestamp 1643678851
transform 1 0 59996 0 1 8298
box 0 0 1 1
use contact_31  contact_31_16
timestamp 1643678851
transform 1 0 59996 0 1 10842
box 0 0 1 1
use contact_31  contact_31_17
timestamp 1643678851
transform 1 0 59572 0 1 10842
box 0 0 1 1
use contact_31  contact_31_18
timestamp 1643678851
transform 1 0 59572 0 1 11690
box 0 0 1 1
use contact_31  contact_31_19
timestamp 1643678851
transform 1 0 56816 0 1 10842
box 0 0 1 1
use contact_31  contact_31_20
timestamp 1643678851
transform 1 0 56816 0 1 11690
box 0 0 1 1
use contact_31  contact_31_21
timestamp 1643678851
transform 1 0 56392 0 1 10842
box 0 0 1 1
use contact_31  contact_31_22
timestamp 1643678851
transform 1 0 56392 0 1 11266
box 0 0 1 1
use contact_31  contact_31_23
timestamp 1643678851
transform 1 0 55756 0 1 11266
box 0 0 1 1
use contact_31  contact_31_24
timestamp 1643678851
transform 1 0 55756 0 1 8298
box 0 0 1 1
use contact_31  contact_31_25
timestamp 1643678851
transform 1 0 53212 0 1 10842
box 0 0 1 1
use contact_31  contact_31_26
timestamp 1643678851
transform 1 0 53212 0 1 11690
box 0 0 1 1
use contact_31  contact_31_27
timestamp 1643678851
transform 1 0 53424 0 1 10842
box 0 0 1 1
use contact_31  contact_31_28
timestamp 1643678851
transform 1 0 53424 0 1 8510
box 0 0 1 1
use contact_31  contact_31_29
timestamp 1643678851
transform 1 0 50456 0 1 10842
box 0 0 1 1
use contact_31  contact_31_30
timestamp 1643678851
transform 1 0 50456 0 1 11690
box 0 0 1 1
use contact_31  contact_31_31
timestamp 1643678851
transform 1 0 50244 0 1 10842
box 0 0 1 1
use contact_31  contact_31_32
timestamp 1643678851
transform 1 0 50244 0 1 11266
box 0 0 1 1
use contact_31  contact_31_33
timestamp 1643678851
transform 1 0 49608 0 1 11266
box 0 0 1 1
use contact_31  contact_31_34
timestamp 1643678851
transform 1 0 49608 0 1 8298
box 0 0 1 1
use contact_31  contact_31_35
timestamp 1643678851
transform 1 0 47488 0 1 8298
box 0 0 1 1
use contact_31  contact_31_36
timestamp 1643678851
transform 1 0 47488 0 1 10842
box 0 0 1 1
use contact_31  contact_31_37
timestamp 1643678851
transform 1 0 47064 0 1 10842
box 0 0 1 1
use contact_31  contact_31_38
timestamp 1643678851
transform 1 0 47064 0 1 11690
box 0 0 1 1
use contact_31  contact_31_39
timestamp 1643678851
transform 1 0 44732 0 1 8298
box 0 0 1 1
use contact_31  contact_31_40
timestamp 1643678851
transform 1 0 44732 0 1 10842
box 0 0 1 1
use contact_31  contact_31_41
timestamp 1643678851
transform 1 0 43884 0 1 10842
box 0 0 1 1
use contact_31  contact_31_42
timestamp 1643678851
transform 1 0 43884 0 1 11690
box 0 0 1 1
use contact_31  contact_31_43
timestamp 1643678851
transform 1 0 41128 0 1 8298
box 0 0 1 1
use contact_31  contact_31_44
timestamp 1643678851
transform 1 0 41128 0 1 10842
box 0 0 1 1
use contact_31  contact_31_45
timestamp 1643678851
transform 1 0 40704 0 1 10842
box 0 0 1 1
use contact_31  contact_31_46
timestamp 1643678851
transform 1 0 40704 0 1 11690
box 0 0 1 1
use contact_31  contact_31_47
timestamp 1643678851
transform 1 0 38584 0 1 8298
box 0 0 1 1
use contact_31  contact_31_48
timestamp 1643678851
transform 1 0 38584 0 1 10842
box 0 0 1 1
use contact_31  contact_31_49
timestamp 1643678851
transform 1 0 37948 0 1 10842
box 0 0 1 1
use contact_31  contact_31_50
timestamp 1643678851
transform 1 0 37948 0 1 11690
box 0 0 1 1
use contact_31  contact_31_51
timestamp 1643678851
transform 1 0 34556 0 1 10842
box 0 0 1 1
use contact_31  contact_31_52
timestamp 1643678851
transform 1 0 34556 0 1 11690
box 0 0 1 1
use contact_31  contact_31_53
timestamp 1643678851
transform 1 0 34980 0 1 10842
box 0 0 1 1
use contact_31  contact_31_54
timestamp 1643678851
transform 1 0 34980 0 1 8510
box 0 0 1 1
use contact_31  contact_31_55
timestamp 1643678851
transform 1 0 32224 0 1 8298
box 0 0 1 1
use contact_31  contact_31_56
timestamp 1643678851
transform 1 0 32224 0 1 10842
box 0 0 1 1
use contact_31  contact_31_57
timestamp 1643678851
transform 1 0 31376 0 1 10842
box 0 0 1 1
use contact_31  contact_31_58
timestamp 1643678851
transform 1 0 31376 0 1 11690
box 0 0 1 1
use contact_31  contact_31_59
timestamp 1643678851
transform 1 0 28408 0 1 11054
box 0 0 1 1
use contact_31  contact_31_60
timestamp 1643678851
transform 1 0 28408 0 1 11690
box 0 0 1 1
use contact_31  contact_31_61
timestamp 1643678851
transform 1 0 28408 0 1 10842
box 0 0 1 1
use contact_31  contact_31_62
timestamp 1643678851
transform 1 0 28196 0 1 8298
box 0 0 1 1
use contact_31  contact_31_63
timestamp 1643678851
transform 1 0 25864 0 1 8298
box 0 0 1 1
use contact_31  contact_31_64
timestamp 1643678851
transform 1 0 25864 0 1 10842
box 0 0 1 1
use contact_31  contact_31_65
timestamp 1643678851
transform 1 0 25228 0 1 10842
box 0 0 1 1
use contact_31  contact_31_66
timestamp 1643678851
transform 1 0 25228 0 1 11690
box 0 0 1 1
use contact_31  contact_31_67
timestamp 1643678851
transform 1 0 22896 0 1 8298
box 0 0 1 1
use contact_31  contact_31_68
timestamp 1643678851
transform 1 0 22896 0 1 10842
box 0 0 1 1
use contact_31  contact_31_69
timestamp 1643678851
transform 1 0 22260 0 1 10842
box 0 0 1 1
use contact_31  contact_31_70
timestamp 1643678851
transform 1 0 22260 0 1 11690
box 0 0 1 1
use contact_31  contact_31_71
timestamp 1643678851
transform 1 0 21412 0 1 62994
box 0 0 1 1
use contact_31  contact_31_72
timestamp 1643678851
transform 1 0 21412 0 1 61298
box 0 0 1 1
use contact_31  contact_31_73
timestamp 1643678851
transform 1 0 21200 0 1 24198
box 0 0 1 1
use contact_31  contact_31_74
timestamp 1643678851
transform 1 0 20988 0 1 21230
box 0 0 1 1
use contact_31  contact_31_75
timestamp 1643678851
transform 1 0 21412 0 1 18262
box 0 0 1 1
use contact_31  contact_31_76
timestamp 1643678851
transform 1 0 21412 0 1 21230
box 0 0 1 1
use contact_31  contact_31_77
timestamp 1643678851
transform 1 0 20140 0 1 15294
box 0 0 1 1
use contact_31  contact_31_78
timestamp 1643678851
transform 1 0 20140 0 1 18050
box 0 0 1 1
use contact_31  contact_31_79
timestamp 1643678851
transform 1 0 20988 0 1 55150
box 0 0 1 1
use contact_31  contact_31_80
timestamp 1643678851
transform 1 0 20988 0 1 57270
box 0 0 1 1
use contact_31  contact_31_81
timestamp 1643678851
transform 1 0 19928 0 1 49002
box 0 0 1 1
use contact_31  contact_31_82
timestamp 1643678851
transform 1 0 19928 0 1 51334
box 0 0 1 1
use contact_31  contact_31_83
timestamp 1643678851
transform 1 0 20988 0 1 51970
box 0 0 1 1
use contact_31  contact_31_84
timestamp 1643678851
transform 1 0 20988 0 1 54302
box 0 0 1 1
use contact_31  contact_31_85
timestamp 1643678851
transform 1 0 21200 0 1 12114
box 0 0 1 1
use contact_31  contact_31_86
timestamp 1643678851
transform 1 0 21200 0 1 14870
box 0 0 1 1
use contact_31  contact_31_87
timestamp 1643678851
transform 1 0 20140 0 1 36706
box 0 0 1 1
use contact_31  contact_31_88
timestamp 1643678851
transform 1 0 20140 0 1 39250
box 0 0 1 1
use contact_31  contact_31_89
timestamp 1643678851
transform 1 0 20988 0 1 30558
box 0 0 1 1
use contact_31  contact_31_90
timestamp 1643678851
transform 1 0 20988 0 1 33102
box 0 0 1 1
use contact_31  contact_31_91
timestamp 1643678851
transform 1 0 19928 0 1 39674
box 0 0 1 1
use contact_31  contact_31_92
timestamp 1643678851
transform 1 0 19928 0 1 42218
box 0 0 1 1
use contact_31  contact_31_93
timestamp 1643678851
transform 1 0 20140 0 1 61086
box 0 0 1 1
use contact_31  contact_31_94
timestamp 1643678851
transform 1 0 20140 0 1 60450
box 0 0 1 1
use contact_31  contact_31_95
timestamp 1643678851
transform 1 0 20988 0 1 58118
box 0 0 1 1
use contact_31  contact_31_96
timestamp 1643678851
transform 1 0 20988 0 1 60450
box 0 0 1 1
use contact_31  contact_31_97
timestamp 1643678851
transform 1 0 21200 0 1 24410
box 0 0 1 1
use contact_31  contact_31_98
timestamp 1643678851
transform 1 0 21200 0 1 26954
box 0 0 1 1
use contact_31  contact_31_99
timestamp 1643678851
transform 1 0 21200 0 1 48790
box 0 0 1 1
use contact_31  contact_31_100
timestamp 1643678851
transform 1 0 21200 0 1 48366
box 0 0 1 1
use contact_31  contact_31_101
timestamp 1643678851
transform 1 0 20988 0 1 45822
box 0 0 1 1
use contact_31  contact_31_102
timestamp 1643678851
transform 1 0 20988 0 1 48154
box 0 0 1 1
use contact_31  contact_31_103
timestamp 1643678851
transform 1 0 20988 0 1 42854
box 0 0 1 1
use contact_31  contact_31_104
timestamp 1643678851
transform 1 0 20988 0 1 45186
box 0 0 1 1
use contact_31  contact_31_105
timestamp 1643678851
transform 1 0 20988 0 1 27378
box 0 0 1 1
use contact_31  contact_31_106
timestamp 1643678851
transform 1 0 20988 0 1 30134
box 0 0 1 1
use contact_31  contact_31_107
timestamp 1643678851
transform 1 0 20988 0 1 33526
box 0 0 1 1
use contact_31  contact_31_108
timestamp 1643678851
transform 1 0 20988 0 1 36070
box 0 0 1 1
use contact_31  contact_31_109
timestamp 1643678851
transform 1 0 19928 0 1 11902
box 0 0 1 1
use contact_31  contact_31_110
timestamp 1643678851
transform 1 0 19928 0 1 11054
box 0 0 1 1
use contact_31  contact_31_111
timestamp 1643678851
transform 1 0 19080 0 1 9146
box 0 0 1 1
use contact_31  contact_31_112
timestamp 1643678851
transform 1 0 19080 0 1 7662
box 0 0 1 1
use contact_31  contact_31_113
timestamp 1643678851
transform 1 0 18020 0 1 9358
box 0 0 1 1
use contact_31  contact_31_114
timestamp 1643678851
transform 1 0 18020 0 1 10842
box 0 0 1 1
use contact_31  contact_31_115
timestamp 1643678851
transform 1 0 16748 0 1 878
box 0 0 1 1
use contact_31  contact_31_116
timestamp 1643678851
transform 1 0 16748 0 1 2574
box 0 0 1 1
use contact_31  contact_31_117
timestamp 1643678851
transform 1 0 16960 0 1 11054
box 0 0 1 1
use contact_31  contact_31_118
timestamp 1643678851
transform 1 0 16960 0 1 11902
box 0 0 1 1
use contact_31  contact_31_119
timestamp 1643678851
transform 1 0 16324 0 1 24198
box 0 0 1 1
use contact_31  contact_31_120
timestamp 1643678851
transform 1 0 16324 0 1 21230
box 0 0 1 1
use contact_31  contact_31_121
timestamp 1643678851
transform 1 0 16112 0 1 18262
box 0 0 1 1
use contact_31  contact_31_122
timestamp 1643678851
transform 1 0 16112 0 1 21230
box 0 0 1 1
use contact_31  contact_31_123
timestamp 1643678851
transform 1 0 16324 0 1 24410
box 0 0 1 1
use contact_31  contact_31_124
timestamp 1643678851
transform 1 0 16324 0 1 27166
box 0 0 1 1
use contact_31  contact_31_125
timestamp 1643678851
transform 1 0 16324 0 1 36494
box 0 0 1 1
use contact_31  contact_31_126
timestamp 1643678851
transform 1 0 16324 0 1 34798
box 0 0 1 1
use contact_31  contact_31_127
timestamp 1643678851
transform 1 0 15476 0 1 34798
box 0 0 1 1
use contact_31  contact_31_128
timestamp 1643678851
transform 1 0 15476 0 1 33526
box 0 0 1 1
use contact_31  contact_31_129
timestamp 1643678851
transform 1 0 16324 0 1 30558
box 0 0 1 1
use contact_31  contact_31_130
timestamp 1643678851
transform 1 0 16112 0 1 33526
box 0 0 1 1
use contact_31  contact_31_131
timestamp 1643678851
transform 1 0 16324 0 1 39674
box 0 0 1 1
use contact_31  contact_31_132
timestamp 1643678851
transform 1 0 16112 0 1 36706
box 0 0 1 1
use contact_31  contact_31_133
timestamp 1643678851
transform 1 0 16112 0 1 42642
box 0 0 1 1
use contact_31  contact_31_134
timestamp 1643678851
transform 1 0 16112 0 1 39674
box 0 0 1 1
use contact_31  contact_31_135
timestamp 1643678851
transform 1 0 16112 0 1 27378
box 0 0 1 1
use contact_31  contact_31_136
timestamp 1643678851
transform 1 0 16112 0 1 30346
box 0 0 1 1
use contact_31  contact_31_137
timestamp 1643678851
transform 1 0 13992 0 1 16990
box 0 0 1 1
use contact_31  contact_31_138
timestamp 1643678851
transform 1 0 13992 0 1 15506
box 0 0 1 1
use contact_31  contact_31_139
timestamp 1643678851
transform 1 0 15688 0 1 18262
box 0 0 1 1
use contact_31  contact_31_140
timestamp 1643678851
transform 1 0 15688 0 1 18686
box 0 0 1 1
use contact_31  contact_31_141
timestamp 1643678851
transform 1 0 13780 0 1 17202
box 0 0 1 1
use contact_31  contact_31_142
timestamp 1643678851
transform 1 0 13780 0 1 18686
box 0 0 1 1
use contact_31  contact_31_143
timestamp 1643678851
transform 1 0 13992 0 1 15294
box 0 0 1 1
use contact_31  contact_31_144
timestamp 1643678851
transform 1 0 13992 0 1 13810
box 0 0 1 1
use contact_31  contact_31_145
timestamp 1643678851
transform 1 0 13780 0 1 12114
box 0 0 1 1
use contact_31  contact_31_146
timestamp 1643678851
transform 1 0 13780 0 1 13810
box 0 0 1 1
use contact_31  contact_31_147
timestamp 1643678851
transform 1 0 848 0 1 7662
box 0 0 1 1
use contact_31  contact_31_148
timestamp 1643678851
transform 1 0 2544 0 1 5966
box 0 0 1 1
use contact_31  contact_31_149
timestamp 1643678851
transform 1 0 2544 0 1 7662
box 0 0 1 1
use contact_31  contact_31_150
timestamp 1643678851
transform 1 0 119568 0 1 9782
box 0 0 1 1
use contact_31  contact_31_151
timestamp 1643678851
transform 1 0 68264 0 1 9994
box 0 0 1 1
use contact_31  contact_31_152
timestamp 1643678851
transform 1 0 68264 0 1 10842
box 0 0 1 1
use contact_31  contact_31_153
timestamp 1643678851
transform 1 0 68476 0 1 10842
box 0 0 1 1
use contact_31  contact_31_154
timestamp 1643678851
transform 1 0 68476 0 1 9782
box 0 0 1 1
use contact_31  contact_31_155
timestamp 1643678851
transform 1 0 65932 0 1 9782
box 0 0 1 1
use contact_31  contact_31_156
timestamp 1643678851
transform 1 0 65932 0 1 11054
box 0 0 1 1
use contact_31  contact_31_157
timestamp 1643678851
transform 1 0 65296 0 1 10842
box 0 0 1 1
use contact_31  contact_31_158
timestamp 1643678851
transform 1 0 65296 0 1 9782
box 0 0 1 1
use contact_31  contact_31_159
timestamp 1643678851
transform 1 0 62752 0 1 9782
box 0 0 1 1
use contact_31  contact_31_160
timestamp 1643678851
transform 1 0 62752 0 1 11054
box 0 0 1 1
use contact_31  contact_31_161
timestamp 1643678851
transform 1 0 62116 0 1 10842
box 0 0 1 1
use contact_31  contact_31_162
timestamp 1643678851
transform 1 0 62116 0 1 9782
box 0 0 1 1
use contact_31  contact_31_163
timestamp 1643678851
transform 1 0 59360 0 1 9782
box 0 0 1 1
use contact_31  contact_31_164
timestamp 1643678851
transform 1 0 59360 0 1 11054
box 0 0 1 1
use contact_31  contact_31_165
timestamp 1643678851
transform 1 0 56604 0 1 9782
box 0 0 1 1
use contact_31  contact_31_166
timestamp 1643678851
transform 1 0 56604 0 1 11054
box 0 0 1 1
use contact_31  contact_31_167
timestamp 1643678851
transform 1 0 55968 0 1 10842
box 0 0 1 1
use contact_31  contact_31_168
timestamp 1643678851
transform 1 0 55968 0 1 9782
box 0 0 1 1
use contact_31  contact_31_169
timestamp 1643678851
transform 1 0 53000 0 1 9782
box 0 0 1 1
use contact_31  contact_31_170
timestamp 1643678851
transform 1 0 53000 0 1 10842
box 0 0 1 1
use contact_31  contact_31_171
timestamp 1643678851
transform 1 0 52788 0 1 10842
box 0 0 1 1
use contact_31  contact_31_172
timestamp 1643678851
transform 1 0 52788 0 1 9782
box 0 0 1 1
use contact_31  contact_31_173
timestamp 1643678851
transform 1 0 50032 0 1 9782
box 0 0 1 1
use contact_31  contact_31_174
timestamp 1643678851
transform 1 0 50032 0 1 11054
box 0 0 1 1
use contact_31  contact_31_175
timestamp 1643678851
transform 1 0 49820 0 1 10842
box 0 0 1 1
use contact_31  contact_31_176
timestamp 1643678851
transform 1 0 49820 0 1 9782
box 0 0 1 1
use contact_31  contact_31_177
timestamp 1643678851
transform 1 0 46428 0 1 9994
box 0 0 1 1
use contact_31  contact_31_178
timestamp 1643678851
transform 1 0 46428 0 1 10842
box 0 0 1 1
use contact_31  contact_31_179
timestamp 1643678851
transform 1 0 46640 0 1 10842
box 0 0 1 1
use contact_31  contact_31_180
timestamp 1643678851
transform 1 0 46640 0 1 9782
box 0 0 1 1
use contact_31  contact_31_181
timestamp 1643678851
transform 1 0 44096 0 1 9782
box 0 0 1 1
use contact_31  contact_31_182
timestamp 1643678851
transform 1 0 44096 0 1 11054
box 0 0 1 1
use contact_31  contact_31_183
timestamp 1643678851
transform 1 0 43460 0 1 10842
box 0 0 1 1
use contact_31  contact_31_184
timestamp 1643678851
transform 1 0 43460 0 1 9782
box 0 0 1 1
use contact_31  contact_31_185
timestamp 1643678851
transform 1 0 40280 0 1 9994
box 0 0 1 1
use contact_31  contact_31_186
timestamp 1643678851
transform 1 0 40280 0 1 10842
box 0 0 1 1
use contact_31  contact_31_187
timestamp 1643678851
transform 1 0 40280 0 1 1938
box 0 0 1 1
use contact_31  contact_31_188
timestamp 1643678851
transform 1 0 40280 0 1 3422
box 0 0 1 1
use contact_31  contact_31_189
timestamp 1643678851
transform 1 0 40492 0 1 10842
box 0 0 1 1
use contact_31  contact_31_190
timestamp 1643678851
transform 1 0 40492 0 1 9782
box 0 0 1 1
use contact_31  contact_31_191
timestamp 1643678851
transform 1 0 37312 0 1 1938
box 0 0 1 1
use contact_31  contact_31_192
timestamp 1643678851
transform 1 0 37312 0 1 3422
box 0 0 1 1
use contact_31  contact_31_193
timestamp 1643678851
transform 1 0 37736 0 1 9782
box 0 0 1 1
use contact_31  contact_31_194
timestamp 1643678851
transform 1 0 37736 0 1 11054
box 0 0 1 1
use contact_31  contact_31_195
timestamp 1643678851
transform 1 0 37312 0 1 10842
box 0 0 1 1
use contact_31  contact_31_196
timestamp 1643678851
transform 1 0 37312 0 1 9782
box 0 0 1 1
use contact_31  contact_31_197
timestamp 1643678851
transform 1 0 34768 0 1 9782
box 0 0 1 1
use contact_31  contact_31_198
timestamp 1643678851
transform 1 0 34768 0 1 11054
box 0 0 1 1
use contact_31  contact_31_199
timestamp 1643678851
transform 1 0 34132 0 1 10842
box 0 0 1 1
use contact_31  contact_31_200
timestamp 1643678851
transform 1 0 34132 0 1 9782
box 0 0 1 1
use contact_31  contact_31_201
timestamp 1643678851
transform 1 0 30952 0 1 9994
box 0 0 1 1
use contact_31  contact_31_202
timestamp 1643678851
transform 1 0 30952 0 1 10842
box 0 0 1 1
use contact_31  contact_31_203
timestamp 1643678851
transform 1 0 30104 0 1 1938
box 0 0 1 1
use contact_31  contact_31_204
timestamp 1643678851
transform 1 0 30104 0 1 3422
box 0 0 1 1
use contact_31  contact_31_205
timestamp 1643678851
transform 1 0 28832 0 1 6390
box 0 0 1 1
use contact_31  contact_31_206
timestamp 1643678851
transform 1 0 28832 0 1 3634
box 0 0 1 1
use contact_31  contact_31_207
timestamp 1643678851
transform 1 0 31164 0 1 10842
box 0 0 1 1
use contact_31  contact_31_208
timestamp 1643678851
transform 1 0 31164 0 1 9782
box 0 0 1 1
use contact_31  contact_31_209
timestamp 1643678851
transform 1 0 28196 0 1 9782
box 0 0 1 1
use contact_31  contact_31_210
timestamp 1643678851
transform 1 0 28196 0 1 11054
box 0 0 1 1
use contact_31  contact_31_211
timestamp 1643678851
transform 1 0 27984 0 1 10842
box 0 0 1 1
use contact_31  contact_31_212
timestamp 1643678851
transform 1 0 27984 0 1 9782
box 0 0 1 1
use contact_31  contact_31_213
timestamp 1643678851
transform 1 0 25016 0 1 9782
box 0 0 1 1
use contact_31  contact_31_214
timestamp 1643678851
transform 1 0 25016 0 1 10842
box 0 0 1 1
use contact_31  contact_31_215
timestamp 1643678851
transform 1 0 24168 0 1 1938
box 0 0 1 1
use contact_31  contact_31_216
timestamp 1643678851
transform 1 0 24168 0 1 3422
box 0 0 1 1
use contact_31  contact_31_217
timestamp 1643678851
transform 1 0 24804 0 1 10842
box 0 0 1 1
use contact_31  contact_31_218
timestamp 1643678851
transform 1 0 24804 0 1 9782
box 0 0 1 1
use contact_31  contact_31_219
timestamp 1643678851
transform 1 0 22048 0 1 9782
box 0 0 1 1
use contact_31  contact_31_220
timestamp 1643678851
transform 1 0 22048 0 1 11054
box 0 0 1 1
use contact_31  contact_31_221
timestamp 1643678851
transform 1 0 21836 0 1 11054
box 0 0 1 1
use contact_31  contact_31_222
timestamp 1643678851
transform 1 0 21836 0 1 13386
box 0 0 1 1
use contact_31  contact_31_223
timestamp 1643678851
transform 1 0 21200 0 1 61934
box 0 0 1 1
use contact_31  contact_31_224
timestamp 1643678851
transform 1 0 21200 0 1 59814
box 0 0 1 1
use contact_31  contact_31_225
timestamp 1643678851
transform 1 0 21200 0 1 19746
box 0 0 1 1
use contact_31  contact_31_226
timestamp 1643678851
transform 1 0 21200 0 1 22714
box 0 0 1 1
use contact_31  contact_31_227
timestamp 1643678851
transform 1 0 21200 0 1 16566
box 0 0 1 1
use contact_31  contact_31_228
timestamp 1643678851
transform 1 0 21200 0 1 19322
box 0 0 1 1
use contact_31  contact_31_229
timestamp 1643678851
transform 1 0 20140 0 1 25894
box 0 0 1 1
use contact_31  contact_31_230
timestamp 1643678851
transform 1 0 20140 0 1 28650
box 0 0 1 1
use contact_31  contact_31_231
timestamp 1643678851
transform 1 0 21200 0 1 47306
box 0 0 1 1
use contact_31  contact_31_232
timestamp 1643678851
transform 1 0 21200 0 1 46882
box 0 0 1 1
use contact_31  contact_31_233
timestamp 1643678851
transform 1 0 21200 0 1 44338
box 0 0 1 1
use contact_31  contact_31_234
timestamp 1643678851
transform 1 0 21200 0 1 46670
box 0 0 1 1
use contact_31  contact_31_235
timestamp 1643678851
transform 1 0 21200 0 1 35010
box 0 0 1 1
use contact_31  contact_31_236
timestamp 1643678851
transform 1 0 21200 0 1 37554
box 0 0 1 1
use contact_31  contact_31_237
timestamp 1643678851
transform 1 0 21200 0 1 53454
box 0 0 1 1
use contact_31  contact_31_238
timestamp 1643678851
transform 1 0 21200 0 1 55786
box 0 0 1 1
use contact_31  contact_31_239
timestamp 1643678851
transform 1 0 21200 0 1 56422
box 0 0 1 1
use contact_31  contact_31_240
timestamp 1643678851
transform 1 0 21200 0 1 55998
box 0 0 1 1
use contact_31  contact_31_241
timestamp 1643678851
transform 1 0 21200 0 1 28862
box 0 0 1 1
use contact_31  contact_31_242
timestamp 1643678851
transform 1 0 21200 0 1 31618
box 0 0 1 1
use contact_31  contact_31_243
timestamp 1643678851
transform 1 0 19928 0 1 13598
box 0 0 1 1
use contact_31  contact_31_244
timestamp 1643678851
transform 1 0 19928 0 1 16354
box 0 0 1 1
use contact_31  contact_31_245
timestamp 1643678851
transform 1 0 21200 0 1 32042
box 0 0 1 1
use contact_31  contact_31_246
timestamp 1643678851
transform 1 0 21200 0 1 34586
box 0 0 1 1
use contact_31  contact_31_247
timestamp 1643678851
transform 1 0 20140 0 1 47306
box 0 0 1 1
use contact_31  contact_31_248
timestamp 1643678851
transform 1 0 20140 0 1 49850
box 0 0 1 1
use contact_31  contact_31_249
timestamp 1643678851
transform 1 0 21200 0 1 50274
box 0 0 1 1
use contact_31  contact_31_250
timestamp 1643678851
transform 1 0 21200 0 1 49850
box 0 0 1 1
use contact_31  contact_31_251
timestamp 1643678851
transform 1 0 20140 0 1 53454
box 0 0 1 1
use contact_31  contact_31_252
timestamp 1643678851
transform 1 0 20140 0 1 52818
box 0 0 1 1
use contact_31  contact_31_253
timestamp 1643678851
transform 1 0 21200 0 1 50486
box 0 0 1 1
use contact_31  contact_31_254
timestamp 1643678851
transform 1 0 21200 0 1 52818
box 0 0 1 1
use contact_31  contact_31_255
timestamp 1643678851
transform 1 0 21200 0 1 41158
box 0 0 1 1
use contact_31  contact_31_256
timestamp 1643678851
transform 1 0 21200 0 1 43702
box 0 0 1 1
use contact_31  contact_31_257
timestamp 1643678851
transform 1 0 20140 0 1 41158
box 0 0 1 1
use contact_31  contact_31_258
timestamp 1643678851
transform 1 0 20140 0 1 40734
box 0 0 1 1
use contact_31  contact_31_259
timestamp 1643678851
transform 1 0 21200 0 1 38190
box 0 0 1 1
use contact_31  contact_31_260
timestamp 1643678851
transform 1 0 21200 0 1 40734
box 0 0 1 1
use contact_31  contact_31_261
timestamp 1643678851
transform 1 0 21200 0 1 56634
box 0 0 1 1
use contact_31  contact_31_262
timestamp 1643678851
transform 1 0 21200 0 1 58754
box 0 0 1 1
use contact_31  contact_31_263
timestamp 1643678851
transform 1 0 21200 0 1 59602
box 0 0 1 1
use contact_31  contact_31_264
timestamp 1643678851
transform 1 0 21200 0 1 58966
box 0 0 1 1
use contact_31  contact_31_265
timestamp 1643678851
transform 1 0 19928 0 1 25470
box 0 0 1 1
use contact_31  contact_31_266
timestamp 1643678851
transform 1 0 19928 0 1 22714
box 0 0 1 1
use contact_31  contact_31_267
timestamp 1643678851
transform 1 0 21836 0 1 10842
box 0 0 1 1
use contact_31  contact_31_268
timestamp 1643678851
transform 1 0 21836 0 1 10206
box 0 0 1 1
use contact_31  contact_31_269
timestamp 1643678851
transform 1 0 18868 0 1 9994
box 0 0 1 1
use contact_31  contact_31_270
timestamp 1643678851
transform 1 0 18868 0 1 8510
box 0 0 1 1
use contact_31  contact_31_271
timestamp 1643678851
transform 1 0 18020 0 1 1938
box 0 0 1 1
use contact_31  contact_31_272
timestamp 1643678851
transform 1 0 18020 0 1 3422
box 0 0 1 1
use contact_31  contact_31_273
timestamp 1643678851
transform 1 0 16112 0 1 25682
box 0 0 1 1
use contact_31  contact_31_274
timestamp 1643678851
transform 1 0 16112 0 1 22714
box 0 0 1 1
use contact_31  contact_31_275
timestamp 1643678851
transform 1 0 15476 0 1 35222
box 0 0 1 1
use contact_31  contact_31_276
timestamp 1643678851
transform 1 0 15476 0 1 37978
box 0 0 1 1
use contact_31  contact_31_277
timestamp 1643678851
transform 1 0 15264 0 1 38190
box 0 0 1 1
use contact_31  contact_31_278
timestamp 1643678851
transform 1 0 15264 0 1 41158
box 0 0 1 1
use contact_31  contact_31_279
timestamp 1643678851
transform 1 0 15264 0 1 35010
box 0 0 1 1
use contact_31  contact_31_280
timestamp 1643678851
transform 1 0 15264 0 1 32042
box 0 0 1 1
use contact_31  contact_31_281
timestamp 1643678851
transform 1 0 15688 0 1 16566
box 0 0 1 1
use contact_31  contact_31_282
timestamp 1643678851
transform 1 0 15688 0 1 17838
box 0 0 1 1
use contact_31  contact_31_283
timestamp 1643678851
transform 1 0 15688 0 1 13386
box 0 0 1 1
use contact_31  contact_31_284
timestamp 1643678851
transform 1 0 15688 0 1 12962
box 0 0 1 1
use contact_31  contact_31_285
timestamp 1643678851
transform 1 0 13568 0 1 12962
box 0 0 1 1
use contact_31  contact_31_286
timestamp 1643678851
transform 1 0 13568 0 1 14658
box 0 0 1 1
use contact_31  contact_31_287
timestamp 1643678851
transform 1 0 13568 0 1 17838
box 0 0 1 1
use contact_31  contact_31_288
timestamp 1643678851
transform 1 0 13568 0 1 16354
box 0 0 1 1
use contact_31  contact_31_289
timestamp 1643678851
transform 1 0 13780 0 1 14658
box 0 0 1 1
use contact_31  contact_31_290
timestamp 1643678851
transform 1 0 13780 0 1 16142
box 0 0 1 1
use contact_31  contact_31_291
timestamp 1643678851
transform 1 0 13568 0 1 18050
box 0 0 1 1
use contact_31  contact_31_292
timestamp 1643678851
transform 1 0 13568 0 1 19534
box 0 0 1 1
use contact_31  contact_31_293
timestamp 1643678851
transform 1 0 1908 0 1 6814
box 0 0 1 1
use contact_33  contact_33_0
timestamp 1643678851
transform 1 0 424 0 1 62994
box 0 0 1 1
use contact_33  contact_33_1
timestamp 1643678851
transform 1 0 120840 0 1 878
box 0 0 1 1
use contact_33  contact_33_2
timestamp 1643678851
transform 1 0 120840 0 1 63418
box 0 0 1 1
use contact_33  contact_33_3
timestamp 1643678851
transform 1 0 121052 0 1 666
box 0 0 1 1
use contact_33  contact_33_4
timestamp 1643678851
transform 1 0 121052 0 1 63206
box 0 0 1 1
use contact_33  contact_33_5
timestamp 1643678851
transform 1 0 120840 0 1 454
box 0 0 1 1
use contact_33  contact_33_6
timestamp 1643678851
transform 1 0 120840 0 1 62994
box 0 0 1 1
use contact_33  contact_33_7
timestamp 1643678851
transform 1 0 636 0 1 666
box 0 0 1 1
use contact_33  contact_33_8
timestamp 1643678851
transform 1 0 424 0 1 666
box 0 0 1 1
use contact_33  contact_33_9
timestamp 1643678851
transform 1 0 848 0 1 666
box 0 0 1 1
use contact_33  contact_33_10
timestamp 1643678851
transform 1 0 120628 0 1 666
box 0 0 1 1
use contact_33  contact_33_11
timestamp 1643678851
transform 1 0 120628 0 1 63206
box 0 0 1 1
use contact_33  contact_33_12
timestamp 1643678851
transform 1 0 848 0 1 63206
box 0 0 1 1
use contact_33  contact_33_13
timestamp 1643678851
transform 1 0 636 0 1 63206
box 0 0 1 1
use contact_33  contact_33_14
timestamp 1643678851
transform 1 0 424 0 1 63206
box 0 0 1 1
use contact_33  contact_33_15
timestamp 1643678851
transform 1 0 120840 0 1 666
box 0 0 1 1
use contact_33  contact_33_16
timestamp 1643678851
transform 1 0 848 0 1 63418
box 0 0 1 1
use contact_33  contact_33_17
timestamp 1643678851
transform 1 0 121052 0 1 878
box 0 0 1 1
use contact_33  contact_33_18
timestamp 1643678851
transform 1 0 121052 0 1 63418
box 0 0 1 1
use contact_33  contact_33_19
timestamp 1643678851
transform 1 0 120628 0 1 63418
box 0 0 1 1
use contact_33  contact_33_20
timestamp 1643678851
transform 1 0 121052 0 1 454
box 0 0 1 1
use contact_33  contact_33_21
timestamp 1643678851
transform 1 0 120840 0 1 63206
box 0 0 1 1
use contact_33  contact_33_22
timestamp 1643678851
transform 1 0 121052 0 1 62994
box 0 0 1 1
use contact_33  contact_33_23
timestamp 1643678851
transform 1 0 636 0 1 63418
box 0 0 1 1
use contact_33  contact_33_24
timestamp 1643678851
transform 1 0 424 0 1 63418
box 0 0 1 1
use contact_33  contact_33_25
timestamp 1643678851
transform 1 0 848 0 1 454
box 0 0 1 1
use contact_33  contact_33_26
timestamp 1643678851
transform 1 0 848 0 1 878
box 0 0 1 1
use contact_33  contact_33_27
timestamp 1643678851
transform 1 0 120628 0 1 878
box 0 0 1 1
use contact_33  contact_33_28
timestamp 1643678851
transform 1 0 848 0 1 62994
box 0 0 1 1
use contact_33  contact_33_29
timestamp 1643678851
transform 1 0 120628 0 1 454
box 0 0 1 1
use contact_33  contact_33_30
timestamp 1643678851
transform 1 0 636 0 1 878
box 0 0 1 1
use contact_33  contact_33_31
timestamp 1643678851
transform 1 0 120628 0 1 62994
box 0 0 1 1
use contact_33  contact_33_32
timestamp 1643678851
transform 1 0 636 0 1 454
box 0 0 1 1
use contact_33  contact_33_33
timestamp 1643678851
transform 1 0 424 0 1 878
box 0 0 1 1
use contact_33  contact_33_34
timestamp 1643678851
transform 1 0 636 0 1 62994
box 0 0 1 1
use contact_33  contact_33_35
timestamp 1643678851
transform 1 0 424 0 1 454
box 0 0 1 1
use contact_33  contact_33_36
timestamp 1643678851
transform 1 0 1908 0 1 1726
box 0 0 1 1
use contact_33  contact_33_37
timestamp 1643678851
transform 1 0 119992 0 1 1514
box 0 0 1 1
use contact_33  contact_33_38
timestamp 1643678851
transform 1 0 1908 0 1 61934
box 0 0 1 1
use contact_33  contact_33_39
timestamp 1643678851
transform 1 0 119568 0 1 1726
box 0 0 1 1
use contact_33  contact_33_40
timestamp 1643678851
transform 1 0 119568 0 1 62358
box 0 0 1 1
use contact_33  contact_33_41
timestamp 1643678851
transform 1 0 119568 0 1 61934
box 0 0 1 1
use contact_33  contact_33_42
timestamp 1643678851
transform 1 0 1696 0 1 62358
box 0 0 1 1
use contact_33  contact_33_43
timestamp 1643678851
transform 1 0 1696 0 1 1726
box 0 0 1 1
use contact_33  contact_33_44
timestamp 1643678851
transform 1 0 1696 0 1 61934
box 0 0 1 1
use contact_33  contact_33_45
timestamp 1643678851
transform 1 0 1484 0 1 1726
box 0 0 1 1
use contact_33  contact_33_46
timestamp 1643678851
transform 1 0 1908 0 1 62358
box 0 0 1 1
use contact_33  contact_33_47
timestamp 1643678851
transform 1 0 1484 0 1 61934
box 0 0 1 1
use contact_33  contact_33_48
timestamp 1643678851
transform 1 0 119780 0 1 62358
box 0 0 1 1
use contact_33  contact_33_49
timestamp 1643678851
transform 1 0 1484 0 1 62358
box 0 0 1 1
use contact_33  contact_33_50
timestamp 1643678851
transform 1 0 119992 0 1 62358
box 0 0 1 1
use contact_33  contact_33_51
timestamp 1643678851
transform 1 0 119992 0 1 1726
box 0 0 1 1
use contact_33  contact_33_52
timestamp 1643678851
transform 1 0 119992 0 1 61934
box 0 0 1 1
use contact_33  contact_33_53
timestamp 1643678851
transform 1 0 119780 0 1 1726
box 0 0 1 1
use contact_33  contact_33_54
timestamp 1643678851
transform 1 0 119780 0 1 61934
box 0 0 1 1
use contact_33  contact_33_55
timestamp 1643678851
transform 1 0 119568 0 1 1938
box 0 0 1 1
use contact_33  contact_33_56
timestamp 1643678851
transform 1 0 119568 0 1 62146
box 0 0 1 1
use contact_33  contact_33_57
timestamp 1643678851
transform 1 0 1696 0 1 1938
box 0 0 1 1
use contact_33  contact_33_58
timestamp 1643678851
transform 1 0 1696 0 1 62146
box 0 0 1 1
use contact_33  contact_33_59
timestamp 1643678851
transform 1 0 1696 0 1 1514
box 0 0 1 1
use contact_33  contact_33_60
timestamp 1643678851
transform 1 0 1908 0 1 1514
box 0 0 1 1
use contact_33  contact_33_61
timestamp 1643678851
transform 1 0 1908 0 1 1938
box 0 0 1 1
use contact_33  contact_33_62
timestamp 1643678851
transform 1 0 119568 0 1 1514
box 0 0 1 1
use contact_33  contact_33_63
timestamp 1643678851
transform 1 0 1908 0 1 62146
box 0 0 1 1
use contact_33  contact_33_64
timestamp 1643678851
transform 1 0 1484 0 1 1938
box 0 0 1 1
use contact_33  contact_33_65
timestamp 1643678851
transform 1 0 1484 0 1 62146
box 0 0 1 1
use contact_33  contact_33_66
timestamp 1643678851
transform 1 0 1484 0 1 1514
box 0 0 1 1
use contact_33  contact_33_67
timestamp 1643678851
transform 1 0 119992 0 1 1938
box 0 0 1 1
use contact_33  contact_33_68
timestamp 1643678851
transform 1 0 119992 0 1 62146
box 0 0 1 1
use contact_33  contact_33_69
timestamp 1643678851
transform 1 0 119780 0 1 62146
box 0 0 1 1
use contact_33  contact_33_70
timestamp 1643678851
transform 1 0 119780 0 1 1514
box 0 0 1 1
use contact_33  contact_33_71
timestamp 1643678851
transform 1 0 119780 0 1 1938
box 0 0 1 1
use contact_31  contact_31_294
timestamp 1643678851
transform 1 0 13144 0 1 12326
box 0 0 1 1
use contact_31  contact_31_295
timestamp 1643678851
transform 1 0 68900 0 1 10630
box 0 0 1 1
use contact_31  contact_31_296
timestamp 1643678851
transform 1 0 65720 0 1 10630
box 0 0 1 1
use contact_31  contact_31_297
timestamp 1643678851
transform 1 0 62540 0 1 10630
box 0 0 1 1
use contact_31  contact_31_298
timestamp 1643678851
transform 1 0 59784 0 1 10630
box 0 0 1 1
use contact_31  contact_31_299
timestamp 1643678851
transform 1 0 56392 0 1 10630
box 0 0 1 1
use contact_31  contact_31_300
timestamp 1643678851
transform 1 0 53212 0 1 10630
box 0 0 1 1
use contact_31  contact_31_301
timestamp 1643678851
transform 1 0 50456 0 1 10630
box 0 0 1 1
use contact_31  contact_31_302
timestamp 1643678851
transform 1 0 47064 0 1 10630
box 0 0 1 1
use contact_31  contact_31_303
timestamp 1643678851
transform 1 0 43884 0 1 10630
box 0 0 1 1
use contact_31  contact_31_304
timestamp 1643678851
transform 1 0 40916 0 1 10630
box 0 0 1 1
use contact_31  contact_31_305
timestamp 1643678851
transform 1 0 37948 0 1 10630
box 0 0 1 1
use contact_31  contact_31_306
timestamp 1643678851
transform 1 0 34556 0 1 10630
box 0 0 1 1
use contact_31  contact_31_307
timestamp 1643678851
transform 1 0 31588 0 1 10630
box 0 0 1 1
use contact_31  contact_31_308
timestamp 1643678851
transform 1 0 28620 0 1 10630
box 0 0 1 1
use contact_31  contact_31_309
timestamp 1643678851
transform 1 0 25440 0 1 10630
box 0 0 1 1
use contact_31  contact_31_310
timestamp 1643678851
transform 1 0 22260 0 1 10630
box 0 0 1 1
use contact_31  contact_31_311
timestamp 1643678851
transform 1 0 6148 0 1 7026
box 0 0 1 1
use contact_31  contact_31_312
timestamp 1643678851
transform 1 0 17596 0 1 2786
box 0 0 1 1
use contact_31  contact_31_313
timestamp 1643678851
transform 1 0 16112 0 1 2786
box 0 0 1 1
use contact_31  contact_31_314
timestamp 1643678851
transform 1 0 41552 0 1 2786
box 0 0 1 1
use contact_31  contact_31_315
timestamp 1643678851
transform 1 0 39856 0 1 2786
box 0 0 1 1
use contact_31  contact_31_316
timestamp 1643678851
transform 1 0 38584 0 1 2786
box 0 0 1 1
use contact_31  contact_31_317
timestamp 1643678851
transform 1 0 36888 0 1 2786
box 0 0 1 1
use contact_31  contact_31_318
timestamp 1643678851
transform 1 0 35616 0 1 2786
box 0 0 1 1
use contact_31  contact_31_319
timestamp 1643678851
transform 1 0 33920 0 1 2786
box 0 0 1 1
use contact_31  contact_31_320
timestamp 1643678851
transform 1 0 32436 0 1 2786
box 0 0 1 1
use contact_31  contact_31_321
timestamp 1643678851
transform 1 0 30952 0 1 2786
box 0 0 1 1
use contact_31  contact_31_322
timestamp 1643678851
transform 1 0 29468 0 1 2786
box 0 0 1 1
use contact_31  contact_31_323
timestamp 1643678851
transform 1 0 28196 0 1 2786
box 0 0 1 1
use contact_31  contact_31_324
timestamp 1643678851
transform 1 0 26712 0 1 2786
box 0 0 1 1
use contact_31  contact_31_325
timestamp 1643678851
transform 1 0 25228 0 1 2786
box 0 0 1 1
use contact_31  contact_31_326
timestamp 1643678851
transform 1 0 23744 0 1 2786
box 0 0 1 1
use contact_31  contact_31_327
timestamp 1643678851
transform 1 0 22048 0 1 2786
box 0 0 1 1
use contact_31  contact_31_328
timestamp 1643678851
transform 1 0 20564 0 1 2786
box 0 0 1 1
use contact_31  contact_31_329
timestamp 1643678851
transform 1 0 19292 0 1 2786
box 0 0 1 1
use contact_18  contact_18_0
timestamp 1643678851
transform 1 0 13227 0 1 17391
box 0 0 1 1
use contact_18  contact_18_1
timestamp 1643678851
transform 1 0 13227 0 1 16899
box 0 0 1 1
use contact_18  contact_18_2
timestamp 1643678851
transform 1 0 13227 0 1 15715
box 0 0 1 1
use contact_18  contact_18_3
timestamp 1643678851
transform 1 0 13227 0 1 15223
box 0 0 1 1
use contact_18  contact_18_4
timestamp 1643678851
transform 1 0 13227 0 1 14039
box 0 0 1 1
use contact_18  contact_18_5
timestamp 1643678851
transform 1 0 13227 0 1 13547
box 0 0 1 1
use contact_18  contact_18_6
timestamp 1643678851
transform 1 0 13227 0 1 12363
box 0 0 1 1
use contact_18  contact_18_7
timestamp 1643678851
transform 1 0 17673 0 1 2915
box 0 0 1 1
use contact_18  contact_18_8
timestamp 1643678851
transform 1 0 16191 0 1 2915
box 0 0 1 1
use contact_18  contact_18_9
timestamp 1643678851
transform 1 0 68940 0 1 10637
box 0 0 1 1
use contact_18  contact_18_10
timestamp 1643678851
transform 1 0 68940 0 1 10637
box 0 0 1 1
use contact_18  contact_18_11
timestamp 1643678851
transform 1 0 65828 0 1 10637
box 0 0 1 1
use contact_18  contact_18_12
timestamp 1643678851
transform 1 0 65828 0 1 10637
box 0 0 1 1
use contact_18  contact_18_13
timestamp 1643678851
transform 1 0 62716 0 1 10637
box 0 0 1 1
use contact_18  contact_18_14
timestamp 1643678851
transform 1 0 62716 0 1 10637
box 0 0 1 1
use contact_18  contact_18_15
timestamp 1643678851
transform 1 0 59604 0 1 10637
box 0 0 1 1
use contact_18  contact_18_16
timestamp 1643678851
transform 1 0 59604 0 1 10637
box 0 0 1 1
use contact_18  contact_18_17
timestamp 1643678851
transform 1 0 56492 0 1 10637
box 0 0 1 1
use contact_18  contact_18_18
timestamp 1643678851
transform 1 0 56492 0 1 10637
box 0 0 1 1
use contact_18  contact_18_19
timestamp 1643678851
transform 1 0 53380 0 1 10637
box 0 0 1 1
use contact_18  contact_18_20
timestamp 1643678851
transform 1 0 53380 0 1 10637
box 0 0 1 1
use contact_18  contact_18_21
timestamp 1643678851
transform 1 0 50268 0 1 10637
box 0 0 1 1
use contact_18  contact_18_22
timestamp 1643678851
transform 1 0 50268 0 1 10637
box 0 0 1 1
use contact_18  contact_18_23
timestamp 1643678851
transform 1 0 47156 0 1 10637
box 0 0 1 1
use contact_18  contact_18_24
timestamp 1643678851
transform 1 0 47156 0 1 10637
box 0 0 1 1
use contact_18  contact_18_25
timestamp 1643678851
transform 1 0 44044 0 1 10637
box 0 0 1 1
use contact_18  contact_18_26
timestamp 1643678851
transform 1 0 44044 0 1 10637
box 0 0 1 1
use contact_18  contact_18_27
timestamp 1643678851
transform 1 0 40932 0 1 10637
box 0 0 1 1
use contact_18  contact_18_28
timestamp 1643678851
transform 1 0 40932 0 1 10637
box 0 0 1 1
use contact_18  contact_18_29
timestamp 1643678851
transform 1 0 37820 0 1 10637
box 0 0 1 1
use contact_18  contact_18_30
timestamp 1643678851
transform 1 0 37820 0 1 10637
box 0 0 1 1
use contact_18  contact_18_31
timestamp 1643678851
transform 1 0 34708 0 1 10637
box 0 0 1 1
use contact_18  contact_18_32
timestamp 1643678851
transform 1 0 34708 0 1 10637
box 0 0 1 1
use contact_18  contact_18_33
timestamp 1643678851
transform 1 0 31596 0 1 10637
box 0 0 1 1
use contact_18  contact_18_34
timestamp 1643678851
transform 1 0 31596 0 1 10637
box 0 0 1 1
use contact_18  contact_18_35
timestamp 1643678851
transform 1 0 28484 0 1 10637
box 0 0 1 1
use contact_18  contact_18_36
timestamp 1643678851
transform 1 0 28484 0 1 10637
box 0 0 1 1
use contact_18  contact_18_37
timestamp 1643678851
transform 1 0 25372 0 1 10637
box 0 0 1 1
use contact_18  contact_18_38
timestamp 1643678851
transform 1 0 25372 0 1 10637
box 0 0 1 1
use contact_18  contact_18_39
timestamp 1643678851
transform 1 0 22260 0 1 10637
box 0 0 1 1
use contact_18  contact_18_40
timestamp 1643678851
transform 1 0 22260 0 1 10637
box 0 0 1 1
use contact_18  contact_18_41
timestamp 1643678851
transform 1 0 41385 0 1 2915
box 0 0 1 1
use contact_18  contact_18_42
timestamp 1643678851
transform 1 0 39903 0 1 2915
box 0 0 1 1
use contact_18  contact_18_43
timestamp 1643678851
transform 1 0 38421 0 1 2915
box 0 0 1 1
use contact_18  contact_18_44
timestamp 1643678851
transform 1 0 36939 0 1 2915
box 0 0 1 1
use contact_18  contact_18_45
timestamp 1643678851
transform 1 0 35457 0 1 2915
box 0 0 1 1
use contact_18  contact_18_46
timestamp 1643678851
transform 1 0 33975 0 1 2915
box 0 0 1 1
use contact_18  contact_18_47
timestamp 1643678851
transform 1 0 32493 0 1 2915
box 0 0 1 1
use contact_18  contact_18_48
timestamp 1643678851
transform 1 0 31011 0 1 2915
box 0 0 1 1
use contact_18  contact_18_49
timestamp 1643678851
transform 1 0 29529 0 1 2915
box 0 0 1 1
use contact_18  contact_18_50
timestamp 1643678851
transform 1 0 28047 0 1 2915
box 0 0 1 1
use contact_18  contact_18_51
timestamp 1643678851
transform 1 0 26565 0 1 2915
box 0 0 1 1
use contact_18  contact_18_52
timestamp 1643678851
transform 1 0 25083 0 1 2915
box 0 0 1 1
use contact_18  contact_18_53
timestamp 1643678851
transform 1 0 23601 0 1 2915
box 0 0 1 1
use contact_18  contact_18_54
timestamp 1643678851
transform 1 0 22119 0 1 2915
box 0 0 1 1
use contact_18  contact_18_55
timestamp 1643678851
transform 1 0 20637 0 1 2915
box 0 0 1 1
use contact_18  contact_18_56
timestamp 1643678851
transform 1 0 19155 0 1 2915
box 0 0 1 1
use contact_18  contact_18_57
timestamp 1643678851
transform 1 0 6185 0 1 7206
box 0 0 1 1
use contact_18  contact_18_58
timestamp 1643678851
transform 1 0 2825 0 1 7421
box 0 0 1 1
use contact_18  contact_18_59
timestamp 1643678851
transform 1 0 2825 0 1 6237
box 0 0 1 1
use contact_18  contact_18_60
timestamp 1643678851
transform 1 0 15061 0 1 17387
box 0 0 1 1
use contact_18  contact_18_61
timestamp 1643678851
transform 1 0 14307 0 1 17387
box 0 0 1 1
use contact_18  contact_18_62
timestamp 1643678851
transform 1 0 14993 0 1 16903
box 0 0 1 1
use contact_18  contact_18_63
timestamp 1643678851
transform 1 0 14307 0 1 16903
box 0 0 1 1
use contact_18  contact_18_64
timestamp 1643678851
transform 1 0 14925 0 1 15711
box 0 0 1 1
use contact_18  contact_18_65
timestamp 1643678851
transform 1 0 14307 0 1 15711
box 0 0 1 1
use contact_18  contact_18_66
timestamp 1643678851
transform 1 0 14857 0 1 15227
box 0 0 1 1
use contact_18  contact_18_67
timestamp 1643678851
transform 1 0 14307 0 1 15227
box 0 0 1 1
use contact_18  contact_18_68
timestamp 1643678851
transform 1 0 14789 0 1 14035
box 0 0 1 1
use contact_18  contact_18_69
timestamp 1643678851
transform 1 0 14307 0 1 14035
box 0 0 1 1
use contact_18  contact_18_70
timestamp 1643678851
transform 1 0 14721 0 1 13551
box 0 0 1 1
use contact_18  contact_18_71
timestamp 1643678851
transform 1 0 14307 0 1 13551
box 0 0 1 1
use contact_18  contact_18_72
timestamp 1643678851
transform 1 0 14653 0 1 12359
box 0 0 1 1
use contact_18  contact_18_73
timestamp 1643678851
transform 1 0 14307 0 1 12359
box 0 0 1 1
use contact_18  contact_18_74
timestamp 1643678851
transform 1 0 20016 0 1 11484
box 0 0 1 1
use contact_18  contact_18_75
timestamp 1643678851
transform 1 0 14502 0 1 11484
box 0 0 1 1
use contact_18  contact_18_76
timestamp 1643678851
transform 1 0 71612 0 1 10551
box 0 0 1 1
use contact_18  contact_18_77
timestamp 1643678851
transform 1 0 14502 0 1 10551
box 0 0 1 1
use contact_18  contact_18_78
timestamp 1643678851
transform 1 0 21138 0 1 9810
box 0 0 1 1
use contact_18  contact_18_79
timestamp 1643678851
transform 1 0 14502 0 1 9810
box 0 0 1 1
use contact_29  contact_29_0
timestamp 1643678851
transform 1 0 12952 0 1 2977
box 0 0 1 1
use contact_29  contact_29_1
timestamp 1643678851
transform 1 0 12952 0 1 2977
box 0 0 1 1
use contact_29  contact_29_2
timestamp 1643678851
transform 1 0 12952 0 1 12425
box 0 0 1 1
use data_dff  data_dff_0
timestamp 1643678851
transform 1 0 19014 0 1 2702
box -39 -42 23712 916
use col_addr_dff  col_addr_dff_0
timestamp 1643678851
transform 1 0 16050 0 1 2702
box -39 -42 2964 916
use row_addr_dff  row_addr_dff_0
timestamp 1643678851
transform 1 0 13086 0 1 12150
box -39 -42 1482 7620
use control_logic_multiport  control_logic_multiport_0
timestamp 1643678851
transform 1 0 2684 0 1 6024
box -66 -42 11884 5922
use bank  bank_0
timestamp 1643678851
transform 1 0 14704 0 1 6224
box -11 0 104150 55154
<< labels >>
rlabel metal3 s 2824 6236 2956 6302 4 web
rlabel metal3 s 2824 7420 2956 7486 4 csb
rlabel metal4 s 6148 0 6300 364 4 clk
rlabel metal4 s 19292 0 19444 364 4 din0[0]
rlabel metal4 s 20564 0 20716 364 4 din0[1]
rlabel metal4 s 22048 0 22200 364 4 din0[2]
rlabel metal4 s 23744 0 23896 364 4 din0[3]
rlabel metal4 s 25228 0 25380 364 4 din0[4]
rlabel metal4 s 26712 0 26864 364 4 din0[5]
rlabel metal4 s 28196 0 28348 364 4 din0[6]
rlabel metal4 s 29468 0 29620 364 4 din0[7]
rlabel metal4 s 30952 0 31104 364 4 din0[8]
rlabel metal4 s 32436 0 32588 364 4 din0[9]
rlabel metal4 s 33920 0 34072 364 4 din0[10]
rlabel metal4 s 35616 0 35768 364 4 din0[11]
rlabel metal4 s 36888 0 37040 364 4 din0[12]
rlabel metal4 s 38584 0 38736 364 4 din0[13]
rlabel metal4 s 39856 0 40008 364 4 din0[14]
rlabel metal4 s 41552 0 41704 364 4 din0[15]
rlabel metal4 s 22260 0 22412 364 4 dout0[0]
rlabel metal3 s 22260 10636 22392 10702 4 dout1[0]
rlabel metal4 s 25440 0 25592 364 4 dout0[1]
rlabel metal3 s 25372 10636 25504 10702 4 dout1[1]
rlabel metal4 s 28620 0 28772 364 4 dout0[2]
rlabel metal3 s 28484 10636 28616 10702 4 dout1[2]
rlabel metal4 s 31588 0 31740 364 4 dout0[3]
rlabel metal3 s 31596 10636 31728 10702 4 dout1[3]
rlabel metal4 s 34556 0 34708 364 4 dout0[4]
rlabel metal3 s 34708 10636 34840 10702 4 dout1[4]
rlabel metal4 s 37948 0 38100 364 4 dout0[5]
rlabel metal3 s 37820 10636 37952 10702 4 dout1[5]
rlabel metal4 s 40916 0 41068 364 4 dout0[6]
rlabel metal3 s 40932 10636 41064 10702 4 dout1[6]
rlabel metal4 s 43884 0 44036 364 4 dout0[7]
rlabel metal3 s 44044 10636 44176 10702 4 dout1[7]
rlabel metal4 s 47064 0 47216 364 4 dout0[8]
rlabel metal3 s 47156 10636 47288 10702 4 dout1[8]
rlabel metal4 s 50456 0 50608 364 4 dout0[9]
rlabel metal3 s 50268 10636 50400 10702 4 dout1[9]
rlabel metal4 s 53212 0 53364 364 4 dout0[10]
rlabel metal3 s 53380 10636 53512 10702 4 dout1[10]
rlabel metal4 s 56392 0 56544 364 4 dout0[11]
rlabel metal3 s 56492 10636 56624 10702 4 dout1[11]
rlabel metal4 s 59784 0 59936 364 4 dout0[12]
rlabel metal3 s 59604 10636 59736 10702 4 dout1[12]
rlabel metal4 s 62540 0 62692 364 4 dout0[13]
rlabel metal3 s 62716 10636 62848 10702 4 dout1[13]
rlabel metal4 s 65720 0 65872 364 4 dout0[14]
rlabel metal3 s 65828 10636 65960 10702 4 dout1[14]
rlabel metal4 s 68900 0 69052 364 4 dout0[15]
rlabel metal3 s 68940 10636 69072 10702 4 dout1[15]
rlabel metal4 s 16112 0 16264 364 4 addr0
rlabel metal4 s 17596 0 17748 364 4 addr1
rlabel metal4 s 13144 0 13296 364 4 addr1[2]
rlabel metal3 s 0 13568 364 13720 4 addr1[3]
rlabel metal3 s 0 13992 364 14144 4 addr1[4]
rlabel metal3 s 0 15264 364 15416 4 addr1[5]
rlabel metal3 s 0 15688 364 15840 4 addr1[6]
rlabel metal3 s 0 16748 364 16900 4 addr1[7]
rlabel metal3 s 0 17384 364 17536 4 addr1[8]
rlabel metal3 s 1484 1484 120144 2060 4 vdd
rlabel metal3 s 1484 61904 120144 62480 4 vdd
rlabel metal4 s 1484 1484 2060 62480 4 vdd
rlabel metal4 s 119568 1484 120144 62480 4 vdd
rlabel metal4 s 120628 424 121204 63540 4 gnd
rlabel metal4 s 424 424 1000 63540 4 gnd
rlabel metal3 s 424 62964 121204 63540 4 gnd
rlabel metal3 s 424 424 121204 1000 4 gnd
<< properties >>
string FIXED_BBOX 0 0 121204 63540
string GDS_FILE sram_0rw2r1w_16_128_sky130A.gds
string GDS_END 232702
string GDS_START 128
<< end >>
