* NGSPICE file created from sram_0rw2r1w_32_128_sky130A.ext - technology: sky130A

.subckt dff clk vdd gnd D Q
X0 net3 net2 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.35e+06u l=150000u
X1 gnd net7 a_922_96# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 vdd clk clkb vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.35e+06u l=150000u
X3 net3 net2 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 vdd net3 net4 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.35e+06u l=150000u
X5 gnd net3 a_474_96# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 gnd clk clkb gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_922_96# clkb net6 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_474_96# clk net2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 net4 clkb net2 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.35e+06u l=150000u
X10 net6 clk net3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 net2 clkb net1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 net7 net6 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.35e+06u l=150000u
X13 net8 clk net6 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.35e+06u l=150000u
X14 net2 clk net1 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.35e+06u l=150000u
X15 net1 D gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 vdd net7 net8 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.35e+06u l=150000u
X17 net1 D vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.35e+06u l=150000u
X18 net6 clkb net3 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.35e+06u l=150000u
X19 Q net7 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.35e+06u l=150000u
X20 net7 net6 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 Q net7 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt nmos_m2_w0_420_sli_dli_da_p S S_uq0 gnd D G
X0 D G S gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 S_uq0 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt pmos_m2_w1_260_sli_dli_da_p w_n59_42# S S_uq0 gnd D G
X0 S_uq0 G D w_n59_42# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.26e+06u l=150000u
X1 D G S w_n59_42# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.26e+06u l=150000u
.ends

.subckt pinv_1 Z gnd vdd A
Xnmos_m2_w0_420_sli_dli_da_p_0 gnd gnd gnd Z A nmos_m2_w0_420_sli_dli_da_p
Xpmos_m2_w1_260_sli_dli_da_p_0 vdd vdd vdd gnd Z A pmos_m2_w1_260_sli_dli_da_p
.ends

.subckt nmos_m4_w0_420_sli_dli_da_p S S_uq0 S_uq1 gnd D G
X0 D G S_uq1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 D G S gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 S G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 S_uq0 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt pmos_m4_w1_260_sli_dli_da_p w_n59_42# S S_uq0 S_uq1 gnd D G
X0 D G S w_n59_42# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.26e+06u l=150000u
X1 S G D w_n59_42# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.26e+06u l=150000u
X2 S_uq0 G D w_n59_42# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.26e+06u l=150000u
X3 D G S_uq1 w_n59_42# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.26e+06u l=150000u
.ends

.subckt pinv_2 Z gnd vdd A
Xnmos_m4_w0_420_sli_dli_da_p_0 gnd gnd gnd gnd Z A nmos_m4_w0_420_sli_dli_da_p
Xpmos_m4_w1_260_sli_dli_da_p_0 vdd vdd vdd vdd gnd Z A pmos_m4_w1_260_sli_dli_da_p
.ends

.subckt dff_buf_0 pinv_2_0/vdd clk Q Qb gnd vdd D
Xdff_0 clk vdd gnd D dff_0/Q dff
Xpinv_1_0 Qb gnd pinv_2_0/vdd dff_0/Q pinv_1
Xpinv_2_0 Q gnd pinv_2_0/vdd Qb pinv_2
.ends

.subckt dff_buf_array vdd dout_0 dout_1 dout_bar_0 dout_bar_1 din_0 din_1
Xdff_buf_0_1 dff_buf_0_1/pinv_2_0/vdd vdd dout_0 dout_bar_0 vdd vdd din_0 dff_buf_0
Xdff_buf_0_0 dff_buf_0_1/pinv_2_0/vdd vdd dout_1 dout_bar_1 vdd vdd din_1 dff_buf_0
.ends

.subckt pmos_m1_w1_260_sli_dli w_n59_42# S gnd D G
X0 D G S w_n59_42# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.26e+06u l=150000u
.ends

.subckt nmos_m1_w0_840_sli_dactive S gnd G a_90_0#
X0 a_90_0# G S gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
.ends

.subckt nmos_m1_w0_840_sactive_dli a_0_0# gnd D G
X0 D G a_0_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
.ends

.subckt pnand2_0 w_n36_402# Z gnd A vdd B
Xpmos_m1_w1_260_sli_dli_0 w_n36_402# Z gnd vdd B pmos_m1_w1_260_sli_dli
Xpmos_m1_w1_260_sli_dli_1 w_n36_402# vdd gnd Z A pmos_m1_w1_260_sli_dli
Xnmos_m1_w0_840_sli_dactive_0 gnd gnd A nmos_m1_w0_840_sactive_dli_0/a_0_0# nmos_m1_w0_840_sli_dactive
Xnmos_m1_w0_840_sactive_dli_0 nmos_m1_w0_840_sactive_dli_0/a_0_0# gnd Z B nmos_m1_w0_840_sactive_dli
.ends

.subckt nmos_m34_w0_495_sli_dli_da_p S S_uq0 S_uq1 S_uq3 S_uq2 S_uq4 S_uq10 S_uq5
+ S_uq11 S_uq6 S_uq13 S_uq12 S_uq7 S_uq14 S_uq8 S_uq15 S_uq9 S_uq16 gnd D G
X0 S_uq13 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X1 S_uq1 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X2 D G S_uq16 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X3 S_uq10 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X4 S_uq5 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X5 S G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X6 S_uq8 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X7 S_uq3 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X8 D G S_uq15 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X9 D G S_uq12 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X10 D G S_uq2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X11 S_uq15 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X12 D G S_uq11 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X13 D G S_uq9 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X14 D G S_uq6 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X15 D G S_uq4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X16 D G S_uq1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X17 S_uq12 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X18 S_uq7 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X19 S_uq4 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X20 S_uq2 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X21 S_uq0 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X22 S_uq11 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X23 S_uq9 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X24 S_uq6 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X25 D G S_uq14 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X26 D G S_uq13 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X27 D G S_uq10 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X28 D G S_uq8 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X29 D G S_uq7 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X30 D G S_uq5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X31 D G S_uq3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X32 D G S gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X33 S_uq14 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
.ends

.subckt pmos_m34_w1_480_sli_dli_da_p w_n59_64# S S_uq0 S_uq1 S_uq3 S_uq2 S_uq4 S_uq10
+ S_uq5 S_uq11 S_uq6 S_uq13 S_uq12 S_uq7 S_uq14 S_uq8 S_uq15 S_uq9 S_uq16 gnd D G
X0 D G S_uq15 w_n59_64# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.48e+06u l=150000u
X1 S_uq8 G D w_n59_64# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.48e+06u l=150000u
X2 S_uq3 G D w_n59_64# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.48e+06u l=150000u
X3 D G S_uq12 w_n59_64# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.48e+06u l=150000u
X4 D G S_uq2 w_n59_64# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.48e+06u l=150000u
X5 S_uq15 G D w_n59_64# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.48e+06u l=150000u
X6 D G S_uq11 w_n59_64# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.48e+06u l=150000u
X7 D G S_uq9 w_n59_64# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.48e+06u l=150000u
X8 D G S_uq6 w_n59_64# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.48e+06u l=150000u
X9 D G S_uq4 w_n59_64# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.48e+06u l=150000u
X10 D G S_uq1 w_n59_64# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.48e+06u l=150000u
X11 S_uq12 G D w_n59_64# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.48e+06u l=150000u
X12 S_uq9 G D w_n59_64# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.48e+06u l=150000u
X13 S_uq7 G D w_n59_64# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.48e+06u l=150000u
X14 S_uq4 G D w_n59_64# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.48e+06u l=150000u
X15 S_uq2 G D w_n59_64# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.48e+06u l=150000u
X16 S_uq0 G D w_n59_64# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.48e+06u l=150000u
X17 S_uq11 G D w_n59_64# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.48e+06u l=150000u
X18 S_uq6 G D w_n59_64# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.48e+06u l=150000u
X19 D G S_uq14 w_n59_64# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.48e+06u l=150000u
X20 D G S_uq13 w_n59_64# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.48e+06u l=150000u
X21 D G S_uq10 w_n59_64# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.48e+06u l=150000u
X22 D G S_uq8 w_n59_64# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.48e+06u l=150000u
X23 D G S_uq7 w_n59_64# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.48e+06u l=150000u
X24 D G S_uq5 w_n59_64# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.48e+06u l=150000u
X25 D G S_uq3 w_n59_64# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.48e+06u l=150000u
X26 D G S w_n59_64# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.48e+06u l=150000u
X27 S_uq14 G D w_n59_64# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.48e+06u l=150000u
X28 S_uq13 G D w_n59_64# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.48e+06u l=150000u
X29 S_uq1 G D w_n59_64# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.48e+06u l=150000u
X30 S G D w_n59_64# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.48e+06u l=150000u
X31 D G S_uq16 w_n59_64# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.48e+06u l=150000u
X32 S_uq10 G D w_n59_64# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.48e+06u l=150000u
X33 S_uq5 G D w_n59_64# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.48e+06u l=150000u
.ends

.subckt pinv_14 gnd vdd Z A
Xnmos_m34_w0_495_sli_dli_da_p_0 gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd
+ gnd gnd gnd gnd gnd gnd Z A nmos_m34_w0_495_sli_dli_da_p
Xpmos_m34_w1_480_sli_dli_da_p_0 vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd
+ vdd vdd vdd vdd vdd vdd gnd Z A pmos_m34_w1_480_sli_dli_da_p
.ends

.subckt pdriver_2 vdd Z gnd A
Xpinv_14_0 gnd vdd Z A pinv_14
.ends

.subckt pand2_0 vdd Z gnd A B
Xpnand2_0_0 vdd pnand2_0_0/Z gnd A vdd B pnand2_0
Xpdriver_2_0 vdd Z gnd pnand2_0_0/Z pdriver_2
.ends

.subckt nmos_m18_w0_490_sli_dli_da_p S S_uq0 S_uq1 S_uq3 S_uq2 S_uq4 S_uq5 S_uq6 S_uq7
+ S_uq8 gnd D G
X0 S_uq5 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=490000u l=150000u
X1 D G S_uq8 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=490000u l=150000u
X2 S_uq2 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=490000u l=150000u
X3 S G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=490000u l=150000u
X4 D G S_uq7 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=490000u l=150000u
X5 D G S_uq4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=490000u l=150000u
X6 S_uq7 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=490000u l=150000u
X7 D G S_uq3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=490000u l=150000u
X8 D G S_uq1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=490000u l=150000u
X9 S_uq4 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=490000u l=150000u
X10 S_uq0 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=490000u l=150000u
X11 S_uq3 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=490000u l=150000u
X12 S_uq1 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=490000u l=150000u
X13 D G S_uq6 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=490000u l=150000u
X14 D G S_uq5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=490000u l=150000u
X15 D G S_uq2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=490000u l=150000u
X16 D G S gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=490000u l=150000u
X17 S_uq6 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=490000u l=150000u
.ends

.subckt pmos_m18_w1_470_sli_dli_da_p w_n59_63# S S_uq0 S_uq1 S_uq3 S_uq2 S_uq4 S_uq5
+ S_uq6 S_uq7 S_uq8 gnd D G
X0 D G S_uq7 w_n59_63# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.47e+06u l=150000u
X1 S G D w_n59_63# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.47e+06u l=150000u
X2 D G S_uq4 w_n59_63# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.47e+06u l=150000u
X3 S_uq7 G D w_n59_63# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.47e+06u l=150000u
X4 D G S_uq3 w_n59_63# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.47e+06u l=150000u
X5 D G S_uq1 w_n59_63# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.47e+06u l=150000u
X6 S_uq4 G D w_n59_63# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.47e+06u l=150000u
X7 S_uq1 G D w_n59_63# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.47e+06u l=150000u
X8 S_uq0 G D w_n59_63# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.47e+06u l=150000u
X9 S_uq3 G D w_n59_63# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.47e+06u l=150000u
X10 D G S_uq6 w_n59_63# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.47e+06u l=150000u
X11 D G S_uq5 w_n59_63# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.47e+06u l=150000u
X12 D G S_uq2 w_n59_63# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.47e+06u l=150000u
X13 D G S w_n59_63# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.47e+06u l=150000u
X14 S_uq6 G D w_n59_63# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.47e+06u l=150000u
X15 S_uq5 G D w_n59_63# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.47e+06u l=150000u
X16 D G S_uq8 w_n59_63# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.47e+06u l=150000u
X17 S_uq2 G D w_n59_63# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.47e+06u l=150000u
.ends

.subckt pinv_13 vdd Z gnd A
Xnmos_m18_w0_490_sli_dli_da_p_0 gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd Z A nmos_m18_w0_490_sli_dli_da_p
Xpmos_m18_w1_470_sli_dli_da_p_0 vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd gnd Z
+ A pmos_m18_w1_470_sli_dli_da_p
.ends

.subckt pinv_11 Z gnd vdd A
Xnmos_m2_w0_420_sli_dli_da_p_0 gnd gnd gnd Z A nmos_m2_w0_420_sli_dli_da_p
Xpmos_m2_w1_260_sli_dli_da_p_0 vdd vdd vdd gnd Z A pmos_m2_w1_260_sli_dli_da_p
.ends

.subckt nmos_m1_w0_420_sli_dli_da_p S gnd D G
X0 D G S gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt pmos_m1_w1_260_sli_dli_da_p w_n59_42# S gnd D G
X0 D G S w_n59_42# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.26e+06u l=150000u
.ends

.subckt pinv_6 A Z gnd vdd
Xnmos_m1_w0_420_sli_dli_da_p_0 gnd gnd Z A nmos_m1_w0_420_sli_dli_da_p
Xpmos_m1_w1_260_sli_dli_da_p_0 vdd vdd gnd Z A pmos_m1_w1_260_sli_dli_da_p
.ends

.subckt pmos_m6_w1_470_sli_dli_da_p w_n59_63# S S_uq0 S_uq1 S_uq2 gnd D G
X0 D G S_uq1 w_n59_63# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.47e+06u l=150000u
X1 S_uq1 G D w_n59_63# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.47e+06u l=150000u
X2 D G S w_n59_63# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.47e+06u l=150000u
X3 S G D w_n59_63# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.47e+06u l=150000u
X4 S_uq0 G D w_n59_63# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.47e+06u l=150000u
X5 D G S_uq2 w_n59_63# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.47e+06u l=150000u
.ends

.subckt nmos_m6_w0_490_sli_dli_da_p S S_uq0 S_uq1 S_uq2 gnd D G
X0 S_uq0 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=490000u l=150000u
X1 D G S_uq2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=490000u l=150000u
X2 D G S_uq1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=490000u l=150000u
X3 S_uq1 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=490000u l=150000u
X4 D G S gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=490000u l=150000u
X5 S G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=490000u l=150000u
.ends

.subckt pinv_12 Z gnd vdd A
Xpmos_m6_w1_470_sli_dli_da_p_0 vdd vdd vdd vdd vdd gnd Z A pmos_m6_w1_470_sli_dli_da_p
Xnmos_m6_w0_490_sli_dli_da_p_0 gnd gnd gnd gnd gnd Z A nmos_m6_w0_490_sli_dli_da_p
.ends

.subckt pdriver_1 gnd A vdd Z
Xpinv_13_0 vdd Z gnd pinv_13_0/A pinv_13
Xpinv_11_0 pinv_12_0/A gnd vdd pinv_6_0/Z pinv_11
Xpinv_6_0 A pinv_6_0/Z gnd vdd pinv_6
Xpinv_12_0 pinv_13_0/A gnd vdd pinv_12_0/A pinv_12
.ends

.subckt pmos_m11_w1_375_sli_dli_da_p S S_uq0 S_uq1 S_uq3 S_uq2 S_uq4 gnd w_n59_53#
+ D G
X0 D G S_uq3 w_n59_53# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=150000u
X1 D G S w_n59_53# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=150000u
X2 S_uq3 G D w_n59_53# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=150000u
X3 D G S_uq0 w_n59_53# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=150000u
X4 S G D w_n59_53# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=150000u
X5 S_uq0 G D w_n59_53# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=150000u
X6 D G S_uq2 w_n59_53# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=150000u
X7 D G S_uq1 w_n59_53# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=150000u
X8 S_uq2 G D w_n59_53# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=150000u
X9 S_uq1 G D w_n59_53# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=150000u
X10 D G S_uq4 w_n59_53# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=150000u
.ends

.subckt nmos_m11_w0_460_sli_dli_da_p S S_uq0 S_uq1 S_uq3 S_uq2 S_uq4 gnd D G
X0 S_uq1 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=460000u l=150000u
X1 D G S_uq4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=460000u l=150000u
X2 D G S_uq3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=460000u l=150000u
X3 D G S gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=460000u l=150000u
X4 S_uq3 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=460000u l=150000u
X5 D G S_uq0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=460000u l=150000u
X6 S G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=460000u l=150000u
X7 S_uq0 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=460000u l=150000u
X8 D G S_uq2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=460000u l=150000u
X9 D G S_uq1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=460000u l=150000u
X10 S_uq2 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=460000u l=150000u
.ends

.subckt pinv_3 gnd vdd Z A
Xpmos_m11_w1_375_sli_dli_da_p_0 vdd vdd vdd vdd vdd vdd gnd vdd Z A pmos_m11_w1_375_sli_dli_da_p
Xnmos_m11_w0_460_sli_dli_da_p_0 gnd gnd gnd gnd gnd gnd gnd Z A nmos_m11_w0_460_sli_dli_da_p
.ends

.subckt pdriver gnd vdd Z A
Xpinv_3_0 gnd vdd Z A pinv_3
.ends

.subckt pand2 vdd gnd Z A B
Xpnand2_0_0 vdd pdriver_0/A gnd A vdd B pnand2_0
Xpdriver_0 gnd vdd Z pdriver_0/A pdriver
.ends

.subckt pnand2_1 Z gnd vdd A
Xpmos_m1_w1_260_sli_dli_0 vdd Z gnd vdd B pmos_m1_w1_260_sli_dli
Xpmos_m1_w1_260_sli_dli_1 vdd vdd gnd Z A pmos_m1_w1_260_sli_dli
Xnmos_m1_w0_840_sli_dactive_0 gnd gnd A nmos_m1_w0_840_sactive_dli_0/a_0_0# nmos_m1_w0_840_sli_dactive
Xnmos_m1_w0_840_sactive_dli_0 nmos_m1_w0_840_sactive_dli_0/a_0_0# gnd Z B nmos_m1_w0_840_sactive_dli
.ends

.subckt pmos_m21_w1_440_sli_dli_da_p w_n59_60# S S_uq0 S_uq1 S_uq3 S_uq2 S_uq4 S_uq5
+ S_uq6 S_uq7 S_uq8 S_uq9 gnd D G
X0 D G S_uq8 w_n59_60# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.44e+06u l=150000u
X1 S_uq1 G D w_n59_60# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.44e+06u l=150000u
X2 D G S_uq5 w_n59_60# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.44e+06u l=150000u
X3 S_uq8 G D w_n59_60# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.44e+06u l=150000u
X4 D G S_uq4 w_n59_60# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.44e+06u l=150000u
X5 D G S_uq2 w_n59_60# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.44e+06u l=150000u
X6 D G S_uq0 w_n59_60# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.44e+06u l=150000u
X7 S_uq5 G D w_n59_60# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.44e+06u l=150000u
X8 S_uq2 G D w_n59_60# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.44e+06u l=150000u
X9 S G D w_n59_60# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.44e+06u l=150000u
X10 S_uq4 G D w_n59_60# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.44e+06u l=150000u
X11 S_uq0 G D w_n59_60# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.44e+06u l=150000u
X12 D G S_uq7 w_n59_60# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.44e+06u l=150000u
X13 D G S_uq6 w_n59_60# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.44e+06u l=150000u
X14 D G S_uq3 w_n59_60# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.44e+06u l=150000u
X15 D G S_uq1 w_n59_60# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.44e+06u l=150000u
X16 D G S w_n59_60# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.44e+06u l=150000u
X17 S_uq7 G D w_n59_60# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.44e+06u l=150000u
X18 S_uq6 G D w_n59_60# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.44e+06u l=150000u
X19 D G S_uq9 w_n59_60# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.44e+06u l=150000u
X20 S_uq3 G D w_n59_60# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.44e+06u l=150000u
.ends

.subckt nmos_m21_w0_480_sli_dli_da_p S S_uq0 S_uq1 S_uq3 S_uq2 S_uq4 S_uq5 S_uq6 S_uq7
+ S_uq8 S_uq9 gnd D G
X0 S_uq6 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=480000u l=150000u
X1 D G S_uq9 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=480000u l=150000u
X2 S_uq3 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=480000u l=150000u
X3 S_uq1 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=480000u l=150000u
X4 D G S_uq8 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=480000u l=150000u
X5 D G S_uq5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=480000u l=150000u
X6 S_uq8 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=480000u l=150000u
X7 D G S_uq4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=480000u l=150000u
X8 D G S_uq2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=480000u l=150000u
X9 D G S_uq0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=480000u l=150000u
X10 S_uq5 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=480000u l=150000u
X11 S G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=480000u l=150000u
X12 S_uq4 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=480000u l=150000u
X13 S_uq2 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=480000u l=150000u
X14 S_uq0 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=480000u l=150000u
X15 D G S_uq7 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=480000u l=150000u
X16 D G S_uq6 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=480000u l=150000u
X17 D G S_uq3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=480000u l=150000u
X18 D G S_uq1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=480000u l=150000u
X19 D G S gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=480000u l=150000u
X20 S_uq7 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=480000u l=150000u
.ends

.subckt pinv_9 gnd Z vdd A
Xpmos_m21_w1_440_sli_dli_da_p_0 vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd gnd
+ Z A pmos_m21_w1_440_sli_dli_da_p
Xnmos_m21_w0_480_sli_dli_da_p_0 gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd Z
+ A nmos_m21_w0_480_sli_dli_da_p
.ends

.subckt nmos_m3_w0_420_sli_dli_da_p S S_uq0 gnd D G
X0 D G S gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 D G S_uq0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 S_uq0 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt pmos_m3_w1_260_sli_dli_da_p w_n59_42# S S_uq0 gnd D G
X0 D G S_uq0 w_n59_42# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.26e+06u l=150000u
X1 S_uq0 G D w_n59_42# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.26e+06u l=150000u
X2 D G S w_n59_42# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.26e+06u l=150000u
.ends

.subckt pinv_7 Z gnd vdd A
Xnmos_m3_w0_420_sli_dli_da_p_0 gnd gnd gnd Z A nmos_m3_w0_420_sli_dli_da_p
Xpmos_m3_w1_260_sli_dli_da_p_0 vdd vdd vdd gnd Z A pmos_m3_w1_260_sli_dli_da_p
.ends

.subckt pmos_m7_w1_440_sli_dli_da_p w_n59_60# S S_uq0 S_uq1 S_uq2 gnd D G
X0 D G S_uq1 w_n59_60# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.44e+06u l=150000u
X1 S_uq1 G D w_n59_60# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.44e+06u l=150000u
X2 D G S w_n59_60# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.44e+06u l=150000u
X3 D G S_uq0 w_n59_60# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.44e+06u l=150000u
X4 S G D w_n59_60# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.44e+06u l=150000u
X5 S_uq0 G D w_n59_60# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.44e+06u l=150000u
X6 D G S_uq2 w_n59_60# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.44e+06u l=150000u
.ends

.subckt nmos_m7_w0_480_sli_dli_da_p S S_uq0 S_uq1 S_uq2 gnd D G
X0 S_uq0 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=480000u l=150000u
X1 D G S_uq2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=480000u l=150000u
X2 D G S_uq1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=480000u l=150000u
X3 S_uq1 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=480000u l=150000u
X4 D G S gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=480000u l=150000u
X5 D G S_uq0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=480000u l=150000u
X6 S G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=480000u l=150000u
.ends

.subckt pinv_8 vdd Z gnd A
Xpmos_m7_w1_440_sli_dli_da_p_0 vdd vdd vdd vdd vdd gnd Z A pmos_m7_w1_440_sli_dli_da_p
Xnmos_m7_w0_480_sli_dli_da_p_0 gnd gnd gnd gnd gnd Z A nmos_m7_w0_480_sli_dli_da_p
.ends

.subckt nmos_m61_w0_495_sli_dli_da_p S S_uq0 S_uq1 S_uq3 S_uq2 S_uq20 S_uq4 S_uq21
+ S_uq10 S_uq5 S_uq22 S_uq11 S_uq6 S_uq24 S_uq23 S_uq13 S_uq12 S_uq7 S_uq25 S_uq14
+ S_uq8 S_uq26 S_uq15 S_uq9 S_uq27 S_uq16 S_uq28 S_uq17 gnd S_uq29 S_uq18 S_uq19 D
+ G
X0 S_uq26 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X1 S_uq14 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X2 S_uq9 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X3 S_uq4 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X4 S_uq2 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X5 S_uq1 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X6 S_uq0 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X7 D G S_uq29 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X8 S_uq23 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X9 S_uq18 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X10 S_uq13 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X11 S_uq21 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X12 S_uq16 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X13 S_uq11 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X14 S_uq6 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X15 D G S_uq28 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X16 D G S_uq25 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X17 D G S_uq3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X18 D G S_uq15 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X19 D G S_uq10 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X20 D G S_uq8 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X21 D G S_uq5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X22 D G S gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X23 D G S_uq7 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X24 S_uq28 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X25 D G S_uq24 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X26 D G S_uq22 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X27 D G S_uq19 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X28 D G S_uq17 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X29 D G S_uq14 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X30 D G S_uq12 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X31 S_uq25 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X32 S_uq8 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X33 S_uq5 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X34 S_uq3 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X35 S G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X36 S_uq10 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X37 S_uq20 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X38 S_uq17 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X39 S_uq15 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X40 S_uq12 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X41 S_uq7 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X42 S_uq24 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X43 S_uq22 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X44 S_uq19 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X45 D G S_uq27 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X46 D G S_uq26 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X47 D G S_uq6 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X48 D G S_uq1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X49 D G S_uq4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X50 D G S_uq2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X51 D G S_uq0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X52 D G S_uq23 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X53 D G S_uq21 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X54 D G S_uq20 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X55 D G S_uq18 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X56 D G S_uq16 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X57 D G S_uq13 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X58 D G S_uq11 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X59 D G S_uq9 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
X60 S_uq27 G D gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=495000u l=150000u
.ends

.subckt pmos_m61_w1_485_sli_dli_da_p w_n59_65# S S_uq0 S_uq1 S_uq3 S_uq2 S_uq20 S_uq4
+ S_uq21 S_uq10 S_uq5 S_uq22 S_uq11 S_uq6 S_uq24 S_uq23 S_uq13 S_uq12 S_uq7 S_uq25
+ S_uq14 S_uq8 S_uq26 S_uq15 S_uq9 S_uq27 S_uq16 S_uq28 S_uq17 gnd S_uq29 S_uq18 S_uq19
+ D G
X0 D G S_uq28 w_n59_65# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.485e+06u l=150000u
X1 S_uq21 G D w_n59_65# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.485e+06u l=150000u
X2 S_uq16 G D w_n59_65# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.485e+06u l=150000u
X3 S_uq11 G D w_n59_65# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.485e+06u l=150000u
X4 D G S_uq25 w_n59_65# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.485e+06u l=150000u
X5 D G S_uq8 w_n59_65# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.485e+06u l=150000u
X6 D G S_uq3 w_n59_65# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.485e+06u l=150000u
X7 D G S w_n59_65# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.485e+06u l=150000u
X8 D G S_uq15 w_n59_65# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.485e+06u l=150000u
X9 D G S_uq10 w_n59_65# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.485e+06u l=150000u
X10 D G S_uq5 w_n59_65# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.485e+06u l=150000u
X11 D G S_uq12 w_n59_65# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.485e+06u l=150000u
X12 D G S_uq7 w_n59_65# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.485e+06u l=150000u
X13 S_uq28 G D w_n59_65# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.485e+06u l=150000u
X14 D G S_uq24 w_n59_65# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.485e+06u l=150000u
X15 D G S_uq22 w_n59_65# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.485e+06u l=150000u
X16 D G S_uq19 w_n59_65# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.485e+06u l=150000u
X17 D G S_uq17 w_n59_65# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.485e+06u l=150000u
X18 D G S_uq14 w_n59_65# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.485e+06u l=150000u
X19 S_uq25 G D w_n59_65# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.485e+06u l=150000u
X20 S_uq10 G D w_n59_65# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.485e+06u l=150000u
X21 S_uq8 G D w_n59_65# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.485e+06u l=150000u
X22 S_uq5 G D w_n59_65# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.485e+06u l=150000u
X23 S_uq3 G D w_n59_65# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.485e+06u l=150000u
X24 S G D w_n59_65# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.485e+06u l=150000u
X25 S_uq22 G D w_n59_65# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.485e+06u l=150000u
X26 S_uq20 G D w_n59_65# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.485e+06u l=150000u
X27 S_uq17 G D w_n59_65# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.485e+06u l=150000u
X28 S_uq15 G D w_n59_65# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.485e+06u l=150000u
X29 S_uq12 G D w_n59_65# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.485e+06u l=150000u
X30 S_uq7 G D w_n59_65# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.485e+06u l=150000u
X31 S_uq24 G D w_n59_65# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.485e+06u l=150000u
X32 S_uq19 G D w_n59_65# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.485e+06u l=150000u
X33 D G S_uq27 w_n59_65# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.485e+06u l=150000u
X34 D G S_uq26 w_n59_65# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.485e+06u l=150000u
X35 D G S_uq6 w_n59_65# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.485e+06u l=150000u
X36 D G S_uq1 w_n59_65# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.485e+06u l=150000u
X37 D G S_uq11 w_n59_65# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.485e+06u l=150000u
X38 D G S_uq9 w_n59_65# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.485e+06u l=150000u
X39 D G S_uq4 w_n59_65# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.485e+06u l=150000u
X40 D G S_uq2 w_n59_65# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.485e+06u l=150000u
X41 D G S_uq0 w_n59_65# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.485e+06u l=150000u
X42 D G S_uq23 w_n59_65# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.485e+06u l=150000u
X43 D G S_uq21 w_n59_65# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.485e+06u l=150000u
X44 D G S_uq20 w_n59_65# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.485e+06u l=150000u
X45 D G S_uq18 w_n59_65# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.485e+06u l=150000u
X46 D G S_uq16 w_n59_65# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.485e+06u l=150000u
X47 D G S_uq13 w_n59_65# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.485e+06u l=150000u
X48 S_uq27 G D w_n59_65# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.485e+06u l=150000u
X49 S_uq26 G D w_n59_65# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.485e+06u l=150000u
X50 S_uq14 G D w_n59_65# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.485e+06u l=150000u
X51 S_uq13 G D w_n59_65# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.485e+06u l=150000u
X52 S_uq9 G D w_n59_65# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.485e+06u l=150000u
X53 S_uq4 G D w_n59_65# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.485e+06u l=150000u
X54 S_uq2 G D w_n59_65# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.485e+06u l=150000u
X55 S_uq1 G D w_n59_65# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.485e+06u l=150000u
X56 S_uq0 G D w_n59_65# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.485e+06u l=150000u
X57 D G S_uq29 w_n59_65# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.485e+06u l=150000u
X58 S_uq23 G D w_n59_65# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.485e+06u l=150000u
X59 S_uq18 G D w_n59_65# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.485e+06u l=150000u
X60 S_uq6 G D w_n59_65# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.485e+06u l=150000u
.ends

.subckt pinv_10 Z gnd vdd A
Xnmos_m61_w0_495_sli_dli_da_p_0 gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd
+ gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd Z A
+ nmos_m61_w0_495_sli_dli_da_p
Xpmos_m61_w1_485_sli_dli_da_p_0 vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd
+ vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd gnd vdd vdd vdd
+ Z A pmos_m61_w1_485_sli_dli_da_p
.ends

.subckt pdriver_0 A vdd Z gnd
Xpinv_9_0 gnd pinv_9_0/Z vdd pinv_9_0/A pinv_9
Xpinv_7_0 pinv_8_0/A gnd vdd pinv_7_0/A pinv_7
Xpinv_8_0 vdd pinv_9_0/A gnd pinv_8_0/A pinv_8
Xpinv_6_0 pinv_6_1/Z pinv_7_0/A gnd vdd pinv_6
Xpinv_6_1 A pinv_6_1/Z gnd vdd pinv_6
Xpinv_10_0 Z gnd vdd pinv_9_0/Z pinv_10
.ends

.subckt pinv_0 A Z gnd vdd
Xnmos_m1_w0_420_sli_dli_da_p_0 gnd gnd Z A nmos_m1_w0_420_sli_dli_da_p
Xpmos_m1_w1_260_sli_dli_da_p_0 vdd vdd gnd Z A pmos_m1_w1_260_sli_dli_da_p
.ends

.subckt control_logic_multiport p_en_bar clk web vdd csb wl_en w_en
Xdff_buf_array_0 vdd dff_buf_array_0/dout_0 dff_buf_array_0/dout_1 pand2_0_0/A pand2_1/B
+ web csb dff_buf_array
Xpand2_0_0 pand2_0/vdd w_en vdd pand2_0_0/A pand2_1/Z pand2_0
Xpdriver_1_0 vdd pnand2_1_0/Z pnand2_1_0/vdd p_en_bar pdriver_1
Xpdriver_1_1 vdd pand2_1/Z pnand2_1_0/vdd wl_en pdriver_1
Xpand2_0 pand2_0/vdd vdd pand2_0/Z vdd pand2_1/B pand2
Xpand2_1 pand2_1/vdd vdd pand2_1/Z pand2_1/A pand2_1/B pand2
Xpnand2_1_0 pnand2_1_0/Z vdd pnand2_1_0/vdd pand2_0/Z pnand2_1
Xpdriver_0_0 clk pand2_1/vdd vdd vdd pdriver_0
Xpinv_0_0 vdd pand2_1/A vdd pand2_1/vdd pinv_0
.ends

.subckt data_dff din_7 clk din_8 vdd din_9 din_30 gnd din_31 din_20 din_21 din_10
+ din_22 din_11 din_23 din_12 din_24 din_13 din_25 din_14 din_26 din_15 din_27 din_16
+ din_28 din_17 din_29 din_18 din_19 din_0 din_1 din_2 din_3 din_4 din_5 din_6
Xdff_19 clk vdd gnd din_12 dout_12 dff
Xdff_0 clk vdd gnd din_31 dout_31 dff
Xdff_1 clk vdd gnd din_30 dout_30 dff
Xdff_2 clk vdd gnd din_29 dout_29 dff
Xdff_3 clk vdd gnd din_28 dout_28 dff
Xdff_4 clk vdd gnd din_27 dout_27 dff
Xdff_5 clk vdd gnd din_26 dout_26 dff
Xdff_6 clk vdd gnd din_25 dout_25 dff
Xdff_7 clk vdd gnd din_24 dout_24 dff
Xdff_8 clk vdd gnd din_23 dout_23 dff
Xdff_9 clk vdd gnd din_22 dout_22 dff
Xdff_30 clk vdd gnd din_1 dout_1 dff
Xdff_31 clk vdd gnd din_0 dout_0 dff
Xdff_20 clk vdd gnd din_11 dout_11 dff
Xdff_10 clk vdd gnd din_21 dout_21 dff
Xdff_21 clk vdd gnd din_10 dout_10 dff
Xdff_11 clk vdd gnd din_20 dout_20 dff
Xdff_22 clk vdd gnd din_9 dout_9 dff
Xdff_12 clk vdd gnd din_19 dout_19 dff
Xdff_23 clk vdd gnd din_8 dout_8 dff
Xdff_13 clk vdd gnd din_18 dout_18 dff
Xdff_24 clk vdd gnd din_7 dout_7 dff
Xdff_14 clk vdd gnd din_17 dout_17 dff
Xdff_25 clk vdd gnd din_6 dout_6 dff
Xdff_15 clk vdd gnd din_16 dout_16 dff
Xdff_26 clk vdd gnd din_5 dout_5 dff
Xdff_27 clk vdd gnd din_4 dout_4 dff
Xdff_16 clk vdd gnd din_15 dout_15 dff
Xdff_28 clk vdd gnd din_3 dout_3 dff
Xdff_17 clk vdd gnd din_14 dout_14 dff
Xdff_29 clk vdd gnd din_2 dout_2 dff
Xdff_18 clk vdd gnd din_13 dout_13 dff
.ends

.subckt col_addr_dff clk gnd vdd din_0
Xdff_0 clk vdd gnd din_0 dout_0 dff
.ends

.subckt row_addr_dff din_7 vdd_uq0 vdd_uq1 vdd_uq2 clk vdd_uq3 dout_0 dout_1 dout_3
+ dout_2 gnd dout_4 dout_5 dout_6 dout_7 vdd din_0 din_1 din_2 din_3 din_4 din_5 din_6
Xdff_0 clk vdd_uq3 gnd din_9 dout_9 dff
Xdff_1 clk vdd_uq3 gnd din_8 dout_8 dff
Xdff_2 clk vdd_uq2 gnd din_7 dout_7 dff
Xdff_3 clk vdd_uq2 gnd din_6 dout_6 dff
Xdff_4 clk vdd_uq1 gnd din_5 dout_5 dff
Xdff_5 clk vdd_uq1 gnd din_4 dout_4 dff
Xdff_6 clk vdd gnd din_3 dout_3 dff
Xdff_7 clk vdd gnd din_2 dout_2 dff
Xdff_8 clk vdd_uq0 gnd din_1 dout_1 dff
Xdff_9 clk vdd_uq0 gnd din_0 dout_0 dff
.ends

.subckt sense_amp_multiport vdd gnd rbl dout
X0 dout rbl gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 dout rbl vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.7e+06u l=150000u
.ends

.subckt sense_amp_array vdd vdd_uq2 data_30 data_31 data_20 vdd_uq4 data_10 data_21
+ data_11 data_22 vdd_uq6 data_12 data_23 data_13 data_24 data_14 data_25 vdd_uq8
+ data_15 data_26 data_27 data_16 vdd_uq9 data_28 data_17 data_29 data_18 data_19
+ gnd vdd_uq60 vdd_uq62 vdd_uq52 vdd_uq42 vdd_uq54 vdd_uq32 data_0 vdd_uq44 vdd_uq22
+ data_1 vdd_uq56 vdd_uq34 vdd_uq12 data_2 vdd_uq46 vdd_uq24 data_3 vdd_uq58 vdd_uq36
+ vdd_uq14 data_4 vdd_uq48 vdd_uq26 data_5 vdd_uq38 vdd_uq16 data_6 vdd_uq50 vdd_uq28
+ data_7 vdd_uq40 vdd_uq18 data_8 vdd_uq30 data_9 vdd_uq20
Xsense_amp_multiport_60 vdd_uq60 gnd rbl_3 data_3 sense_amp_multiport
Xsense_amp_multiport_61 vdd_uq60 gnd rbl_2 data_2 sense_amp_multiport
Xsense_amp_multiport_50 vdd_uq50 gnd rbl_13 data_13 sense_amp_multiport
Xsense_amp_multiport_40 vdd_uq40 gnd rbl_23 data_23 sense_amp_multiport
Xsense_amp_multiport_62 vdd_uq62 gnd rbl_1 data_1 sense_amp_multiport
Xsense_amp_multiport_51 vdd_uq50 gnd rbl_12 data_12 sense_amp_multiport
Xsense_amp_multiport_30 vdd_uq30 gnd rbl_33 data_33 sense_amp_multiport
Xsense_amp_multiport_41 vdd_uq40 gnd rbl_22 data_22 sense_amp_multiport
Xsense_amp_multiport_63 vdd_uq62 gnd rbl_0 data_0 sense_amp_multiport
Xsense_amp_multiport_52 vdd_uq52 gnd rbl_11 data_11 sense_amp_multiport
Xsense_amp_multiport_0 vdd gnd rbl_63 data_63 sense_amp_multiport
Xsense_amp_multiport_20 vdd_uq20 gnd rbl_43 data_43 sense_amp_multiport
Xsense_amp_multiport_31 vdd_uq30 gnd rbl_32 data_32 sense_amp_multiport
Xsense_amp_multiport_42 vdd_uq42 gnd rbl_21 data_21 sense_amp_multiport
Xsense_amp_multiport_53 vdd_uq52 gnd rbl_10 data_10 sense_amp_multiport
Xsense_amp_multiport_10 vdd_uq9 gnd rbl_53 data_53 sense_amp_multiport
Xsense_amp_multiport_21 vdd_uq20 gnd rbl_42 data_42 sense_amp_multiport
Xsense_amp_multiport_32 vdd_uq32 gnd rbl_31 data_31 sense_amp_multiport
Xsense_amp_multiport_43 vdd_uq42 gnd rbl_20 data_20 sense_amp_multiport
Xsense_amp_multiport_54 vdd_uq54 gnd rbl_9 data_9 sense_amp_multiport
Xsense_amp_multiport_1 vdd gnd rbl_62 data_62 sense_amp_multiport
Xsense_amp_multiport_2 vdd_uq2 gnd rbl_61 data_61 sense_amp_multiport
Xsense_amp_multiport_11 vdd_uq9 gnd rbl_52 data_52 sense_amp_multiport
Xsense_amp_multiport_22 vdd_uq22 gnd rbl_41 data_41 sense_amp_multiport
Xsense_amp_multiport_33 vdd_uq32 gnd rbl_30 data_30 sense_amp_multiport
Xsense_amp_multiport_55 vdd_uq54 gnd rbl_8 data_8 sense_amp_multiport
Xsense_amp_multiport_44 vdd_uq44 gnd rbl_19 data_19 sense_amp_multiport
Xsense_amp_multiport_12 vdd_uq12 gnd rbl_51 data_51 sense_amp_multiport
Xsense_amp_multiport_23 vdd_uq22 gnd rbl_40 data_40 sense_amp_multiport
Xsense_amp_multiport_34 vdd_uq34 gnd rbl_29 data_29 sense_amp_multiport
Xsense_amp_multiport_56 vdd_uq56 gnd rbl_7 data_7 sense_amp_multiport
Xsense_amp_multiport_45 vdd_uq44 gnd rbl_18 data_18 sense_amp_multiport
Xsense_amp_multiport_3 vdd_uq2 gnd rbl_60 data_60 sense_amp_multiport
Xsense_amp_multiport_13 vdd_uq12 gnd rbl_50 data_50 sense_amp_multiport
Xsense_amp_multiport_24 vdd_uq24 gnd rbl_39 data_39 sense_amp_multiport
Xsense_amp_multiport_35 vdd_uq34 gnd rbl_28 data_28 sense_amp_multiport
Xsense_amp_multiport_57 vdd_uq56 gnd rbl_6 data_6 sense_amp_multiport
Xsense_amp_multiport_46 vdd_uq46 gnd rbl_17 data_17 sense_amp_multiport
Xsense_amp_multiport_4 vdd_uq4 gnd rbl_59 data_59 sense_amp_multiport
Xsense_amp_multiport_14 vdd_uq14 gnd rbl_49 data_49 sense_amp_multiport
Xsense_amp_multiport_25 vdd_uq24 gnd rbl_38 data_38 sense_amp_multiport
Xsense_amp_multiport_36 vdd_uq36 gnd rbl_27 data_27 sense_amp_multiport
Xsense_amp_multiport_58 vdd_uq58 gnd rbl_5 data_5 sense_amp_multiport
Xsense_amp_multiport_47 vdd_uq46 gnd rbl_16 data_16 sense_amp_multiport
Xsense_amp_multiport_5 vdd_uq4 gnd rbl_58 data_58 sense_amp_multiport
Xsense_amp_multiport_15 vdd_uq14 gnd rbl_48 data_48 sense_amp_multiport
Xsense_amp_multiport_26 vdd_uq26 gnd rbl_37 data_37 sense_amp_multiport
Xsense_amp_multiport_37 vdd_uq36 gnd rbl_26 data_26 sense_amp_multiport
Xsense_amp_multiport_59 vdd_uq58 gnd rbl_4 data_4 sense_amp_multiport
Xsense_amp_multiport_48 vdd_uq48 gnd rbl_15 data_15 sense_amp_multiport
Xsense_amp_multiport_6 vdd_uq6 gnd rbl_57 data_57 sense_amp_multiport
Xsense_amp_multiport_7 vdd_uq6 gnd rbl_56 data_56 sense_amp_multiport
Xsense_amp_multiport_16 vdd_uq16 gnd rbl_47 data_47 sense_amp_multiport
Xsense_amp_multiport_27 vdd_uq26 gnd rbl_36 data_36 sense_amp_multiport
Xsense_amp_multiport_38 vdd_uq38 gnd rbl_25 data_25 sense_amp_multiport
Xsense_amp_multiport_49 vdd_uq48 gnd rbl_14 data_14 sense_amp_multiport
Xsense_amp_multiport_17 vdd_uq16 gnd rbl_46 data_46 sense_amp_multiport
Xsense_amp_multiport_28 vdd_uq28 gnd rbl_35 data_35 sense_amp_multiport
Xsense_amp_multiport_39 vdd_uq38 gnd rbl_24 data_24 sense_amp_multiport
Xsense_amp_multiport_8 vdd_uq8 gnd rbl_55 data_55 sense_amp_multiport
Xsense_amp_multiport_9 vdd_uq8 gnd rbl_54 data_54 sense_amp_multiport
Xsense_amp_multiport_18 vdd_uq18 gnd rbl_45 data_45 sense_amp_multiport
Xsense_amp_multiport_29 vdd_uq28 gnd rbl_34 data_34 sense_amp_multiport
Xsense_amp_multiport_19 vdd_uq18 gnd rbl_44 data_44 sense_amp_multiport
.ends

.subckt nmos_m1_w3_360_sli_dli S gnd D G
X0 D G S gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3.36e+06u l=150000u
.ends

.subckt column_mux_multiport rbl1_out sel rbl0_out gnd rbl0 rbl1
Xnmos_m1_w3_360_sli_dli_0 nmos_m1_w3_360_sli_dli_0/S gnd rbl0 sel nmos_m1_w3_360_sli_dli
Xnmos_m1_w3_360_sli_dli_1 rbl1_out gnd nmos_m1_w3_360_sli_dli_1/D sel nmos_m1_w3_360_sli_dli
.ends

.subckt column_mux_array_multiport rbl0_0 rbl0_60 sel_1 rbl0_61 rbl0_50 rbl0_1 sel_0
+ rbl0_2 rbl0_40 rbl0_62 rbl0_51 rbl0_30 rbl0_41 rbl0_63 rbl0_52 rbl0_3 rbl0_4 rbl0_20
+ rbl0_31 rbl0_42 rbl0_53 rbl0_10 rbl0_21 rbl0_32 rbl0_43 rbl0_54 rbl0_5 rbl0_6 rbl0_11
+ rbl0_22 rbl0_33 rbl0_44 rbl0_55 rbl0_12 rbl0_23 rbl0_34 rbl0_45 rbl0_56 rbl0_7 rbl0_8
+ rbl0_13 rbl0_24 rbl0_35 rbl0_46 rbl0_57 rbl0_14 rbl0_25 rbl0_36 rbl0_47 rbl0_58
+ rbl0_9 rbl0_15 rbl0_26 rbl0_37 rbl0_59 rbl0_48 rbl0_16 rbl0_27 rbl0_38 rbl0_49 rbl0_17
+ rbl0_28 rbl0_39 rbl1_60 rbl0_18 rbl0_29 rbl1_61 rbl1_50 rbl0_19 rbl1_40 rbl1_62
+ rbl1_51 rbl1_30 rbl1_41 rbl1_63 rbl1_52 rbl1_20 rbl1_31 rbl1_42 rbl1_53 rbl1_0 rbl1_10
+ rbl1_21 rbl1_32 rbl1_43 rbl1_54 rbl1_1 rbl1_11 rbl1_22 rbl1_33 rbl1_44 rbl1_55 rbl1_2
+ gnd rbl1_12 rbl1_23 rbl1_34 rbl1_45 rbl1_56 rbl1_3 rbl1_13 rbl1_24 rbl1_35 rbl1_46
+ rbl1_57 rbl1_4 rbl1_14 rbl1_25 rbl1_36 rbl1_47 rbl1_58 rbl1_5 rbl1_15 rbl1_26 rbl1_37
+ rbl1_59 rbl1_48 rbl1_6 rbl1_16 rbl1_27 rbl1_38 rbl1_49 rbl1_7 rbl1_17 rbl1_28 rbl1_39
+ rbl1_8 rbl1_18 rbl1_29 rbl1_9 rbl1_19
Xcolumn_mux_multiport_60 rbl1_out_1 sel_1 rbl0_out_1 gnd rbl0_3 rbl1_3 column_mux_multiport
Xcolumn_mux_multiport_0 rbl1_out_31 sel_1 rbl0_out_31 gnd rbl0_63 rbl1_63 column_mux_multiport
Xcolumn_mux_multiport_61 rbl1_out_1 sel_0 rbl0_out_1 gnd rbl0_2 rbl1_2 column_mux_multiport
Xcolumn_mux_multiport_50 rbl1_out_6 sel_1 rbl0_out_6 gnd rbl0_13 rbl1_13 column_mux_multiport
Xcolumn_mux_multiport_1 rbl1_out_31 sel_0 rbl0_out_31 gnd rbl0_62 rbl1_62 column_mux_multiport
Xcolumn_mux_multiport_40 rbl1_out_11 sel_1 rbl0_out_11 gnd rbl0_23 rbl1_23 column_mux_multiport
Xcolumn_mux_multiport_62 rbl1_out_0 sel_1 rbl0_out_0 gnd rbl0_1 rbl1_1 column_mux_multiport
Xcolumn_mux_multiport_51 rbl1_out_6 sel_0 rbl0_out_6 gnd rbl0_12 rbl1_12 column_mux_multiport
Xcolumn_mux_multiport_2 rbl1_out_30 sel_1 rbl0_out_30 gnd rbl0_61 rbl1_61 column_mux_multiport
Xcolumn_mux_multiport_30 rbl1_out_16 sel_1 rbl0_out_16 gnd rbl0_33 rbl1_33 column_mux_multiport
Xcolumn_mux_multiport_41 rbl1_out_11 sel_0 rbl0_out_11 gnd rbl0_22 rbl1_22 column_mux_multiport
Xcolumn_mux_multiport_63 rbl1_out_0 sel_0 rbl0_out_0 gnd rbl0_0 rbl1_0 column_mux_multiport
Xcolumn_mux_multiport_52 rbl1_out_5 sel_1 rbl0_out_5 gnd rbl0_11 rbl1_11 column_mux_multiport
Xcolumn_mux_multiport_3 rbl1_out_30 sel_0 rbl0_out_30 gnd rbl0_60 rbl1_60 column_mux_multiport
Xcolumn_mux_multiport_20 rbl1_out_21 sel_1 rbl0_out_21 gnd rbl0_43 rbl1_43 column_mux_multiport
Xcolumn_mux_multiport_31 rbl1_out_16 sel_0 rbl0_out_16 gnd rbl0_32 rbl1_32 column_mux_multiport
Xcolumn_mux_multiport_42 rbl1_out_10 sel_1 rbl0_out_10 gnd rbl0_21 rbl1_21 column_mux_multiport
Xcolumn_mux_multiport_53 rbl1_out_5 sel_0 rbl0_out_5 gnd rbl0_10 rbl1_10 column_mux_multiport
Xcolumn_mux_multiport_4 rbl1_out_29 sel_1 rbl0_out_29 gnd rbl0_59 rbl1_59 column_mux_multiport
Xcolumn_mux_multiport_10 rbl1_out_26 sel_1 rbl0_out_26 gnd rbl0_53 rbl1_53 column_mux_multiport
Xcolumn_mux_multiport_21 rbl1_out_21 sel_0 rbl0_out_21 gnd rbl0_42 rbl1_42 column_mux_multiport
Xcolumn_mux_multiport_32 rbl1_out_15 sel_1 rbl0_out_15 gnd rbl0_31 rbl1_31 column_mux_multiport
Xcolumn_mux_multiport_43 rbl1_out_10 sel_0 rbl0_out_10 gnd rbl0_20 rbl1_20 column_mux_multiport
Xcolumn_mux_multiport_54 rbl1_out_4 sel_1 rbl0_out_4 gnd rbl0_9 rbl1_9 column_mux_multiport
Xcolumn_mux_multiport_5 rbl1_out_29 sel_0 rbl0_out_29 gnd rbl0_58 rbl1_58 column_mux_multiport
Xcolumn_mux_multiport_11 rbl1_out_26 sel_0 rbl0_out_26 gnd rbl0_52 rbl1_52 column_mux_multiport
Xcolumn_mux_multiport_22 rbl1_out_20 sel_1 rbl0_out_20 gnd rbl0_41 rbl1_41 column_mux_multiport
Xcolumn_mux_multiport_33 rbl1_out_15 sel_0 rbl0_out_15 gnd rbl0_30 rbl1_30 column_mux_multiport
Xcolumn_mux_multiport_55 rbl1_out_4 sel_0 rbl0_out_4 gnd rbl0_8 rbl1_8 column_mux_multiport
Xcolumn_mux_multiport_44 rbl1_out_9 sel_1 rbl0_out_9 gnd rbl0_19 rbl1_19 column_mux_multiport
Xcolumn_mux_multiport_6 rbl1_out_28 sel_1 rbl0_out_28 gnd rbl0_57 rbl1_57 column_mux_multiport
Xcolumn_mux_multiport_12 rbl1_out_25 sel_1 rbl0_out_25 gnd rbl0_51 rbl1_51 column_mux_multiport
Xcolumn_mux_multiport_23 rbl1_out_20 sel_0 rbl0_out_20 gnd rbl0_40 rbl1_40 column_mux_multiport
Xcolumn_mux_multiport_34 rbl1_out_14 sel_1 rbl0_out_14 gnd rbl0_29 rbl1_29 column_mux_multiport
Xcolumn_mux_multiport_56 rbl1_out_3 sel_1 rbl0_out_3 gnd rbl0_7 rbl1_7 column_mux_multiport
Xcolumn_mux_multiport_45 rbl1_out_9 sel_0 rbl0_out_9 gnd rbl0_18 rbl1_18 column_mux_multiport
Xcolumn_mux_multiport_7 rbl1_out_28 sel_0 rbl0_out_28 gnd rbl0_56 rbl1_56 column_mux_multiport
Xcolumn_mux_multiport_13 rbl1_out_25 sel_0 rbl0_out_25 gnd rbl0_50 rbl1_50 column_mux_multiport
Xcolumn_mux_multiport_24 rbl1_out_19 sel_1 rbl0_out_19 gnd rbl0_39 rbl1_39 column_mux_multiport
Xcolumn_mux_multiport_35 rbl1_out_14 sel_0 rbl0_out_14 gnd rbl0_28 rbl1_28 column_mux_multiport
Xcolumn_mux_multiport_57 rbl1_out_3 sel_0 rbl0_out_3 gnd rbl0_6 rbl1_6 column_mux_multiport
Xcolumn_mux_multiport_46 rbl1_out_8 sel_1 rbl0_out_8 gnd rbl0_17 rbl1_17 column_mux_multiport
Xcolumn_mux_multiport_8 rbl1_out_27 sel_1 rbl0_out_27 gnd rbl0_55 rbl1_55 column_mux_multiport
Xcolumn_mux_multiport_14 rbl1_out_24 sel_1 rbl0_out_24 gnd rbl0_49 rbl1_49 column_mux_multiport
Xcolumn_mux_multiport_25 rbl1_out_19 sel_0 rbl0_out_19 gnd rbl0_38 rbl1_38 column_mux_multiport
Xcolumn_mux_multiport_36 rbl1_out_13 sel_1 rbl0_out_13 gnd rbl0_27 rbl1_27 column_mux_multiport
Xcolumn_mux_multiport_58 rbl1_out_2 sel_1 rbl0_out_2 gnd rbl0_5 rbl1_5 column_mux_multiport
Xcolumn_mux_multiport_47 rbl1_out_8 sel_0 rbl0_out_8 gnd rbl0_16 rbl1_16 column_mux_multiport
Xcolumn_mux_multiport_9 rbl1_out_27 sel_0 rbl0_out_27 gnd rbl0_54 rbl1_54 column_mux_multiport
Xcolumn_mux_multiport_15 rbl1_out_24 sel_0 rbl0_out_24 gnd rbl0_48 rbl1_48 column_mux_multiport
Xcolumn_mux_multiport_26 rbl1_out_18 sel_1 rbl0_out_18 gnd rbl0_37 rbl1_37 column_mux_multiport
Xcolumn_mux_multiport_37 rbl1_out_13 sel_0 rbl0_out_13 gnd rbl0_26 rbl1_26 column_mux_multiport
Xcolumn_mux_multiport_59 rbl1_out_2 sel_0 rbl0_out_2 gnd rbl0_4 rbl1_4 column_mux_multiport
Xcolumn_mux_multiport_48 rbl1_out_7 sel_1 rbl0_out_7 gnd rbl0_15 rbl1_15 column_mux_multiport
Xcolumn_mux_multiport_16 rbl1_out_23 sel_1 rbl0_out_23 gnd rbl0_47 rbl1_47 column_mux_multiport
Xcolumn_mux_multiport_27 rbl1_out_18 sel_0 rbl0_out_18 gnd rbl0_36 rbl1_36 column_mux_multiport
Xcolumn_mux_multiport_38 rbl1_out_12 sel_1 rbl0_out_12 gnd rbl0_25 rbl1_25 column_mux_multiport
Xcolumn_mux_multiport_49 rbl1_out_7 sel_0 rbl0_out_7 gnd rbl0_14 rbl1_14 column_mux_multiport
Xcolumn_mux_multiport_17 rbl1_out_23 sel_0 rbl0_out_23 gnd rbl0_46 rbl1_46 column_mux_multiport
Xcolumn_mux_multiport_28 rbl1_out_17 sel_1 rbl0_out_17 gnd rbl0_35 rbl1_35 column_mux_multiport
Xcolumn_mux_multiport_39 rbl1_out_12 sel_0 rbl0_out_12 gnd rbl0_24 rbl1_24 column_mux_multiport
Xcolumn_mux_multiport_18 rbl1_out_22 sel_1 rbl0_out_22 gnd rbl0_45 rbl1_45 column_mux_multiport
Xcolumn_mux_multiport_29 rbl1_out_17 sel_0 rbl0_out_17 gnd rbl0_34 rbl1_34 column_mux_multiport
Xcolumn_mux_multiport_19 rbl1_out_22 sel_0 rbl0_out_22 gnd rbl0_44 rbl1_44 column_mux_multiport
.ends

.subckt write_driver_multiport din vdd gnd en wbl
X0 net2 net1 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.35e+06u l=150000u
X1 net1 din gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 wbl en a_478_138# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 gnd en enb gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_478_138# net1 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 net1 din vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.35e+06u l=150000u
X6 wbl enb net2 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.35e+06u l=150000u
X7 vdd en enb vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.35e+06u l=150000u
.ends

.subckt write_driver_array din_7 din_8 vdd_uq0 din_9 vdd_uq1 en vdd_uq2 vdd_uq3 vdd_uq4
+ vdd_uq5 vdd_uq6 vdd_uq7 vdd_uq8 vdd_uq9 wbl0_0 wbl0_1 din_30 gnd din_31 din_20 din_21
+ din_10 din_22 din_11 din_23 din_12 vdd_uq30 din_24 din_13 din_25 din_14 vdd_uq20
+ vdd_uq21 vdd_uq10 din_26 din_15 din_27 din_16 vdd_uq22 vdd_uq11 vdd_uq23 vdd_uq12
+ din_28 din_17 din_29 din_18 vdd_uq24 vdd_uq13 vdd vdd_uq25 vdd_uq14 din_19 din_0
+ vdd_uq26 vdd_uq15 din_1 vdd_uq16 vdd_uq27 din_2 vdd_uq28 vdd_uq17 din_3 vdd_uq29
+ vdd_uq18 din_4 vdd_uq19 din_5 din_6
Xwrite_driver_multiport_30 din_1 vdd_uq29 gnd en wbl0_1 write_driver_multiport
Xwrite_driver_multiport_31 din_0 vdd_uq30 gnd en wbl0_0 write_driver_multiport
Xwrite_driver_multiport_20 din_11 vdd_uq19 gnd en wbl0_11 write_driver_multiport
Xwrite_driver_multiport_10 din_21 vdd_uq9 gnd en wbl0_21 write_driver_multiport
Xwrite_driver_multiport_21 din_10 vdd_uq20 gnd en wbl0_10 write_driver_multiport
Xwrite_driver_multiport_11 din_20 vdd_uq10 gnd en wbl0_20 write_driver_multiport
Xwrite_driver_multiport_22 din_9 vdd_uq21 gnd en wbl0_9 write_driver_multiport
Xwrite_driver_multiport_23 din_8 vdd_uq22 gnd en wbl0_8 write_driver_multiport
Xwrite_driver_multiport_12 din_19 vdd_uq11 gnd en wbl0_19 write_driver_multiport
Xwrite_driver_multiport_0 din_31 vdd_uq0 gnd en wbl0_31 write_driver_multiport
Xwrite_driver_multiport_24 din_7 vdd_uq23 gnd en wbl0_7 write_driver_multiport
Xwrite_driver_multiport_13 din_18 vdd_uq12 gnd en wbl0_18 write_driver_multiport
Xwrite_driver_multiport_1 din_30 vdd gnd en wbl0_30 write_driver_multiport
Xwrite_driver_multiport_25 din_6 vdd_uq24 gnd en wbl0_6 write_driver_multiport
Xwrite_driver_multiport_14 din_17 vdd_uq13 gnd en wbl0_17 write_driver_multiport
Xwrite_driver_multiport_2 din_29 vdd_uq1 gnd en wbl0_29 write_driver_multiport
Xwrite_driver_multiport_26 din_5 vdd_uq25 gnd en wbl0_5 write_driver_multiport
Xwrite_driver_multiport_15 din_16 vdd_uq14 gnd en wbl0_16 write_driver_multiport
Xwrite_driver_multiport_3 din_28 vdd_uq2 gnd en wbl0_28 write_driver_multiport
Xwrite_driver_multiport_27 din_4 vdd_uq26 gnd en wbl0_4 write_driver_multiport
Xwrite_driver_multiport_16 din_15 vdd_uq15 gnd en wbl0_15 write_driver_multiport
Xwrite_driver_multiport_4 din_27 vdd_uq3 gnd en wbl0_27 write_driver_multiport
Xwrite_driver_multiport_28 din_3 vdd_uq27 gnd en wbl0_3 write_driver_multiport
Xwrite_driver_multiport_17 din_14 vdd_uq16 gnd en wbl0_14 write_driver_multiport
Xwrite_driver_multiport_5 din_26 vdd_uq4 gnd en wbl0_26 write_driver_multiport
Xwrite_driver_multiport_29 din_2 vdd_uq28 gnd en wbl0_2 write_driver_multiport
Xwrite_driver_multiport_18 din_13 vdd_uq17 gnd en wbl0_13 write_driver_multiport
Xwrite_driver_multiport_6 din_25 vdd_uq5 gnd en wbl0_25 write_driver_multiport
Xwrite_driver_multiport_19 din_12 vdd_uq18 gnd en wbl0_12 write_driver_multiport
Xwrite_driver_multiport_7 din_24 vdd_uq6 gnd en wbl0_24 write_driver_multiport
Xwrite_driver_multiport_8 din_23 vdd_uq7 gnd en wbl0_23 write_driver_multiport
Xwrite_driver_multiport_9 din_22 vdd_uq8 gnd en wbl0_22 write_driver_multiport
.ends

.subckt precharge_multiport_0 en_bar rbl1 gnd rbl0 vdd
Xpmos_m1_w1_260_sli_dli_0 vdd vdd gnd rbl1 en_bar pmos_m1_w1_260_sli_dli
Xpmos_m1_w1_260_sli_dli_1 vdd rbl0 gnd vdd en_bar pmos_m1_w1_260_sli_dli
Xpmos_m1_w1_260_sli_dli_2 vdd rbl0 gnd rbl1 en_bar pmos_m1_w1_260_sli_dli
.ends

.subckt precharge_array_multiport rbl0_0 rbl0_60 en_bar rbl0_61 rbl0_50 rbl0_1 vdd
+ rbl0_2 rbl0_40 rbl0_62 rbl0_51 rbl0_30 rbl0_41 rbl0_63 rbl0_52 rbl0_3 rbl0_4 rbl0_20
+ rbl0_31 rbl0_42 rbl0_53 rbl0_10 rbl0_21 rbl0_32 rbl0_43 rbl0_54 rbl0_5 rbl0_6 rbl0_11
+ rbl0_22 rbl0_33 rbl0_44 rbl0_55 rbl0_12 rbl0_23 rbl0_34 rbl0_45 rbl0_56 rbl0_7 rbl0_8
+ rbl0_13 rbl0_24 rbl0_35 rbl0_46 rbl0_57 rbl0_14 rbl0_25 rbl0_36 rbl0_47 rbl0_58
+ rbl0_9 rbl0_15 rbl0_26 rbl0_37 rbl0_48 rbl0_59 rbl0_16 rbl0_27 rbl0_38 rbl0_49 rbl0_17
+ rbl0_28 rbl0_39 rbl1_60 rbl0_18 rbl0_29 rbl1_61 rbl1_50 rbl0_19 rbl1_40 rbl1_62
+ rbl1_51 rbl1_30 rbl1_41 rbl1_63 rbl1_52 rbl1_20 rbl1_31 rbl1_42 rbl1_64 rbl1_53
+ rbl1_0 rbl1_10 rbl1_21 rbl1_32 rbl1_43 rbl1_54 rbl1_1 rbl1_11 rbl1_22 rbl1_33 rbl1_44
+ rbl1_55 rbl1_2 rbl1_12 rbl1_23 rbl1_34 rbl1_45 rbl1_56 rbl1_3 rbl1_13 rbl1_24 rbl1_35
+ rbl1_46 rbl1_57 rbl1_4 rbl1_14 rbl1_25 rbl1_36 rbl1_47 rbl1_58 rbl1_5 rbl1_15 rbl1_26
+ rbl1_37 rbl1_48 rbl1_59 rbl1_6 rbl1_16 rbl1_27 rbl1_38 rbl1_49 rbl1_7 gnd rbl1_17
+ rbl1_28 rbl1_39 rbl1_8 rbl1_18 rbl1_29 rbl1_9 rbl1_19
Xprecharge_multiport_0_1 en_bar rbl1_63 gnd rbl0_63 vdd precharge_multiport_0
Xprecharge_multiport_0_2 en_bar rbl1_62 gnd rbl0_62 vdd precharge_multiport_0
Xprecharge_multiport_0_3 en_bar rbl1_61 gnd rbl0_61 vdd precharge_multiport_0
Xprecharge_multiport_0_4 en_bar rbl1_60 gnd rbl0_60 vdd precharge_multiport_0
Xprecharge_multiport_0_60 en_bar rbl1_4 gnd rbl0_4 vdd precharge_multiport_0
Xprecharge_multiport_0_5 en_bar rbl1_59 gnd rbl0_59 vdd precharge_multiport_0
Xprecharge_multiport_0_50 en_bar rbl1_14 gnd rbl0_14 vdd precharge_multiport_0
Xprecharge_multiport_0_61 en_bar rbl1_3 gnd rbl0_3 vdd precharge_multiport_0
Xprecharge_multiport_0_6 en_bar rbl1_58 gnd rbl0_58 vdd precharge_multiport_0
Xprecharge_multiport_0_7 en_bar rbl1_57 gnd rbl0_57 vdd precharge_multiport_0
Xprecharge_multiport_0_40 en_bar rbl1_24 gnd rbl0_24 vdd precharge_multiport_0
Xprecharge_multiport_0_51 en_bar rbl1_13 gnd rbl0_13 vdd precharge_multiport_0
Xprecharge_multiport_0_62 en_bar rbl1_2 gnd rbl0_2 vdd precharge_multiport_0
Xprecharge_multiport_0_8 en_bar rbl1_56 gnd rbl0_56 vdd precharge_multiport_0
Xprecharge_multiport_0_30 en_bar rbl1_34 gnd rbl0_34 vdd precharge_multiport_0
Xprecharge_multiport_0_41 en_bar rbl1_23 gnd rbl0_23 vdd precharge_multiport_0
Xprecharge_multiport_0_52 en_bar rbl1_12 gnd rbl0_12 vdd precharge_multiport_0
Xprecharge_multiport_0_63 en_bar rbl1_1 gnd rbl0_1 vdd precharge_multiport_0
Xprecharge_multiport_0_9 en_bar rbl1_55 gnd rbl0_55 vdd precharge_multiport_0
Xprecharge_multiport_0_20 en_bar rbl1_44 gnd rbl0_44 vdd precharge_multiport_0
Xprecharge_multiport_0_31 en_bar rbl1_33 gnd rbl0_33 vdd precharge_multiport_0
Xprecharge_multiport_0_42 en_bar rbl1_22 gnd rbl0_22 vdd precharge_multiport_0
Xprecharge_multiport_0_53 en_bar rbl1_11 gnd rbl0_11 vdd precharge_multiport_0
Xprecharge_multiport_0_64 en_bar rbl1_0 gnd rbl0_0 vdd precharge_multiport_0
Xprecharge_multiport_0_10 en_bar rbl1_54 gnd rbl0_54 vdd precharge_multiport_0
Xprecharge_multiport_0_21 en_bar rbl1_43 gnd rbl0_43 vdd precharge_multiport_0
Xprecharge_multiport_0_32 en_bar rbl1_32 gnd rbl0_32 vdd precharge_multiport_0
Xprecharge_multiport_0_43 en_bar rbl1_21 gnd rbl0_21 vdd precharge_multiport_0
Xprecharge_multiport_0_54 en_bar rbl1_10 gnd rbl0_10 vdd precharge_multiport_0
Xprecharge_multiport_0_11 en_bar rbl1_53 gnd rbl0_53 vdd precharge_multiport_0
Xprecharge_multiport_0_22 en_bar rbl1_42 gnd rbl0_42 vdd precharge_multiport_0
Xprecharge_multiport_0_33 en_bar rbl1_31 gnd rbl0_31 vdd precharge_multiport_0
Xprecharge_multiport_0_44 en_bar rbl1_20 gnd rbl0_20 vdd precharge_multiport_0
Xprecharge_multiport_0_55 en_bar rbl1_9 gnd rbl0_9 vdd precharge_multiport_0
Xprecharge_multiport_0_12 en_bar rbl1_52 gnd rbl0_52 vdd precharge_multiport_0
Xprecharge_multiport_0_13 en_bar rbl1_51 gnd rbl0_51 vdd precharge_multiport_0
Xprecharge_multiport_0_23 en_bar rbl1_41 gnd rbl0_41 vdd precharge_multiport_0
Xprecharge_multiport_0_24 en_bar rbl1_40 gnd rbl0_40 vdd precharge_multiport_0
Xprecharge_multiport_0_34 en_bar rbl1_30 gnd rbl0_30 vdd precharge_multiport_0
Xprecharge_multiport_0_35 en_bar rbl1_29 gnd rbl0_29 vdd precharge_multiport_0
Xprecharge_multiport_0_45 en_bar rbl1_19 gnd rbl0_19 vdd precharge_multiport_0
Xprecharge_multiport_0_46 en_bar rbl1_18 gnd rbl0_18 vdd precharge_multiport_0
Xprecharge_multiport_0_56 en_bar rbl1_8 gnd rbl0_8 vdd precharge_multiport_0
Xprecharge_multiport_0_57 en_bar rbl1_7 gnd rbl0_7 vdd precharge_multiport_0
Xprecharge_multiport_0_14 en_bar rbl1_50 gnd rbl0_50 vdd precharge_multiport_0
Xprecharge_multiport_0_25 en_bar rbl1_39 gnd rbl0_39 vdd precharge_multiport_0
Xprecharge_multiport_0_36 en_bar rbl1_28 gnd rbl0_28 vdd precharge_multiport_0
Xprecharge_multiport_0_47 en_bar rbl1_17 gnd rbl0_17 vdd precharge_multiport_0
Xprecharge_multiport_0_58 en_bar rbl1_6 gnd rbl0_6 vdd precharge_multiport_0
Xprecharge_multiport_0_15 en_bar rbl1_49 gnd rbl0_49 vdd precharge_multiport_0
Xprecharge_multiport_0_26 en_bar rbl1_38 gnd rbl0_38 vdd precharge_multiport_0
Xprecharge_multiport_0_37 en_bar rbl1_27 gnd rbl0_27 vdd precharge_multiport_0
Xprecharge_multiport_0_48 en_bar rbl1_16 gnd rbl0_16 vdd precharge_multiport_0
Xprecharge_multiport_0_59 en_bar rbl1_5 gnd rbl0_5 vdd precharge_multiport_0
Xprecharge_multiport_0_16 en_bar rbl1_48 gnd rbl0_48 vdd precharge_multiport_0
Xprecharge_multiport_0_27 en_bar rbl1_37 gnd rbl0_37 vdd precharge_multiport_0
Xprecharge_multiport_0_38 en_bar rbl1_26 gnd rbl0_26 vdd precharge_multiport_0
Xprecharge_multiport_0_49 en_bar rbl1_15 gnd rbl0_15 vdd precharge_multiport_0
Xprecharge_multiport_0_17 en_bar rbl1_47 gnd rbl0_47 vdd precharge_multiport_0
Xprecharge_multiport_0_28 en_bar rbl1_36 gnd rbl0_36 vdd precharge_multiport_0
Xprecharge_multiport_0_39 en_bar rbl1_25 gnd rbl0_25 vdd precharge_multiport_0
Xprecharge_multiport_0_18 en_bar rbl1_46 gnd rbl0_46 vdd precharge_multiport_0
Xprecharge_multiport_0_29 en_bar rbl1_35 gnd rbl0_35 vdd precharge_multiport_0
Xprecharge_multiport_0_19 en_bar rbl1_45 gnd rbl0_45 vdd precharge_multiport_0
Xprecharge_multiport_0_0 en_bar rbl1_64 gnd rbl0_64 vdd precharge_multiport_0
.ends

.subckt port_data din0_15 din0_26 dout1_19 din0_6 din0_16 din0_27 p_en_bar din0_7
+ dout1_30 din0_17 din0_28 gnd sel_1 din0_8 dout1_20 dout1_31 din0_18 din0_29 din0_9
+ vdd dout1_10 dout1_21 din0_19 dout1_11 dout1_22 dout1_12 dout1_23 dout1_13 dout1_24
+ w_en dout1_14 dout1_25 dout1_15 dout1_26 dout1_0 dout1_16 dout1_27 dout1_1 dout1_17
+ dout1_28 dout1_2 dout1_18 dout1_29 dout1_3 dout1_4 dout1_5 dout1_6 vdd_uq150 dout1_7
+ vdd_uq91 vdd_uq140 vdd_uq151 dout1_8 vdd_uq81 vdd_uq130 vdd_uq141 vdd_uq152 dout1_9
+ vdd_uq71 vdd_uq93 vdd_uq121 vdd_uq131 vdd_uq142 vdd_uq153 vdd_uq83 vdd_uq111 vdd_uq132
+ vdd_uq143 vdd_uq154 vdd_uq73 vdd_uq95 vdd_uq101 vdd_uq123 vdd_uq133 vdd_uq144 vdd_uq155
+ vdd_uq85 vdd_uq113 vdd_uq134 vdd_uq145 vdd_uq156 vdd_uq125 vdd_uq75 vdd_uq97 vdd_uq103
+ vdd_uq135 vdd_uq146 vdd_uq157 precharge_array_multiport_0/rbl1_64 vdd_uq65 vdd_uq87
+ vdd_uq115 vdd_uq136 vdd_uq147 vdd_uq158 vdd_uq77 vdd_uq99 vdd_uq105 vdd_uq127 vdd_uq137
+ vdd_uq148 vdd_uq159 din0_21 vdd_uq67 vdd_uq89 vdd_uq117 vdd_uq138 vdd_uq149 vdd_uq107
+ vdd_uq79 vdd_uq128 vdd_uq139 sel_0 vdd_uq69 vdd_uq119 vdd_uq129 vdd_uq109 din0_30
+ din0_20 din0_31 din0_0 din0_10 din0_1 din0_11 din0_22 din0_2 din0_12 din0_23 din0_3
+ din0_13 din0_24 din0_4 din0_14 din0_25 din0_5
Xsense_amp_array_0 vdd_uq65 vdd_uq67 dout1_30 dout1_31 dout1_20 vdd_uq69 dout1_10
+ dout1_21 dout1_11 dout1_22 vdd_uq71 dout1_12 dout1_23 dout1_13 dout1_24 dout1_14
+ dout1_25 vdd_uq73 dout1_15 dout1_26 dout1_27 dout1_16 vdd_uq75 dout1_28 dout1_17
+ dout1_29 dout1_18 dout1_19 gnd vdd_uq125 vdd_uq127 vdd_uq117 vdd_uq107 vdd_uq119
+ vdd_uq97 dout1_0 vdd_uq109 vdd_uq87 dout1_1 vdd_uq121 vdd_uq99 vdd_uq77 dout1_2
+ vdd_uq111 vdd_uq89 dout1_3 vdd_uq123 vdd_uq101 vdd_uq79 dout1_4 vdd_uq113 vdd_uq91
+ dout1_5 vdd_uq103 vdd_uq81 dout1_6 vdd_uq115 vdd_uq93 dout1_7 vdd_uq105 vdd_uq83
+ dout1_8 vdd_uq95 dout1_9 vdd_uq85 sense_amp_array
Xcolumn_mux_array_multiport_0 rbl0_0 rbl0_60 sel_1 rbl0_61 rbl0_50 rbl0_1 sel_0 rbl0_2
+ rbl0_40 rbl0_62 rbl0_51 rbl0_30 rbl0_41 rbl0_63 rbl0_52 rbl0_3 rbl0_4 rbl0_20 rbl0_31
+ rbl0_42 rbl0_53 rbl0_10 rbl0_21 rbl0_32 rbl0_43 rbl0_54 rbl0_5 rbl0_6 rbl0_11 rbl0_22
+ rbl0_33 rbl0_44 rbl0_55 rbl0_12 rbl0_23 rbl0_34 rbl0_45 rbl0_56 rbl0_7 rbl0_8 rbl0_13
+ rbl0_24 rbl0_35 rbl0_46 rbl0_57 rbl0_14 rbl0_25 rbl0_36 rbl0_47 rbl0_58 rbl0_9 rbl0_15
+ rbl0_26 rbl0_37 rbl0_59 rbl0_48 rbl0_16 rbl0_27 rbl0_38 rbl0_49 rbl0_17 rbl0_28
+ rbl0_39 rbl1_60 rbl0_18 rbl0_29 rbl1_61 rbl1_50 rbl0_19 rbl1_40 rbl1_62 rbl1_51
+ rbl1_30 rbl1_41 rbl1_63 rbl1_52 rbl1_20 rbl1_31 rbl1_42 rbl1_53 rbl1_0 rbl1_10 rbl1_21
+ rbl1_32 rbl1_43 rbl1_54 rbl1_1 rbl1_11 rbl1_22 rbl1_33 rbl1_44 rbl1_55 rbl1_2 gnd
+ rbl1_12 rbl1_23 rbl1_34 rbl1_45 rbl1_56 rbl1_3 rbl1_13 rbl1_24 rbl1_35 rbl1_46 rbl1_57
+ rbl1_4 rbl1_14 rbl1_25 rbl1_36 rbl1_47 rbl1_58 rbl1_5 rbl1_15 rbl1_26 rbl1_37 rbl1_59
+ rbl1_48 rbl1_6 rbl1_16 rbl1_27 rbl1_38 rbl1_49 rbl1_7 rbl1_17 rbl1_28 rbl1_39 rbl1_8
+ rbl1_18 rbl1_29 rbl1_9 rbl1_19 column_mux_array_multiport
Xwrite_driver_array_0 din0_7 din0_8 vdd_uq128 din0_9 vdd_uq130 w_en vdd_uq131 vdd_uq132
+ vdd_uq133 vdd_uq134 vdd_uq135 vdd_uq136 vdd_uq137 vdd_uq138 wbl0_0 wbl0_1 din0_30
+ gnd din0_31 din0_20 din0_21 din0_10 din0_22 din0_11 din0_23 din0_12 vdd_uq159 din0_24
+ din0_13 din0_25 din0_14 vdd_uq149 vdd_uq150 vdd_uq139 din0_26 din0_15 din0_27 din0_16
+ vdd_uq151 vdd_uq140 vdd_uq152 vdd_uq141 din0_28 din0_17 din0_29 din0_18 vdd_uq153
+ vdd_uq142 vdd_uq129 vdd_uq154 vdd_uq143 din0_19 din0_0 vdd_uq155 vdd_uq144 din0_1
+ vdd_uq145 vdd_uq156 din0_2 vdd_uq157 vdd_uq146 din0_3 vdd_uq158 vdd_uq147 din0_4
+ vdd_uq148 din0_5 din0_6 write_driver_array
Xprecharge_array_multiport_0 rbl0_0 rbl0_60 p_en_bar rbl0_61 rbl0_50 rbl0_1 vdd rbl0_2
+ rbl0_40 rbl0_62 rbl0_51 rbl0_30 rbl0_41 rbl0_63 rbl0_52 rbl0_3 rbl0_4 rbl0_20 rbl0_31
+ rbl0_42 rbl0_53 rbl0_10 rbl0_21 rbl0_32 rbl0_43 rbl0_54 rbl0_5 rbl0_6 rbl0_11 rbl0_22
+ rbl0_33 rbl0_44 rbl0_55 rbl0_12 rbl0_23 rbl0_34 rbl0_45 rbl0_56 rbl0_7 rbl0_8 rbl0_13
+ rbl0_24 rbl0_35 rbl0_46 rbl0_57 rbl0_14 rbl0_25 rbl0_36 rbl0_47 rbl0_58 rbl0_9 rbl0_15
+ rbl0_26 rbl0_37 rbl0_48 rbl0_59 rbl0_16 rbl0_27 rbl0_38 rbl0_49 rbl0_17 rbl0_28
+ rbl0_39 rbl1_60 rbl0_18 rbl0_29 rbl1_61 rbl1_50 rbl0_19 rbl1_40 rbl1_62 rbl1_51
+ rbl1_30 rbl1_41 rbl1_63 rbl1_52 rbl1_20 rbl1_31 rbl1_42 precharge_array_multiport_0/rbl1_64
+ rbl1_53 rbl1_0 rbl1_10 rbl1_21 rbl1_32 rbl1_43 rbl1_54 rbl1_1 rbl1_11 rbl1_22 rbl1_33
+ rbl1_44 rbl1_55 rbl1_2 rbl1_12 rbl1_23 rbl1_34 rbl1_45 rbl1_56 rbl1_3 rbl1_13 rbl1_24
+ rbl1_35 rbl1_46 rbl1_57 rbl1_4 rbl1_14 rbl1_25 rbl1_36 rbl1_47 rbl1_58 rbl1_5 rbl1_15
+ rbl1_26 rbl1_37 rbl1_48 rbl1_59 rbl1_6 rbl1_16 rbl1_27 rbl1_38 rbl1_49 rbl1_7 gnd
+ rbl1_17 rbl1_28 rbl1_39 rbl1_8 rbl1_18 rbl1_29 rbl1_9 rbl1_19 precharge_array_multiport
.ends

.subckt pinvbuf pinv_2_0/A Zb Z gnd vdd A
Xpinv_1_0 pinv_2_1/A gnd vdd pinv_2_0/A pinv_1
Xpinv_2_0 Z gnd vdd pinv_2_0/A pinv_2
Xpinv_2_1 Zb gnd vdd pinv_2_1/A pinv_2
Xpinv_0_0 A pinv_2_0/A gnd vdd pinv_0
.ends

.subckt pinv Z A gnd vdd
Xnmos_m1_w0_420_sli_dli_da_p_0 gnd gnd Z A nmos_m1_w0_420_sli_dli_da_p
Xpmos_m1_w1_260_sli_dli_da_p_0 vdd vdd gnd Z A pmos_m1_w1_260_sli_dli_da_p
.ends

.subckt pnand2 Z gnd vdd A B
Xpmos_m1_w1_260_sli_dli_0 vdd Z gnd vdd B pmos_m1_w1_260_sli_dli
Xpmos_m1_w1_260_sli_dli_1 vdd vdd gnd Z A pmos_m1_w1_260_sli_dli
Xnmos_m1_w0_840_sli_dactive_0 gnd gnd A nmos_m1_w0_840_sactive_dli_0/a_0_0# nmos_m1_w0_840_sli_dactive
Xnmos_m1_w0_840_sactive_dli_0 nmos_m1_w0_840_sactive_dli_0/a_0_0# gnd Z B nmos_m1_w0_840_sactive_dli
.ends

.subckt and2_dec Z gnd vdd A B
Xpinv_0 Z pinv_0/A gnd vdd pinv
Xpnand2_0 pinv_0/A gnd vdd A B pnand2
.ends

.subckt hierarchical_predecode2x4 in_1 vdd_uq0 out_0 out_1 out_2 out_3 in_0 gnd vdd
Xand2_dec_0 out_3 gnd vdd in_0 in_1 and2_dec
Xand2_dec_1 out_2 gnd vdd pinv_1/Z in_1 and2_dec
Xpinv_0 pinv_0/Z in_1 gnd vdd_uq0 pinv
Xand2_dec_2 out_1 gnd vdd_uq0 in_0 pinv_0/Z and2_dec
Xpinv_1 pinv_1/Z in_0 gnd vdd_uq0 pinv
Xand2_dec_3 out_0 gnd vdd_uq0 pinv_1/Z pinv_0/Z and2_dec
.ends

.subckt dec_cell3_2r1w A0 B0 C0 A1 B1 C1 A2 B2 C2 OUT2 vdd gnd OUT0 OUT1
X0 vdd A2 net9 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_124_132# A0 net3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 net6 A1 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 OUT2 net9 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.35e+06u l=150000u
X4 OUT2 net9 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 vdd C0 net3 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 net6 C1 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 vdd C2 net9 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 OUT0 net6 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.35e+06u l=150000u
X9 a_220_132# B0 a_124_132# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_412_132# A1 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 gnd net3 OUT1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 OUT0 net6 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 gnd C0 a_220_132# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_508_132# B1 a_412_132# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 net6 C1 a_508_132# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 vdd B1 net6 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 vdd A0 net3 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 net9 B2 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 vdd net3 OUT1 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.35e+06u l=150000u
X20 a_808_132# A2 net9 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 a_904_132# B2 a_808_132# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 gnd C2 a_904_132# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 net3 B0 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt pnand3 Z gnd vdd A B C
Xpmos_m1_w1_260_sli_dli_0 vdd vdd gnd Z C pmos_m1_w1_260_sli_dli
Xpmos_m1_w1_260_sli_dli_1 vdd Z gnd vdd B pmos_m1_w1_260_sli_dli
Xpmos_m1_w1_260_sli_dli_2 vdd vdd gnd Z A pmos_m1_w1_260_sli_dli
Xnmos_m1_w0_840_sli_dactive_0 gnd gnd A a_154_51# nmos_m1_w0_840_sli_dactive
Xnmos_m1_w0_840_sactive_dli_0 a_244_51# gnd Z C nmos_m1_w0_840_sactive_dli
X0 a_244_51# B a_154_51# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
.ends

.subckt and3_dec Z gnd vdd A B C
Xpinv_0 Z pinv_0/A gnd vdd pinv
Xpnand3_0 pinv_0/A gnd vdd A B C pnand3
.ends

.subckt hierarchical_predecode3x8 vdd_uq0 vdd_uq1 vdd_uq2 out_5 out_0 out_1 out_2
+ out_3 out_4 out_7 out_6 in_0 gnd in_1 in_2 vdd
Xand3_dec_1 out_6 gnd vdd_uq2 pinv_2/Z in_1 in_2 and3_dec
Xand3_dec_2 out_5 gnd vdd_uq1 in_0 pinv_1/Z in_2 and3_dec
Xpinv_0 pinv_0/Z in_2 gnd vdd pinv
Xand3_dec_3 out_4 gnd vdd_uq1 pinv_2/Z pinv_1/Z in_2 and3_dec
Xpinv_1 pinv_1/Z in_1 gnd vdd_uq0 pinv
Xand3_dec_4 out_3 gnd vdd in_0 in_1 pinv_0/Z and3_dec
Xpinv_2 pinv_2/Z in_0 gnd vdd_uq0 pinv
Xand3_dec_5 out_2 gnd vdd pinv_2/Z in_1 pinv_0/Z and3_dec
Xand3_dec_6 out_1 gnd vdd_uq0 in_0 pinv_1/Z pinv_0/Z and3_dec
Xand3_dec_7 out_0 gnd vdd_uq0 pinv_2/Z pinv_1/Z pinv_0/Z and3_dec
Xand3_dec_0 out_7 gnd vdd_uq2 in_0 in_1 in_2 and3_dec
.ends

.subckt hierarchical_decoder addr_0 decode0_6 decode2_9 addr_2 decode1_54 decode1_43
+ decode1_32 decode1_21 decode1_10 addr_1 gnd addr_3 decode1_55 decode1_44 decode1_33
+ decode1_22 decode1_11 decode0_7 addr_4 decode1_56 decode1_45 decode1_34 decode1_23
+ decode1_12 vdd_uq2 decode0_8 decode1_57 decode1_46 decode1_35 decode1_24 decode1_13
+ decode0_9 decode1_58 decode1_47 decode1_36 decode1_25 decode1_14 vdd_uq4 addr_5
+ decode1_59 decode1_48 decode1_37 decode1_26 decode1_15 addr_6 decode1_49 decode1_38
+ decode1_27 decode1_16 vdd_uq6 addr_7 decode2_60 decode1_39 decode1_28 decode1_17
+ decode1_29 decode1_18 decode2_61 decode2_50 vdd_uq8 decode2_62 decode2_51 decode2_40
+ decode1_19 decode2_63 decode2_52 decode2_41 decode2_30 vdd_uq9 decode1_0 decode2_53
+ decode2_42 decode2_31 decode2_20 decode1_1 decode2_54 decode2_43 decode2_32 decode2_21
+ decode2_10 decode1_2 decode2_55 decode2_44 decode2_33 decode2_22 decode2_11 decode1_3
+ decode2_56 decode2_45 decode2_34 decode2_23 decode2_12 decode1_4 decode2_57 decode2_46
+ decode2_35 decode2_24 decode2_13 decode1_5 decode2_58 decode2_47 decode2_36 decode2_25
+ decode2_14 decode1_6 decode2_59 decode2_48 decode2_37 decode2_26 decode2_15 decode1_7
+ decode2_49 decode2_38 decode2_27 decode2_16 decode1_8 decode0_60 decode2_39 decode2_28
+ decode2_17 decode1_9 decode0_61 decode0_50 vdd_uq50 decode2_29 decode2_18 decode0_62
+ decode0_51 decode0_40 decode2_19 vdd_uq40 decode0_63 decode0_52 decode0_41 decode0_30
+ vdd_uq41 vdd_uq30 decode0_53 decode0_42 decode0_31 decode0_20 vdd_uq42 vdd_uq31
+ vdd_uq20 decode0_54 decode0_43 decode0_32 decode0_21 decode0_10 vdd_uq43 vdd_uq32
+ vdd_uq21 decode0_55 decode0_44 decode0_33 decode0_22 decode0_11 vdd_uq44 vdd_uq33
+ vdd_uq12 vdd_uq22 decode0_56 decode0_45 decode0_34 decode0_23 decode0_12 vdd_uq45
+ vdd_uq34 vdd_uq23 decode0_57 decode0_46 decode0_35 decode0_24 decode0_13 decode2_0
+ vdd_uq46 vdd_uq35 vdd_uq14 vdd_uq24 decode0_58 decode0_47 decode0_36 decode0_25
+ decode0_14 vdd decode2_1 vdd_uq47 vdd_uq36 vdd_uq25 decode0_59 decode0_48 decode0_37
+ decode0_26 decode0_15 decode2_2 vdd_uq48 vdd_uq37 vdd_uq26 vdd_uq16 decode0_27 decode0_16
+ decode0_49 decode0_38 decode0_0 decode2_3 vdd_uq49 vdd_uq38 vdd_uq27 decode0_39
+ decode0_28 decode0_17 decode2_4 decode1_60 decode0_1 vdd_uq39 vdd_uq28 vdd_uq18
+ decode1_61 decode1_50 decode0_29 decode0_18 decode0_2 decode2_5 vdd_uq29 decode0_19
+ decode2_6 decode1_62 decode1_51 decode1_40 decode0_3 vdd_uq19 decode0_4 decode2_7
+ decode1_63 decode1_52 decode1_41 decode1_30 decode2_8 decode1_53 decode1_42 decode1_31
+ decode1_20 decode0_5
Xhierarchical_predecode2x4_0 addr_1 vdd predecode_0 predecode_1 predecode_2 predecode_3
+ addr_0 gnd vdd_uq2 hierarchical_predecode2x4
Xdec_cell3_2r1w_60 predecode_0 predecode_6 predecode_12 predecode_1 predecode_6 predecode_12
+ predecode_2 predecode_6 predecode_12 decode2_3 vdd_uq20 gnd decode0_3 decode1_3
+ dec_cell3_2r1w
Xdec_cell3_2r1w_61 predecode_1 predecode_5 predecode_12 predecode_2 predecode_5 predecode_12
+ predecode_3 predecode_5 predecode_12 decode2_2 vdd_uq20 gnd decode0_2 decode1_2
+ dec_cell3_2r1w
Xdec_cell3_2r1w_50 predecode_2 predecode_5 predecode_13 predecode_3 predecode_5 predecode_13
+ predecode_0 predecode_6 predecode_13 decode2_13 vdd_uq25 gnd decode0_13 decode1_13
+ dec_cell3_2r1w
Xdec_cell3_2r1w_40 predecode_0 predecode_5 predecode_14 predecode_1 predecode_5 predecode_14
+ predecode_2 predecode_5 predecode_14 decode2_23 vdd_uq30 gnd decode0_23 decode1_23
+ dec_cell3_2r1w
Xdec_cell3_2r1w_62 predecode_2 predecode_4 predecode_12 predecode_3 predecode_4 predecode_12
+ predecode_0 predecode_5 predecode_12 decode2_1 vdd_uq19 gnd decode0_1 decode1_1
+ dec_cell3_2r1w
Xdec_cell3_2r1w_51 predecode_3 predecode_4 predecode_13 predecode_0 predecode_5 predecode_13
+ predecode_1 predecode_5 predecode_13 decode2_12 vdd_uq25 gnd decode0_12 decode1_12
+ dec_cell3_2r1w
Xdec_cell3_2r1w_30 predecode_2 predecode_4 predecode_15 predecode_3 predecode_4 predecode_15
+ predecode_0 predecode_5 predecode_15 decode2_33 vdd_uq35 gnd decode0_33 decode1_33
+ dec_cell3_2r1w
Xdec_cell3_2r1w_41 predecode_1 predecode_4 predecode_14 predecode_2 predecode_4 predecode_14
+ predecode_3 predecode_4 predecode_14 decode2_22 vdd_uq30 gnd decode0_22 decode1_22
+ dec_cell3_2r1w
Xdec_cell3_2r1w_63 dec_cell3_2r1w_63/A0 dec_cell3_2r1w_63/B0 dec_cell3_2r1w_63/C0
+ predecode_0 predecode_4 predecode_12 predecode_1 predecode_4 predecode_12 decode2_0
+ vdd_uq19 gnd decode0_0 decode1_0 dec_cell3_2r1w
Xdec_cell3_2r1w_52 predecode_0 predecode_4 predecode_13 predecode_1 predecode_4 predecode_13
+ predecode_2 predecode_4 predecode_13 decode2_11 vdd_uq24 gnd decode0_11 decode1_11
+ dec_cell3_2r1w
Xdec_cell3_2r1w_0 predecode_0 predecode_11 predecode_17 predecode_1 predecode_11 predecode_17
+ predecode_2 predecode_11 predecode_17 decode2_63 vdd_uq50 gnd decode0_63 decode1_63
+ dec_cell3_2r1w
Xdec_cell3_2r1w_20 predecode_0 predecode_4 predecode_16 predecode_1 predecode_4 predecode_16
+ predecode_2 predecode_4 predecode_16 decode2_43 vdd_uq40 gnd decode0_43 decode1_43
+ dec_cell3_2r1w
Xdec_cell3_2r1w_31 predecode_3 predecode_11 predecode_14 predecode_0 predecode_4 predecode_15
+ predecode_1 predecode_4 predecode_15 decode2_32 vdd_uq35 gnd decode0_32 decode1_32
+ dec_cell3_2r1w
Xdec_cell3_2r1w_53 predecode_1 predecode_11 predecode_12 predecode_2 predecode_11
+ predecode_12 predecode_3 predecode_11 predecode_12 decode2_10 vdd_uq24 gnd decode0_10
+ decode1_10 dec_cell3_2r1w
Xdec_cell3_2r1w_42 predecode_2 predecode_11 predecode_13 predecode_3 predecode_11
+ predecode_13 predecode_0 predecode_4 predecode_14 decode2_21 vdd_uq29 gnd decode0_21
+ decode1_21 dec_cell3_2r1w
Xdec_cell3_2r1w_1 predecode_1 predecode_10 predecode_17 predecode_2 predecode_10 predecode_17
+ predecode_3 predecode_10 predecode_17 decode2_62 vdd_uq50 gnd decode0_62 decode1_62
+ dec_cell3_2r1w
Xdec_cell3_2r1w_10 predecode_2 predecode_11 predecode_16 predecode_3 predecode_11
+ predecode_16 predecode_0 predecode_4 predecode_17 decode2_53 vdd_uq45 gnd decode0_53
+ decode1_53 dec_cell3_2r1w
Xdec_cell3_2r1w_21 predecode_1 predecode_11 predecode_15 predecode_2 predecode_11
+ predecode_15 predecode_3 predecode_11 predecode_15 decode2_42 vdd_uq40 gnd decode0_42
+ decode1_42 dec_cell3_2r1w
Xdec_cell3_2r1w_32 predecode_0 predecode_11 predecode_14 predecode_1 predecode_11
+ predecode_14 predecode_2 predecode_11 predecode_14 decode2_31 vdd_uq34 gnd decode0_31
+ decode1_31 dec_cell3_2r1w
Xdec_cell3_2r1w_54 predecode_2 predecode_10 predecode_12 predecode_3 predecode_10
+ predecode_12 predecode_0 predecode_11 predecode_12 decode2_9 vdd_uq23 gnd decode0_9
+ decode1_9 dec_cell3_2r1w
Xdec_cell3_2r1w_43 predecode_3 predecode_10 predecode_13 predecode_0 predecode_11
+ predecode_13 predecode_1 predecode_11 predecode_13 decode2_20 vdd_uq29 gnd decode0_20
+ decode1_20 dec_cell3_2r1w
Xdec_cell3_2r1w_2 predecode_2 predecode_9 predecode_17 predecode_3 predecode_9 predecode_17
+ predecode_0 predecode_10 predecode_17 decode2_61 vdd_uq49 gnd decode0_61 decode1_61
+ dec_cell3_2r1w
Xdec_cell3_2r1w_11 predecode_3 predecode_10 predecode_16 predecode_0 predecode_11
+ predecode_16 predecode_1 predecode_11 predecode_16 decode2_52 vdd_uq45 gnd decode0_52
+ decode1_52 dec_cell3_2r1w
Xdec_cell3_2r1w_22 predecode_2 predecode_10 predecode_15 predecode_3 predecode_10
+ predecode_15 predecode_0 predecode_11 predecode_15 decode2_41 vdd_uq39 gnd decode0_41
+ decode1_41 dec_cell3_2r1w
Xdec_cell3_2r1w_33 predecode_1 predecode_10 predecode_14 predecode_2 predecode_10
+ predecode_14 predecode_3 predecode_10 predecode_14 decode2_30 vdd_uq34 gnd decode0_30
+ decode1_30 dec_cell3_2r1w
Xdec_cell3_2r1w_55 predecode_3 predecode_9 predecode_12 predecode_0 predecode_10 predecode_12
+ predecode_1 predecode_10 predecode_12 decode2_8 vdd_uq23 gnd decode0_8 decode1_8
+ dec_cell3_2r1w
Xdec_cell3_2r1w_44 predecode_0 predecode_10 predecode_13 predecode_1 predecode_10
+ predecode_13 predecode_2 predecode_10 predecode_13 decode2_19 vdd_uq28 gnd decode0_19
+ decode1_19 dec_cell3_2r1w
Xdec_cell3_2r1w_3 predecode_3 predecode_8 predecode_17 predecode_0 predecode_9 predecode_17
+ predecode_1 predecode_9 predecode_17 decode2_60 vdd_uq49 gnd decode0_60 decode1_60
+ dec_cell3_2r1w
Xdec_cell3_2r1w_12 predecode_0 predecode_10 predecode_16 predecode_1 predecode_10
+ predecode_16 predecode_2 predecode_10 predecode_16 decode2_51 vdd_uq44 gnd decode0_51
+ decode1_51 dec_cell3_2r1w
Xdec_cell3_2r1w_23 predecode_3 predecode_9 predecode_15 predecode_0 predecode_10 predecode_15
+ predecode_1 predecode_10 predecode_15 decode2_40 vdd_uq39 gnd decode0_40 decode1_40
+ dec_cell3_2r1w
Xdec_cell3_2r1w_34 predecode_2 predecode_9 predecode_14 predecode_3 predecode_9 predecode_14
+ predecode_0 predecode_10 predecode_14 decode2_29 vdd_uq33 gnd decode0_29 decode1_29
+ dec_cell3_2r1w
Xdec_cell3_2r1w_56 predecode_0 predecode_9 predecode_12 predecode_1 predecode_9 predecode_12
+ predecode_2 predecode_9 predecode_12 decode2_7 vdd_uq22 gnd decode0_7 decode1_7
+ dec_cell3_2r1w
Xdec_cell3_2r1w_45 predecode_1 predecode_9 predecode_13 predecode_2 predecode_9 predecode_13
+ predecode_3 predecode_9 predecode_13 decode2_18 vdd_uq28 gnd decode0_18 decode1_18
+ dec_cell3_2r1w
Xdec_cell3_2r1w_4 predecode_0 predecode_8 predecode_17 predecode_1 predecode_8 predecode_17
+ predecode_2 predecode_8 predecode_17 decode2_59 vdd_uq48 gnd decode0_59 decode1_59
+ dec_cell3_2r1w
Xdec_cell3_2r1w_13 predecode_1 predecode_9 predecode_16 predecode_2 predecode_9 predecode_16
+ predecode_3 predecode_9 predecode_16 decode2_50 vdd_uq44 gnd decode0_50 decode1_50
+ dec_cell3_2r1w
Xdec_cell3_2r1w_24 predecode_0 predecode_9 predecode_15 predecode_1 predecode_9 predecode_15
+ predecode_2 predecode_9 predecode_15 decode2_39 vdd_uq38 gnd decode0_39 decode1_39
+ dec_cell3_2r1w
Xdec_cell3_2r1w_35 predecode_3 predecode_8 predecode_14 predecode_0 predecode_9 predecode_14
+ predecode_1 predecode_9 predecode_14 decode2_28 vdd_uq33 gnd decode0_28 decode1_28
+ dec_cell3_2r1w
Xdec_cell3_2r1w_57 predecode_1 predecode_8 predecode_12 predecode_2 predecode_8 predecode_12
+ predecode_3 predecode_8 predecode_12 decode2_6 vdd_uq22 gnd decode0_6 decode1_6
+ dec_cell3_2r1w
Xdec_cell3_2r1w_46 predecode_2 predecode_8 predecode_13 predecode_3 predecode_8 predecode_13
+ predecode_0 predecode_9 predecode_13 decode2_17 vdd_uq27 gnd decode0_17 decode1_17
+ dec_cell3_2r1w
Xdec_cell3_2r1w_5 predecode_1 predecode_7 predecode_17 predecode_2 predecode_7 predecode_17
+ predecode_3 predecode_7 predecode_17 decode2_58 vdd_uq48 gnd decode0_58 decode1_58
+ dec_cell3_2r1w
Xdec_cell3_2r1w_14 predecode_2 predecode_8 predecode_16 predecode_3 predecode_8 predecode_16
+ predecode_0 predecode_9 predecode_16 decode2_49 vdd_uq43 gnd decode0_49 decode1_49
+ dec_cell3_2r1w
Xdec_cell3_2r1w_25 predecode_1 predecode_8 predecode_15 predecode_2 predecode_8 predecode_15
+ predecode_3 predecode_8 predecode_15 decode2_38 vdd_uq38 gnd decode0_38 decode1_38
+ dec_cell3_2r1w
Xdec_cell3_2r1w_36 predecode_0 predecode_8 predecode_14 predecode_1 predecode_8 predecode_14
+ predecode_2 predecode_8 predecode_14 decode2_27 vdd_uq32 gnd decode0_27 decode1_27
+ dec_cell3_2r1w
Xdec_cell3_2r1w_58 predecode_2 predecode_7 predecode_12 predecode_3 predecode_7 predecode_12
+ predecode_0 predecode_8 predecode_12 decode2_5 vdd_uq21 gnd decode0_5 decode1_5
+ dec_cell3_2r1w
Xdec_cell3_2r1w_47 predecode_3 predecode_7 predecode_13 predecode_0 predecode_8 predecode_13
+ predecode_1 predecode_8 predecode_13 decode2_16 vdd_uq27 gnd decode0_16 decode1_16
+ dec_cell3_2r1w
Xdec_cell3_2r1w_6 predecode_2 predecode_6 predecode_17 predecode_3 predecode_6 predecode_17
+ predecode_0 predecode_7 predecode_17 decode2_57 vdd_uq47 gnd decode0_57 decode1_57
+ dec_cell3_2r1w
Xdec_cell3_2r1w_15 predecode_3 predecode_7 predecode_16 predecode_0 predecode_8 predecode_16
+ predecode_1 predecode_8 predecode_16 decode2_48 vdd_uq43 gnd decode0_48 decode1_48
+ dec_cell3_2r1w
Xdec_cell3_2r1w_26 predecode_2 predecode_7 predecode_15 predecode_3 predecode_7 predecode_15
+ predecode_0 predecode_8 predecode_15 decode2_37 vdd_uq37 gnd decode0_37 decode1_37
+ dec_cell3_2r1w
Xdec_cell3_2r1w_37 predecode_1 predecode_7 predecode_14 predecode_2 predecode_7 predecode_14
+ predecode_3 predecode_7 predecode_14 decode2_26 vdd_uq32 gnd decode0_26 decode1_26
+ dec_cell3_2r1w
Xdec_cell3_2r1w_59 predecode_3 predecode_6 predecode_12 predecode_0 predecode_7 predecode_12
+ predecode_1 predecode_7 predecode_12 decode2_4 vdd_uq21 gnd decode0_4 decode1_4
+ dec_cell3_2r1w
Xdec_cell3_2r1w_48 predecode_0 predecode_7 predecode_13 predecode_1 predecode_7 predecode_13
+ predecode_2 predecode_7 predecode_13 decode2_15 vdd_uq26 gnd decode0_15 decode1_15
+ dec_cell3_2r1w
Xdec_cell3_2r1w_7 predecode_3 predecode_5 predecode_17 predecode_0 predecode_6 predecode_17
+ predecode_1 predecode_6 predecode_17 decode2_56 vdd_uq47 gnd decode0_56 decode1_56
+ dec_cell3_2r1w
Xhierarchical_predecode3x8_0 vdd_uq12 vdd_uq16 vdd_uq18 predecode_17 predecode_12
+ predecode_13 predecode_14 predecode_15 predecode_16 predecode_19 predecode_18 addr_5
+ gnd addr_6 addr_7 vdd_uq14 hierarchical_predecode3x8
Xdec_cell3_2r1w_16 predecode_0 predecode_7 predecode_16 predecode_1 predecode_7 predecode_16
+ predecode_2 predecode_7 predecode_16 decode2_47 vdd_uq42 gnd decode0_47 decode1_47
+ dec_cell3_2r1w
Xdec_cell3_2r1w_27 predecode_3 predecode_6 predecode_15 predecode_0 predecode_7 predecode_15
+ predecode_1 predecode_7 predecode_15 decode2_36 vdd_uq37 gnd decode0_36 decode1_36
+ dec_cell3_2r1w
Xdec_cell3_2r1w_38 predecode_2 predecode_6 predecode_14 predecode_3 predecode_6 predecode_14
+ predecode_0 predecode_7 predecode_14 decode2_25 vdd_uq31 gnd decode0_25 decode1_25
+ dec_cell3_2r1w
Xdec_cell3_2r1w_49 predecode_1 predecode_6 predecode_13 predecode_2 predecode_6 predecode_13
+ predecode_3 predecode_6 predecode_13 decode2_14 vdd_uq26 gnd decode0_14 decode1_14
+ dec_cell3_2r1w
Xdec_cell3_2r1w_8 predecode_0 predecode_5 predecode_17 predecode_1 predecode_5 predecode_17
+ predecode_2 predecode_5 predecode_17 decode2_55 vdd_uq46 gnd decode0_55 decode1_55
+ dec_cell3_2r1w
Xhierarchical_predecode3x8_1 vdd_uq4 vdd_uq8 vdd_uq9 predecode_9 predecode_4 predecode_5
+ predecode_6 predecode_7 predecode_8 predecode_11 predecode_10 addr_2 gnd addr_3
+ addr_4 vdd_uq6 hierarchical_predecode3x8
Xdec_cell3_2r1w_17 predecode_1 predecode_6 predecode_16 predecode_2 predecode_6 predecode_16
+ predecode_3 predecode_6 predecode_16 decode2_46 vdd_uq42 gnd decode0_46 decode1_46
+ dec_cell3_2r1w
Xdec_cell3_2r1w_28 predecode_0 predecode_6 predecode_15 predecode_1 predecode_6 predecode_15
+ predecode_2 predecode_6 predecode_15 decode2_35 vdd_uq36 gnd decode0_35 decode1_35
+ dec_cell3_2r1w
Xdec_cell3_2r1w_39 predecode_3 predecode_5 predecode_14 predecode_0 predecode_6 predecode_14
+ predecode_1 predecode_6 predecode_14 decode2_24 vdd_uq31 gnd decode0_24 decode1_24
+ dec_cell3_2r1w
Xdec_cell3_2r1w_9 predecode_1 predecode_4 predecode_17 predecode_2 predecode_4 predecode_17
+ predecode_3 predecode_4 predecode_17 decode2_54 vdd_uq46 gnd decode0_54 decode1_54
+ dec_cell3_2r1w
Xdec_cell3_2r1w_18 predecode_2 predecode_5 predecode_16 predecode_3 predecode_5 predecode_16
+ predecode_0 predecode_6 predecode_16 decode2_45 vdd_uq41 gnd decode0_45 decode1_45
+ dec_cell3_2r1w
Xdec_cell3_2r1w_29 predecode_1 predecode_5 predecode_15 predecode_2 predecode_5 predecode_15
+ predecode_3 predecode_5 predecode_15 decode2_34 vdd_uq36 gnd decode0_34 decode1_34
+ dec_cell3_2r1w
Xdec_cell3_2r1w_19 predecode_3 predecode_4 predecode_16 predecode_0 predecode_5 predecode_16
+ predecode_1 predecode_5 predecode_16 decode2_44 vdd_uq41 gnd decode0_44 decode1_44
+ dec_cell3_2r1w
.ends

.subckt wordline_driver_cell A0 vdd gnd wl_en A1 A2 rwl0 wwl0 rwl1
X0 gnd wl_en a_124_308# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X1 net4 wl_en a_316_308# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X2 a_316_308# A1 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X3 vdd wl_en net4 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 vdd net4 rwl0 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.35e+06u l=150000u
X5 a_616_308# A2 net6 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X6 gnd wl_en a_616_308# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X7 wwl0 net6 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 net4 A1 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 vdd wl_en net6 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_124_308# A0 net2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X11 net6 A2 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 wwl0 net6 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.35e+06u l=150000u
X13 gnd net4 rwl0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 net2 A0 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 rwl1 net2 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 vdd wl_en net2 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 rwl1 net2 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.35e+06u l=150000u
.ends

.subckt wordline_driver_array wl_en in1_19 rwl1_0 wwl0_0 in2_62 in2_51 in2_40 rwl1_55
+ rwl1_11 rwl1_22 rwl1_33 rwl1_44 rwl1_1 in2_63 in2_52 wwl0_1 in2_30 in2_41 vdd_uq0
+ rwl1_56 rwl1_12 rwl1_23 rwl1_34 rwl1_45 rwl1_2 wwl0_2 in2_53 vdd_uq1 in2_20 in2_31
+ in2_42 rwl1_13 rwl1_24 rwl1_57 rwl1_46 rwl1_35 rwl1_3 wwl0_3 in2_54 in2_10 in2_21
+ in2_32 in2_43 vdd_uq2 rwl1_58 rwl1_47 rwl1_14 rwl1_25 rwl1_36 wwl0_4 rwl1_4 in2_55
+ in2_11 in2_22 in2_33 in2_44 vdd_uq3 rwl1_59 rwl1_48 rwl1_15 rwl1_26 rwl1_37 rwl1_5
+ wwl0_5 in2_56 in2_45 in2_12 in2_23 in2_34 vdd_uq4 rwl1_49 rwl1_16 rwl1_27 rwl1_38
+ in1_0 rwl1_6 in2_57 in2_46 wwl0_6 in2_13 in2_24 in2_35 vdd_uq5 rwl1_17 rwl1_28 rwl1_39
+ in1_1 rwl1_7 wwl0_7 in2_14 in2_58 in2_47 vdd_uq6 in2_25 in2_36 rwl1_18 rwl1_29 in1_2
+ rwl1_8 wwl0_8 in2_59 in2_48 in2_15 in2_26 in2_37 vdd_uq7 in1_3 rwl1_19 rwl1_9 wwl0_9
+ in2_49 in2_16 in2_27 in2_38 vdd_uq8 in1_4 in0_60 in2_17 in2_28 in2_39 vdd_uq9 in1_5
+ in0_61 in0_50 in2_18 in2_29 in1_6 in0_51 in0_40 in0_62 wwl0_60 in2_19 in1_7 in0_63
+ in0_52 in0_30 in0_41 wwl0_61 wwl0_50 in1_8 in0_53 in0_20 in0_31 in0_42 wwl0_62 wwl0_51
+ wwl0_40 in1_9 in0_54 in0_10 in0_21 in0_32 in0_43 wwl0_63 wwl0_52 wwl0_30 wwl0_41
+ in0_55 in0_11 in0_22 in0_33 in0_44 wwl0_53 wwl0_20 wwl0_31 wwl0_42 in0_56 in0_12
+ in0_23 in0_34 in0_45 wwl0_54 wwl0_10 wwl0_21 wwl0_32 wwl0_43 gnd in0_57 in0_46 in0_13
+ in0_24 in0_35 wwl0_55 wwl0_11 wwl0_22 wwl0_33 wwl0_44 rwl0_60 in0_58 in0_47 in0_14
+ in0_25 in0_36 wwl0_56 wwl0_45 wwl0_12 wwl0_23 wwl0_34 rwl0_61 rwl0_50 rwl0_0 in0_59
+ in0_48 in0_15 in0_26 in0_37 wwl0_57 wwl0_46 wwl0_13 wwl0_24 wwl0_35 rwl0_40 rwl0_62
+ rwl0_51 in0_49 rwl0_1 in0_16 in0_27 in0_38 wwl0_58 wwl0_47 wwl0_14 wwl0_25 wwl0_36
+ rwl0_63 rwl0_52 rwl0_30 rwl0_41 rwl0_2 in0_17 in0_28 in0_39 wwl0_59 wwl0_48 wwl0_15
+ wwl0_26 wwl0_37 in2_0 in1_60 rwl0_53 rwl0_20 rwl0_31 rwl0_42 vdd_uq30 rwl0_3 in0_18
+ in0_29 wwl0_49 wwl0_16 wwl0_27 wwl0_38 in2_1 in1_61 in1_50 rwl0_54 rwl0_10 rwl0_21
+ rwl0_32 rwl0_43 vdd_uq20 rwl0_4 in0_19 wwl0_17 wwl0_28 wwl0_39 in2_2 in1_62 in1_51
+ in1_40 rwl0_55 rwl0_11 rwl0_22 rwl0_33 rwl0_44 vdd_uq10 vdd_uq21 rwl0_5 wwl0_18
+ wwl0_29 in2_3 in1_63 in1_52 in1_30 in1_41 in0_0 rwl0_56 rwl0_12 rwl0_23 rwl0_34
+ rwl0_45 vdd_uq11 vdd_uq22 rwl0_6 wwl0_19 in2_4 in1_53 in1_20 in1_31 in1_42 in0_1
+ rwl0_57 rwl0_46 rwl0_13 rwl0_24 rwl0_35 vdd_uq23 vdd_uq12 rwl0_7 in2_5 in1_54 in1_10
+ in1_21 in1_32 in1_43 in0_2 rwl0_58 rwl0_47 rwl0_14 rwl0_25 rwl0_36 vdd_uq24 vdd_uq13
+ rwl0_8 vdd in2_6 in1_55 in1_11 in1_22 in1_33 in1_44 in0_3 rwl0_59 rwl0_48 rwl0_15
+ rwl0_26 rwl0_37 vdd_uq25 vdd_uq14 rwl0_9 in2_7 in1_56 in1_45 in1_12 in1_23 in1_34
+ in0_4 rwl0_49 rwl0_16 rwl0_27 rwl0_38 vdd_uq26 vdd_uq15 in2_8 in1_13 in1_24 in1_35
+ in1_57 in1_46 in0_5 rwl0_17 rwl0_28 rwl0_39 vdd_uq16 rwl1_60 vdd_uq27 in2_9 in1_58
+ in1_47 in1_14 in1_25 in1_36 in0_6 rwl0_18 rwl0_29 rwl1_61 vdd_uq28 rwl1_50 vdd_uq17
+ in1_59 in1_48 in1_15 in1_26 in1_37 in0_7 rwl0_19 rwl1_62 vdd_uq29 rwl1_51 vdd_uq18
+ rwl1_40 in1_49 in1_16 in1_27 in1_38 in0_8 vdd_uq19 rwl1_63 rwl1_52 rwl1_30 rwl1_41
+ in1_17 in1_28 in1_39 in0_9 in2_60 rwl1_53 rwl1_20 rwl1_31 rwl1_42 in1_18 in1_29
+ in2_61 in2_50 rwl1_54 rwl1_10 rwl1_21 rwl1_32 rwl1_43
Xwordline_driver_cell_18 in0_45 vdd_uq21 gnd wl_en in1_45 in2_45 rwl0_45 wwl0_45 rwl1_45
+ wordline_driver_cell
Xwordline_driver_cell_29 in0_34 vdd_uq16 gnd wl_en in1_34 in2_34 rwl0_34 wwl0_34 rwl1_34
+ wordline_driver_cell
Xwordline_driver_cell_19 in0_44 vdd_uq21 gnd wl_en in1_44 in2_44 rwl0_44 wwl0_44 rwl1_44
+ wordline_driver_cell
Xwordline_driver_cell_0 in0_63 vdd_uq30 gnd wl_en in1_63 in2_63 rwl0_63 wwl0_63 rwl1_63
+ wordline_driver_cell
Xwordline_driver_cell_1 in0_62 vdd_uq30 gnd wl_en in1_62 in2_62 rwl0_62 wwl0_62 rwl1_62
+ wordline_driver_cell
Xwordline_driver_cell_60 in0_3 vdd gnd wl_en in1_3 in2_3 rwl0_3 wwl0_3 rwl1_3 wordline_driver_cell
Xwordline_driver_cell_2 in0_61 vdd_uq29 gnd wl_en in1_61 in2_61 rwl0_61 wwl0_61 rwl1_61
+ wordline_driver_cell
Xwordline_driver_cell_61 in0_2 vdd gnd wl_en in1_2 in2_2 rwl0_2 wwl0_2 rwl1_2 wordline_driver_cell
Xwordline_driver_cell_50 in0_13 vdd_uq5 gnd wl_en in1_13 in2_13 rwl0_13 wwl0_13 rwl1_13
+ wordline_driver_cell
Xwordline_driver_cell_3 in0_60 vdd_uq29 gnd wl_en in1_60 in2_60 rwl0_60 wwl0_60 rwl1_60
+ wordline_driver_cell
Xwordline_driver_cell_40 in0_23 vdd_uq10 gnd wl_en in1_23 in2_23 rwl0_23 wwl0_23 rwl1_23
+ wordline_driver_cell
Xwordline_driver_cell_62 in0_1 vdd_uq0 gnd wl_en in1_1 in2_1 rwl0_1 wwl0_1 rwl1_1
+ wordline_driver_cell
Xwordline_driver_cell_51 in0_12 vdd_uq5 gnd wl_en in1_12 in2_12 rwl0_12 wwl0_12 rwl1_12
+ wordline_driver_cell
Xwordline_driver_cell_4 in0_59 vdd_uq28 gnd wl_en in1_59 in2_59 rwl0_59 wwl0_59 rwl1_59
+ wordline_driver_cell
Xwordline_driver_cell_30 in0_33 vdd_uq15 gnd wl_en in1_33 in2_33 rwl0_33 wwl0_33 rwl1_33
+ wordline_driver_cell
Xwordline_driver_cell_41 in0_22 vdd_uq10 gnd wl_en in1_22 in2_22 rwl0_22 wwl0_22 rwl1_22
+ wordline_driver_cell
Xwordline_driver_cell_63 in0_0 vdd_uq0 gnd wl_en in1_0 in2_0 rwl0_0 wwl0_0 rwl1_0
+ wordline_driver_cell
Xwordline_driver_cell_52 in0_11 vdd_uq4 gnd wl_en in1_11 in2_11 rwl0_11 wwl0_11 rwl1_11
+ wordline_driver_cell
Xwordline_driver_cell_5 in0_58 vdd_uq28 gnd wl_en in1_58 in2_58 rwl0_58 wwl0_58 rwl1_58
+ wordline_driver_cell
Xwordline_driver_cell_20 in0_43 vdd_uq20 gnd wl_en in1_43 in2_43 rwl0_43 wwl0_43 rwl1_43
+ wordline_driver_cell
Xwordline_driver_cell_31 in0_32 vdd_uq15 gnd wl_en in1_32 in2_32 rwl0_32 wwl0_32 rwl1_32
+ wordline_driver_cell
Xwordline_driver_cell_42 in0_21 vdd_uq9 gnd wl_en in1_21 in2_21 rwl0_21 wwl0_21 rwl1_21
+ wordline_driver_cell
Xwordline_driver_cell_53 in0_10 vdd_uq4 gnd wl_en in1_10 in2_10 rwl0_10 wwl0_10 rwl1_10
+ wordline_driver_cell
Xwordline_driver_cell_6 in0_57 vdd_uq27 gnd wl_en in1_57 in2_57 rwl0_57 wwl0_57 rwl1_57
+ wordline_driver_cell
Xwordline_driver_cell_10 in0_53 vdd_uq25 gnd wl_en in1_53 in2_53 rwl0_53 wwl0_53 rwl1_53
+ wordline_driver_cell
Xwordline_driver_cell_21 in0_42 vdd_uq20 gnd wl_en in1_42 in2_42 rwl0_42 wwl0_42 rwl1_42
+ wordline_driver_cell
Xwordline_driver_cell_32 in0_31 vdd_uq14 gnd wl_en in1_31 in2_31 rwl0_31 wwl0_31 rwl1_31
+ wordline_driver_cell
Xwordline_driver_cell_43 in0_20 vdd_uq9 gnd wl_en in1_20 in2_20 rwl0_20 wwl0_20 rwl1_20
+ wordline_driver_cell
Xwordline_driver_cell_54 in0_9 vdd_uq3 gnd wl_en in1_9 in2_9 rwl0_9 wwl0_9 rwl1_9
+ wordline_driver_cell
Xwordline_driver_cell_7 in0_56 vdd_uq27 gnd wl_en in1_56 in2_56 rwl0_56 wwl0_56 rwl1_56
+ wordline_driver_cell
Xwordline_driver_cell_11 in0_52 vdd_uq25 gnd wl_en in1_52 in2_52 rwl0_52 wwl0_52 rwl1_52
+ wordline_driver_cell
Xwordline_driver_cell_22 in0_41 vdd_uq19 gnd wl_en in1_41 in2_41 rwl0_41 wwl0_41 rwl1_41
+ wordline_driver_cell
Xwordline_driver_cell_33 in0_30 vdd_uq14 gnd wl_en in1_30 in2_30 rwl0_30 wwl0_30 rwl1_30
+ wordline_driver_cell
Xwordline_driver_cell_55 in0_8 vdd_uq3 gnd wl_en in1_8 in2_8 rwl0_8 wwl0_8 rwl1_8
+ wordline_driver_cell
Xwordline_driver_cell_44 in0_19 vdd_uq8 gnd wl_en in1_19 in2_19 rwl0_19 wwl0_19 rwl1_19
+ wordline_driver_cell
Xwordline_driver_cell_8 in0_55 vdd_uq26 gnd wl_en in1_55 in2_55 rwl0_55 wwl0_55 rwl1_55
+ wordline_driver_cell
Xwordline_driver_cell_12 in0_51 vdd_uq24 gnd wl_en in1_51 in2_51 rwl0_51 wwl0_51 rwl1_51
+ wordline_driver_cell
Xwordline_driver_cell_23 in0_40 vdd_uq19 gnd wl_en in1_40 in2_40 rwl0_40 wwl0_40 rwl1_40
+ wordline_driver_cell
Xwordline_driver_cell_34 in0_29 vdd_uq13 gnd wl_en in1_29 in2_29 rwl0_29 wwl0_29 rwl1_29
+ wordline_driver_cell
Xwordline_driver_cell_56 in0_7 vdd_uq2 gnd wl_en in1_7 in2_7 rwl0_7 wwl0_7 rwl1_7
+ wordline_driver_cell
Xwordline_driver_cell_45 in0_18 vdd_uq8 gnd wl_en in1_18 in2_18 rwl0_18 wwl0_18 rwl1_18
+ wordline_driver_cell
Xwordline_driver_cell_9 in0_54 vdd_uq26 gnd wl_en in1_54 in2_54 rwl0_54 wwl0_54 rwl1_54
+ wordline_driver_cell
Xwordline_driver_cell_13 in0_50 vdd_uq24 gnd wl_en in1_50 in2_50 rwl0_50 wwl0_50 rwl1_50
+ wordline_driver_cell
Xwordline_driver_cell_24 in0_39 vdd_uq18 gnd wl_en in1_39 in2_39 rwl0_39 wwl0_39 rwl1_39
+ wordline_driver_cell
Xwordline_driver_cell_35 in0_28 vdd_uq13 gnd wl_en in1_28 in2_28 rwl0_28 wwl0_28 rwl1_28
+ wordline_driver_cell
Xwordline_driver_cell_57 in0_6 vdd_uq2 gnd wl_en in1_6 in2_6 rwl0_6 wwl0_6 rwl1_6
+ wordline_driver_cell
Xwordline_driver_cell_46 in0_17 vdd_uq7 gnd wl_en in1_17 in2_17 rwl0_17 wwl0_17 rwl1_17
+ wordline_driver_cell
Xwordline_driver_cell_14 in0_49 vdd_uq23 gnd wl_en in1_49 in2_49 rwl0_49 wwl0_49 rwl1_49
+ wordline_driver_cell
Xwordline_driver_cell_25 in0_38 vdd_uq18 gnd wl_en in1_38 in2_38 rwl0_38 wwl0_38 rwl1_38
+ wordline_driver_cell
Xwordline_driver_cell_36 in0_27 vdd_uq12 gnd wl_en in1_27 in2_27 rwl0_27 wwl0_27 rwl1_27
+ wordline_driver_cell
Xwordline_driver_cell_58 in0_5 vdd_uq1 gnd wl_en in1_5 in2_5 rwl0_5 wwl0_5 rwl1_5
+ wordline_driver_cell
Xwordline_driver_cell_47 in0_16 vdd_uq7 gnd wl_en in1_16 in2_16 rwl0_16 wwl0_16 rwl1_16
+ wordline_driver_cell
Xwordline_driver_cell_15 in0_48 vdd_uq23 gnd wl_en in1_48 in2_48 rwl0_48 wwl0_48 rwl1_48
+ wordline_driver_cell
Xwordline_driver_cell_26 in0_37 vdd_uq17 gnd wl_en in1_37 in2_37 rwl0_37 wwl0_37 rwl1_37
+ wordline_driver_cell
Xwordline_driver_cell_37 in0_26 vdd_uq12 gnd wl_en in1_26 in2_26 rwl0_26 wwl0_26 rwl1_26
+ wordline_driver_cell
Xwordline_driver_cell_59 in0_4 vdd_uq1 gnd wl_en in1_4 in2_4 rwl0_4 wwl0_4 rwl1_4
+ wordline_driver_cell
Xwordline_driver_cell_48 in0_15 vdd_uq6 gnd wl_en in1_15 in2_15 rwl0_15 wwl0_15 rwl1_15
+ wordline_driver_cell
Xwordline_driver_cell_16 in0_47 vdd_uq22 gnd wl_en in1_47 in2_47 rwl0_47 wwl0_47 rwl1_47
+ wordline_driver_cell
Xwordline_driver_cell_27 in0_36 vdd_uq17 gnd wl_en in1_36 in2_36 rwl0_36 wwl0_36 rwl1_36
+ wordline_driver_cell
Xwordline_driver_cell_38 in0_25 vdd_uq11 gnd wl_en in1_25 in2_25 rwl0_25 wwl0_25 rwl1_25
+ wordline_driver_cell
Xwordline_driver_cell_49 in0_14 vdd_uq6 gnd wl_en in1_14 in2_14 rwl0_14 wwl0_14 rwl1_14
+ wordline_driver_cell
Xwordline_driver_cell_17 in0_46 vdd_uq22 gnd wl_en in1_46 in2_46 rwl0_46 wwl0_46 rwl1_46
+ wordline_driver_cell
Xwordline_driver_cell_28 in0_35 vdd_uq16 gnd wl_en in1_35 in2_35 rwl0_35 wwl0_35 rwl1_35
+ wordline_driver_cell
Xwordline_driver_cell_39 in0_24 vdd_uq11 gnd wl_en in1_24 in2_24 rwl0_24 wwl0_24 rwl1_24
+ wordline_driver_cell
.ends

.subckt port_address addr2 wl_en wwl0_0 rwl1_0 rwl1_55 rwl1_44 rwl1_11 rwl1_22 rwl1_33
+ addr3 gnd rwl1_1 wwl0_1 vdd_uq0 rwl1_56 rwl1_45 rwl1_34 rwl1_12 rwl1_23 addr4 vdd_uq82
+ rwl1_2 wwl0_2 vdd_uq2 rwl1_13 rwl1_24 rwl1_57 rwl1_46 rwl1_35 addr5 vdd_uq62 rwl1_3
+ wwl0_3 rwl1_58 rwl1_47 rwl1_36 rwl1_14 rwl1_25 addr6 vdd_uq64 vdd_uq40 wwl0_4 rwl1_4
+ vdd_uq3 rwl1_59 rwl1_48 rwl1_37 rwl1_15 rwl1_26 addr7 vdd_uq66 vdd_uq44 vdd_uq4
+ rwl1_5 wwl0_5 rwl1_49 rwl1_38 rwl1_16 rwl1_27 vdd_uq68 vdd_uq46 vdd_uq8 rwl1_6 wwl0_6
+ vdd_uq6 rwl1_39 rwl1_17 rwl1_28 vdd_uq70 vdd_uq48 vdd_uq10 rwl1_7 wwl0_7 rwl1_18
+ rwl1_29 vdd_uq72 vdd_uq50 vdd_uq14 rwl1_8 wwl0_8 vdd_uq7 rwl1_19 vdd_uq74 vdd_uq52
+ vdd_uq18 rwl1_9 wwl0_9 vdd_uq76 vdd_uq54 vdd_uq22 vdd_uq9 vdd_uq78 vdd_uq56 vdd_uq26
+ wwl0_60 vdd_uq80 vdd_uq58 vdd_uq28 wwl0_61 wwl0_50 vdd_uq60 vdd_uq32 wwl0_62 wwl0_51
+ wwl0_40 vdd_uq36 wwl0_63 wwl0_52 wwl0_41 wwl0_30 vdd wwl0_53 wwl0_42 wwl0_20 wwl0_31
+ addr0 wwl0_54 wwl0_43 wwl0_10 wwl0_21 wwl0_32 addr1 wwl0_55 wwl0_44 wwl0_33 wwl0_11
+ wwl0_22 rwl0_60 vdd_uq81 wwl0_56 wwl0_45 wwl0_34 wwl0_12 wwl0_23 rwl0_61 rwl0_50
+ vdd_uq71 rwl0_0 wwl0_57 wwl0_46 wwl0_35 wwl0_13 wwl0_24 vdd_uq79 rwl0_40 rwl0_62
+ rwl0_51 vdd_uq61 rwl0_1 wwl0_58 wwl0_47 wwl0_36 wwl0_14 wwl0_25 rwl0_63 rwl0_52
+ rwl0_41 rwl0_30 vdd_uq51 vdd_uq73 rwl0_2 wwl0_59 wwl0_48 wwl0_37 wwl0_15 wwl0_26
+ rwl0_53 rwl0_42 rwl0_20 rwl0_31 vdd_uq42 vdd_uq30 vdd_uq63 rwl0_3 wwl0_49 wwl0_38
+ wwl0_16 wwl0_27 rwl0_54 rwl0_43 rwl0_10 rwl0_21 rwl0_32 vdd_uq31 vdd_uq20 vdd_uq53
+ vdd_uq75 rwl0_4 wwl0_39 wwl0_17 wwl0_28 rwl0_55 rwl0_44 rwl0_33 rwl0_11 rwl0_22
+ vdd_uq21 vdd_uq43 vdd_uq65 rwl0_5 wwl0_18 wwl0_29 rwl0_56 rwl0_45 rwl0_34 rwl0_12
+ rwl0_23 vdd_uq12 vdd_uq34 vdd_uq55 vdd_uq77 rwl0_6 wwl0_19 rwl0_57 rwl0_46 rwl0_35
+ rwl0_13 rwl0_24 vdd_uq24 vdd_uq45 vdd_uq67 rwl0_7 rwl0_58 rwl0_47 rwl0_36 rwl0_14
+ rwl0_25 vdd_uq35 vdd_uq13 vdd_uq57 rwl0_8 rwl0_59 rwl0_48 rwl0_37 rwl0_15 rwl0_26
+ vdd_uq25 vdd_uq47 vdd_uq69 rwl0_9 rwl0_49 rwl0_38 rwl0_16 rwl0_27 vdd_uq38 vdd_uq16
+ vdd_uq59 rwl0_39 rwl0_17 rwl0_28 rwl1_60 vdd_uq27 vdd_uq49 rwl0_18 rwl0_29 rwl1_61
+ rwl1_50 vdd_uq39 vdd_uq17 rwl0_19 rwl1_62 rwl1_51 rwl1_40 rwl1_63 rwl1_52 rwl1_41
+ rwl1_30 rwl1_53 rwl1_42 rwl1_20 rwl1_31 rwl1_54 rwl1_43 rwl1_10 rwl1_21 rwl1_32
Xhierarchical_decoder_0 addr0 wordline_driver_array_0/in0_6 wordline_driver_array_0/in2_9
+ addr2 wordline_driver_array_0/in1_54 wordline_driver_array_0/in1_43 wordline_driver_array_0/in1_32
+ wordline_driver_array_0/in1_21 wordline_driver_array_0/in1_10 addr1 gnd addr3 wordline_driver_array_0/in1_55
+ wordline_driver_array_0/in1_44 wordline_driver_array_0/in1_33 wordline_driver_array_0/in1_22
+ wordline_driver_array_0/in1_11 wordline_driver_array_0/in0_7 addr4 wordline_driver_array_0/in1_56
+ wordline_driver_array_0/in1_45 wordline_driver_array_0/in1_34 wordline_driver_array_0/in1_23
+ wordline_driver_array_0/in1_12 vdd_uq6 wordline_driver_array_0/in0_8 wordline_driver_array_0/in1_57
+ wordline_driver_array_0/in1_46 wordline_driver_array_0/in1_35 wordline_driver_array_0/in1_24
+ wordline_driver_array_0/in1_13 wordline_driver_array_0/in0_9 wordline_driver_array_0/in1_58
+ wordline_driver_array_0/in1_47 wordline_driver_array_0/in1_36 wordline_driver_array_0/in1_25
+ wordline_driver_array_0/in1_14 vdd_uq12 addr5 wordline_driver_array_0/in1_59 wordline_driver_array_0/in1_48
+ wordline_driver_array_0/in1_37 wordline_driver_array_0/in1_26 wordline_driver_array_0/in1_15
+ addr6 wordline_driver_array_0/in1_49 wordline_driver_array_0/in1_38 wordline_driver_array_0/in1_27
+ wordline_driver_array_0/in1_16 vdd_uq16 addr7 wordline_driver_array_0/in2_60 wordline_driver_array_0/in1_39
+ wordline_driver_array_0/in1_28 wordline_driver_array_0/in1_17 wordline_driver_array_0/in1_29
+ wordline_driver_array_0/in1_18 wordline_driver_array_0/in2_61 wordline_driver_array_0/in2_50
+ vdd_uq20 wordline_driver_array_0/in2_62 wordline_driver_array_0/in2_51 wordline_driver_array_0/in2_40
+ wordline_driver_array_0/in1_19 wordline_driver_array_0/in2_63 wordline_driver_array_0/in2_52
+ wordline_driver_array_0/in2_41 wordline_driver_array_0/in2_30 vdd_uq24 wordline_driver_array_0/in1_0
+ wordline_driver_array_0/in2_53 wordline_driver_array_0/in2_42 wordline_driver_array_0/in2_31
+ wordline_driver_array_0/in2_20 wordline_driver_array_0/in1_1 wordline_driver_array_0/in2_54
+ wordline_driver_array_0/in2_43 wordline_driver_array_0/in2_32 wordline_driver_array_0/in2_21
+ wordline_driver_array_0/in2_10 wordline_driver_array_0/in1_2 wordline_driver_array_0/in2_55
+ wordline_driver_array_0/in2_44 wordline_driver_array_0/in2_33 wordline_driver_array_0/in2_22
+ wordline_driver_array_0/in2_11 wordline_driver_array_0/in1_3 wordline_driver_array_0/in2_56
+ wordline_driver_array_0/in2_45 wordline_driver_array_0/in2_34 wordline_driver_array_0/in2_23
+ wordline_driver_array_0/in2_12 wordline_driver_array_0/in1_4 wordline_driver_array_0/in2_57
+ wordline_driver_array_0/in2_46 wordline_driver_array_0/in2_35 wordline_driver_array_0/in2_24
+ wordline_driver_array_0/in2_13 wordline_driver_array_0/in1_5 wordline_driver_array_0/in2_58
+ wordline_driver_array_0/in2_47 wordline_driver_array_0/in2_36 wordline_driver_array_0/in2_25
+ wordline_driver_array_0/in2_14 wordline_driver_array_0/in1_6 wordline_driver_array_0/in2_59
+ wordline_driver_array_0/in2_48 wordline_driver_array_0/in2_37 wordline_driver_array_0/in2_26
+ wordline_driver_array_0/in2_15 wordline_driver_array_0/in1_7 wordline_driver_array_0/in2_49
+ wordline_driver_array_0/in2_38 wordline_driver_array_0/in2_27 wordline_driver_array_0/in2_16
+ wordline_driver_array_0/in1_8 wordline_driver_array_0/in0_60 wordline_driver_array_0/in2_39
+ wordline_driver_array_0/in2_28 wordline_driver_array_0/in2_17 wordline_driver_array_0/in1_9
+ wordline_driver_array_0/in0_61 wordline_driver_array_0/in0_50 vdd_uq82 wordline_driver_array_0/in2_29
+ wordline_driver_array_0/in2_18 wordline_driver_array_0/in0_62 wordline_driver_array_0/in0_51
+ wordline_driver_array_0/in0_40 wordline_driver_array_0/in2_19 vdd_uq62 wordline_driver_array_0/in0_63
+ wordline_driver_array_0/in0_52 wordline_driver_array_0/in0_41 wordline_driver_array_0/in0_30
+ vdd_uq64 vdd_uq40 wordline_driver_array_0/in0_53 wordline_driver_array_0/in0_42
+ wordline_driver_array_0/in0_31 wordline_driver_array_0/in0_20 vdd_uq66 vdd_uq44
+ vdd_uq4 wordline_driver_array_0/in0_54 wordline_driver_array_0/in0_43 wordline_driver_array_0/in0_32
+ wordline_driver_array_0/in0_21 wordline_driver_array_0/in0_10 vdd_uq68 vdd_uq46
+ vdd_uq8 wordline_driver_array_0/in0_55 wordline_driver_array_0/in0_44 wordline_driver_array_0/in0_33
+ wordline_driver_array_0/in0_22 wordline_driver_array_0/in0_11 vdd_uq70 vdd_uq48
+ vdd_uq30 vdd_uq10 wordline_driver_array_0/in0_56 wordline_driver_array_0/in0_45
+ wordline_driver_array_0/in0_34 wordline_driver_array_0/in0_23 wordline_driver_array_0/in0_12
+ vdd_uq72 vdd_uq50 vdd_uq14 wordline_driver_array_0/in0_57 wordline_driver_array_0/in0_46
+ wordline_driver_array_0/in0_35 wordline_driver_array_0/in0_24 wordline_driver_array_0/in0_13
+ wordline_driver_array_0/in2_0 vdd_uq74 vdd_uq52 vdd_uq34 vdd_uq18 wordline_driver_array_0/in0_58
+ wordline_driver_array_0/in0_47 wordline_driver_array_0/in0_36 wordline_driver_array_0/in0_25
+ wordline_driver_array_0/in0_14 vdd_uq2 wordline_driver_array_0/in2_1 vdd_uq76 vdd_uq54
+ vdd_uq22 wordline_driver_array_0/in0_59 wordline_driver_array_0/in0_48 wordline_driver_array_0/in0_37
+ wordline_driver_array_0/in0_26 wordline_driver_array_0/in0_15 wordline_driver_array_0/in2_2
+ vdd_uq78 vdd_uq56 vdd_uq26 vdd_uq38 wordline_driver_array_0/in0_27 wordline_driver_array_0/in0_16
+ wordline_driver_array_0/in0_49 wordline_driver_array_0/in0_38 wordline_driver_array_0/in0_0
+ wordline_driver_array_0/in2_3 vdd_uq80 vdd_uq58 vdd_uq28 wordline_driver_array_0/in0_39
+ wordline_driver_array_0/in0_28 wordline_driver_array_0/in0_17 wordline_driver_array_0/in2_4
+ wordline_driver_array_0/in1_60 wordline_driver_array_0/in0_1 vdd_uq60 vdd_uq32 vdd_uq42
+ wordline_driver_array_0/in1_61 wordline_driver_array_0/in1_50 wordline_driver_array_0/in0_29
+ wordline_driver_array_0/in0_18 wordline_driver_array_0/in0_2 wordline_driver_array_0/in2_5
+ vdd_uq36 wordline_driver_array_0/in0_19 wordline_driver_array_0/in2_6 wordline_driver_array_0/in1_62
+ wordline_driver_array_0/in1_51 wordline_driver_array_0/in1_40 wordline_driver_array_0/in0_3
+ vdd wordline_driver_array_0/in0_4 wordline_driver_array_0/in2_7 wordline_driver_array_0/in1_63
+ wordline_driver_array_0/in1_52 wordline_driver_array_0/in1_41 wordline_driver_array_0/in1_30
+ wordline_driver_array_0/in2_8 wordline_driver_array_0/in1_53 wordline_driver_array_0/in1_42
+ wordline_driver_array_0/in1_31 wordline_driver_array_0/in1_20 wordline_driver_array_0/in0_5
+ hierarchical_decoder
Xwordline_driver_array_0 wl_en wordline_driver_array_0/in1_19 rwl1_0 wwl0_0 wordline_driver_array_0/in2_62
+ wordline_driver_array_0/in2_51 wordline_driver_array_0/in2_40 rwl1_55 rwl1_11 rwl1_22
+ rwl1_33 rwl1_44 rwl1_1 wordline_driver_array_0/in2_63 wordline_driver_array_0/in2_52
+ wwl0_1 wordline_driver_array_0/in2_30 wordline_driver_array_0/in2_41 vdd_uq0 rwl1_56
+ rwl1_12 rwl1_23 rwl1_34 rwl1_45 rwl1_2 wwl0_2 wordline_driver_array_0/in2_53 vdd_uq7
+ wordline_driver_array_0/in2_20 wordline_driver_array_0/in2_31 wordline_driver_array_0/in2_42
+ rwl1_13 rwl1_24 rwl1_57 rwl1_46 rwl1_35 rwl1_3 wwl0_3 wordline_driver_array_0/in2_54
+ wordline_driver_array_0/in2_10 wordline_driver_array_0/in2_21 wordline_driver_array_0/in2_32
+ wordline_driver_array_0/in2_43 vdd_uq9 rwl1_58 rwl1_47 rwl1_14 rwl1_25 rwl1_36 wwl0_4
+ rwl1_4 wordline_driver_array_0/in2_55 wordline_driver_array_0/in2_11 wordline_driver_array_0/in2_22
+ wordline_driver_array_0/in2_33 wordline_driver_array_0/in2_44 vdd_uq13 rwl1_59 rwl1_48
+ rwl1_15 rwl1_26 rwl1_37 rwl1_5 wwl0_5 wordline_driver_array_0/in2_56 wordline_driver_array_0/in2_45
+ wordline_driver_array_0/in2_12 wordline_driver_array_0/in2_23 wordline_driver_array_0/in2_34
+ vdd_uq17 rwl1_49 rwl1_16 rwl1_27 rwl1_38 wordline_driver_array_0/in1_0 rwl1_6 wordline_driver_array_0/in2_57
+ wordline_driver_array_0/in2_46 wwl0_6 wordline_driver_array_0/in2_13 wordline_driver_array_0/in2_24
+ wordline_driver_array_0/in2_35 vdd_uq21 rwl1_17 rwl1_28 rwl1_39 wordline_driver_array_0/in1_1
+ rwl1_7 wwl0_7 wordline_driver_array_0/in2_14 wordline_driver_array_0/in2_58 wordline_driver_array_0/in2_47
+ vdd_uq25 wordline_driver_array_0/in2_25 wordline_driver_array_0/in2_36 rwl1_18 rwl1_29
+ wordline_driver_array_0/in1_2 rwl1_8 wwl0_8 wordline_driver_array_0/in2_59 wordline_driver_array_0/in2_48
+ wordline_driver_array_0/in2_15 wordline_driver_array_0/in2_26 wordline_driver_array_0/in2_37
+ vdd_uq27 wordline_driver_array_0/in1_3 rwl1_19 rwl1_9 wwl0_9 wordline_driver_array_0/in2_49
+ wordline_driver_array_0/in2_16 wordline_driver_array_0/in2_27 wordline_driver_array_0/in2_38
+ vdd_uq31 wordline_driver_array_0/in1_4 wordline_driver_array_0/in0_60 wordline_driver_array_0/in2_17
+ wordline_driver_array_0/in2_28 wordline_driver_array_0/in2_39 vdd_uq35 wordline_driver_array_0/in1_5
+ wordline_driver_array_0/in0_61 wordline_driver_array_0/in0_50 wordline_driver_array_0/in2_18
+ wordline_driver_array_0/in2_29 wordline_driver_array_0/in1_6 wordline_driver_array_0/in0_51
+ wordline_driver_array_0/in0_40 wordline_driver_array_0/in0_62 wwl0_60 wordline_driver_array_0/in2_19
+ wordline_driver_array_0/in1_7 wordline_driver_array_0/in0_63 wordline_driver_array_0/in0_52
+ wordline_driver_array_0/in0_30 wordline_driver_array_0/in0_41 wwl0_61 wwl0_50 wordline_driver_array_0/in1_8
+ wordline_driver_array_0/in0_53 wordline_driver_array_0/in0_20 wordline_driver_array_0/in0_31
+ wordline_driver_array_0/in0_42 wwl0_62 wwl0_51 wwl0_40 wordline_driver_array_0/in1_9
+ wordline_driver_array_0/in0_54 wordline_driver_array_0/in0_10 wordline_driver_array_0/in0_21
+ wordline_driver_array_0/in0_32 wordline_driver_array_0/in0_43 wwl0_63 wwl0_52 wwl0_30
+ wwl0_41 wordline_driver_array_0/in0_55 wordline_driver_array_0/in0_11 wordline_driver_array_0/in0_22
+ wordline_driver_array_0/in0_33 wordline_driver_array_0/in0_44 wwl0_53 wwl0_20 wwl0_31
+ wwl0_42 wordline_driver_array_0/in0_56 wordline_driver_array_0/in0_12 wordline_driver_array_0/in0_23
+ wordline_driver_array_0/in0_34 wordline_driver_array_0/in0_45 wwl0_54 wwl0_10 wwl0_21
+ wwl0_32 wwl0_43 gnd wordline_driver_array_0/in0_57 wordline_driver_array_0/in0_46
+ wordline_driver_array_0/in0_13 wordline_driver_array_0/in0_24 wordline_driver_array_0/in0_35
+ wwl0_55 wwl0_11 wwl0_22 wwl0_33 wwl0_44 rwl0_60 wordline_driver_array_0/in0_58 wordline_driver_array_0/in0_47
+ wordline_driver_array_0/in0_14 wordline_driver_array_0/in0_25 wordline_driver_array_0/in0_36
+ wwl0_56 wwl0_45 wwl0_12 wwl0_23 wwl0_34 rwl0_61 rwl0_50 rwl0_0 wordline_driver_array_0/in0_59
+ wordline_driver_array_0/in0_48 wordline_driver_array_0/in0_15 wordline_driver_array_0/in0_26
+ wordline_driver_array_0/in0_37 wwl0_57 wwl0_46 wwl0_13 wwl0_24 wwl0_35 rwl0_40 rwl0_62
+ rwl0_51 wordline_driver_array_0/in0_49 rwl0_1 wordline_driver_array_0/in0_16 wordline_driver_array_0/in0_27
+ wordline_driver_array_0/in0_38 wwl0_58 wwl0_47 wwl0_14 wwl0_25 wwl0_36 rwl0_63 rwl0_52
+ rwl0_30 rwl0_41 rwl0_2 wordline_driver_array_0/in0_17 wordline_driver_array_0/in0_28
+ wordline_driver_array_0/in0_39 wwl0_59 wwl0_48 wwl0_15 wwl0_26 wwl0_37 wordline_driver_array_0/in2_0
+ wordline_driver_array_0/in1_60 rwl0_53 rwl0_20 rwl0_31 rwl0_42 vdd_uq81 rwl0_3 wordline_driver_array_0/in0_18
+ wordline_driver_array_0/in0_29 wwl0_49 wwl0_16 wwl0_27 wwl0_38 wordline_driver_array_0/in2_1
+ wordline_driver_array_0/in1_61 wordline_driver_array_0/in1_50 rwl0_54 rwl0_10 rwl0_21
+ rwl0_32 rwl0_43 vdd_uq61 rwl0_4 wordline_driver_array_0/in0_19 wwl0_17 wwl0_28 wwl0_39
+ wordline_driver_array_0/in2_2 wordline_driver_array_0/in1_62 wordline_driver_array_0/in1_51
+ wordline_driver_array_0/in1_40 rwl0_55 rwl0_11 rwl0_22 rwl0_33 rwl0_44 vdd_uq39
+ vdd_uq63 rwl0_5 wwl0_18 wwl0_29 wordline_driver_array_0/in2_3 wordline_driver_array_0/in1_63
+ wordline_driver_array_0/in1_52 wordline_driver_array_0/in1_30 wordline_driver_array_0/in1_41
+ wordline_driver_array_0/in0_0 rwl0_56 rwl0_12 rwl0_23 rwl0_34 rwl0_45 vdd_uq43 vdd_uq65
+ rwl0_6 wwl0_19 wordline_driver_array_0/in2_4 wordline_driver_array_0/in1_53 wordline_driver_array_0/in1_20
+ wordline_driver_array_0/in1_31 wordline_driver_array_0/in1_42 wordline_driver_array_0/in0_1
+ rwl0_57 rwl0_46 rwl0_13 rwl0_24 rwl0_35 vdd_uq67 vdd_uq45 rwl0_7 wordline_driver_array_0/in2_5
+ wordline_driver_array_0/in1_54 wordline_driver_array_0/in1_10 wordline_driver_array_0/in1_21
+ wordline_driver_array_0/in1_32 wordline_driver_array_0/in1_43 wordline_driver_array_0/in0_2
+ rwl0_58 rwl0_47 rwl0_14 rwl0_25 rwl0_36 vdd_uq69 vdd_uq47 rwl0_8 vdd_uq3 wordline_driver_array_0/in2_6
+ wordline_driver_array_0/in1_55 wordline_driver_array_0/in1_11 wordline_driver_array_0/in1_22
+ wordline_driver_array_0/in1_33 wordline_driver_array_0/in1_44 wordline_driver_array_0/in0_3
+ rwl0_59 rwl0_48 rwl0_15 rwl0_26 rwl0_37 vdd_uq71 vdd_uq49 rwl0_9 wordline_driver_array_0/in2_7
+ wordline_driver_array_0/in1_56 wordline_driver_array_0/in1_45 wordline_driver_array_0/in1_12
+ wordline_driver_array_0/in1_23 wordline_driver_array_0/in1_34 wordline_driver_array_0/in0_4
+ rwl0_49 rwl0_16 rwl0_27 rwl0_38 vdd_uq73 vdd_uq51 wordline_driver_array_0/in2_8
+ wordline_driver_array_0/in1_13 wordline_driver_array_0/in1_24 wordline_driver_array_0/in1_35
+ wordline_driver_array_0/in1_57 wordline_driver_array_0/in1_46 wordline_driver_array_0/in0_5
+ rwl0_17 rwl0_28 rwl0_39 vdd_uq53 rwl1_60 vdd_uq75 wordline_driver_array_0/in2_9
+ wordline_driver_array_0/in1_58 wordline_driver_array_0/in1_47 wordline_driver_array_0/in1_14
+ wordline_driver_array_0/in1_25 wordline_driver_array_0/in1_36 wordline_driver_array_0/in0_6
+ rwl0_18 rwl0_29 rwl1_61 vdd_uq77 rwl1_50 vdd_uq55 wordline_driver_array_0/in1_59
+ wordline_driver_array_0/in1_48 wordline_driver_array_0/in1_15 wordline_driver_array_0/in1_26
+ wordline_driver_array_0/in1_37 wordline_driver_array_0/in0_7 rwl0_19 rwl1_62 vdd_uq79
+ rwl1_51 vdd_uq57 rwl1_40 wordline_driver_array_0/in1_49 wordline_driver_array_0/in1_16
+ wordline_driver_array_0/in1_27 wordline_driver_array_0/in1_38 wordline_driver_array_0/in0_8
+ vdd_uq59 rwl1_63 rwl1_52 rwl1_30 rwl1_41 wordline_driver_array_0/in1_17 wordline_driver_array_0/in1_28
+ wordline_driver_array_0/in1_39 wordline_driver_array_0/in0_9 wordline_driver_array_0/in2_60
+ rwl1_53 rwl1_20 rwl1_31 rwl1_42 wordline_driver_array_0/in1_18 wordline_driver_array_0/in1_29
+ wordline_driver_array_0/in2_61 wordline_driver_array_0/in2_50 rwl1_54 rwl1_10 rwl1_21
+ rwl1_32 rwl1_43 wordline_driver_array
.ends

.subckt cell_2r1w vdd gnd rbl0 rbl1 wbl0 wwl0 rwl1 rwl0
X0 q qbar vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X1 net2 q gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X2 gnd qbar q gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 wbl0 wwl0 q gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X4 net1 wwl0 qbar gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X5 rbl1 rwl1 net3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X6 vdd q qbar vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X7 rbl0 rwl0 net2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X8 gnd q net3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X9 net1 wbl0 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X10 qbar q gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 net1 wbl0 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt bitcell_array write_bl_0_56 wwl_0_1 read_bl_1_29 read_bl_0_0 rwl_0_0 write_bl_0_44
+ read_bl_0_24 wwl_0_57 rwl_0_47 write_bl_0_53 wwl_0_43 read_bl_0_51 read_bl_1_26
+ read_bl_0_22 write_bl_0_5 wwl_0_35 read_bl_0_39 read_bl_0_2 read_bl_0_48 wwl_0_56
+ wwl_0_37 write_bl_0_3 read_bl_0_37 write_bl_0_20 rwl_1_12 read_bl_0_60 rwl_0_11
+ wwl_0_20 write_bl_0_15 read_bl_0_31 write_bl_0_32 read_bl_0_58 write_bl_0_61 read_bl_0_63
+ read_bl_0_47 rwl_0_24 write_bl_0_12 read_bl_1_21 write_bl_0_30 read_bl_0_29 read_bl_0_10
+ write_bl_0_37 rwl_0_2 read_bl_1_19 read_bl_1_36 read_bl_0_7 write_bl_0_34 read_bl_1_34
+ read_bl_1_57 rwl_1_43 rwl_1_5 wwl_0_42 rwl_0_46 read_bl_1_28 rwl_1_35 write_bl_0_0
+ read_bl_1_55 rwl_1_21 read_bl_0_41 rwl_1_47 read_bl_1_44 read_bl_1_7 wwl_0_55 read_bl_0_50
+ rwl_1_13 write_bl_0_22 write_bl_0_42 read_bl_0_20 rwl_1_15 rwl_1_60 write_bl_0_49
+ wwl_0_33 read_bl_1_4 rwl_0_3 rwl_0_40 read_bl_0_17 rwl_1_57 read_bl_0_12 write_bl_0_58
+ write_bl_0_63 read_bl_1_14 rwl_0_1 read_bl_0_46 read_bl_0_27 read_bl_0_9 read_bl_0_34
+ read_bl_0_25 read_bl_1_30 rwl_0_45 rwl_1_20 read_bl_1_46 rwl_1_46 rwl_0_23 read_bl_1_9
+ rwl_1_24 rwl_1_59 write_bl_0_51 wwl_0_6 wwl_0_32 read_bl_1_6 write_bl_0_39 write_bl_0_2
+ read_bl_0_19 rwl_1_37 write_bl_0_48 rwl_1_56 wwl_0_10 read_bl_1_16 wwl_0_50 rwl_1_34
+ wwl_0_28 read_bl_1_49 wwl_0_54 rwl_1_39 write_bl_0_47 read_bl_1_38 write_bl_0_10
+ wwl_0_3 rwl_0_58 write_bl_0_7 read_bl_1_48 rwl_0_22 wwl_0_5 read_bl_1_56 wwl_0_47
+ read_bl_1_45 rwl_1_58 read_bl_1_8 read_bl_1_54 write_bl_0_41 rwl_1_10 read_bl_0_21
+ rwl_1_36 rwl_0_9 write_bl_0_50 read_bl_0_36 rwl_1_33 wwl_0_40 wwl_0_62 wwl_0_51
+ wwl_0_41 write_bl_0_60 wwl_0_27 read_bl_1_40 rwl_1_32 wwl_0_19 read_bl_0_55 rwl_1_16
+ write_bl_0_46 rwl_0_57 rwl_0_31 read_bl_1_18 read_bl_0_26 write_bl_0_9 read_bl_0_44
+ read_bl_0_53 rwl_0_6 read_bl_0_4 rwl_1_9 read_bl_1_47 wwl_0_24 read_bl_1_25 rwl_0_50
+ write_bl_0_52 read_bl_0_14 rwl_0_34 read_bl_0_42 read_bl_1_52 read_bl_1_23 rwl_0_28
+ write_bl_0_19 read_bl_1_50 rwl_1_19 read_bl_1_62 wwl_0_18 write_bl_0_17 wwl_0_4
+ rwl_0_30 rwl_0_56 write_bl_0_29 read_bl_0_28 write_bl_0_11 read_bl_1_59 write_bl_0_57
+ rwl_0_8 wwl_0_17 write_bl_0_62 write_bl_0_27 read_bl_0_6 wwl_0_59 rwl_1_50 read_bl_0_16
+ rwl_0_44 rwl_0_27 read_bl_0_49 write_bl_0_21 read_bl_0_38 read_bl_1_3 read_bl_1_61
+ rwl_0_21 read_bl_0_57 rwl_0_7 read_bl_0_45 wwl_0_16 read_bl_0_8 write_bl_0_55 read_bl_1_11
+ wwl_0_58 read_bl_0_54 write_bl_0_26 rwl_0_20 rwl_0_62 read_bl_1_33 write_bl_0_4
+ rwl_0_43 wwl_0_26 rwl_1_27 write_bl_0_16 read_bl_1_42 rwl_0_4 write_bl_0_14 write_bl_0_38
+ read_bl_1_51 wwl_0_46 read_bl_0_35 write_bl_0_36 write_bl_0_31 read_bl_1_13 write_bl_0_28
+ rwl_0_19 rwl_1_62 read_bl_0_52 wwl_0_9 read_bl_1_35 rwl_0_61 write_bl_0_43 write_bl_0_6
+ read_bl_0_23 wwl_0_48 read_bl_0_62 read_bl_1_1 wwl_0_45 rwl_1_42 read_bl_0_59 read_bl_1_5
+ rwl_0_49 read_bl_0_18 rwl_1_55 read_bl_1_20 read_bl_1_32 read_bl_1_15 rwl_0_60 read_bl_1_12
+ write_bl_0_45 write_bl_0_8 wwl_0_21 rwl_0_38 rwl_0_12 write_bl_0_24 read_bl_0_3
+ read_bl_0_1 read_bl_0_61 wwl_0_22 read_bl_0_13 rwl_0_48 rwl_1_54 read_bl_0_11 write_bl_0_35
+ read_bl_0_33 rwl_0_37 wwl_0_49 read_bl_1_10 rwl_1_25 write_bl_0_23 read_bl_0_40
+ read_bl_1_0 rwl_0_33 rwl_1_0 read_bl_1_24 rwl_0_25 rwl_1_31 read_bl_1_22 read_bl_1_39
+ write_bl_0_18 read_bl_1_37 read_bl_1_60 write_bl_0_33 rwl_1_49 read_bl_1_31 wwl_0_61
+ rwl_1_41 rwl_1_53 read_bl_1_63 read_bl_1_58 rwl_0_52 write_bl_0_54 write_bl_0_25
+ read_bl_0_5 rwl_1_2 rwl_1_4 write_bl_0_1 read_bl_0_15 wwl_0_7 rwl_0_10 read_bl_1_41
+ read_bl_0_30 write_bl_0_59 read_bl_1_17 rwl_1_40 rwl_1_26 wwl_0_38 rwl_1_18 read_bl_1_27
+ rwl_1_1 rwl_1_45 rwl_1_23 wwl_0_31 write_bl_0_13 rwl_0_35 read_bl_1_2 rwl_0_13 rwl_1_3
+ wwl_0_53 rwl_1_22 read_bl_0_32 wwl_0_8 read_bl_0_56 wwl_0_30 wwl_0_63 wwl_0_52 read_bl_1_53
+ read_bl_0_43 rwl_0_55 rwl_1_30 rwl_1_8 write_bl_0_40 rwl_1_44 wwl_0_13 rwl_0_32
+ rwl_1_7 wwl_0_29 wwl_0_15 rwl_0_41 rwl_0_16 wwl_0_34 wwl_0_14 rwl_0_18 rwl_0_54
+ wwl_0_11 rwl_1_6 rwl_0_17 rwl_0_53 rwl_0_14 rwl_1_52 rwl_0_59 rwl_0_5 rwl_1_51 rwl_1_63
+ rwl_1_29 rwl_1_28 rwl_1_14 rwl_1_11 wwl_0_23 rwl_0_42 rwl_1_17 read_bl_1_43 wwl_0_39
+ wwl_0_25 rwl_0_51 rwl_0_29 wwl_0_0 rwl_0_26 wwl_0_2 wwl_0_44 rwl_0_63 rwl_1_61 rwl_1_38
+ wwl_0_36 rwl_0_39 rwl_0_36 wwl_0_12 rwl_0_15 rwl_1_48 wwl_0_60 gnd
Xcell_2r1w_1924 vdd_uq28 gnd read_bl_0_33 read_bl_1_33 write_bl_0_33 wwl_0_59 rwl_1_59
+ rwl_0_59 cell_2r1w
Xcell_2r1w_1935 vdd_uq23 gnd read_bl_0_33 read_bl_1_33 write_bl_0_33 wwl_0_48 rwl_1_48
+ rwl_0_48 cell_2r1w
Xcell_2r1w_1946 vdd_uq17 gnd read_bl_0_33 read_bl_1_33 write_bl_0_33 wwl_0_37 rwl_1_37
+ rwl_0_37 cell_2r1w
Xcell_2r1w_2658 vdd_uq13 gnd read_bl_0_22 read_bl_1_22 write_bl_0_22 wwl_0_29 rwl_1_29
+ rwl_0_29 cell_2r1w
Xcell_2r1w_1957 vdd_uq12 gnd read_bl_0_33 read_bl_1_33 write_bl_0_33 wwl_0_26 rwl_1_26
+ rwl_0_26 cell_2r1w
Xcell_2r1w_1979 vdd_uq1 gnd read_bl_0_33 read_bl_1_33 write_bl_0_33 wwl_0_4 rwl_1_4
+ rwl_0_4 cell_2r1w
Xcell_2r1w_1968 vdd_uq6 gnd read_bl_0_33 read_bl_1_33 write_bl_0_33 wwl_0_15 rwl_1_15
+ rwl_0_15 cell_2r1w
Xcell_2r1w_2669 vdd_uq8 gnd read_bl_0_22 read_bl_1_22 write_bl_0_22 wwl_0_18 rwl_1_18
+ rwl_0_18 cell_2r1w
Xcell_2r1w_3860 vdd_uq20 gnd read_bl_0_3 read_bl_1_3 write_bl_0_3 wwl_0_43 rwl_1_43
+ rwl_0_43 cell_2r1w
Xcell_2r1w_3871 vdd_uq15 gnd read_bl_0_3 read_bl_1_3 write_bl_0_3 wwl_0_32 rwl_1_32
+ rwl_0_32 cell_2r1w
Xcell_2r1w_3893 vdd_uq4 gnd read_bl_0_3 read_bl_1_3 write_bl_0_3 wwl_0_10 rwl_1_10
+ rwl_0_10 cell_2r1w
Xcell_2r1w_3882 vdd_uq9 gnd read_bl_0_3 read_bl_1_3 write_bl_0_3 wwl_0_21 rwl_1_21
+ rwl_0_21 cell_2r1w
Xcell_2r1w_458 vdd_uq25 gnd read_bl_0_56 read_bl_1_56 write_bl_0_56 wwl_0_53 rwl_1_53
+ rwl_0_53 cell_2r1w
Xcell_2r1w_403 vdd_uq21 gnd read_bl_0_57 read_bl_1_57 write_bl_0_57 wwl_0_44 rwl_1_44
+ rwl_0_44 cell_2r1w
Xcell_2r1w_469 vdd_uq20 gnd read_bl_0_56 read_bl_1_56 write_bl_0_56 wwl_0_42 rwl_1_42
+ rwl_0_42 cell_2r1w
Xcell_2r1w_414 vdd_uq15 gnd read_bl_0_57 read_bl_1_57 write_bl_0_57 wwl_0_33 rwl_1_33
+ rwl_0_33 cell_2r1w
Xcell_2r1w_447 vdd_uq0 gnd read_bl_0_57 read_bl_1_57 write_bl_0_57 wwl_0_0 rwl_1_0
+ rwl_0_0 cell_2r1w
Xcell_2r1w_1209 vdd_uq2 gnd read_bl_0_45 read_bl_1_45 write_bl_0_45 wwl_0_6 rwl_1_6
+ rwl_0_6 cell_2r1w
Xcell_2r1w_436 vdd_uq4 gnd read_bl_0_57 read_bl_1_57 write_bl_0_57 wwl_0_11 rwl_1_11
+ rwl_0_11 cell_2r1w
Xcell_2r1w_425 vdd_uq10 gnd read_bl_0_57 read_bl_1_57 write_bl_0_57 wwl_0_22 rwl_1_22
+ rwl_0_22 cell_2r1w
Xcell_2r1w_3101 vdd_uq16 gnd read_bl_0_15 read_bl_1_15 write_bl_0_15 wwl_0_34 rwl_1_34
+ rwl_0_34 cell_2r1w
Xcell_2r1w_2433 vdd_uq30 gnd read_bl_0_25 read_bl_1_25 write_bl_0_25 wwl_0_62 rwl_1_62
+ rwl_0_62 cell_2r1w
Xcell_2r1w_2499 vdd_uq29 gnd read_bl_0_24 read_bl_1_24 write_bl_0_24 wwl_0_60 rwl_1_60
+ rwl_0_60 cell_2r1w
Xcell_2r1w_1732 vdd_uq28 gnd read_bl_0_36 read_bl_1_36 write_bl_0_36 wwl_0_59 rwl_1_59
+ rwl_0_59 cell_2r1w
Xcell_2r1w_3145 vdd_uq26 gnd read_bl_0_14 read_bl_1_14 write_bl_0_14 wwl_0_54 rwl_1_54
+ rwl_0_54 cell_2r1w
Xcell_2r1w_2444 vdd_uq24 gnd read_bl_0_25 read_bl_1_25 write_bl_0_25 wwl_0_51 rwl_1_51
+ rwl_0_51 cell_2r1w
Xcell_2r1w_1743 vdd_uq23 gnd read_bl_0_36 read_bl_1_36 write_bl_0_36 wwl_0_48 rwl_1_48
+ rwl_0_48 cell_2r1w
Xcell_2r1w_3156 vdd_uq20 gnd read_bl_0_14 read_bl_1_14 write_bl_0_14 wwl_0_43 rwl_1_43
+ rwl_0_43 cell_2r1w
Xcell_2r1w_2455 vdd_uq19 gnd read_bl_0_25 read_bl_1_25 write_bl_0_25 wwl_0_40 rwl_1_40
+ rwl_0_40 cell_2r1w
Xcell_2r1w_1754 vdd_uq17 gnd read_bl_0_36 read_bl_1_36 write_bl_0_36 wwl_0_37 rwl_1_37
+ rwl_0_37 cell_2r1w
Xcell_2r1w_3167 vdd_uq15 gnd read_bl_0_14 read_bl_1_14 write_bl_0_14 wwl_0_32 rwl_1_32
+ rwl_0_32 cell_2r1w
Xcell_2r1w_2400 vdd_uq14 gnd read_bl_0_26 read_bl_1_26 write_bl_0_26 wwl_0_31 rwl_1_31
+ rwl_0_31 cell_2r1w
Xcell_2r1w_2466 vdd_uq13 gnd read_bl_0_25 read_bl_1_25 write_bl_0_25 wwl_0_29 rwl_1_29
+ rwl_0_29 cell_2r1w
Xcell_2r1w_3134 vdd_uq0 gnd read_bl_0_15 read_bl_1_15 write_bl_0_15 wwl_0_1 rwl_1_1
+ rwl_0_1 cell_2r1w
Xcell_2r1w_1721 vdd_uq2 gnd read_bl_0_37 read_bl_1_37 write_bl_0_37 wwl_0_6 rwl_1_6
+ rwl_0_6 cell_2r1w
Xcell_2r1w_2488 vdd_uq2 gnd read_bl_0_25 read_bl_1_25 write_bl_0_25 wwl_0_7 rwl_1_7
+ rwl_0_7 cell_2r1w
Xcell_2r1w_2422 vdd_uq3 gnd read_bl_0_26 read_bl_1_26 write_bl_0_26 wwl_0_9 rwl_1_9
+ rwl_0_9 cell_2r1w
Xcell_2r1w_3189 vdd_uq4 gnd read_bl_0_14 read_bl_1_14 write_bl_0_14 wwl_0_10 rwl_1_10
+ rwl_0_10 cell_2r1w
Xcell_2r1w_3123 vdd_uq5 gnd read_bl_0_15 read_bl_1_15 write_bl_0_15 wwl_0_12 rwl_1_12
+ rwl_0_12 cell_2r1w
Xcell_2r1w_1710 vdd_uq7 gnd read_bl_0_37 read_bl_1_37 write_bl_0_37 wwl_0_17 rwl_1_17
+ rwl_0_17 cell_2r1w
Xcell_2r1w_2477 vdd_uq8 gnd read_bl_0_25 read_bl_1_25 write_bl_0_25 wwl_0_18 rwl_1_18
+ rwl_0_18 cell_2r1w
Xcell_2r1w_2411 vdd_uq9 gnd read_bl_0_26 read_bl_1_26 write_bl_0_26 wwl_0_20 rwl_1_20
+ rwl_0_20 cell_2r1w
Xcell_2r1w_3178 vdd_uq9 gnd read_bl_0_14 read_bl_1_14 write_bl_0_14 wwl_0_21 rwl_1_21
+ rwl_0_21 cell_2r1w
Xcell_2r1w_3112 vdd_uq10 gnd read_bl_0_15 read_bl_1_15 write_bl_0_15 wwl_0_23 rwl_1_23
+ rwl_0_23 cell_2r1w
Xcell_2r1w_1798 vdd_uq27 gnd read_bl_0_35 read_bl_1_35 write_bl_0_35 wwl_0_57 rwl_1_57
+ rwl_0_57 cell_2r1w
Xcell_2r1w_970 vdd_uq25 gnd read_bl_0_48 read_bl_1_48 write_bl_0_48 wwl_0_53 rwl_1_53
+ rwl_0_53 cell_2r1w
Xcell_2r1w_981 vdd_uq20 gnd read_bl_0_48 read_bl_1_48 write_bl_0_48 wwl_0_42 rwl_1_42
+ rwl_0_42 cell_2r1w
Xcell_2r1w_992 vdd_uq14 gnd read_bl_0_48 read_bl_1_48 write_bl_0_48 wwl_0_31 rwl_1_31
+ rwl_0_31 cell_2r1w
Xcell_2r1w_1765 vdd_uq12 gnd read_bl_0_36 read_bl_1_36 write_bl_0_36 wwl_0_26 rwl_1_26
+ rwl_0_26 cell_2r1w
Xcell_2r1w_1787 vdd_uq1 gnd read_bl_0_36 read_bl_1_36 write_bl_0_36 wwl_0_4 rwl_1_4
+ rwl_0_4 cell_2r1w
Xcell_2r1w_1776 vdd_uq6 gnd read_bl_0_36 read_bl_1_36 write_bl_0_36 wwl_0_15 rwl_1_15
+ rwl_0_15 cell_2r1w
Xcell_2r1w_3690 vdd_uq9 gnd read_bl_0_6 read_bl_1_6 write_bl_0_6 wwl_0_21 rwl_1_21
+ rwl_0_21 cell_2r1w
Xcell_2r1w_71 vdd_uq27 gnd read_bl_0_62 read_bl_1_62 write_bl_0_62 wwl_0_56 rwl_1_56
+ rwl_0_56 cell_2r1w
Xcell_2r1w_82 vdd_uq21 gnd read_bl_0_62 read_bl_1_62 write_bl_0_62 wwl_0_45 rwl_1_45
+ rwl_0_45 cell_2r1w
Xcell_2r1w_60 vdd gnd read_bl_0_63 read_bl_1_63 write_bl_0_63 wwl_0_3 rwl_1_3 rwl_0_3
+ cell_2r1w
Xcell_2r1w_93 vdd_uq16 gnd read_bl_0_62 read_bl_1_62 write_bl_0_62 wwl_0_34 rwl_1_34
+ rwl_0_34 cell_2r1w
Xcell_2r1w_1028 vdd_uq28 gnd read_bl_0_47 read_bl_1_47 write_bl_0_47 wwl_0_59 rwl_1_59
+ rwl_0_59 cell_2r1w
Xcell_2r1w_200 vdd_uq26 gnd read_bl_0_60 read_bl_1_60 write_bl_0_60 wwl_0_55 rwl_1_55
+ rwl_0_55 cell_2r1w
Xcell_2r1w_1039 vdd_uq23 gnd read_bl_0_47 read_bl_1_47 write_bl_0_47 wwl_0_48 rwl_1_48
+ rwl_0_48 cell_2r1w
Xcell_2r1w_211 vdd_uq21 gnd read_bl_0_60 read_bl_1_60 write_bl_0_60 wwl_0_44 rwl_1_44
+ rwl_0_44 cell_2r1w
Xcell_2r1w_1017 vdd_uq2 gnd read_bl_0_48 read_bl_1_48 write_bl_0_48 wwl_0_6 rwl_1_6
+ rwl_0_6 cell_2r1w
Xcell_2r1w_1006 vdd_uq7 gnd read_bl_0_48 read_bl_1_48 write_bl_0_48 wwl_0_17 rwl_1_17
+ rwl_0_17 cell_2r1w
Xcell_2r1w_266 vdd_uq25 gnd read_bl_0_59 read_bl_1_59 write_bl_0_59 wwl_0_53 rwl_1_53
+ rwl_0_53 cell_2r1w
Xcell_2r1w_277 vdd_uq20 gnd read_bl_0_59 read_bl_1_59 write_bl_0_59 wwl_0_42 rwl_1_42
+ rwl_0_42 cell_2r1w
Xcell_2r1w_222 vdd_uq15 gnd read_bl_0_60 read_bl_1_60 write_bl_0_60 wwl_0_33 rwl_1_33
+ rwl_0_33 cell_2r1w
Xcell_2r1w_288 vdd_uq14 gnd read_bl_0_59 read_bl_1_59 write_bl_0_59 wwl_0_31 rwl_1_31
+ rwl_0_31 cell_2r1w
Xcell_2r1w_255 vdd_uq0 gnd read_bl_0_60 read_bl_1_60 write_bl_0_60 wwl_0_0 rwl_1_0
+ rwl_0_0 cell_2r1w
Xcell_2r1w_244 vdd_uq4 gnd read_bl_0_60 read_bl_1_60 write_bl_0_60 wwl_0_11 rwl_1_11
+ rwl_0_11 cell_2r1w
Xcell_2r1w_299 vdd_uq9 gnd read_bl_0_59 read_bl_1_59 write_bl_0_59 wwl_0_20 rwl_1_20
+ rwl_0_20 cell_2r1w
Xcell_2r1w_233 vdd_uq10 gnd read_bl_0_60 read_bl_1_60 write_bl_0_60 wwl_0_22 rwl_1_22
+ rwl_0_22 cell_2r1w
Xcell_2r1w_2241 vdd_uq30 gnd read_bl_0_28 read_bl_1_28 write_bl_0_28 wwl_0_62 rwl_1_62
+ rwl_0_62 cell_2r1w
Xcell_2r1w_1540 vdd_uq28 gnd read_bl_0_39 read_bl_1_39 write_bl_0_39 wwl_0_59 rwl_1_59
+ rwl_0_59 cell_2r1w
Xcell_2r1w_2252 vdd_uq24 gnd read_bl_0_28 read_bl_1_28 write_bl_0_28 wwl_0_51 rwl_1_51
+ rwl_0_51 cell_2r1w
Xcell_2r1w_1551 vdd_uq23 gnd read_bl_0_39 read_bl_1_39 write_bl_0_39 wwl_0_48 rwl_1_48
+ rwl_0_48 cell_2r1w
Xcell_2r1w_2263 vdd_uq19 gnd read_bl_0_28 read_bl_1_28 write_bl_0_28 wwl_0_40 rwl_1_40
+ rwl_0_40 cell_2r1w
Xcell_2r1w_1562 vdd_uq17 gnd read_bl_0_39 read_bl_1_39 write_bl_0_39 wwl_0_37 rwl_1_37
+ rwl_0_37 cell_2r1w
Xcell_2r1w_2274 vdd_uq13 gnd read_bl_0_28 read_bl_1_28 write_bl_0_28 wwl_0_29 rwl_1_29
+ rwl_0_29 cell_2r1w
Xcell_2r1w_1573 vdd_uq12 gnd read_bl_0_39 read_bl_1_39 write_bl_0_39 wwl_0_26 rwl_1_26
+ rwl_0_26 cell_2r1w
Xcell_2r1w_1595 vdd_uq1 gnd read_bl_0_39 read_bl_1_39 write_bl_0_39 wwl_0_4 rwl_1_4
+ rwl_0_4 cell_2r1w
Xcell_2r1w_2296 vdd_uq2 gnd read_bl_0_28 read_bl_1_28 write_bl_0_28 wwl_0_7 rwl_1_7
+ rwl_0_7 cell_2r1w
Xcell_2r1w_2230 vdd_uq3 gnd read_bl_0_29 read_bl_1_29 write_bl_0_29 wwl_0_9 rwl_1_9
+ rwl_0_9 cell_2r1w
Xcell_2r1w_1584 vdd_uq6 gnd read_bl_0_39 read_bl_1_39 write_bl_0_39 wwl_0_15 rwl_1_15
+ rwl_0_15 cell_2r1w
Xcell_2r1w_2285 vdd_uq8 gnd read_bl_0_28 read_bl_1_28 write_bl_0_28 wwl_0_18 rwl_1_18
+ rwl_0_18 cell_2r1w
Xcell_2r1w_2060 vdd_uq24 gnd read_bl_0_31 read_bl_1_31 write_bl_0_31 wwl_0_51 rwl_1_51
+ rwl_0_51 cell_2r1w
Xcell_2r1w_2071 vdd_uq19 gnd read_bl_0_31 read_bl_1_31 write_bl_0_31 wwl_0_40 rwl_1_40
+ rwl_0_40 cell_2r1w
Xcell_2r1w_1370 vdd_uq17 gnd read_bl_0_42 read_bl_1_42 write_bl_0_42 wwl_0_37 rwl_1_37
+ rwl_0_37 cell_2r1w
Xcell_2r1w_2082 vdd_uq13 gnd read_bl_0_31 read_bl_1_31 write_bl_0_31 wwl_0_29 rwl_1_29
+ rwl_0_29 cell_2r1w
Xcell_2r1w_1381 vdd_uq12 gnd read_bl_0_42 read_bl_1_42 write_bl_0_42 wwl_0_26 rwl_1_26
+ rwl_0_26 cell_2r1w
Xcell_2r1w_1392 vdd_uq6 gnd read_bl_0_42 read_bl_1_42 write_bl_0_42 wwl_0_15 rwl_1_15
+ rwl_0_15 cell_2r1w
Xcell_2r1w_2093 vdd_uq8 gnd read_bl_0_31 read_bl_1_31 write_bl_0_31 wwl_0_18 rwl_1_18
+ rwl_0_18 cell_2r1w
Xcell_2r1w_2818 vdd_uq29 gnd read_bl_0_19 read_bl_1_19 write_bl_0_19 wwl_0_61 rwl_1_61
+ rwl_0_61 cell_2r1w
Xcell_2r1w_2829 vdd_uq24 gnd read_bl_0_19 read_bl_1_19 write_bl_0_19 wwl_0_50 rwl_1_50
+ rwl_0_50 cell_2r1w
Xcell_2r1w_3519 vdd_uq0 gnd read_bl_0_9 read_bl_1_9 write_bl_0_9 wwl_0_0 rwl_1_0 rwl_0_0
+ cell_2r1w
Xcell_2r1w_2807 vdd_uq3 gnd read_bl_0_20 read_bl_1_20 write_bl_0_20 wwl_0_8 rwl_1_8
+ rwl_0_8 cell_2r1w
Xcell_2r1w_3508 vdd_uq4 gnd read_bl_0_9 read_bl_1_9 write_bl_0_9 wwl_0_11 rwl_1_11
+ rwl_0_11 cell_2r1w
Xcell_2r1w_607 vdd_uq15 gnd read_bl_0_54 read_bl_1_54 write_bl_0_54 wwl_0_32 rwl_1_32
+ rwl_0_32 cell_2r1w
Xcell_2r1w_629 vdd_uq4 gnd read_bl_0_54 read_bl_1_54 write_bl_0_54 wwl_0_10 rwl_1_10
+ rwl_0_10 cell_2r1w
Xcell_2r1w_618 vdd_uq9 gnd read_bl_0_54 read_bl_1_54 write_bl_0_54 wwl_0_21 rwl_1_21
+ rwl_0_21 cell_2r1w
Xcell_2r1w_4006 vdd_uq11 gnd read_bl_0_1 read_bl_1_1 write_bl_0_1 wwl_0_25 rwl_1_25
+ rwl_0_25 cell_2r1w
Xcell_2r1w_4028 vdd gnd read_bl_0_1 read_bl_1_1 write_bl_0_1 wwl_0_3 rwl_1_3 rwl_0_3
+ cell_2r1w
Xcell_2r1w_4017 vdd_uq6 gnd read_bl_0_1 read_bl_1_1 write_bl_0_1 wwl_0_14 rwl_1_14
+ rwl_0_14 cell_2r1w
Xcell_2r1w_2626 vdd_uq29 gnd read_bl_0_22 read_bl_1_22 write_bl_0_22 wwl_0_61 rwl_1_61
+ rwl_0_61 cell_2r1w
Xcell_2r1w_1925 vdd_uq28 gnd read_bl_0_33 read_bl_1_33 write_bl_0_33 wwl_0_58 rwl_1_58
+ rwl_0_58 cell_2r1w
Xcell_2r1w_4039 vdd_uq27 gnd read_bl_0_0 read_bl_1_0 write_bl_0_0 wwl_0_56 rwl_1_56
+ rwl_0_56 cell_2r1w
Xcell_2r1w_3338 vdd_uq25 gnd read_bl_0_11 read_bl_1_11 write_bl_0_11 wwl_0_53 rwl_1_53
+ rwl_0_53 cell_2r1w
Xcell_2r1w_2637 vdd_uq24 gnd read_bl_0_22 read_bl_1_22 write_bl_0_22 wwl_0_50 rwl_1_50
+ rwl_0_50 cell_2r1w
Xcell_2r1w_1936 vdd_uq22 gnd read_bl_0_33 read_bl_1_33 write_bl_0_33 wwl_0_47 rwl_1_47
+ rwl_0_47 cell_2r1w
Xcell_2r1w_3349 vdd_uq20 gnd read_bl_0_11 read_bl_1_11 write_bl_0_11 wwl_0_42 rwl_1_42
+ rwl_0_42 cell_2r1w
Xcell_2r1w_2648 vdd_uq18 gnd read_bl_0_22 read_bl_1_22 write_bl_0_22 wwl_0_39 rwl_1_39
+ rwl_0_39 cell_2r1w
Xcell_2r1w_2659 vdd_uq13 gnd read_bl_0_22 read_bl_1_22 write_bl_0_22 wwl_0_28 rwl_1_28
+ rwl_0_28 cell_2r1w
Xcell_2r1w_1914 vdd_uq1 gnd read_bl_0_34 read_bl_1_34 write_bl_0_34 wwl_0_5 rwl_1_5
+ rwl_0_5 cell_2r1w
Xcell_2r1w_3327 vdd_uq0 gnd read_bl_0_12 read_bl_1_12 write_bl_0_12 wwl_0_0 rwl_1_0
+ rwl_0_0 cell_2r1w
Xcell_2r1w_2615 vdd_uq3 gnd read_bl_0_23 read_bl_1_23 write_bl_0_23 wwl_0_8 rwl_1_8
+ rwl_0_8 cell_2r1w
Xcell_2r1w_3316 vdd_uq4 gnd read_bl_0_12 read_bl_1_12 write_bl_0_12 wwl_0_11 rwl_1_11
+ rwl_0_11 cell_2r1w
Xcell_2r1w_1903 vdd_uq7 gnd read_bl_0_34 read_bl_1_34 write_bl_0_34 wwl_0_16 rwl_1_16
+ rwl_0_16 cell_2r1w
Xcell_2r1w_2604 vdd_uq8 gnd read_bl_0_23 read_bl_1_23 write_bl_0_23 wwl_0_19 rwl_1_19
+ rwl_0_19 cell_2r1w
Xcell_2r1w_3305 vdd_uq10 gnd read_bl_0_12 read_bl_1_12 write_bl_0_12 wwl_0_22 rwl_1_22
+ rwl_0_22 cell_2r1w
Xcell_2r1w_1947 vdd_uq17 gnd read_bl_0_33 read_bl_1_33 write_bl_0_33 wwl_0_36 rwl_1_36
+ rwl_0_36 cell_2r1w
Xcell_2r1w_1958 vdd_uq11 gnd read_bl_0_33 read_bl_1_33 write_bl_0_33 wwl_0_25 rwl_1_25
+ rwl_0_25 cell_2r1w
Xcell_2r1w_1969 vdd_uq6 gnd read_bl_0_33 read_bl_1_33 write_bl_0_33 wwl_0_14 rwl_1_14
+ rwl_0_14 cell_2r1w
Xcell_2r1w_3850 vdd_uq25 gnd read_bl_0_3 read_bl_1_3 write_bl_0_3 wwl_0_53 rwl_1_53
+ rwl_0_53 cell_2r1w
Xcell_2r1w_3861 vdd_uq20 gnd read_bl_0_3 read_bl_1_3 write_bl_0_3 wwl_0_42 rwl_1_42
+ rwl_0_42 cell_2r1w
Xcell_2r1w_3872 vdd_uq14 gnd read_bl_0_3 read_bl_1_3 write_bl_0_3 wwl_0_31 rwl_1_31
+ rwl_0_31 cell_2r1w
Xcell_2r1w_3894 vdd_uq3 gnd read_bl_0_3 read_bl_1_3 write_bl_0_3 wwl_0_9 rwl_1_9 rwl_0_9
+ cell_2r1w
Xcell_2r1w_3883 vdd_uq9 gnd read_bl_0_3 read_bl_1_3 write_bl_0_3 wwl_0_20 rwl_1_20
+ rwl_0_20 cell_2r1w
Xcell_2r1w_448 vdd_uq30 gnd read_bl_0_56 read_bl_1_56 write_bl_0_56 wwl_0_63 rwl_1_63
+ rwl_0_63 cell_2r1w
Xcell_2r1w_459 vdd_uq25 gnd read_bl_0_56 read_bl_1_56 write_bl_0_56 wwl_0_52 rwl_1_52
+ rwl_0_52 cell_2r1w
Xcell_2r1w_404 vdd_uq20 gnd read_bl_0_57 read_bl_1_57 write_bl_0_57 wwl_0_43 rwl_1_43
+ rwl_0_43 cell_2r1w
Xcell_2r1w_415 vdd_uq15 gnd read_bl_0_57 read_bl_1_57 write_bl_0_57 wwl_0_32 rwl_1_32
+ rwl_0_32 cell_2r1w
Xcell_2r1w_437 vdd_uq4 gnd read_bl_0_57 read_bl_1_57 write_bl_0_57 wwl_0_10 rwl_1_10
+ rwl_0_10 cell_2r1w
Xcell_2r1w_426 vdd_uq9 gnd read_bl_0_57 read_bl_1_57 write_bl_0_57 wwl_0_21 rwl_1_21
+ rwl_0_21 cell_2r1w
Xcell_2r1w_3102 vdd_uq15 gnd read_bl_0_15 read_bl_1_15 write_bl_0_15 wwl_0_33 rwl_1_33
+ rwl_0_33 cell_2r1w
Xcell_2r1w_3124 vdd_uq4 gnd read_bl_0_15 read_bl_1_15 write_bl_0_15 wwl_0_11 rwl_1_11
+ rwl_0_11 cell_2r1w
Xcell_2r1w_3113 vdd_uq10 gnd read_bl_0_15 read_bl_1_15 write_bl_0_15 wwl_0_22 rwl_1_22
+ rwl_0_22 cell_2r1w
Xcell_2r1w_2434 vdd_uq29 gnd read_bl_0_25 read_bl_1_25 write_bl_0_25 wwl_0_61 rwl_1_61
+ rwl_0_61 cell_2r1w
Xcell_2r1w_1733 vdd_uq28 gnd read_bl_0_36 read_bl_1_36 write_bl_0_36 wwl_0_58 rwl_1_58
+ rwl_0_58 cell_2r1w
Xcell_2r1w_3146 vdd_uq25 gnd read_bl_0_14 read_bl_1_14 write_bl_0_14 wwl_0_53 rwl_1_53
+ rwl_0_53 cell_2r1w
Xcell_2r1w_2445 vdd_uq24 gnd read_bl_0_25 read_bl_1_25 write_bl_0_25 wwl_0_50 rwl_1_50
+ rwl_0_50 cell_2r1w
Xcell_2r1w_1744 vdd_uq22 gnd read_bl_0_36 read_bl_1_36 write_bl_0_36 wwl_0_47 rwl_1_47
+ rwl_0_47 cell_2r1w
Xcell_2r1w_3157 vdd_uq20 gnd read_bl_0_14 read_bl_1_14 write_bl_0_14 wwl_0_42 rwl_1_42
+ rwl_0_42 cell_2r1w
Xcell_2r1w_2456 vdd_uq18 gnd read_bl_0_25 read_bl_1_25 write_bl_0_25 wwl_0_39 rwl_1_39
+ rwl_0_39 cell_2r1w
Xcell_2r1w_1755 vdd_uq17 gnd read_bl_0_36 read_bl_1_36 write_bl_0_36 wwl_0_36 rwl_1_36
+ rwl_0_36 cell_2r1w
Xcell_2r1w_3168 vdd_uq14 gnd read_bl_0_14 read_bl_1_14 write_bl_0_14 wwl_0_31 rwl_1_31
+ rwl_0_31 cell_2r1w
Xcell_2r1w_2401 vdd_uq14 gnd read_bl_0_26 read_bl_1_26 write_bl_0_26 wwl_0_30 rwl_1_30
+ rwl_0_30 cell_2r1w
Xcell_2r1w_1700 vdd_uq12 gnd read_bl_0_37 read_bl_1_37 write_bl_0_37 wwl_0_27 rwl_1_27
+ rwl_0_27 cell_2r1w
Xcell_2r1w_2467 vdd_uq13 gnd read_bl_0_25 read_bl_1_25 write_bl_0_25 wwl_0_28 rwl_1_28
+ rwl_0_28 cell_2r1w
Xcell_2r1w_1766 vdd_uq11 gnd read_bl_0_36 read_bl_1_36 write_bl_0_36 wwl_0_25 rwl_1_25
+ rwl_0_25 cell_2r1w
Xcell_2r1w_1722 vdd_uq1 gnd read_bl_0_37 read_bl_1_37 write_bl_0_37 wwl_0_5 rwl_1_5
+ rwl_0_5 cell_2r1w
Xcell_2r1w_1788 vdd gnd read_bl_0_36 read_bl_1_36 write_bl_0_36 wwl_0_3 rwl_1_3 rwl_0_3
+ cell_2r1w
Xcell_2r1w_3135 vdd_uq0 gnd read_bl_0_15 read_bl_1_15 write_bl_0_15 wwl_0_0 rwl_1_0
+ rwl_0_0 cell_2r1w
Xcell_2r1w_2489 vdd_uq2 gnd read_bl_0_25 read_bl_1_25 write_bl_0_25 wwl_0_6 rwl_1_6
+ rwl_0_6 cell_2r1w
Xcell_2r1w_2423 vdd_uq3 gnd read_bl_0_26 read_bl_1_26 write_bl_0_26 wwl_0_8 rwl_1_8
+ rwl_0_8 cell_2r1w
Xcell_2r1w_1777 vdd_uq6 gnd read_bl_0_36 read_bl_1_36 write_bl_0_36 wwl_0_14 rwl_1_14
+ rwl_0_14 cell_2r1w
Xcell_2r1w_1711 vdd_uq7 gnd read_bl_0_37 read_bl_1_37 write_bl_0_37 wwl_0_16 rwl_1_16
+ rwl_0_16 cell_2r1w
Xcell_2r1w_2478 vdd_uq7 gnd read_bl_0_25 read_bl_1_25 write_bl_0_25 wwl_0_17 rwl_1_17
+ rwl_0_17 cell_2r1w
Xcell_2r1w_2412 vdd_uq8 gnd read_bl_0_26 read_bl_1_26 write_bl_0_26 wwl_0_19 rwl_1_19
+ rwl_0_19 cell_2r1w
Xcell_2r1w_3179 vdd_uq9 gnd read_bl_0_14 read_bl_1_14 write_bl_0_14 wwl_0_20 rwl_1_20
+ rwl_0_20 cell_2r1w
Xcell_2r1w_960 vdd_uq30 gnd read_bl_0_48 read_bl_1_48 write_bl_0_48 wwl_0_63 rwl_1_63
+ rwl_0_63 cell_2r1w
Xcell_2r1w_1799 vdd_uq27 gnd read_bl_0_35 read_bl_1_35 write_bl_0_35 wwl_0_56 rwl_1_56
+ rwl_0_56 cell_2r1w
Xcell_2r1w_971 vdd_uq25 gnd read_bl_0_48 read_bl_1_48 write_bl_0_48 wwl_0_52 rwl_1_52
+ rwl_0_52 cell_2r1w
Xcell_2r1w_982 vdd_uq19 gnd read_bl_0_48 read_bl_1_48 write_bl_0_48 wwl_0_41 rwl_1_41
+ rwl_0_41 cell_2r1w
Xcell_2r1w_993 vdd_uq14 gnd read_bl_0_48 read_bl_1_48 write_bl_0_48 wwl_0_30 rwl_1_30
+ rwl_0_30 cell_2r1w
Xcell_2r1w_3680 vdd_uq14 gnd read_bl_0_6 read_bl_1_6 write_bl_0_6 wwl_0_31 rwl_1_31
+ rwl_0_31 cell_2r1w
Xcell_2r1w_2990 vdd_uq7 gnd read_bl_0_17 read_bl_1_17 write_bl_0_17 wwl_0_17 rwl_1_17
+ rwl_0_17 cell_2r1w
Xcell_2r1w_3691 vdd_uq9 gnd read_bl_0_6 read_bl_1_6 write_bl_0_6 wwl_0_20 rwl_1_20
+ rwl_0_20 cell_2r1w
Xcell_2r1w_72 vdd_uq26 gnd read_bl_0_62 read_bl_1_62 write_bl_0_62 wwl_0_55 rwl_1_55
+ rwl_0_55 cell_2r1w
Xcell_2r1w_83 vdd_uq21 gnd read_bl_0_62 read_bl_1_62 write_bl_0_62 wwl_0_44 rwl_1_44
+ rwl_0_44 cell_2r1w
Xcell_2r1w_94 vdd_uq15 gnd read_bl_0_62 read_bl_1_62 write_bl_0_62 wwl_0_33 rwl_1_33
+ rwl_0_33 cell_2r1w
Xcell_2r1w_61 vdd gnd read_bl_0_63 read_bl_1_63 write_bl_0_63 wwl_0_2 rwl_1_2 rwl_0_2
+ cell_2r1w
Xcell_2r1w_50 vdd_uq5 gnd read_bl_0_63 read_bl_1_63 write_bl_0_63 wwl_0_13 rwl_1_13
+ rwl_0_13 cell_2r1w
Xcell_2r1w_1029 vdd_uq28 gnd read_bl_0_47 read_bl_1_47 write_bl_0_47 wwl_0_58 rwl_1_58
+ rwl_0_58 cell_2r1w
Xcell_2r1w_201 vdd_uq26 gnd read_bl_0_60 read_bl_1_60 write_bl_0_60 wwl_0_54 rwl_1_54
+ rwl_0_54 cell_2r1w
Xcell_2r1w_212 vdd_uq20 gnd read_bl_0_60 read_bl_1_60 write_bl_0_60 wwl_0_43 rwl_1_43
+ rwl_0_43 cell_2r1w
Xcell_2r1w_223 vdd_uq15 gnd read_bl_0_60 read_bl_1_60 write_bl_0_60 wwl_0_32 rwl_1_32
+ rwl_0_32 cell_2r1w
Xcell_2r1w_1018 vdd_uq1 gnd read_bl_0_48 read_bl_1_48 write_bl_0_48 wwl_0_5 rwl_1_5
+ rwl_0_5 cell_2r1w
Xcell_2r1w_245 vdd_uq4 gnd read_bl_0_60 read_bl_1_60 write_bl_0_60 wwl_0_10 rwl_1_10
+ rwl_0_10 cell_2r1w
Xcell_2r1w_1007 vdd_uq7 gnd read_bl_0_48 read_bl_1_48 write_bl_0_48 wwl_0_16 rwl_1_16
+ rwl_0_16 cell_2r1w
Xcell_2r1w_234 vdd_uq9 gnd read_bl_0_60 read_bl_1_60 write_bl_0_60 wwl_0_21 rwl_1_21
+ rwl_0_21 cell_2r1w
Xcell_2r1w_256 vdd_uq30 gnd read_bl_0_59 read_bl_1_59 write_bl_0_59 wwl_0_63 rwl_1_63
+ rwl_0_63 cell_2r1w
Xcell_2r1w_267 vdd_uq25 gnd read_bl_0_59 read_bl_1_59 write_bl_0_59 wwl_0_52 rwl_1_52
+ rwl_0_52 cell_2r1w
Xcell_2r1w_278 vdd_uq19 gnd read_bl_0_59 read_bl_1_59 write_bl_0_59 wwl_0_41 rwl_1_41
+ rwl_0_41 cell_2r1w
Xcell_2r1w_289 vdd_uq14 gnd read_bl_0_59 read_bl_1_59 write_bl_0_59 wwl_0_30 rwl_1_30
+ rwl_0_30 cell_2r1w
Xcell_2r1w_2231 vdd_uq3 gnd read_bl_0_29 read_bl_1_29 write_bl_0_29 wwl_0_8 rwl_1_8
+ rwl_0_8 cell_2r1w
Xcell_2r1w_2220 vdd_uq8 gnd read_bl_0_29 read_bl_1_29 write_bl_0_29 wwl_0_19 rwl_1_19
+ rwl_0_19 cell_2r1w
Xcell_2r1w_2242 vdd_uq29 gnd read_bl_0_28 read_bl_1_28 write_bl_0_28 wwl_0_61 rwl_1_61
+ rwl_0_61 cell_2r1w
Xcell_2r1w_1541 vdd_uq28 gnd read_bl_0_39 read_bl_1_39 write_bl_0_39 wwl_0_58 rwl_1_58
+ rwl_0_58 cell_2r1w
Xcell_2r1w_2253 vdd_uq24 gnd read_bl_0_28 read_bl_1_28 write_bl_0_28 wwl_0_50 rwl_1_50
+ rwl_0_50 cell_2r1w
Xcell_2r1w_1552 vdd_uq22 gnd read_bl_0_39 read_bl_1_39 write_bl_0_39 wwl_0_47 rwl_1_47
+ rwl_0_47 cell_2r1w
Xcell_2r1w_790 vdd_uq19 gnd read_bl_0_51 read_bl_1_51 write_bl_0_51 wwl_0_41 rwl_1_41
+ rwl_0_41 cell_2r1w
Xcell_2r1w_2264 vdd_uq18 gnd read_bl_0_28 read_bl_1_28 write_bl_0_28 wwl_0_39 rwl_1_39
+ rwl_0_39 cell_2r1w
Xcell_2r1w_1563 vdd_uq17 gnd read_bl_0_39 read_bl_1_39 write_bl_0_39 wwl_0_36 rwl_1_36
+ rwl_0_36 cell_2r1w
Xcell_2r1w_2275 vdd_uq13 gnd read_bl_0_28 read_bl_1_28 write_bl_0_28 wwl_0_28 rwl_1_28
+ rwl_0_28 cell_2r1w
Xcell_2r1w_1574 vdd_uq11 gnd read_bl_0_39 read_bl_1_39 write_bl_0_39 wwl_0_25 rwl_1_25
+ rwl_0_25 cell_2r1w
Xcell_2r1w_1530 vdd_uq1 gnd read_bl_0_40 read_bl_1_40 write_bl_0_40 wwl_0_5 rwl_1_5
+ rwl_0_5 cell_2r1w
Xcell_2r1w_1596 vdd gnd read_bl_0_39 read_bl_1_39 write_bl_0_39 wwl_0_3 rwl_1_3 rwl_0_3
+ cell_2r1w
Xcell_2r1w_2297 vdd_uq2 gnd read_bl_0_28 read_bl_1_28 write_bl_0_28 wwl_0_6 rwl_1_6
+ rwl_0_6 cell_2r1w
Xcell_2r1w_1585 vdd_uq6 gnd read_bl_0_39 read_bl_1_39 write_bl_0_39 wwl_0_14 rwl_1_14
+ rwl_0_14 cell_2r1w
Xcell_2r1w_2286 vdd_uq7 gnd read_bl_0_28 read_bl_1_28 write_bl_0_28 wwl_0_17 rwl_1_17
+ rwl_0_17 cell_2r1w
Xcell_2r1w_2050 vdd_uq29 gnd read_bl_0_31 read_bl_1_31 write_bl_0_31 wwl_0_61 rwl_1_61
+ rwl_0_61 cell_2r1w
Xcell_2r1w_2061 vdd_uq24 gnd read_bl_0_31 read_bl_1_31 write_bl_0_31 wwl_0_50 rwl_1_50
+ rwl_0_50 cell_2r1w
Xcell_2r1w_2072 vdd_uq18 gnd read_bl_0_31 read_bl_1_31 write_bl_0_31 wwl_0_39 rwl_1_39
+ rwl_0_39 cell_2r1w
Xcell_2r1w_2083 vdd_uq13 gnd read_bl_0_31 read_bl_1_31 write_bl_0_31 wwl_0_28 rwl_1_28
+ rwl_0_28 cell_2r1w
Xcell_2r1w_1360 vdd_uq22 gnd read_bl_0_42 read_bl_1_42 write_bl_0_42 wwl_0_47 rwl_1_47
+ rwl_0_47 cell_2r1w
Xcell_2r1w_1371 vdd_uq17 gnd read_bl_0_42 read_bl_1_42 write_bl_0_42 wwl_0_36 rwl_1_36
+ rwl_0_36 cell_2r1w
Xcell_2r1w_1382 vdd_uq11 gnd read_bl_0_42 read_bl_1_42 write_bl_0_42 wwl_0_25 rwl_1_25
+ rwl_0_25 cell_2r1w
Xcell_2r1w_1393 vdd_uq6 gnd read_bl_0_42 read_bl_1_42 write_bl_0_42 wwl_0_14 rwl_1_14
+ rwl_0_14 cell_2r1w
Xcell_2r1w_2094 vdd_uq7 gnd read_bl_0_31 read_bl_1_31 write_bl_0_31 wwl_0_17 rwl_1_17
+ rwl_0_17 cell_2r1w
Xcell_2r1w_1190 vdd_uq11 gnd read_bl_0_45 read_bl_1_45 write_bl_0_45 wwl_0_25 rwl_1_25
+ rwl_0_25 cell_2r1w
Xcell_2r1w_2819 vdd_uq29 gnd read_bl_0_19 read_bl_1_19 write_bl_0_19 wwl_0_60 rwl_1_60
+ rwl_0_60 cell_2r1w
Xcell_2r1w_2808 vdd_uq2 gnd read_bl_0_20 read_bl_1_20 write_bl_0_20 wwl_0_7 rwl_1_7
+ rwl_0_7 cell_2r1w
Xcell_2r1w_3509 vdd_uq4 gnd read_bl_0_9 read_bl_1_9 write_bl_0_9 wwl_0_10 rwl_1_10
+ rwl_0_10 cell_2r1w
Xcell_2r1w_608 vdd_uq14 gnd read_bl_0_54 read_bl_1_54 write_bl_0_54 wwl_0_31 rwl_1_31
+ rwl_0_31 cell_2r1w
Xcell_2r1w_619 vdd_uq9 gnd read_bl_0_54 read_bl_1_54 write_bl_0_54 wwl_0_20 rwl_1_20
+ rwl_0_20 cell_2r1w
Xcell_2r1w_4007 vdd_uq11 gnd read_bl_0_1 read_bl_1_1 write_bl_0_1 wwl_0_24 rwl_1_24
+ rwl_0_24 cell_2r1w
Xcell_2r1w_4029 vdd gnd read_bl_0_1 read_bl_1_1 write_bl_0_1 wwl_0_2 rwl_1_2 rwl_0_2
+ cell_2r1w
Xcell_2r1w_3317 vdd_uq4 gnd read_bl_0_12 read_bl_1_12 write_bl_0_12 wwl_0_10 rwl_1_10
+ rwl_0_10 cell_2r1w
Xcell_2r1w_4018 vdd_uq5 gnd read_bl_0_1 read_bl_1_1 write_bl_0_1 wwl_0_13 rwl_1_13
+ rwl_0_13 cell_2r1w
Xcell_2r1w_3306 vdd_uq9 gnd read_bl_0_12 read_bl_1_12 write_bl_0_12 wwl_0_21 rwl_1_21
+ rwl_0_21 cell_2r1w
Xcell_2r1w_3328 vdd_uq30 gnd read_bl_0_11 read_bl_1_11 write_bl_0_11 wwl_0_63 rwl_1_63
+ rwl_0_63 cell_2r1w
Xcell_2r1w_2627 vdd_uq29 gnd read_bl_0_22 read_bl_1_22 write_bl_0_22 wwl_0_60 rwl_1_60
+ rwl_0_60 cell_2r1w
Xcell_2r1w_1926 vdd_uq27 gnd read_bl_0_33 read_bl_1_33 write_bl_0_33 wwl_0_57 rwl_1_57
+ rwl_0_57 cell_2r1w
Xcell_2r1w_3339 vdd_uq25 gnd read_bl_0_11 read_bl_1_11 write_bl_0_11 wwl_0_52 rwl_1_52
+ rwl_0_52 cell_2r1w
Xcell_2r1w_2638 vdd_uq23 gnd read_bl_0_22 read_bl_1_22 write_bl_0_22 wwl_0_49 rwl_1_49
+ rwl_0_49 cell_2r1w
Xcell_2r1w_1937 vdd_uq22 gnd read_bl_0_33 read_bl_1_33 write_bl_0_33 wwl_0_46 rwl_1_46
+ rwl_0_46 cell_2r1w
Xcell_2r1w_2649 vdd_uq18 gnd read_bl_0_22 read_bl_1_22 write_bl_0_22 wwl_0_38 rwl_1_38
+ rwl_0_38 cell_2r1w
Xcell_2r1w_1948 vdd_uq16 gnd read_bl_0_33 read_bl_1_33 write_bl_0_33 wwl_0_35 rwl_1_35
+ rwl_0_35 cell_2r1w
Xcell_2r1w_1959 vdd_uq11 gnd read_bl_0_33 read_bl_1_33 write_bl_0_33 wwl_0_24 rwl_1_24
+ rwl_0_24 cell_2r1w
Xcell_2r1w_1915 vdd_uq1 gnd read_bl_0_34 read_bl_1_34 write_bl_0_34 wwl_0_4 rwl_1_4
+ rwl_0_4 cell_2r1w
Xcell_2r1w_2616 vdd_uq2 gnd read_bl_0_23 read_bl_1_23 write_bl_0_23 wwl_0_7 rwl_1_7
+ rwl_0_7 cell_2r1w
Xcell_2r1w_1904 vdd_uq6 gnd read_bl_0_34 read_bl_1_34 write_bl_0_34 wwl_0_15 rwl_1_15
+ rwl_0_15 cell_2r1w
Xcell_2r1w_2605 vdd_uq8 gnd read_bl_0_23 read_bl_1_23 write_bl_0_23 wwl_0_18 rwl_1_18
+ rwl_0_18 cell_2r1w
Xcell_2r1w_3840 vdd_uq30 gnd read_bl_0_3 read_bl_1_3 write_bl_0_3 wwl_0_63 rwl_1_63
+ rwl_0_63 cell_2r1w
Xcell_2r1w_3851 vdd_uq25 gnd read_bl_0_3 read_bl_1_3 write_bl_0_3 wwl_0_52 rwl_1_52
+ rwl_0_52 cell_2r1w
Xcell_2r1w_3862 vdd_uq19 gnd read_bl_0_3 read_bl_1_3 write_bl_0_3 wwl_0_41 rwl_1_41
+ rwl_0_41 cell_2r1w
Xcell_2r1w_3873 vdd_uq14 gnd read_bl_0_3 read_bl_1_3 write_bl_0_3 wwl_0_30 rwl_1_30
+ rwl_0_30 cell_2r1w
Xcell_2r1w_3895 vdd_uq3 gnd read_bl_0_3 read_bl_1_3 write_bl_0_3 wwl_0_8 rwl_1_8 rwl_0_8
+ cell_2r1w
Xcell_2r1w_3884 vdd_uq8 gnd read_bl_0_3 read_bl_1_3 write_bl_0_3 wwl_0_19 rwl_1_19
+ rwl_0_19 cell_2r1w
Xcell_2r1w_405 vdd_uq20 gnd read_bl_0_57 read_bl_1_57 write_bl_0_57 wwl_0_42 rwl_1_42
+ rwl_0_42 cell_2r1w
Xcell_2r1w_416 vdd_uq14 gnd read_bl_0_57 read_bl_1_57 write_bl_0_57 wwl_0_31 rwl_1_31
+ rwl_0_31 cell_2r1w
Xcell_2r1w_427 vdd_uq9 gnd read_bl_0_57 read_bl_1_57 write_bl_0_57 wwl_0_20 rwl_1_20
+ rwl_0_20 cell_2r1w
Xcell_2r1w_449 vdd_uq30 gnd read_bl_0_56 read_bl_1_56 write_bl_0_56 wwl_0_62 rwl_1_62
+ rwl_0_62 cell_2r1w
Xcell_2r1w_438 vdd_uq3 gnd read_bl_0_57 read_bl_1_57 write_bl_0_57 wwl_0_9 rwl_1_9
+ rwl_0_9 cell_2r1w
Xcell_2r1w_3136 vdd_uq30 gnd read_bl_0_14 read_bl_1_14 write_bl_0_14 wwl_0_63 rwl_1_63
+ rwl_0_63 cell_2r1w
Xcell_2r1w_3147 vdd_uq25 gnd read_bl_0_14 read_bl_1_14 write_bl_0_14 wwl_0_52 rwl_1_52
+ rwl_0_52 cell_2r1w
Xcell_2r1w_3158 vdd_uq19 gnd read_bl_0_14 read_bl_1_14 write_bl_0_14 wwl_0_41 rwl_1_41
+ rwl_0_41 cell_2r1w
Xcell_2r1w_3103 vdd_uq15 gnd read_bl_0_15 read_bl_1_15 write_bl_0_15 wwl_0_32 rwl_1_32
+ rwl_0_32 cell_2r1w
Xcell_2r1w_2402 vdd_uq13 gnd read_bl_0_26 read_bl_1_26 write_bl_0_26 wwl_0_29 rwl_1_29
+ rwl_0_29 cell_2r1w
Xcell_2r1w_3125 vdd_uq4 gnd read_bl_0_15 read_bl_1_15 write_bl_0_15 wwl_0_10 rwl_1_10
+ rwl_0_10 cell_2r1w
Xcell_2r1w_2413 vdd_uq8 gnd read_bl_0_26 read_bl_1_26 write_bl_0_26 wwl_0_18 rwl_1_18
+ rwl_0_18 cell_2r1w
Xcell_2r1w_3114 vdd_uq9 gnd read_bl_0_15 read_bl_1_15 write_bl_0_15 wwl_0_21 rwl_1_21
+ rwl_0_21 cell_2r1w
Xcell_2r1w_961 vdd_uq30 gnd read_bl_0_48 read_bl_1_48 write_bl_0_48 wwl_0_62 rwl_1_62
+ rwl_0_62 cell_2r1w
Xcell_2r1w_2435 vdd_uq29 gnd read_bl_0_25 read_bl_1_25 write_bl_0_25 wwl_0_60 rwl_1_60
+ rwl_0_60 cell_2r1w
Xcell_2r1w_1734 vdd_uq27 gnd read_bl_0_36 read_bl_1_36 write_bl_0_36 wwl_0_57 rwl_1_57
+ rwl_0_57 cell_2r1w
Xcell_2r1w_972 vdd_uq24 gnd read_bl_0_48 read_bl_1_48 write_bl_0_48 wwl_0_51 rwl_1_51
+ rwl_0_51 cell_2r1w
Xcell_2r1w_2446 vdd_uq23 gnd read_bl_0_25 read_bl_1_25 write_bl_0_25 wwl_0_49 rwl_1_49
+ rwl_0_49 cell_2r1w
Xcell_2r1w_1745 vdd_uq22 gnd read_bl_0_36 read_bl_1_36 write_bl_0_36 wwl_0_46 rwl_1_46
+ rwl_0_46 cell_2r1w
Xcell_2r1w_983 vdd_uq19 gnd read_bl_0_48 read_bl_1_48 write_bl_0_48 wwl_0_40 rwl_1_40
+ rwl_0_40 cell_2r1w
Xcell_2r1w_2457 vdd_uq18 gnd read_bl_0_25 read_bl_1_25 write_bl_0_25 wwl_0_38 rwl_1_38
+ rwl_0_38 cell_2r1w
Xcell_2r1w_1756 vdd_uq16 gnd read_bl_0_36 read_bl_1_36 write_bl_0_36 wwl_0_35 rwl_1_35
+ rwl_0_35 cell_2r1w
Xcell_2r1w_3169 vdd_uq14 gnd read_bl_0_14 read_bl_1_14 write_bl_0_14 wwl_0_30 rwl_1_30
+ rwl_0_30 cell_2r1w
Xcell_2r1w_2468 vdd_uq12 gnd read_bl_0_25 read_bl_1_25 write_bl_0_25 wwl_0_27 rwl_1_27
+ rwl_0_27 cell_2r1w
Xcell_2r1w_1701 vdd_uq12 gnd read_bl_0_37 read_bl_1_37 write_bl_0_37 wwl_0_26 rwl_1_26
+ rwl_0_26 cell_2r1w
Xcell_2r1w_1767 vdd_uq11 gnd read_bl_0_36 read_bl_1_36 write_bl_0_36 wwl_0_24 rwl_1_24
+ rwl_0_24 cell_2r1w
Xcell_2r1w_1723 vdd_uq1 gnd read_bl_0_37 read_bl_1_37 write_bl_0_37 wwl_0_4 rwl_1_4
+ rwl_0_4 cell_2r1w
Xcell_2r1w_1789 vdd gnd read_bl_0_36 read_bl_1_36 write_bl_0_36 wwl_0_2 rwl_1_2 rwl_0_2
+ cell_2r1w
Xcell_2r1w_2424 vdd_uq2 gnd read_bl_0_26 read_bl_1_26 write_bl_0_26 wwl_0_7 rwl_1_7
+ rwl_0_7 cell_2r1w
Xcell_2r1w_950 vdd_uq3 gnd read_bl_0_49 read_bl_1_49 write_bl_0_49 wwl_0_9 rwl_1_9
+ rwl_0_9 cell_2r1w
Xcell_2r1w_1778 vdd_uq5 gnd read_bl_0_36 read_bl_1_36 write_bl_0_36 wwl_0_13 rwl_1_13
+ rwl_0_13 cell_2r1w
Xcell_2r1w_1712 vdd_uq6 gnd read_bl_0_37 read_bl_1_37 write_bl_0_37 wwl_0_15 rwl_1_15
+ rwl_0_15 cell_2r1w
Xcell_2r1w_2479 vdd_uq7 gnd read_bl_0_25 read_bl_1_25 write_bl_0_25 wwl_0_16 rwl_1_16
+ rwl_0_16 cell_2r1w
Xcell_2r1w_994 vdd_uq13 gnd read_bl_0_48 read_bl_1_48 write_bl_0_48 wwl_0_29 rwl_1_29
+ rwl_0_29 cell_2r1w
Xcell_2r1w_3670 vdd_uq19 gnd read_bl_0_6 read_bl_1_6 write_bl_0_6 wwl_0_41 rwl_1_41
+ rwl_0_41 cell_2r1w
Xcell_2r1w_3681 vdd_uq14 gnd read_bl_0_6 read_bl_1_6 write_bl_0_6 wwl_0_30 rwl_1_30
+ rwl_0_30 cell_2r1w
Xcell_2r1w_3692 vdd_uq8 gnd read_bl_0_6 read_bl_1_6 write_bl_0_6 wwl_0_19 rwl_1_19
+ rwl_0_19 cell_2r1w
Xcell_2r1w_2980 vdd_uq12 gnd read_bl_0_17 read_bl_1_17 write_bl_0_17 wwl_0_27 rwl_1_27
+ rwl_0_27 cell_2r1w
Xcell_2r1w_2991 vdd_uq7 gnd read_bl_0_17 read_bl_1_17 write_bl_0_17 wwl_0_16 rwl_1_16
+ rwl_0_16 cell_2r1w
Xcell_2r1w_73 vdd_uq26 gnd read_bl_0_62 read_bl_1_62 write_bl_0_62 wwl_0_54 rwl_1_54
+ rwl_0_54 cell_2r1w
Xcell_2r1w_84 vdd_uq20 gnd read_bl_0_62 read_bl_1_62 write_bl_0_62 wwl_0_43 rwl_1_43
+ rwl_0_43 cell_2r1w
Xcell_2r1w_95 vdd_uq15 gnd read_bl_0_62 read_bl_1_62 write_bl_0_62 wwl_0_32 rwl_1_32
+ rwl_0_32 cell_2r1w
Xcell_2r1w_62 vdd_uq0 gnd read_bl_0_63 read_bl_1_63 write_bl_0_63 wwl_0_1 rwl_1_1
+ rwl_0_1 cell_2r1w
Xcell_2r1w_51 vdd_uq5 gnd read_bl_0_63 read_bl_1_63 write_bl_0_63 wwl_0_12 rwl_1_12
+ rwl_0_12 cell_2r1w
Xcell_2r1w_40 vdd_uq10 gnd read_bl_0_63 read_bl_1_63 write_bl_0_63 wwl_0_23 rwl_1_23
+ rwl_0_23 cell_2r1w
Xcell_2r1w_257 vdd_uq30 gnd read_bl_0_59 read_bl_1_59 write_bl_0_59 wwl_0_62 rwl_1_62
+ rwl_0_62 cell_2r1w
Xcell_2r1w_202 vdd_uq25 gnd read_bl_0_60 read_bl_1_60 write_bl_0_60 wwl_0_53 rwl_1_53
+ rwl_0_53 cell_2r1w
Xcell_2r1w_268 vdd_uq24 gnd read_bl_0_59 read_bl_1_59 write_bl_0_59 wwl_0_51 rwl_1_51
+ rwl_0_51 cell_2r1w
Xcell_2r1w_213 vdd_uq20 gnd read_bl_0_60 read_bl_1_60 write_bl_0_60 wwl_0_42 rwl_1_42
+ rwl_0_42 cell_2r1w
Xcell_2r1w_224 vdd_uq14 gnd read_bl_0_60 read_bl_1_60 write_bl_0_60 wwl_0_31 rwl_1_31
+ rwl_0_31 cell_2r1w
Xcell_2r1w_1019 vdd_uq1 gnd read_bl_0_48 read_bl_1_48 write_bl_0_48 wwl_0_4 rwl_1_4
+ rwl_0_4 cell_2r1w
Xcell_2r1w_246 vdd_uq3 gnd read_bl_0_60 read_bl_1_60 write_bl_0_60 wwl_0_9 rwl_1_9
+ rwl_0_9 cell_2r1w
Xcell_2r1w_1008 vdd_uq6 gnd read_bl_0_48 read_bl_1_48 write_bl_0_48 wwl_0_15 rwl_1_15
+ rwl_0_15 cell_2r1w
Xcell_2r1w_235 vdd_uq9 gnd read_bl_0_60 read_bl_1_60 write_bl_0_60 wwl_0_20 rwl_1_20
+ rwl_0_20 cell_2r1w
Xcell_2r1w_279 vdd_uq19 gnd read_bl_0_59 read_bl_1_59 write_bl_0_59 wwl_0_40 rwl_1_40
+ rwl_0_40 cell_2r1w
Xcell_2r1w_2243 vdd_uq29 gnd read_bl_0_28 read_bl_1_28 write_bl_0_28 wwl_0_60 rwl_1_60
+ rwl_0_60 cell_2r1w
Xcell_2r1w_2254 vdd_uq23 gnd read_bl_0_28 read_bl_1_28 write_bl_0_28 wwl_0_49 rwl_1_49
+ rwl_0_49 cell_2r1w
Xcell_2r1w_2265 vdd_uq18 gnd read_bl_0_28 read_bl_1_28 write_bl_0_28 wwl_0_38 rwl_1_38
+ rwl_0_38 cell_2r1w
Xcell_2r1w_2210 vdd_uq13 gnd read_bl_0_29 read_bl_1_29 write_bl_0_29 wwl_0_29 rwl_1_29
+ rwl_0_29 cell_2r1w
Xcell_2r1w_2232 vdd_uq2 gnd read_bl_0_29 read_bl_1_29 write_bl_0_29 wwl_0_7 rwl_1_7
+ rwl_0_7 cell_2r1w
Xcell_2r1w_1520 vdd_uq6 gnd read_bl_0_40 read_bl_1_40 write_bl_0_40 wwl_0_15 rwl_1_15
+ rwl_0_15 cell_2r1w
Xcell_2r1w_2221 vdd_uq8 gnd read_bl_0_29 read_bl_1_29 write_bl_0_29 wwl_0_18 rwl_1_18
+ rwl_0_18 cell_2r1w
Xcell_2r1w_1542 vdd_uq27 gnd read_bl_0_39 read_bl_1_39 write_bl_0_39 wwl_0_57 rwl_1_57
+ rwl_0_57 cell_2r1w
Xcell_2r1w_780 vdd_uq24 gnd read_bl_0_51 read_bl_1_51 write_bl_0_51 wwl_0_51 rwl_1_51
+ rwl_0_51 cell_2r1w
Xcell_2r1w_1553 vdd_uq22 gnd read_bl_0_39 read_bl_1_39 write_bl_0_39 wwl_0_46 rwl_1_46
+ rwl_0_46 cell_2r1w
Xcell_2r1w_791 vdd_uq19 gnd read_bl_0_51 read_bl_1_51 write_bl_0_51 wwl_0_40 rwl_1_40
+ rwl_0_40 cell_2r1w
Xcell_2r1w_1564 vdd_uq16 gnd read_bl_0_39 read_bl_1_39 write_bl_0_39 wwl_0_35 rwl_1_35
+ rwl_0_35 cell_2r1w
Xcell_2r1w_2276 vdd_uq12 gnd read_bl_0_28 read_bl_1_28 write_bl_0_28 wwl_0_27 rwl_1_27
+ rwl_0_27 cell_2r1w
Xcell_2r1w_1575 vdd_uq11 gnd read_bl_0_39 read_bl_1_39 write_bl_0_39 wwl_0_24 rwl_1_24
+ rwl_0_24 cell_2r1w
Xcell_2r1w_2298 vdd_uq1 gnd read_bl_0_28 read_bl_1_28 write_bl_0_28 wwl_0_5 rwl_1_5
+ rwl_0_5 cell_2r1w
Xcell_2r1w_1531 vdd_uq1 gnd read_bl_0_40 read_bl_1_40 write_bl_0_40 wwl_0_4 rwl_1_4
+ rwl_0_4 cell_2r1w
Xcell_2r1w_1597 vdd gnd read_bl_0_39 read_bl_1_39 write_bl_0_39 wwl_0_2 rwl_1_2 rwl_0_2
+ cell_2r1w
Xcell_2r1w_1586 vdd_uq5 gnd read_bl_0_39 read_bl_1_39 write_bl_0_39 wwl_0_13 rwl_1_13
+ rwl_0_13 cell_2r1w
Xcell_2r1w_2287 vdd_uq7 gnd read_bl_0_28 read_bl_1_28 write_bl_0_28 wwl_0_16 rwl_1_16
+ rwl_0_16 cell_2r1w
Xcell_2r1w_2051 vdd_uq29 gnd read_bl_0_31 read_bl_1_31 write_bl_0_31 wwl_0_60 rwl_1_60
+ rwl_0_60 cell_2r1w
Xcell_2r1w_1350 vdd_uq27 gnd read_bl_0_42 read_bl_1_42 write_bl_0_42 wwl_0_57 rwl_1_57
+ rwl_0_57 cell_2r1w
Xcell_2r1w_2062 vdd_uq23 gnd read_bl_0_31 read_bl_1_31 write_bl_0_31 wwl_0_49 rwl_1_49
+ rwl_0_49 cell_2r1w
Xcell_2r1w_1361 vdd_uq22 gnd read_bl_0_42 read_bl_1_42 write_bl_0_42 wwl_0_46 rwl_1_46
+ rwl_0_46 cell_2r1w
Xcell_2r1w_2073 vdd_uq18 gnd read_bl_0_31 read_bl_1_31 write_bl_0_31 wwl_0_38 rwl_1_38
+ rwl_0_38 cell_2r1w
Xcell_2r1w_1372 vdd_uq16 gnd read_bl_0_42 read_bl_1_42 write_bl_0_42 wwl_0_35 rwl_1_35
+ rwl_0_35 cell_2r1w
Xcell_2r1w_2084 vdd_uq12 gnd read_bl_0_31 read_bl_1_31 write_bl_0_31 wwl_0_27 rwl_1_27
+ rwl_0_27 cell_2r1w
Xcell_2r1w_2040 vdd_uq2 gnd read_bl_0_32 read_bl_1_32 write_bl_0_32 wwl_0_7 rwl_1_7
+ rwl_0_7 cell_2r1w
Xcell_2r1w_2095 vdd_uq7 gnd read_bl_0_31 read_bl_1_31 write_bl_0_31 wwl_0_16 rwl_1_16
+ rwl_0_16 cell_2r1w
Xcell_2r1w_1383 vdd_uq11 gnd read_bl_0_42 read_bl_1_42 write_bl_0_42 wwl_0_24 rwl_1_24
+ rwl_0_24 cell_2r1w
Xcell_2r1w_1394 vdd_uq5 gnd read_bl_0_42 read_bl_1_42 write_bl_0_42 wwl_0_13 rwl_1_13
+ rwl_0_13 cell_2r1w
Xcell_2r1w_1180 vdd_uq16 gnd read_bl_0_45 read_bl_1_45 write_bl_0_45 wwl_0_35 rwl_1_35
+ rwl_0_35 cell_2r1w
Xcell_2r1w_1191 vdd_uq11 gnd read_bl_0_45 read_bl_1_45 write_bl_0_45 wwl_0_24 rwl_1_24
+ rwl_0_24 cell_2r1w
Xcell_2r1w_2809 vdd_uq2 gnd read_bl_0_20 read_bl_1_20 write_bl_0_20 wwl_0_6 rwl_1_6
+ rwl_0_6 cell_2r1w
Xcell_2r1w_609 vdd_uq14 gnd read_bl_0_54 read_bl_1_54 write_bl_0_54 wwl_0_30 rwl_1_30
+ rwl_0_30 cell_2r1w
Xcell_2r1w_3329 vdd_uq30 gnd read_bl_0_11 read_bl_1_11 write_bl_0_11 wwl_0_62 rwl_1_62
+ rwl_0_62 cell_2r1w
Xcell_2r1w_3318 vdd_uq3 gnd read_bl_0_12 read_bl_1_12 write_bl_0_12 wwl_0_9 rwl_1_9
+ rwl_0_9 cell_2r1w
Xcell_2r1w_4019 vdd_uq5 gnd read_bl_0_1 read_bl_1_1 write_bl_0_1 wwl_0_12 rwl_1_12
+ rwl_0_12 cell_2r1w
Xcell_2r1w_2606 vdd_uq7 gnd read_bl_0_23 read_bl_1_23 write_bl_0_23 wwl_0_17 rwl_1_17
+ rwl_0_17 cell_2r1w
Xcell_2r1w_3307 vdd_uq9 gnd read_bl_0_12 read_bl_1_12 write_bl_0_12 wwl_0_20 rwl_1_20
+ rwl_0_20 cell_2r1w
Xcell_2r1w_4008 vdd_uq10 gnd read_bl_0_1 read_bl_1_1 write_bl_0_1 wwl_0_23 rwl_1_23
+ rwl_0_23 cell_2r1w
Xcell_2r1w_2628 vdd_uq28 gnd read_bl_0_22 read_bl_1_22 write_bl_0_22 wwl_0_59 rwl_1_59
+ rwl_0_59 cell_2r1w
Xcell_2r1w_1927 vdd_uq27 gnd read_bl_0_33 read_bl_1_33 write_bl_0_33 wwl_0_56 rwl_1_56
+ rwl_0_56 cell_2r1w
Xcell_2r1w_2639 vdd_uq23 gnd read_bl_0_22 read_bl_1_22 write_bl_0_22 wwl_0_48 rwl_1_48
+ rwl_0_48 cell_2r1w
Xcell_2r1w_1938 vdd_uq21 gnd read_bl_0_33 read_bl_1_33 write_bl_0_33 wwl_0_45 rwl_1_45
+ rwl_0_45 cell_2r1w
Xcell_2r1w_1949 vdd_uq16 gnd read_bl_0_33 read_bl_1_33 write_bl_0_33 wwl_0_34 rwl_1_34
+ rwl_0_34 cell_2r1w
Xcell_2r1w_1916 vdd gnd read_bl_0_34 read_bl_1_34 write_bl_0_34 wwl_0_3 rwl_1_3 rwl_0_3
+ cell_2r1w
Xcell_2r1w_2617 vdd_uq2 gnd read_bl_0_23 read_bl_1_23 write_bl_0_23 wwl_0_6 rwl_1_6
+ rwl_0_6 cell_2r1w
Xcell_2r1w_1905 vdd_uq6 gnd read_bl_0_34 read_bl_1_34 write_bl_0_34 wwl_0_14 rwl_1_14
+ rwl_0_14 cell_2r1w
Xcell_2r1w_3841 vdd_uq30 gnd read_bl_0_3 read_bl_1_3 write_bl_0_3 wwl_0_62 rwl_1_62
+ rwl_0_62 cell_2r1w
Xcell_2r1w_3852 vdd_uq24 gnd read_bl_0_3 read_bl_1_3 write_bl_0_3 wwl_0_51 rwl_1_51
+ rwl_0_51 cell_2r1w
Xcell_2r1w_3863 vdd_uq19 gnd read_bl_0_3 read_bl_1_3 write_bl_0_3 wwl_0_40 rwl_1_40
+ rwl_0_40 cell_2r1w
Xcell_2r1w_3874 vdd_uq13 gnd read_bl_0_3 read_bl_1_3 write_bl_0_3 wwl_0_29 rwl_1_29
+ rwl_0_29 cell_2r1w
Xcell_2r1w_3896 vdd_uq2 gnd read_bl_0_3 read_bl_1_3 write_bl_0_3 wwl_0_7 rwl_1_7 rwl_0_7
+ cell_2r1w
Xcell_2r1w_3830 vdd_uq3 gnd read_bl_0_4 read_bl_1_4 write_bl_0_4 wwl_0_9 rwl_1_9 rwl_0_9
+ cell_2r1w
Xcell_2r1w_3885 vdd_uq8 gnd read_bl_0_3 read_bl_1_3 write_bl_0_3 wwl_0_18 rwl_1_18
+ rwl_0_18 cell_2r1w
Xcell_2r1w_406 vdd_uq19 gnd read_bl_0_57 read_bl_1_57 write_bl_0_57 wwl_0_41 rwl_1_41
+ rwl_0_41 cell_2r1w
Xcell_2r1w_417 vdd_uq14 gnd read_bl_0_57 read_bl_1_57 write_bl_0_57 wwl_0_30 rwl_1_30
+ rwl_0_30 cell_2r1w
Xcell_2r1w_439 vdd_uq3 gnd read_bl_0_57 read_bl_1_57 write_bl_0_57 wwl_0_8 rwl_1_8
+ rwl_0_8 cell_2r1w
Xcell_2r1w_428 vdd_uq8 gnd read_bl_0_57 read_bl_1_57 write_bl_0_57 wwl_0_19 rwl_1_19
+ rwl_0_19 cell_2r1w
Xcell_2r1w_3137 vdd_uq30 gnd read_bl_0_14 read_bl_1_14 write_bl_0_14 wwl_0_62 rwl_1_62
+ rwl_0_62 cell_2r1w
Xcell_2r1w_2436 vdd_uq28 gnd read_bl_0_25 read_bl_1_25 write_bl_0_25 wwl_0_59 rwl_1_59
+ rwl_0_59 cell_2r1w
Xcell_2r1w_3148 vdd_uq24 gnd read_bl_0_14 read_bl_1_14 write_bl_0_14 wwl_0_51 rwl_1_51
+ rwl_0_51 cell_2r1w
Xcell_2r1w_2447 vdd_uq23 gnd read_bl_0_25 read_bl_1_25 write_bl_0_25 wwl_0_48 rwl_1_48
+ rwl_0_48 cell_2r1w
Xcell_2r1w_3159 vdd_uq19 gnd read_bl_0_14 read_bl_1_14 write_bl_0_14 wwl_0_40 rwl_1_40
+ rwl_0_40 cell_2r1w
Xcell_2r1w_3104 vdd_uq14 gnd read_bl_0_15 read_bl_1_15 write_bl_0_15 wwl_0_31 rwl_1_31
+ rwl_0_31 cell_2r1w
Xcell_2r1w_2403 vdd_uq13 gnd read_bl_0_26 read_bl_1_26 write_bl_0_26 wwl_0_28 rwl_1_28
+ rwl_0_28 cell_2r1w
Xcell_2r1w_1702 vdd_uq11 gnd read_bl_0_37 read_bl_1_37 write_bl_0_37 wwl_0_25 rwl_1_25
+ rwl_0_25 cell_2r1w
Xcell_2r1w_2425 vdd_uq2 gnd read_bl_0_26 read_bl_1_26 write_bl_0_26 wwl_0_6 rwl_1_6
+ rwl_0_6 cell_2r1w
Xcell_2r1w_3126 vdd_uq3 gnd read_bl_0_15 read_bl_1_15 write_bl_0_15 wwl_0_9 rwl_1_9
+ rwl_0_9 cell_2r1w
Xcell_2r1w_2414 vdd_uq7 gnd read_bl_0_26 read_bl_1_26 write_bl_0_26 wwl_0_17 rwl_1_17
+ rwl_0_17 cell_2r1w
Xcell_2r1w_3115 vdd_uq9 gnd read_bl_0_15 read_bl_1_15 write_bl_0_15 wwl_0_20 rwl_1_20
+ rwl_0_20 cell_2r1w
Xcell_2r1w_962 vdd_uq29 gnd read_bl_0_48 read_bl_1_48 write_bl_0_48 wwl_0_61 rwl_1_61
+ rwl_0_61 cell_2r1w
Xcell_2r1w_1735 vdd_uq27 gnd read_bl_0_36 read_bl_1_36 write_bl_0_36 wwl_0_56 rwl_1_56
+ rwl_0_56 cell_2r1w
Xcell_2r1w_973 vdd_uq24 gnd read_bl_0_48 read_bl_1_48 write_bl_0_48 wwl_0_50 rwl_1_50
+ rwl_0_50 cell_2r1w
Xcell_2r1w_1746 vdd_uq21 gnd read_bl_0_36 read_bl_1_36 write_bl_0_36 wwl_0_45 rwl_1_45
+ rwl_0_45 cell_2r1w
Xcell_2r1w_984 vdd_uq18 gnd read_bl_0_48 read_bl_1_48 write_bl_0_48 wwl_0_39 rwl_1_39
+ rwl_0_39 cell_2r1w
Xcell_2r1w_2458 vdd_uq17 gnd read_bl_0_25 read_bl_1_25 write_bl_0_25 wwl_0_37 rwl_1_37
+ rwl_0_37 cell_2r1w
Xcell_2r1w_1757 vdd_uq16 gnd read_bl_0_36 read_bl_1_36 write_bl_0_36 wwl_0_34 rwl_1_34
+ rwl_0_34 cell_2r1w
Xcell_2r1w_995 vdd_uq13 gnd read_bl_0_48 read_bl_1_48 write_bl_0_48 wwl_0_28 rwl_1_28
+ rwl_0_28 cell_2r1w
Xcell_2r1w_2469 vdd_uq12 gnd read_bl_0_25 read_bl_1_25 write_bl_0_25 wwl_0_26 rwl_1_26
+ rwl_0_26 cell_2r1w
Xcell_2r1w_1724 vdd gnd read_bl_0_37 read_bl_1_37 write_bl_0_37 wwl_0_3 rwl_1_3 rwl_0_3
+ cell_2r1w
Xcell_2r1w_951 vdd_uq3 gnd read_bl_0_49 read_bl_1_49 write_bl_0_49 wwl_0_8 rwl_1_8
+ rwl_0_8 cell_2r1w
Xcell_2r1w_1779 vdd_uq5 gnd read_bl_0_36 read_bl_1_36 write_bl_0_36 wwl_0_12 rwl_1_12
+ rwl_0_12 cell_2r1w
Xcell_2r1w_1713 vdd_uq6 gnd read_bl_0_37 read_bl_1_37 write_bl_0_37 wwl_0_14 rwl_1_14
+ rwl_0_14 cell_2r1w
Xcell_2r1w_940 vdd_uq8 gnd read_bl_0_49 read_bl_1_49 write_bl_0_49 wwl_0_19 rwl_1_19
+ rwl_0_19 cell_2r1w
Xcell_2r1w_1768 vdd_uq10 gnd read_bl_0_36 read_bl_1_36 write_bl_0_36 wwl_0_23 rwl_1_23
+ rwl_0_23 cell_2r1w
Xcell_2r1w_3660 vdd_uq24 gnd read_bl_0_6 read_bl_1_6 write_bl_0_6 wwl_0_51 rwl_1_51
+ rwl_0_51 cell_2r1w
Xcell_2r1w_3671 vdd_uq19 gnd read_bl_0_6 read_bl_1_6 write_bl_0_6 wwl_0_40 rwl_1_40
+ rwl_0_40 cell_2r1w
Xcell_2r1w_2970 vdd_uq17 gnd read_bl_0_17 read_bl_1_17 write_bl_0_17 wwl_0_37 rwl_1_37
+ rwl_0_37 cell_2r1w
Xcell_2r1w_3682 vdd_uq13 gnd read_bl_0_6 read_bl_1_6 write_bl_0_6 wwl_0_29 rwl_1_29
+ rwl_0_29 cell_2r1w
Xcell_2r1w_2981 vdd_uq12 gnd read_bl_0_17 read_bl_1_17 write_bl_0_17 wwl_0_26 rwl_1_26
+ rwl_0_26 cell_2r1w
Xcell_2r1w_2992 vdd_uq6 gnd read_bl_0_17 read_bl_1_17 write_bl_0_17 wwl_0_15 rwl_1_15
+ rwl_0_15 cell_2r1w
Xcell_2r1w_3693 vdd_uq8 gnd read_bl_0_6 read_bl_1_6 write_bl_0_6 wwl_0_18 rwl_1_18
+ rwl_0_18 cell_2r1w
Xcell_2r1w_30 vdd_uq15 gnd read_bl_0_63 read_bl_1_63 write_bl_0_63 wwl_0_33 rwl_1_33
+ rwl_0_33 cell_2r1w
Xcell_2r1w_74 vdd_uq25 gnd read_bl_0_62 read_bl_1_62 write_bl_0_62 wwl_0_53 rwl_1_53
+ rwl_0_53 cell_2r1w
Xcell_2r1w_85 vdd_uq20 gnd read_bl_0_62 read_bl_1_62 write_bl_0_62 wwl_0_42 rwl_1_42
+ rwl_0_42 cell_2r1w
Xcell_2r1w_96 vdd_uq14 gnd read_bl_0_62 read_bl_1_62 write_bl_0_62 wwl_0_31 rwl_1_31
+ rwl_0_31 cell_2r1w
Xcell_2r1w_63 vdd_uq0 gnd read_bl_0_63 read_bl_1_63 write_bl_0_63 wwl_0_0 rwl_1_0
+ rwl_0_0 cell_2r1w
Xcell_2r1w_52 vdd_uq4 gnd read_bl_0_63 read_bl_1_63 write_bl_0_63 wwl_0_11 rwl_1_11
+ rwl_0_11 cell_2r1w
Xcell_2r1w_41 vdd_uq10 gnd read_bl_0_63 read_bl_1_63 write_bl_0_63 wwl_0_22 rwl_1_22
+ rwl_0_22 cell_2r1w
Xcell_2r1w_258 vdd_uq29 gnd read_bl_0_59 read_bl_1_59 write_bl_0_59 wwl_0_61 rwl_1_61
+ rwl_0_61 cell_2r1w
Xcell_2r1w_203 vdd_uq25 gnd read_bl_0_60 read_bl_1_60 write_bl_0_60 wwl_0_52 rwl_1_52
+ rwl_0_52 cell_2r1w
Xcell_2r1w_269 vdd_uq24 gnd read_bl_0_59 read_bl_1_59 write_bl_0_59 wwl_0_50 rwl_1_50
+ rwl_0_50 cell_2r1w
Xcell_2r1w_214 vdd_uq19 gnd read_bl_0_60 read_bl_1_60 write_bl_0_60 wwl_0_41 rwl_1_41
+ rwl_0_41 cell_2r1w
Xcell_2r1w_225 vdd_uq14 gnd read_bl_0_60 read_bl_1_60 write_bl_0_60 wwl_0_30 rwl_1_30
+ rwl_0_30 cell_2r1w
Xcell_2r1w_247 vdd_uq3 gnd read_bl_0_60 read_bl_1_60 write_bl_0_60 wwl_0_8 rwl_1_8
+ rwl_0_8 cell_2r1w
Xcell_2r1w_1009 vdd_uq6 gnd read_bl_0_48 read_bl_1_48 write_bl_0_48 wwl_0_14 rwl_1_14
+ rwl_0_14 cell_2r1w
Xcell_2r1w_236 vdd_uq8 gnd read_bl_0_60 read_bl_1_60 write_bl_0_60 wwl_0_19 rwl_1_19
+ rwl_0_19 cell_2r1w
Xcell_2r1w_2244 vdd_uq28 gnd read_bl_0_28 read_bl_1_28 write_bl_0_28 wwl_0_59 rwl_1_59
+ rwl_0_59 cell_2r1w
Xcell_2r1w_1543 vdd_uq27 gnd read_bl_0_39 read_bl_1_39 write_bl_0_39 wwl_0_56 rwl_1_56
+ rwl_0_56 cell_2r1w
Xcell_2r1w_2255 vdd_uq23 gnd read_bl_0_28 read_bl_1_28 write_bl_0_28 wwl_0_48 rwl_1_48
+ rwl_0_48 cell_2r1w
Xcell_2r1w_1554 vdd_uq21 gnd read_bl_0_39 read_bl_1_39 write_bl_0_39 wwl_0_45 rwl_1_45
+ rwl_0_45 cell_2r1w
Xcell_2r1w_2200 vdd_uq18 gnd read_bl_0_29 read_bl_1_29 write_bl_0_29 wwl_0_39 rwl_1_39
+ rwl_0_39 cell_2r1w
Xcell_2r1w_2266 vdd_uq17 gnd read_bl_0_28 read_bl_1_28 write_bl_0_28 wwl_0_37 rwl_1_37
+ rwl_0_37 cell_2r1w
Xcell_2r1w_2211 vdd_uq13 gnd read_bl_0_29 read_bl_1_29 write_bl_0_29 wwl_0_28 rwl_1_28
+ rwl_0_28 cell_2r1w
Xcell_2r1w_2277 vdd_uq12 gnd read_bl_0_28 read_bl_1_28 write_bl_0_28 wwl_0_26 rwl_1_26
+ rwl_0_26 cell_2r1w
Xcell_2r1w_1510 vdd_uq11 gnd read_bl_0_40 read_bl_1_40 write_bl_0_40 wwl_0_25 rwl_1_25
+ rwl_0_25 cell_2r1w
Xcell_2r1w_2299 vdd_uq1 gnd read_bl_0_28 read_bl_1_28 write_bl_0_28 wwl_0_4 rwl_1_4
+ rwl_0_4 cell_2r1w
Xcell_2r1w_1532 vdd gnd read_bl_0_40 read_bl_1_40 write_bl_0_40 wwl_0_3 rwl_1_3 rwl_0_3
+ cell_2r1w
Xcell_2r1w_2233 vdd_uq2 gnd read_bl_0_29 read_bl_1_29 write_bl_0_29 wwl_0_6 rwl_1_6
+ rwl_0_6 cell_2r1w
Xcell_2r1w_1521 vdd_uq6 gnd read_bl_0_40 read_bl_1_40 write_bl_0_40 wwl_0_14 rwl_1_14
+ rwl_0_14 cell_2r1w
Xcell_2r1w_2288 vdd_uq6 gnd read_bl_0_28 read_bl_1_28 write_bl_0_28 wwl_0_15 rwl_1_15
+ rwl_0_15 cell_2r1w
Xcell_2r1w_2222 vdd_uq7 gnd read_bl_0_29 read_bl_1_29 write_bl_0_29 wwl_0_17 rwl_1_17
+ rwl_0_17 cell_2r1w
Xcell_2r1w_770 vdd_uq29 gnd read_bl_0_51 read_bl_1_51 write_bl_0_51 wwl_0_61 rwl_1_61
+ rwl_0_61 cell_2r1w
Xcell_2r1w_781 vdd_uq24 gnd read_bl_0_51 read_bl_1_51 write_bl_0_51 wwl_0_50 rwl_1_50
+ rwl_0_50 cell_2r1w
Xcell_2r1w_792 vdd_uq18 gnd read_bl_0_51 read_bl_1_51 write_bl_0_51 wwl_0_39 rwl_1_39
+ rwl_0_39 cell_2r1w
Xcell_2r1w_1565 vdd_uq16 gnd read_bl_0_39 read_bl_1_39 write_bl_0_39 wwl_0_34 rwl_1_34
+ rwl_0_34 cell_2r1w
Xcell_2r1w_1598 vdd_uq0 gnd read_bl_0_39 read_bl_1_39 write_bl_0_39 wwl_0_1 rwl_1_1
+ rwl_0_1 cell_2r1w
Xcell_2r1w_1587 vdd_uq5 gnd read_bl_0_39 read_bl_1_39 write_bl_0_39 wwl_0_12 rwl_1_12
+ rwl_0_12 cell_2r1w
Xcell_2r1w_1576 vdd_uq10 gnd read_bl_0_39 read_bl_1_39 write_bl_0_39 wwl_0_23 rwl_1_23
+ rwl_0_23 cell_2r1w
Xcell_2r1w_3490 vdd_uq13 gnd read_bl_0_9 read_bl_1_9 write_bl_0_9 wwl_0_29 rwl_1_29
+ rwl_0_29 cell_2r1w
Xcell_2r1w_2052 vdd_uq28 gnd read_bl_0_31 read_bl_1_31 write_bl_0_31 wwl_0_59 rwl_1_59
+ rwl_0_59 cell_2r1w
Xcell_2r1w_1351 vdd_uq27 gnd read_bl_0_42 read_bl_1_42 write_bl_0_42 wwl_0_56 rwl_1_56
+ rwl_0_56 cell_2r1w
Xcell_2r1w_2063 vdd_uq23 gnd read_bl_0_31 read_bl_1_31 write_bl_0_31 wwl_0_48 rwl_1_48
+ rwl_0_48 cell_2r1w
Xcell_2r1w_1362 vdd_uq21 gnd read_bl_0_42 read_bl_1_42 write_bl_0_42 wwl_0_45 rwl_1_45
+ rwl_0_45 cell_2r1w
Xcell_2r1w_2074 vdd_uq17 gnd read_bl_0_31 read_bl_1_31 write_bl_0_31 wwl_0_37 rwl_1_37
+ rwl_0_37 cell_2r1w
Xcell_2r1w_1373 vdd_uq16 gnd read_bl_0_42 read_bl_1_42 write_bl_0_42 wwl_0_34 rwl_1_34
+ rwl_0_34 cell_2r1w
Xcell_2r1w_2085 vdd_uq12 gnd read_bl_0_31 read_bl_1_31 write_bl_0_31 wwl_0_26 rwl_1_26
+ rwl_0_26 cell_2r1w
Xcell_2r1w_1340 vdd gnd read_bl_0_43 read_bl_1_43 write_bl_0_43 wwl_0_3 rwl_1_3 rwl_0_3
+ cell_2r1w
Xcell_2r1w_2041 vdd_uq2 gnd read_bl_0_32 read_bl_1_32 write_bl_0_32 wwl_0_6 rwl_1_6
+ rwl_0_6 cell_2r1w
Xcell_2r1w_1395 vdd_uq5 gnd read_bl_0_42 read_bl_1_42 write_bl_0_42 wwl_0_12 rwl_1_12
+ rwl_0_12 cell_2r1w
Xcell_2r1w_2096 vdd_uq6 gnd read_bl_0_31 read_bl_1_31 write_bl_0_31 wwl_0_15 rwl_1_15
+ rwl_0_15 cell_2r1w
Xcell_2r1w_2030 vdd_uq7 gnd read_bl_0_32 read_bl_1_32 write_bl_0_32 wwl_0_17 rwl_1_17
+ rwl_0_17 cell_2r1w
Xcell_2r1w_1384 vdd_uq10 gnd read_bl_0_42 read_bl_1_42 write_bl_0_42 wwl_0_23 rwl_1_23
+ rwl_0_23 cell_2r1w
Xcell_2r1w_1170 vdd_uq21 gnd read_bl_0_45 read_bl_1_45 write_bl_0_45 wwl_0_45 rwl_1_45
+ rwl_0_45 cell_2r1w
Xcell_2r1w_1181 vdd_uq16 gnd read_bl_0_45 read_bl_1_45 write_bl_0_45 wwl_0_34 rwl_1_34
+ rwl_0_34 cell_2r1w
Xcell_2r1w_1192 vdd_uq10 gnd read_bl_0_45 read_bl_1_45 write_bl_0_45 wwl_0_23 rwl_1_23
+ rwl_0_23 cell_2r1w
Xcell_2r1w_2629 vdd_uq28 gnd read_bl_0_22 read_bl_1_22 write_bl_0_22 wwl_0_58 rwl_1_58
+ rwl_0_58 cell_2r1w
Xcell_2r1w_2618 vdd_uq1 gnd read_bl_0_23 read_bl_1_23 write_bl_0_23 wwl_0_5 rwl_1_5
+ rwl_0_5 cell_2r1w
Xcell_2r1w_3319 vdd_uq3 gnd read_bl_0_12 read_bl_1_12 write_bl_0_12 wwl_0_8 rwl_1_8
+ rwl_0_8 cell_2r1w
Xcell_2r1w_2607 vdd_uq7 gnd read_bl_0_23 read_bl_1_23 write_bl_0_23 wwl_0_16 rwl_1_16
+ rwl_0_16 cell_2r1w
Xcell_2r1w_3308 vdd_uq8 gnd read_bl_0_12 read_bl_1_12 write_bl_0_12 wwl_0_19 rwl_1_19
+ rwl_0_19 cell_2r1w
Xcell_2r1w_4009 vdd_uq10 gnd read_bl_0_1 read_bl_1_1 write_bl_0_1 wwl_0_22 rwl_1_22
+ rwl_0_22 cell_2r1w
Xcell_2r1w_1928 vdd_uq26 gnd read_bl_0_33 read_bl_1_33 write_bl_0_33 wwl_0_55 rwl_1_55
+ rwl_0_55 cell_2r1w
Xcell_2r1w_1939 vdd_uq21 gnd read_bl_0_33 read_bl_1_33 write_bl_0_33 wwl_0_44 rwl_1_44
+ rwl_0_44 cell_2r1w
Xcell_2r1w_1917 vdd gnd read_bl_0_34 read_bl_1_34 write_bl_0_34 wwl_0_2 rwl_1_2 rwl_0_2
+ cell_2r1w
Xcell_2r1w_1906 vdd_uq5 gnd read_bl_0_34 read_bl_1_34 write_bl_0_34 wwl_0_13 rwl_1_13
+ rwl_0_13 cell_2r1w
Xcell_2r1w_3842 vdd_uq29 gnd read_bl_0_3 read_bl_1_3 write_bl_0_3 wwl_0_61 rwl_1_61
+ rwl_0_61 cell_2r1w
Xcell_2r1w_3853 vdd_uq24 gnd read_bl_0_3 read_bl_1_3 write_bl_0_3 wwl_0_50 rwl_1_50
+ rwl_0_50 cell_2r1w
Xcell_2r1w_3864 vdd_uq18 gnd read_bl_0_3 read_bl_1_3 write_bl_0_3 wwl_0_39 rwl_1_39
+ rwl_0_39 cell_2r1w
Xcell_2r1w_3875 vdd_uq13 gnd read_bl_0_3 read_bl_1_3 write_bl_0_3 wwl_0_28 rwl_1_28
+ rwl_0_28 cell_2r1w
Xcell_2r1w_3897 vdd_uq2 gnd read_bl_0_3 read_bl_1_3 write_bl_0_3 wwl_0_6 rwl_1_6 rwl_0_6
+ cell_2r1w
Xcell_2r1w_3831 vdd_uq3 gnd read_bl_0_4 read_bl_1_4 write_bl_0_4 wwl_0_8 rwl_1_8 rwl_0_8
+ cell_2r1w
Xcell_2r1w_3886 vdd_uq7 gnd read_bl_0_3 read_bl_1_3 write_bl_0_3 wwl_0_17 rwl_1_17
+ rwl_0_17 cell_2r1w
Xcell_2r1w_3820 vdd_uq8 gnd read_bl_0_4 read_bl_1_4 write_bl_0_4 wwl_0_19 rwl_1_19
+ rwl_0_19 cell_2r1w
Xcell_2r1w_407 vdd_uq19 gnd read_bl_0_57 read_bl_1_57 write_bl_0_57 wwl_0_40 rwl_1_40
+ rwl_0_40 cell_2r1w
Xcell_2r1w_418 vdd_uq13 gnd read_bl_0_57 read_bl_1_57 write_bl_0_57 wwl_0_29 rwl_1_29
+ rwl_0_29 cell_2r1w
Xcell_2r1w_429 vdd_uq8 gnd read_bl_0_57 read_bl_1_57 write_bl_0_57 wwl_0_18 rwl_1_18
+ rwl_0_18 cell_2r1w
Xcell_2r1w_3138 vdd_uq29 gnd read_bl_0_14 read_bl_1_14 write_bl_0_14 wwl_0_61 rwl_1_61
+ rwl_0_61 cell_2r1w
Xcell_2r1w_2437 vdd_uq28 gnd read_bl_0_25 read_bl_1_25 write_bl_0_25 wwl_0_58 rwl_1_58
+ rwl_0_58 cell_2r1w
Xcell_2r1w_1736 vdd_uq26 gnd read_bl_0_36 read_bl_1_36 write_bl_0_36 wwl_0_55 rwl_1_55
+ rwl_0_55 cell_2r1w
Xcell_2r1w_3149 vdd_uq24 gnd read_bl_0_14 read_bl_1_14 write_bl_0_14 wwl_0_50 rwl_1_50
+ rwl_0_50 cell_2r1w
Xcell_2r1w_2448 vdd_uq22 gnd read_bl_0_25 read_bl_1_25 write_bl_0_25 wwl_0_47 rwl_1_47
+ rwl_0_47 cell_2r1w
Xcell_2r1w_2459 vdd_uq17 gnd read_bl_0_25 read_bl_1_25 write_bl_0_25 wwl_0_36 rwl_1_36
+ rwl_0_36 cell_2r1w
Xcell_2r1w_3105 vdd_uq14 gnd read_bl_0_15 read_bl_1_15 write_bl_0_15 wwl_0_30 rwl_1_30
+ rwl_0_30 cell_2r1w
Xcell_2r1w_2404 vdd_uq12 gnd read_bl_0_26 read_bl_1_26 write_bl_0_26 wwl_0_27 rwl_1_27
+ rwl_0_27 cell_2r1w
Xcell_2r1w_1703 vdd_uq11 gnd read_bl_0_37 read_bl_1_37 write_bl_0_37 wwl_0_24 rwl_1_24
+ rwl_0_24 cell_2r1w
Xcell_2r1w_2426 vdd_uq1 gnd read_bl_0_26 read_bl_1_26 write_bl_0_26 wwl_0_5 rwl_1_5
+ rwl_0_5 cell_2r1w
Xcell_2r1w_1725 vdd gnd read_bl_0_37 read_bl_1_37 write_bl_0_37 wwl_0_2 rwl_1_2 rwl_0_2
+ cell_2r1w
Xcell_2r1w_3127 vdd_uq3 gnd read_bl_0_15 read_bl_1_15 write_bl_0_15 wwl_0_8 rwl_1_8
+ rwl_0_8 cell_2r1w
Xcell_2r1w_1714 vdd_uq5 gnd read_bl_0_37 read_bl_1_37 write_bl_0_37 wwl_0_13 rwl_1_13
+ rwl_0_13 cell_2r1w
Xcell_2r1w_2415 vdd_uq7 gnd read_bl_0_26 read_bl_1_26 write_bl_0_26 wwl_0_16 rwl_1_16
+ rwl_0_16 cell_2r1w
Xcell_2r1w_3116 vdd_uq8 gnd read_bl_0_15 read_bl_1_15 write_bl_0_15 wwl_0_19 rwl_1_19
+ rwl_0_19 cell_2r1w
Xcell_2r1w_963 vdd_uq29 gnd read_bl_0_48 read_bl_1_48 write_bl_0_48 wwl_0_60 rwl_1_60
+ rwl_0_60 cell_2r1w
Xcell_2r1w_974 vdd_uq23 gnd read_bl_0_48 read_bl_1_48 write_bl_0_48 wwl_0_49 rwl_1_49
+ rwl_0_49 cell_2r1w
Xcell_2r1w_1747 vdd_uq21 gnd read_bl_0_36 read_bl_1_36 write_bl_0_36 wwl_0_44 rwl_1_44
+ rwl_0_44 cell_2r1w
Xcell_2r1w_985 vdd_uq18 gnd read_bl_0_48 read_bl_1_48 write_bl_0_48 wwl_0_38 rwl_1_38
+ rwl_0_38 cell_2r1w
Xcell_2r1w_1758 vdd_uq15 gnd read_bl_0_36 read_bl_1_36 write_bl_0_36 wwl_0_33 rwl_1_33
+ rwl_0_33 cell_2r1w
Xcell_2r1w_930 vdd_uq13 gnd read_bl_0_49 read_bl_1_49 write_bl_0_49 wwl_0_29 rwl_1_29
+ rwl_0_29 cell_2r1w
Xcell_2r1w_996 vdd_uq12 gnd read_bl_0_48 read_bl_1_48 write_bl_0_48 wwl_0_27 rwl_1_27
+ rwl_0_27 cell_2r1w
Xcell_2r1w_952 vdd_uq2 gnd read_bl_0_49 read_bl_1_49 write_bl_0_49 wwl_0_7 rwl_1_7
+ rwl_0_7 cell_2r1w
Xcell_2r1w_941 vdd_uq8 gnd read_bl_0_49 read_bl_1_49 write_bl_0_49 wwl_0_18 rwl_1_18
+ rwl_0_18 cell_2r1w
Xcell_2r1w_1769 vdd_uq10 gnd read_bl_0_36 read_bl_1_36 write_bl_0_36 wwl_0_22 rwl_1_22
+ rwl_0_22 cell_2r1w
Xcell_2r1w_3650 vdd_uq29 gnd read_bl_0_6 read_bl_1_6 write_bl_0_6 wwl_0_61 rwl_1_61
+ rwl_0_61 cell_2r1w
Xcell_2r1w_3661 vdd_uq24 gnd read_bl_0_6 read_bl_1_6 write_bl_0_6 wwl_0_50 rwl_1_50
+ rwl_0_50 cell_2r1w
Xcell_2r1w_2960 vdd_uq22 gnd read_bl_0_17 read_bl_1_17 write_bl_0_17 wwl_0_47 rwl_1_47
+ rwl_0_47 cell_2r1w
Xcell_2r1w_3672 vdd_uq18 gnd read_bl_0_6 read_bl_1_6 write_bl_0_6 wwl_0_39 rwl_1_39
+ rwl_0_39 cell_2r1w
Xcell_2r1w_2971 vdd_uq17 gnd read_bl_0_17 read_bl_1_17 write_bl_0_17 wwl_0_36 rwl_1_36
+ rwl_0_36 cell_2r1w
Xcell_2r1w_3683 vdd_uq13 gnd read_bl_0_6 read_bl_1_6 write_bl_0_6 wwl_0_28 rwl_1_28
+ rwl_0_28 cell_2r1w
Xcell_2r1w_2982 vdd_uq11 gnd read_bl_0_17 read_bl_1_17 write_bl_0_17 wwl_0_25 rwl_1_25
+ rwl_0_25 cell_2r1w
Xcell_2r1w_2993 vdd_uq6 gnd read_bl_0_17 read_bl_1_17 write_bl_0_17 wwl_0_14 rwl_1_14
+ rwl_0_14 cell_2r1w
Xcell_2r1w_3694 vdd_uq7 gnd read_bl_0_6 read_bl_1_6 write_bl_0_6 wwl_0_17 rwl_1_17
+ rwl_0_17 cell_2r1w
Xcell_2r1w_64 vdd_uq30 gnd read_bl_0_62 read_bl_1_62 write_bl_0_62 wwl_0_63 rwl_1_63
+ rwl_0_63 cell_2r1w
Xcell_2r1w_20 vdd_uq20 gnd read_bl_0_63 read_bl_1_63 write_bl_0_63 wwl_0_43 rwl_1_43
+ rwl_0_43 cell_2r1w
Xcell_2r1w_31 vdd_uq15 gnd read_bl_0_63 read_bl_1_63 write_bl_0_63 wwl_0_32 rwl_1_32
+ rwl_0_32 cell_2r1w
Xcell_2r1w_53 vdd_uq4 gnd read_bl_0_63 read_bl_1_63 write_bl_0_63 wwl_0_10 rwl_1_10
+ rwl_0_10 cell_2r1w
Xcell_2r1w_42 vdd_uq9 gnd read_bl_0_63 read_bl_1_63 write_bl_0_63 wwl_0_21 rwl_1_21
+ rwl_0_21 cell_2r1w
Xcell_2r1w_75 vdd_uq25 gnd read_bl_0_62 read_bl_1_62 write_bl_0_62 wwl_0_52 rwl_1_52
+ rwl_0_52 cell_2r1w
Xcell_2r1w_86 vdd_uq19 gnd read_bl_0_62 read_bl_1_62 write_bl_0_62 wwl_0_41 rwl_1_41
+ rwl_0_41 cell_2r1w
Xcell_2r1w_97 vdd_uq14 gnd read_bl_0_62 read_bl_1_62 write_bl_0_62 wwl_0_30 rwl_1_30
+ rwl_0_30 cell_2r1w
Xcell_2r1w_259 vdd_uq29 gnd read_bl_0_59 read_bl_1_59 write_bl_0_59 wwl_0_60 rwl_1_60
+ rwl_0_60 cell_2r1w
Xcell_2r1w_204 vdd_uq24 gnd read_bl_0_60 read_bl_1_60 write_bl_0_60 wwl_0_51 rwl_1_51
+ rwl_0_51 cell_2r1w
Xcell_2r1w_215 vdd_uq19 gnd read_bl_0_60 read_bl_1_60 write_bl_0_60 wwl_0_40 rwl_1_40
+ rwl_0_40 cell_2r1w
Xcell_2r1w_226 vdd_uq13 gnd read_bl_0_60 read_bl_1_60 write_bl_0_60 wwl_0_29 rwl_1_29
+ rwl_0_29 cell_2r1w
Xcell_2r1w_248 vdd_uq2 gnd read_bl_0_60 read_bl_1_60 write_bl_0_60 wwl_0_7 rwl_1_7
+ rwl_0_7 cell_2r1w
Xcell_2r1w_237 vdd_uq8 gnd read_bl_0_60 read_bl_1_60 write_bl_0_60 wwl_0_18 rwl_1_18
+ rwl_0_18 cell_2r1w
Xcell_2r1w_2245 vdd_uq28 gnd read_bl_0_28 read_bl_1_28 write_bl_0_28 wwl_0_58 rwl_1_58
+ rwl_0_58 cell_2r1w
Xcell_2r1w_1544 vdd_uq26 gnd read_bl_0_39 read_bl_1_39 write_bl_0_39 wwl_0_55 rwl_1_55
+ rwl_0_55 cell_2r1w
Xcell_2r1w_2256 vdd_uq22 gnd read_bl_0_28 read_bl_1_28 write_bl_0_28 wwl_0_47 rwl_1_47
+ rwl_0_47 cell_2r1w
Xcell_2r1w_1555 vdd_uq21 gnd read_bl_0_39 read_bl_1_39 write_bl_0_39 wwl_0_44 rwl_1_44
+ rwl_0_44 cell_2r1w
Xcell_2r1w_2201 vdd_uq18 gnd read_bl_0_29 read_bl_1_29 write_bl_0_29 wwl_0_38 rwl_1_38
+ rwl_0_38 cell_2r1w
Xcell_2r1w_2267 vdd_uq17 gnd read_bl_0_28 read_bl_1_28 write_bl_0_28 wwl_0_36 rwl_1_36
+ rwl_0_36 cell_2r1w
Xcell_2r1w_1500 vdd_uq16 gnd read_bl_0_40 read_bl_1_40 write_bl_0_40 wwl_0_35 rwl_1_35
+ rwl_0_35 cell_2r1w
Xcell_2r1w_1566 vdd_uq15 gnd read_bl_0_39 read_bl_1_39 write_bl_0_39 wwl_0_33 rwl_1_33
+ rwl_0_33 cell_2r1w
Xcell_2r1w_2212 vdd_uq12 gnd read_bl_0_29 read_bl_1_29 write_bl_0_29 wwl_0_27 rwl_1_27
+ rwl_0_27 cell_2r1w
Xcell_2r1w_2278 vdd_uq11 gnd read_bl_0_28 read_bl_1_28 write_bl_0_28 wwl_0_25 rwl_1_25
+ rwl_0_25 cell_2r1w
Xcell_2r1w_1511 vdd_uq11 gnd read_bl_0_40 read_bl_1_40 write_bl_0_40 wwl_0_24 rwl_1_24
+ rwl_0_24 cell_2r1w
Xcell_2r1w_2234 vdd_uq1 gnd read_bl_0_29 read_bl_1_29 write_bl_0_29 wwl_0_5 rwl_1_5
+ rwl_0_5 cell_2r1w
Xcell_2r1w_1533 vdd gnd read_bl_0_40 read_bl_1_40 write_bl_0_40 wwl_0_2 rwl_1_2 rwl_0_2
+ cell_2r1w
Xcell_2r1w_1588 vdd_uq4 gnd read_bl_0_39 read_bl_1_39 write_bl_0_39 wwl_0_11 rwl_1_11
+ rwl_0_11 cell_2r1w
Xcell_2r1w_2289 vdd_uq6 gnd read_bl_0_28 read_bl_1_28 write_bl_0_28 wwl_0_14 rwl_1_14
+ rwl_0_14 cell_2r1w
Xcell_2r1w_1522 vdd_uq5 gnd read_bl_0_40 read_bl_1_40 write_bl_0_40 wwl_0_13 rwl_1_13
+ rwl_0_13 cell_2r1w
Xcell_2r1w_2223 vdd_uq7 gnd read_bl_0_29 read_bl_1_29 write_bl_0_29 wwl_0_16 rwl_1_16
+ rwl_0_16 cell_2r1w
Xcell_2r1w_1577 vdd_uq10 gnd read_bl_0_39 read_bl_1_39 write_bl_0_39 wwl_0_22 rwl_1_22
+ rwl_0_22 cell_2r1w
Xcell_2r1w_771 vdd_uq29 gnd read_bl_0_51 read_bl_1_51 write_bl_0_51 wwl_0_60 rwl_1_60
+ rwl_0_60 cell_2r1w
Xcell_2r1w_782 vdd_uq23 gnd read_bl_0_51 read_bl_1_51 write_bl_0_51 wwl_0_49 rwl_1_49
+ rwl_0_49 cell_2r1w
Xcell_2r1w_793 vdd_uq18 gnd read_bl_0_51 read_bl_1_51 write_bl_0_51 wwl_0_38 rwl_1_38
+ rwl_0_38 cell_2r1w
Xcell_2r1w_1599 vdd_uq0 gnd read_bl_0_39 read_bl_1_39 write_bl_0_39 wwl_0_0 rwl_1_0
+ rwl_0_0 cell_2r1w
Xcell_2r1w_760 vdd_uq2 gnd read_bl_0_52 read_bl_1_52 write_bl_0_52 wwl_0_7 rwl_1_7
+ rwl_0_7 cell_2r1w
Xcell_2r1w_3480 vdd_uq18 gnd read_bl_0_9 read_bl_1_9 write_bl_0_9 wwl_0_39 rwl_1_39
+ rwl_0_39 cell_2r1w
Xcell_2r1w_3491 vdd_uq13 gnd read_bl_0_9 read_bl_1_9 write_bl_0_9 wwl_0_28 rwl_1_28
+ rwl_0_28 cell_2r1w
Xcell_2r1w_2790 vdd_uq11 gnd read_bl_0_20 read_bl_1_20 write_bl_0_20 wwl_0_25 rwl_1_25
+ rwl_0_25 cell_2r1w
Xcell_2r1w_2020 vdd_uq12 gnd read_bl_0_32 read_bl_1_32 write_bl_0_32 wwl_0_27 rwl_1_27
+ rwl_0_27 cell_2r1w
Xcell_2r1w_2031 vdd_uq7 gnd read_bl_0_32 read_bl_1_32 write_bl_0_32 wwl_0_16 rwl_1_16
+ rwl_0_16 cell_2r1w
Xcell_2r1w_2053 vdd_uq28 gnd read_bl_0_31 read_bl_1_31 write_bl_0_31 wwl_0_58 rwl_1_58
+ rwl_0_58 cell_2r1w
Xcell_2r1w_1352 vdd_uq26 gnd read_bl_0_42 read_bl_1_42 write_bl_0_42 wwl_0_55 rwl_1_55
+ rwl_0_55 cell_2r1w
Xcell_2r1w_590 vdd_uq23 gnd read_bl_0_54 read_bl_1_54 write_bl_0_54 wwl_0_49 rwl_1_49
+ rwl_0_49 cell_2r1w
Xcell_2r1w_2064 vdd_uq22 gnd read_bl_0_31 read_bl_1_31 write_bl_0_31 wwl_0_47 rwl_1_47
+ rwl_0_47 cell_2r1w
Xcell_2r1w_1363 vdd_uq21 gnd read_bl_0_42 read_bl_1_42 write_bl_0_42 wwl_0_44 rwl_1_44
+ rwl_0_44 cell_2r1w
Xcell_2r1w_2075 vdd_uq17 gnd read_bl_0_31 read_bl_1_31 write_bl_0_31 wwl_0_36 rwl_1_36
+ rwl_0_36 cell_2r1w
Xcell_2r1w_1374 vdd_uq15 gnd read_bl_0_42 read_bl_1_42 write_bl_0_42 wwl_0_33 rwl_1_33
+ rwl_0_33 cell_2r1w
Xcell_2r1w_2086 vdd_uq11 gnd read_bl_0_31 read_bl_1_31 write_bl_0_31 wwl_0_25 rwl_1_25
+ rwl_0_25 cell_2r1w
Xcell_2r1w_2042 vdd_uq1 gnd read_bl_0_32 read_bl_1_32 write_bl_0_32 wwl_0_5 rwl_1_5
+ rwl_0_5 cell_2r1w
Xcell_2r1w_1341 vdd gnd read_bl_0_43 read_bl_1_43 write_bl_0_43 wwl_0_2 rwl_1_2 rwl_0_2
+ cell_2r1w
Xcell_2r1w_1396 vdd_uq4 gnd read_bl_0_42 read_bl_1_42 write_bl_0_42 wwl_0_11 rwl_1_11
+ rwl_0_11 cell_2r1w
Xcell_2r1w_2097 vdd_uq6 gnd read_bl_0_31 read_bl_1_31 write_bl_0_31 wwl_0_14 rwl_1_14
+ rwl_0_14 cell_2r1w
Xcell_2r1w_1330 vdd_uq5 gnd read_bl_0_43 read_bl_1_43 write_bl_0_43 wwl_0_13 rwl_1_13
+ rwl_0_13 cell_2r1w
Xcell_2r1w_1385 vdd_uq10 gnd read_bl_0_42 read_bl_1_42 write_bl_0_42 wwl_0_22 rwl_1_22
+ rwl_0_22 cell_2r1w
Xcell_2r1w_1160 vdd_uq26 gnd read_bl_0_45 read_bl_1_45 write_bl_0_45 wwl_0_55 rwl_1_55
+ rwl_0_55 cell_2r1w
Xcell_2r1w_1171 vdd_uq21 gnd read_bl_0_45 read_bl_1_45 write_bl_0_45 wwl_0_44 rwl_1_44
+ rwl_0_44 cell_2r1w
Xcell_2r1w_1182 vdd_uq15 gnd read_bl_0_45 read_bl_1_45 write_bl_0_45 wwl_0_33 rwl_1_33
+ rwl_0_33 cell_2r1w
Xcell_2r1w_1193 vdd_uq10 gnd read_bl_0_45 read_bl_1_45 write_bl_0_45 wwl_0_22 rwl_1_22
+ rwl_0_22 cell_2r1w
Xcell_2r1w_2619 vdd_uq1 gnd read_bl_0_23 read_bl_1_23 write_bl_0_23 wwl_0_4 rwl_1_4
+ rwl_0_4 cell_2r1w
Xcell_2r1w_1918 vdd_uq0 gnd read_bl_0_34 read_bl_1_34 write_bl_0_34 wwl_0_1 rwl_1_1
+ rwl_0_1 cell_2r1w
Xcell_2r1w_1907 vdd_uq5 gnd read_bl_0_34 read_bl_1_34 write_bl_0_34 wwl_0_12 rwl_1_12
+ rwl_0_12 cell_2r1w
Xcell_2r1w_2608 vdd_uq6 gnd read_bl_0_23 read_bl_1_23 write_bl_0_23 wwl_0_15 rwl_1_15
+ rwl_0_15 cell_2r1w
Xcell_2r1w_3309 vdd_uq8 gnd read_bl_0_12 read_bl_1_12 write_bl_0_12 wwl_0_18 rwl_1_18
+ rwl_0_18 cell_2r1w
Xcell_2r1w_1929 vdd_uq26 gnd read_bl_0_33 read_bl_1_33 write_bl_0_33 wwl_0_54 rwl_1_54
+ rwl_0_54 cell_2r1w
Xcell_2r1w_3810 vdd_uq13 gnd read_bl_0_4 read_bl_1_4 write_bl_0_4 wwl_0_29 rwl_1_29
+ rwl_0_29 cell_2r1w
Xcell_2r1w_3821 vdd_uq8 gnd read_bl_0_4 read_bl_1_4 write_bl_0_4 wwl_0_18 rwl_1_18
+ rwl_0_18 cell_2r1w
Xcell_2r1w_3843 vdd_uq29 gnd read_bl_0_3 read_bl_1_3 write_bl_0_3 wwl_0_60 rwl_1_60
+ rwl_0_60 cell_2r1w
Xcell_2r1w_3854 vdd_uq23 gnd read_bl_0_3 read_bl_1_3 write_bl_0_3 wwl_0_49 rwl_1_49
+ rwl_0_49 cell_2r1w
Xcell_2r1w_3865 vdd_uq18 gnd read_bl_0_3 read_bl_1_3 write_bl_0_3 wwl_0_38 rwl_1_38
+ rwl_0_38 cell_2r1w
Xcell_2r1w_3876 vdd_uq12 gnd read_bl_0_3 read_bl_1_3 write_bl_0_3 wwl_0_27 rwl_1_27
+ rwl_0_27 cell_2r1w
Xcell_2r1w_3898 vdd_uq1 gnd read_bl_0_3 read_bl_1_3 write_bl_0_3 wwl_0_5 rwl_1_5 rwl_0_5
+ cell_2r1w
Xcell_2r1w_3832 vdd_uq2 gnd read_bl_0_4 read_bl_1_4 write_bl_0_4 wwl_0_7 rwl_1_7 rwl_0_7
+ cell_2r1w
Xcell_2r1w_3887 vdd_uq7 gnd read_bl_0_3 read_bl_1_3 write_bl_0_3 wwl_0_16 rwl_1_16
+ rwl_0_16 cell_2r1w
Xcell_2r1w_408 vdd_uq18 gnd read_bl_0_57 read_bl_1_57 write_bl_0_57 wwl_0_39 rwl_1_39
+ rwl_0_39 cell_2r1w
Xcell_2r1w_419 vdd_uq13 gnd read_bl_0_57 read_bl_1_57 write_bl_0_57 wwl_0_28 rwl_1_28
+ rwl_0_28 cell_2r1w
Xcell_2r1w_3106 vdd_uq13 gnd read_bl_0_15 read_bl_1_15 write_bl_0_15 wwl_0_29 rwl_1_29
+ rwl_0_29 cell_2r1w
Xcell_2r1w_3139 vdd_uq29 gnd read_bl_0_14 read_bl_1_14 write_bl_0_14 wwl_0_60 rwl_1_60
+ rwl_0_60 cell_2r1w
Xcell_2r1w_2438 vdd_uq27 gnd read_bl_0_25 read_bl_1_25 write_bl_0_25 wwl_0_57 rwl_1_57
+ rwl_0_57 cell_2r1w
Xcell_2r1w_1737 vdd_uq26 gnd read_bl_0_36 read_bl_1_36 write_bl_0_36 wwl_0_54 rwl_1_54
+ rwl_0_54 cell_2r1w
Xcell_2r1w_2449 vdd_uq22 gnd read_bl_0_25 read_bl_1_25 write_bl_0_25 wwl_0_46 rwl_1_46
+ rwl_0_46 cell_2r1w
Xcell_2r1w_1748 vdd_uq20 gnd read_bl_0_36 read_bl_1_36 write_bl_0_36 wwl_0_43 rwl_1_43
+ rwl_0_43 cell_2r1w
Xcell_2r1w_920 vdd_uq18 gnd read_bl_0_49 read_bl_1_49 write_bl_0_49 wwl_0_39 rwl_1_39
+ rwl_0_39 cell_2r1w
Xcell_2r1w_1759 vdd_uq15 gnd read_bl_0_36 read_bl_1_36 write_bl_0_36 wwl_0_32 rwl_1_32
+ rwl_0_32 cell_2r1w
Xcell_2r1w_931 vdd_uq13 gnd read_bl_0_49 read_bl_1_49 write_bl_0_49 wwl_0_28 rwl_1_28
+ rwl_0_28 cell_2r1w
Xcell_2r1w_2405 vdd_uq12 gnd read_bl_0_26 read_bl_1_26 write_bl_0_26 wwl_0_26 rwl_1_26
+ rwl_0_26 cell_2r1w
Xcell_2r1w_2427 vdd_uq1 gnd read_bl_0_26 read_bl_1_26 write_bl_0_26 wwl_0_4 rwl_1_4
+ rwl_0_4 cell_2r1w
Xcell_2r1w_1726 vdd_uq0 gnd read_bl_0_37 read_bl_1_37 write_bl_0_37 wwl_0_1 rwl_1_1
+ rwl_0_1 cell_2r1w
Xcell_2r1w_3128 vdd_uq2 gnd read_bl_0_15 read_bl_1_15 write_bl_0_15 wwl_0_7 rwl_1_7
+ rwl_0_7 cell_2r1w
Xcell_2r1w_1715 vdd_uq5 gnd read_bl_0_37 read_bl_1_37 write_bl_0_37 wwl_0_12 rwl_1_12
+ rwl_0_12 cell_2r1w
Xcell_2r1w_2416 vdd_uq6 gnd read_bl_0_26 read_bl_1_26 write_bl_0_26 wwl_0_15 rwl_1_15
+ rwl_0_15 cell_2r1w
Xcell_2r1w_3117 vdd_uq8 gnd read_bl_0_15 read_bl_1_15 write_bl_0_15 wwl_0_18 rwl_1_18
+ rwl_0_18 cell_2r1w
Xcell_2r1w_1704 vdd_uq10 gnd read_bl_0_37 read_bl_1_37 write_bl_0_37 wwl_0_23 rwl_1_23
+ rwl_0_23 cell_2r1w
Xcell_2r1w_964 vdd_uq28 gnd read_bl_0_48 read_bl_1_48 write_bl_0_48 wwl_0_59 rwl_1_59
+ rwl_0_59 cell_2r1w
Xcell_2r1w_975 vdd_uq23 gnd read_bl_0_48 read_bl_1_48 write_bl_0_48 wwl_0_48 rwl_1_48
+ rwl_0_48 cell_2r1w
Xcell_2r1w_986 vdd_uq17 gnd read_bl_0_48 read_bl_1_48 write_bl_0_48 wwl_0_37 rwl_1_37
+ rwl_0_37 cell_2r1w
Xcell_2r1w_997 vdd_uq12 gnd read_bl_0_48 read_bl_1_48 write_bl_0_48 wwl_0_26 rwl_1_26
+ rwl_0_26 cell_2r1w
Xcell_2r1w_953 vdd_uq2 gnd read_bl_0_49 read_bl_1_49 write_bl_0_49 wwl_0_6 rwl_1_6
+ rwl_0_6 cell_2r1w
Xcell_2r1w_942 vdd_uq7 gnd read_bl_0_49 read_bl_1_49 write_bl_0_49 wwl_0_17 rwl_1_17
+ rwl_0_17 cell_2r1w
Xcell_2r1w_3651 vdd_uq29 gnd read_bl_0_6 read_bl_1_6 write_bl_0_6 wwl_0_60 rwl_1_60
+ rwl_0_60 cell_2r1w
Xcell_2r1w_3662 vdd_uq23 gnd read_bl_0_6 read_bl_1_6 write_bl_0_6 wwl_0_49 rwl_1_49
+ rwl_0_49 cell_2r1w
Xcell_2r1w_3640 vdd_uq2 gnd read_bl_0_7 read_bl_1_7 write_bl_0_7 wwl_0_7 rwl_1_7 rwl_0_7
+ cell_2r1w
Xcell_2r1w_2950 vdd_uq27 gnd read_bl_0_17 read_bl_1_17 write_bl_0_17 wwl_0_57 rwl_1_57
+ rwl_0_57 cell_2r1w
Xcell_2r1w_2961 vdd_uq22 gnd read_bl_0_17 read_bl_1_17 write_bl_0_17 wwl_0_46 rwl_1_46
+ rwl_0_46 cell_2r1w
Xcell_2r1w_3673 vdd_uq18 gnd read_bl_0_6 read_bl_1_6 write_bl_0_6 wwl_0_38 rwl_1_38
+ rwl_0_38 cell_2r1w
Xcell_2r1w_2972 vdd_uq16 gnd read_bl_0_17 read_bl_1_17 write_bl_0_17 wwl_0_35 rwl_1_35
+ rwl_0_35 cell_2r1w
Xcell_2r1w_3684 vdd_uq12 gnd read_bl_0_6 read_bl_1_6 write_bl_0_6 wwl_0_27 rwl_1_27
+ rwl_0_27 cell_2r1w
Xcell_2r1w_2983 vdd_uq11 gnd read_bl_0_17 read_bl_1_17 write_bl_0_17 wwl_0_24 rwl_1_24
+ rwl_0_24 cell_2r1w
Xcell_2r1w_2994 vdd_uq5 gnd read_bl_0_17 read_bl_1_17 write_bl_0_17 wwl_0_13 rwl_1_13
+ rwl_0_13 cell_2r1w
Xcell_2r1w_3695 vdd_uq7 gnd read_bl_0_6 read_bl_1_6 write_bl_0_6 wwl_0_16 rwl_1_16
+ rwl_0_16 cell_2r1w
Xcell_2r1w_65 vdd_uq30 gnd read_bl_0_62 read_bl_1_62 write_bl_0_62 wwl_0_62 rwl_1_62
+ rwl_0_62 cell_2r1w
Xcell_2r1w_10 vdd_uq25 gnd read_bl_0_63 read_bl_1_63 write_bl_0_63 wwl_0_53 rwl_1_53
+ rwl_0_53 cell_2r1w
Xcell_2r1w_76 vdd_uq24 gnd read_bl_0_62 read_bl_1_62 write_bl_0_62 wwl_0_51 rwl_1_51
+ rwl_0_51 cell_2r1w
Xcell_2r1w_21 vdd_uq20 gnd read_bl_0_63 read_bl_1_63 write_bl_0_63 wwl_0_42 rwl_1_42
+ rwl_0_42 cell_2r1w
Xcell_2r1w_87 vdd_uq19 gnd read_bl_0_62 read_bl_1_62 write_bl_0_62 wwl_0_40 rwl_1_40
+ rwl_0_40 cell_2r1w
Xcell_2r1w_32 vdd_uq14 gnd read_bl_0_63 read_bl_1_63 write_bl_0_63 wwl_0_31 rwl_1_31
+ rwl_0_31 cell_2r1w
Xcell_2r1w_98 vdd_uq13 gnd read_bl_0_62 read_bl_1_62 write_bl_0_62 wwl_0_29 rwl_1_29
+ rwl_0_29 cell_2r1w
Xcell_2r1w_54 vdd_uq3 gnd read_bl_0_63 read_bl_1_63 write_bl_0_63 wwl_0_9 rwl_1_9
+ rwl_0_9 cell_2r1w
Xcell_2r1w_43 vdd_uq9 gnd read_bl_0_63 read_bl_1_63 write_bl_0_63 wwl_0_20 rwl_1_20
+ rwl_0_20 cell_2r1w
Xcell_2r1w_205 vdd_uq24 gnd read_bl_0_60 read_bl_1_60 write_bl_0_60 wwl_0_50 rwl_1_50
+ rwl_0_50 cell_2r1w
Xcell_2r1w_216 vdd_uq18 gnd read_bl_0_60 read_bl_1_60 write_bl_0_60 wwl_0_39 rwl_1_39
+ rwl_0_39 cell_2r1w
Xcell_2r1w_227 vdd_uq13 gnd read_bl_0_60 read_bl_1_60 write_bl_0_60 wwl_0_28 rwl_1_28
+ rwl_0_28 cell_2r1w
Xcell_2r1w_249 vdd_uq2 gnd read_bl_0_60 read_bl_1_60 write_bl_0_60 wwl_0_6 rwl_1_6
+ rwl_0_6 cell_2r1w
Xcell_2r1w_238 vdd_uq7 gnd read_bl_0_60 read_bl_1_60 write_bl_0_60 wwl_0_17 rwl_1_17
+ rwl_0_17 cell_2r1w
Xcell_2r1w_2202 vdd_uq17 gnd read_bl_0_29 read_bl_1_29 write_bl_0_29 wwl_0_37 rwl_1_37
+ rwl_0_37 cell_2r1w
Xcell_2r1w_2213 vdd_uq12 gnd read_bl_0_29 read_bl_1_29 write_bl_0_29 wwl_0_26 rwl_1_26
+ rwl_0_26 cell_2r1w
Xcell_2r1w_772 vdd_uq28 gnd read_bl_0_51 read_bl_1_51 write_bl_0_51 wwl_0_59 rwl_1_59
+ rwl_0_59 cell_2r1w
Xcell_2r1w_2246 vdd_uq27 gnd read_bl_0_28 read_bl_1_28 write_bl_0_28 wwl_0_57 rwl_1_57
+ rwl_0_57 cell_2r1w
Xcell_2r1w_1545 vdd_uq26 gnd read_bl_0_39 read_bl_1_39 write_bl_0_39 wwl_0_54 rwl_1_54
+ rwl_0_54 cell_2r1w
Xcell_2r1w_2257 vdd_uq22 gnd read_bl_0_28 read_bl_1_28 write_bl_0_28 wwl_0_46 rwl_1_46
+ rwl_0_46 cell_2r1w
Xcell_2r1w_1556 vdd_uq20 gnd read_bl_0_39 read_bl_1_39 write_bl_0_39 wwl_0_43 rwl_1_43
+ rwl_0_43 cell_2r1w
Xcell_2r1w_2268 vdd_uq16 gnd read_bl_0_28 read_bl_1_28 write_bl_0_28 wwl_0_35 rwl_1_35
+ rwl_0_35 cell_2r1w
Xcell_2r1w_1501 vdd_uq16 gnd read_bl_0_40 read_bl_1_40 write_bl_0_40 wwl_0_34 rwl_1_34
+ rwl_0_34 cell_2r1w
Xcell_2r1w_1567 vdd_uq15 gnd read_bl_0_39 read_bl_1_39 write_bl_0_39 wwl_0_32 rwl_1_32
+ rwl_0_32 cell_2r1w
Xcell_2r1w_2279 vdd_uq11 gnd read_bl_0_28 read_bl_1_28 write_bl_0_28 wwl_0_24 rwl_1_24
+ rwl_0_24 cell_2r1w
Xcell_2r1w_2235 vdd_uq1 gnd read_bl_0_29 read_bl_1_29 write_bl_0_29 wwl_0_4 rwl_1_4
+ rwl_0_4 cell_2r1w
Xcell_2r1w_1534 vdd_uq0 gnd read_bl_0_40 read_bl_1_40 write_bl_0_40 wwl_0_1 rwl_1_1
+ rwl_0_1 cell_2r1w
Xcell_2r1w_761 vdd_uq2 gnd read_bl_0_52 read_bl_1_52 write_bl_0_52 wwl_0_6 rwl_1_6
+ rwl_0_6 cell_2r1w
Xcell_2r1w_1589 vdd_uq4 gnd read_bl_0_39 read_bl_1_39 write_bl_0_39 wwl_0_10 rwl_1_10
+ rwl_0_10 cell_2r1w
Xcell_2r1w_1523 vdd_uq5 gnd read_bl_0_40 read_bl_1_40 write_bl_0_40 wwl_0_12 rwl_1_12
+ rwl_0_12 cell_2r1w
Xcell_2r1w_2224 vdd_uq6 gnd read_bl_0_29 read_bl_1_29 write_bl_0_29 wwl_0_15 rwl_1_15
+ rwl_0_15 cell_2r1w
Xcell_2r1w_750 vdd_uq7 gnd read_bl_0_52 read_bl_1_52 write_bl_0_52 wwl_0_17 rwl_1_17
+ rwl_0_17 cell_2r1w
Xcell_2r1w_1578 vdd_uq9 gnd read_bl_0_39 read_bl_1_39 write_bl_0_39 wwl_0_21 rwl_1_21
+ rwl_0_21 cell_2r1w
Xcell_2r1w_1512 vdd_uq10 gnd read_bl_0_40 read_bl_1_40 write_bl_0_40 wwl_0_23 rwl_1_23
+ rwl_0_23 cell_2r1w
Xcell_2r1w_783 vdd_uq23 gnd read_bl_0_51 read_bl_1_51 write_bl_0_51 wwl_0_48 rwl_1_48
+ rwl_0_48 cell_2r1w
Xcell_2r1w_794 vdd_uq17 gnd read_bl_0_51 read_bl_1_51 write_bl_0_51 wwl_0_37 rwl_1_37
+ rwl_0_37 cell_2r1w
Xcell_2r1w_0 vdd_uq30 gnd read_bl_0_63 read_bl_1_63 write_bl_0_63 wwl_0_63 rwl_1_63
+ rwl_0_63 cell_2r1w
Xcell_2r1w_3470 vdd_uq23 gnd read_bl_0_9 read_bl_1_9 write_bl_0_9 wwl_0_49 rwl_1_49
+ rwl_0_49 cell_2r1w
Xcell_2r1w_3481 vdd_uq18 gnd read_bl_0_9 read_bl_1_9 write_bl_0_9 wwl_0_38 rwl_1_38
+ rwl_0_38 cell_2r1w
Xcell_2r1w_3492 vdd_uq12 gnd read_bl_0_9 read_bl_1_9 write_bl_0_9 wwl_0_27 rwl_1_27
+ rwl_0_27 cell_2r1w
Xcell_2r1w_2780 vdd_uq16 gnd read_bl_0_20 read_bl_1_20 write_bl_0_20 wwl_0_35 rwl_1_35
+ rwl_0_35 cell_2r1w
Xcell_2r1w_2791 vdd_uq11 gnd read_bl_0_20 read_bl_1_20 write_bl_0_20 wwl_0_24 rwl_1_24
+ rwl_0_24 cell_2r1w
Xcell_2r1w_2054 vdd_uq27 gnd read_bl_0_31 read_bl_1_31 write_bl_0_31 wwl_0_57 rwl_1_57
+ rwl_0_57 cell_2r1w
Xcell_2r1w_2065 vdd_uq22 gnd read_bl_0_31 read_bl_1_31 write_bl_0_31 wwl_0_46 rwl_1_46
+ rwl_0_46 cell_2r1w
Xcell_2r1w_2010 vdd_uq17 gnd read_bl_0_32 read_bl_1_32 write_bl_0_32 wwl_0_37 rwl_1_37
+ rwl_0_37 cell_2r1w
Xcell_2r1w_2021 vdd_uq12 gnd read_bl_0_32 read_bl_1_32 write_bl_0_32 wwl_0_26 rwl_1_26
+ rwl_0_26 cell_2r1w
Xcell_2r1w_2043 vdd_uq1 gnd read_bl_0_32 read_bl_1_32 write_bl_0_32 wwl_0_4 rwl_1_4
+ rwl_0_4 cell_2r1w
Xcell_2r1w_2032 vdd_uq6 gnd read_bl_0_32 read_bl_1_32 write_bl_0_32 wwl_0_15 rwl_1_15
+ rwl_0_15 cell_2r1w
Xcell_2r1w_1320 vdd_uq10 gnd read_bl_0_43 read_bl_1_43 write_bl_0_43 wwl_0_23 rwl_1_23
+ rwl_0_23 cell_2r1w
Xcell_2r1w_580 vdd_uq28 gnd read_bl_0_54 read_bl_1_54 write_bl_0_54 wwl_0_59 rwl_1_59
+ rwl_0_59 cell_2r1w
Xcell_2r1w_1353 vdd_uq26 gnd read_bl_0_42 read_bl_1_42 write_bl_0_42 wwl_0_54 rwl_1_54
+ rwl_0_54 cell_2r1w
Xcell_2r1w_591 vdd_uq23 gnd read_bl_0_54 read_bl_1_54 write_bl_0_54 wwl_0_48 rwl_1_48
+ rwl_0_48 cell_2r1w
Xcell_2r1w_1364 vdd_uq20 gnd read_bl_0_42 read_bl_1_42 write_bl_0_42 wwl_0_43 rwl_1_43
+ rwl_0_43 cell_2r1w
Xcell_2r1w_2076 vdd_uq16 gnd read_bl_0_31 read_bl_1_31 write_bl_0_31 wwl_0_35 rwl_1_35
+ rwl_0_35 cell_2r1w
Xcell_2r1w_1375 vdd_uq15 gnd read_bl_0_42 read_bl_1_42 write_bl_0_42 wwl_0_32 rwl_1_32
+ rwl_0_32 cell_2r1w
Xcell_2r1w_2087 vdd_uq11 gnd read_bl_0_31 read_bl_1_31 write_bl_0_31 wwl_0_24 rwl_1_24
+ rwl_0_24 cell_2r1w
Xcell_2r1w_1342 vdd_uq0 gnd read_bl_0_43 read_bl_1_43 write_bl_0_43 wwl_0_1 rwl_1_1
+ rwl_0_1 cell_2r1w
Xcell_2r1w_1397 vdd_uq4 gnd read_bl_0_42 read_bl_1_42 write_bl_0_42 wwl_0_10 rwl_1_10
+ rwl_0_10 cell_2r1w
Xcell_2r1w_1331 vdd_uq5 gnd read_bl_0_43 read_bl_1_43 write_bl_0_43 wwl_0_12 rwl_1_12
+ rwl_0_12 cell_2r1w
Xcell_2r1w_2098 vdd_uq5 gnd read_bl_0_31 read_bl_1_31 write_bl_0_31 wwl_0_13 rwl_1_13
+ rwl_0_13 cell_2r1w
Xcell_2r1w_1386 vdd_uq9 gnd read_bl_0_42 read_bl_1_42 write_bl_0_42 wwl_0_21 rwl_1_21
+ rwl_0_21 cell_2r1w
Xcell_2r1w_1161 vdd_uq26 gnd read_bl_0_45 read_bl_1_45 write_bl_0_45 wwl_0_54 rwl_1_54
+ rwl_0_54 cell_2r1w
Xcell_2r1w_1150 vdd_uq0 gnd read_bl_0_46 read_bl_1_46 write_bl_0_46 wwl_0_1 rwl_1_1
+ rwl_0_1 cell_2r1w
Xcell_2r1w_1172 vdd_uq20 gnd read_bl_0_45 read_bl_1_45 write_bl_0_45 wwl_0_43 rwl_1_43
+ rwl_0_43 cell_2r1w
Xcell_2r1w_1183 vdd_uq15 gnd read_bl_0_45 read_bl_1_45 write_bl_0_45 wwl_0_32 rwl_1_32
+ rwl_0_32 cell_2r1w
Xcell_2r1w_1194 vdd_uq9 gnd read_bl_0_45 read_bl_1_45 write_bl_0_45 wwl_0_21 rwl_1_21
+ rwl_0_21 cell_2r1w
Xcell_2r1w_1919 vdd_uq0 gnd read_bl_0_34 read_bl_1_34 write_bl_0_34 wwl_0_0 rwl_1_0
+ rwl_0_0 cell_2r1w
Xcell_2r1w_1908 vdd_uq4 gnd read_bl_0_34 read_bl_1_34 write_bl_0_34 wwl_0_11 rwl_1_11
+ rwl_0_11 cell_2r1w
Xcell_2r1w_2609 vdd_uq6 gnd read_bl_0_23 read_bl_1_23 write_bl_0_23 wwl_0_14 rwl_1_14
+ rwl_0_14 cell_2r1w
Xcell_2r1w_3844 vdd_uq28 gnd read_bl_0_3 read_bl_1_3 write_bl_0_3 wwl_0_59 rwl_1_59
+ rwl_0_59 cell_2r1w
Xcell_2r1w_3855 vdd_uq23 gnd read_bl_0_3 read_bl_1_3 write_bl_0_3 wwl_0_48 rwl_1_48
+ rwl_0_48 cell_2r1w
Xcell_2r1w_3800 vdd_uq18 gnd read_bl_0_4 read_bl_1_4 write_bl_0_4 wwl_0_39 rwl_1_39
+ rwl_0_39 cell_2r1w
Xcell_2r1w_3811 vdd_uq13 gnd read_bl_0_4 read_bl_1_4 write_bl_0_4 wwl_0_28 rwl_1_28
+ rwl_0_28 cell_2r1w
Xcell_2r1w_3833 vdd_uq2 gnd read_bl_0_4 read_bl_1_4 write_bl_0_4 wwl_0_6 rwl_1_6 rwl_0_6
+ cell_2r1w
Xcell_2r1w_3822 vdd_uq7 gnd read_bl_0_4 read_bl_1_4 write_bl_0_4 wwl_0_17 rwl_1_17
+ rwl_0_17 cell_2r1w
Xcell_2r1w_3866 vdd_uq17 gnd read_bl_0_3 read_bl_1_3 write_bl_0_3 wwl_0_37 rwl_1_37
+ rwl_0_37 cell_2r1w
Xcell_2r1w_3877 vdd_uq12 gnd read_bl_0_3 read_bl_1_3 write_bl_0_3 wwl_0_26 rwl_1_26
+ rwl_0_26 cell_2r1w
Xcell_2r1w_3899 vdd_uq1 gnd read_bl_0_3 read_bl_1_3 write_bl_0_3 wwl_0_4 rwl_1_4 rwl_0_4
+ cell_2r1w
Xcell_2r1w_3888 vdd_uq6 gnd read_bl_0_3 read_bl_1_3 write_bl_0_3 wwl_0_15 rwl_1_15
+ rwl_0_15 cell_2r1w
Xcell_2r1w_409 vdd_uq18 gnd read_bl_0_57 read_bl_1_57 write_bl_0_57 wwl_0_38 rwl_1_38
+ rwl_0_38 cell_2r1w
Xcell_2r1w_3107 vdd_uq13 gnd read_bl_0_15 read_bl_1_15 write_bl_0_15 wwl_0_28 rwl_1_28
+ rwl_0_28 cell_2r1w
Xcell_2r1w_3129 vdd_uq2 gnd read_bl_0_15 read_bl_1_15 write_bl_0_15 wwl_0_6 rwl_1_6
+ rwl_0_6 cell_2r1w
Xcell_2r1w_3118 vdd_uq7 gnd read_bl_0_15 read_bl_1_15 write_bl_0_15 wwl_0_17 rwl_1_17
+ rwl_0_17 cell_2r1w
Xcell_2r1w_965 vdd_uq28 gnd read_bl_0_48 read_bl_1_48 write_bl_0_48 wwl_0_58 rwl_1_58
+ rwl_0_58 cell_2r1w
Xcell_2r1w_2439 vdd_uq27 gnd read_bl_0_25 read_bl_1_25 write_bl_0_25 wwl_0_56 rwl_1_56
+ rwl_0_56 cell_2r1w
Xcell_2r1w_1738 vdd_uq25 gnd read_bl_0_36 read_bl_1_36 write_bl_0_36 wwl_0_53 rwl_1_53
+ rwl_0_53 cell_2r1w
Xcell_2r1w_910 vdd_uq23 gnd read_bl_0_49 read_bl_1_49 write_bl_0_49 wwl_0_49 rwl_1_49
+ rwl_0_49 cell_2r1w
Xcell_2r1w_1749 vdd_uq20 gnd read_bl_0_36 read_bl_1_36 write_bl_0_36 wwl_0_42 rwl_1_42
+ rwl_0_42 cell_2r1w
Xcell_2r1w_921 vdd_uq18 gnd read_bl_0_49 read_bl_1_49 write_bl_0_49 wwl_0_38 rwl_1_38
+ rwl_0_38 cell_2r1w
Xcell_2r1w_932 vdd_uq12 gnd read_bl_0_49 read_bl_1_49 write_bl_0_49 wwl_0_27 rwl_1_27
+ rwl_0_27 cell_2r1w
Xcell_2r1w_2406 vdd_uq11 gnd read_bl_0_26 read_bl_1_26 write_bl_0_26 wwl_0_25 rwl_1_25
+ rwl_0_25 cell_2r1w
Xcell_2r1w_954 vdd_uq1 gnd read_bl_0_49 read_bl_1_49 write_bl_0_49 wwl_0_5 rwl_1_5
+ rwl_0_5 cell_2r1w
Xcell_2r1w_2428 vdd gnd read_bl_0_26 read_bl_1_26 write_bl_0_26 wwl_0_3 rwl_1_3 rwl_0_3
+ cell_2r1w
Xcell_2r1w_1727 vdd_uq0 gnd read_bl_0_37 read_bl_1_37 write_bl_0_37 wwl_0_0 rwl_1_0
+ rwl_0_0 cell_2r1w
Xcell_2r1w_1716 vdd_uq4 gnd read_bl_0_37 read_bl_1_37 write_bl_0_37 wwl_0_11 rwl_1_11
+ rwl_0_11 cell_2r1w
Xcell_2r1w_2417 vdd_uq6 gnd read_bl_0_26 read_bl_1_26 write_bl_0_26 wwl_0_14 rwl_1_14
+ rwl_0_14 cell_2r1w
Xcell_2r1w_943 vdd_uq7 gnd read_bl_0_49 read_bl_1_49 write_bl_0_49 wwl_0_16 rwl_1_16
+ rwl_0_16 cell_2r1w
Xcell_2r1w_1705 vdd_uq10 gnd read_bl_0_37 read_bl_1_37 write_bl_0_37 wwl_0_22 rwl_1_22
+ rwl_0_22 cell_2r1w
Xcell_2r1w_976 vdd_uq22 gnd read_bl_0_48 read_bl_1_48 write_bl_0_48 wwl_0_47 rwl_1_47
+ rwl_0_47 cell_2r1w
Xcell_2r1w_987 vdd_uq17 gnd read_bl_0_48 read_bl_1_48 write_bl_0_48 wwl_0_36 rwl_1_36
+ rwl_0_36 cell_2r1w
Xcell_2r1w_998 vdd_uq11 gnd read_bl_0_48 read_bl_1_48 write_bl_0_48 wwl_0_25 rwl_1_25
+ rwl_0_25 cell_2r1w
Xcell_2r1w_3652 vdd_uq28 gnd read_bl_0_6 read_bl_1_6 write_bl_0_6 wwl_0_59 rwl_1_59
+ rwl_0_59 cell_2r1w
Xcell_2r1w_2951 vdd_uq27 gnd read_bl_0_17 read_bl_1_17 write_bl_0_17 wwl_0_56 rwl_1_56
+ rwl_0_56 cell_2r1w
Xcell_2r1w_3663 vdd_uq23 gnd read_bl_0_6 read_bl_1_6 write_bl_0_6 wwl_0_48 rwl_1_48
+ rwl_0_48 cell_2r1w
Xcell_2r1w_3674 vdd_uq17 gnd read_bl_0_6 read_bl_1_6 write_bl_0_6 wwl_0_37 rwl_1_37
+ rwl_0_37 cell_2r1w
Xcell_2r1w_3685 vdd_uq12 gnd read_bl_0_6 read_bl_1_6 write_bl_0_6 wwl_0_26 rwl_1_26
+ rwl_0_26 cell_2r1w
Xcell_2r1w_2940 vdd gnd read_bl_0_18 read_bl_1_18 write_bl_0_18 wwl_0_3 rwl_1_3 rwl_0_3
+ cell_2r1w
Xcell_2r1w_3641 vdd_uq2 gnd read_bl_0_7 read_bl_1_7 write_bl_0_7 wwl_0_6 rwl_1_6 rwl_0_6
+ cell_2r1w
Xcell_2r1w_3696 vdd_uq6 gnd read_bl_0_6 read_bl_1_6 write_bl_0_6 wwl_0_15 rwl_1_15
+ rwl_0_15 cell_2r1w
Xcell_2r1w_3630 vdd_uq7 gnd read_bl_0_7 read_bl_1_7 write_bl_0_7 wwl_0_17 rwl_1_17
+ rwl_0_17 cell_2r1w
Xcell_2r1w_2962 vdd_uq21 gnd read_bl_0_17 read_bl_1_17 write_bl_0_17 wwl_0_45 rwl_1_45
+ rwl_0_45 cell_2r1w
Xcell_2r1w_2973 vdd_uq16 gnd read_bl_0_17 read_bl_1_17 write_bl_0_17 wwl_0_34 rwl_1_34
+ rwl_0_34 cell_2r1w
Xcell_2r1w_2995 vdd_uq5 gnd read_bl_0_17 read_bl_1_17 write_bl_0_17 wwl_0_12 rwl_1_12
+ rwl_0_12 cell_2r1w
Xcell_2r1w_2984 vdd_uq10 gnd read_bl_0_17 read_bl_1_17 write_bl_0_17 wwl_0_23 rwl_1_23
+ rwl_0_23 cell_2r1w
Xcell_2r1w_66 vdd_uq29 gnd read_bl_0_62 read_bl_1_62 write_bl_0_62 wwl_0_61 rwl_1_61
+ rwl_0_61 cell_2r1w
Xcell_2r1w_11 vdd_uq25 gnd read_bl_0_63 read_bl_1_63 write_bl_0_63 wwl_0_52 rwl_1_52
+ rwl_0_52 cell_2r1w
Xcell_2r1w_77 vdd_uq24 gnd read_bl_0_62 read_bl_1_62 write_bl_0_62 wwl_0_50 rwl_1_50
+ rwl_0_50 cell_2r1w
Xcell_2r1w_22 vdd_uq19 gnd read_bl_0_63 read_bl_1_63 write_bl_0_63 wwl_0_41 rwl_1_41
+ rwl_0_41 cell_2r1w
Xcell_2r1w_88 vdd_uq18 gnd read_bl_0_62 read_bl_1_62 write_bl_0_62 wwl_0_39 rwl_1_39
+ rwl_0_39 cell_2r1w
Xcell_2r1w_33 vdd_uq14 gnd read_bl_0_63 read_bl_1_63 write_bl_0_63 wwl_0_30 rwl_1_30
+ rwl_0_30 cell_2r1w
Xcell_2r1w_99 vdd_uq13 gnd read_bl_0_62 read_bl_1_62 write_bl_0_62 wwl_0_28 rwl_1_28
+ rwl_0_28 cell_2r1w
Xcell_2r1w_55 vdd_uq3 gnd read_bl_0_63 read_bl_1_63 write_bl_0_63 wwl_0_8 rwl_1_8
+ rwl_0_8 cell_2r1w
Xcell_2r1w_44 vdd_uq8 gnd read_bl_0_63 read_bl_1_63 write_bl_0_63 wwl_0_19 rwl_1_19
+ rwl_0_19 cell_2r1w
Xcell_2r1w_206 vdd_uq23 gnd read_bl_0_60 read_bl_1_60 write_bl_0_60 wwl_0_49 rwl_1_49
+ rwl_0_49 cell_2r1w
Xcell_2r1w_217 vdd_uq18 gnd read_bl_0_60 read_bl_1_60 write_bl_0_60 wwl_0_38 rwl_1_38
+ rwl_0_38 cell_2r1w
Xcell_2r1w_228 vdd_uq12 gnd read_bl_0_60 read_bl_1_60 write_bl_0_60 wwl_0_27 rwl_1_27
+ rwl_0_27 cell_2r1w
Xcell_2r1w_239 vdd_uq7 gnd read_bl_0_60 read_bl_1_60 write_bl_0_60 wwl_0_16 rwl_1_16
+ rwl_0_16 cell_2r1w
Xcell_2r1w_2247 vdd_uq27 gnd read_bl_0_28 read_bl_1_28 write_bl_0_28 wwl_0_56 rwl_1_56
+ rwl_0_56 cell_2r1w
Xcell_2r1w_2203 vdd_uq17 gnd read_bl_0_29 read_bl_1_29 write_bl_0_29 wwl_0_36 rwl_1_36
+ rwl_0_36 cell_2r1w
Xcell_2r1w_1502 vdd_uq15 gnd read_bl_0_40 read_bl_1_40 write_bl_0_40 wwl_0_33 rwl_1_33
+ rwl_0_33 cell_2r1w
Xcell_2r1w_2214 vdd_uq11 gnd read_bl_0_29 read_bl_1_29 write_bl_0_29 wwl_0_25 rwl_1_25
+ rwl_0_25 cell_2r1w
Xcell_2r1w_2236 vdd gnd read_bl_0_29 read_bl_1_29 write_bl_0_29 wwl_0_3 rwl_1_3 rwl_0_3
+ cell_2r1w
Xcell_2r1w_2225 vdd_uq6 gnd read_bl_0_29 read_bl_1_29 write_bl_0_29 wwl_0_14 rwl_1_14
+ rwl_0_14 cell_2r1w
Xcell_2r1w_773 vdd_uq28 gnd read_bl_0_51 read_bl_1_51 write_bl_0_51 wwl_0_58 rwl_1_58
+ rwl_0_58 cell_2r1w
Xcell_2r1w_1546 vdd_uq25 gnd read_bl_0_39 read_bl_1_39 write_bl_0_39 wwl_0_53 rwl_1_53
+ rwl_0_53 cell_2r1w
Xcell_2r1w_784 vdd_uq22 gnd read_bl_0_51 read_bl_1_51 write_bl_0_51 wwl_0_47 rwl_1_47
+ rwl_0_47 cell_2r1w
Xcell_2r1w_2258 vdd_uq21 gnd read_bl_0_28 read_bl_1_28 write_bl_0_28 wwl_0_45 rwl_1_45
+ rwl_0_45 cell_2r1w
Xcell_2r1w_1557 vdd_uq20 gnd read_bl_0_39 read_bl_1_39 write_bl_0_39 wwl_0_42 rwl_1_42
+ rwl_0_42 cell_2r1w
Xcell_2r1w_795 vdd_uq17 gnd read_bl_0_51 read_bl_1_51 write_bl_0_51 wwl_0_36 rwl_1_36
+ rwl_0_36 cell_2r1w
Xcell_2r1w_2269 vdd_uq16 gnd read_bl_0_28 read_bl_1_28 write_bl_0_28 wwl_0_34 rwl_1_34
+ rwl_0_34 cell_2r1w
Xcell_2r1w_1568 vdd_uq14 gnd read_bl_0_39 read_bl_1_39 write_bl_0_39 wwl_0_31 rwl_1_31
+ rwl_0_31 cell_2r1w
Xcell_2r1w_740 vdd_uq12 gnd read_bl_0_52 read_bl_1_52 write_bl_0_52 wwl_0_27 rwl_1_27
+ rwl_0_27 cell_2r1w
Xcell_2r1w_762 vdd_uq1 gnd read_bl_0_52 read_bl_1_52 write_bl_0_52 wwl_0_5 rwl_1_5
+ rwl_0_5 cell_2r1w
Xcell_2r1w_1535 vdd_uq0 gnd read_bl_0_40 read_bl_1_40 write_bl_0_40 wwl_0_0 rwl_1_0
+ rwl_0_0 cell_2r1w
Xcell_2r1w_1524 vdd_uq4 gnd read_bl_0_40 read_bl_1_40 write_bl_0_40 wwl_0_11 rwl_1_11
+ rwl_0_11 cell_2r1w
Xcell_2r1w_751 vdd_uq7 gnd read_bl_0_52 read_bl_1_52 write_bl_0_52 wwl_0_16 rwl_1_16
+ rwl_0_16 cell_2r1w
Xcell_2r1w_1579 vdd_uq9 gnd read_bl_0_39 read_bl_1_39 write_bl_0_39 wwl_0_20 rwl_1_20
+ rwl_0_20 cell_2r1w
Xcell_2r1w_1513 vdd_uq10 gnd read_bl_0_40 read_bl_1_40 write_bl_0_40 wwl_0_22 rwl_1_22
+ rwl_0_22 cell_2r1w
Xcell_2r1w_1 vdd_uq30 gnd read_bl_0_63 read_bl_1_63 write_bl_0_63 wwl_0_62 rwl_1_62
+ rwl_0_62 cell_2r1w
Xcell_2r1w_3460 vdd_uq28 gnd read_bl_0_9 read_bl_1_9 write_bl_0_9 wwl_0_59 rwl_1_59
+ rwl_0_59 cell_2r1w
Xcell_2r1w_3471 vdd_uq23 gnd read_bl_0_9 read_bl_1_9 write_bl_0_9 wwl_0_48 rwl_1_48
+ rwl_0_48 cell_2r1w
Xcell_2r1w_2770 vdd_uq21 gnd read_bl_0_20 read_bl_1_20 write_bl_0_20 wwl_0_45 rwl_1_45
+ rwl_0_45 cell_2r1w
Xcell_2r1w_3482 vdd_uq17 gnd read_bl_0_9 read_bl_1_9 write_bl_0_9 wwl_0_37 rwl_1_37
+ rwl_0_37 cell_2r1w
Xcell_2r1w_2781 vdd_uq16 gnd read_bl_0_20 read_bl_1_20 write_bl_0_20 wwl_0_34 rwl_1_34
+ rwl_0_34 cell_2r1w
Xcell_2r1w_3493 vdd_uq12 gnd read_bl_0_9 read_bl_1_9 write_bl_0_9 wwl_0_26 rwl_1_26
+ rwl_0_26 cell_2r1w
Xcell_2r1w_2792 vdd_uq10 gnd read_bl_0_20 read_bl_1_20 write_bl_0_20 wwl_0_23 rwl_1_23
+ rwl_0_23 cell_2r1w
Xcell_2r1w_2055 vdd_uq27 gnd read_bl_0_31 read_bl_1_31 write_bl_0_31 wwl_0_56 rwl_1_56
+ rwl_0_56 cell_2r1w
Xcell_2r1w_1354 vdd_uq25 gnd read_bl_0_42 read_bl_1_42 write_bl_0_42 wwl_0_53 rwl_1_53
+ rwl_0_53 cell_2r1w
Xcell_2r1w_2000 vdd_uq22 gnd read_bl_0_32 read_bl_1_32 write_bl_0_32 wwl_0_47 rwl_1_47
+ rwl_0_47 cell_2r1w
Xcell_2r1w_2066 vdd_uq21 gnd read_bl_0_31 read_bl_1_31 write_bl_0_31 wwl_0_45 rwl_1_45
+ rwl_0_45 cell_2r1w
Xcell_2r1w_2011 vdd_uq17 gnd read_bl_0_32 read_bl_1_32 write_bl_0_32 wwl_0_36 rwl_1_36
+ rwl_0_36 cell_2r1w
Xcell_2r1w_2077 vdd_uq16 gnd read_bl_0_31 read_bl_1_31 write_bl_0_31 wwl_0_34 rwl_1_34
+ rwl_0_34 cell_2r1w
Xcell_2r1w_1310 vdd_uq15 gnd read_bl_0_43 read_bl_1_43 write_bl_0_43 wwl_0_33 rwl_1_33
+ rwl_0_33 cell_2r1w
Xcell_2r1w_2022 vdd_uq11 gnd read_bl_0_32 read_bl_1_32 write_bl_0_32 wwl_0_25 rwl_1_25
+ rwl_0_25 cell_2r1w
Xcell_2r1w_2044 vdd gnd read_bl_0_32 read_bl_1_32 write_bl_0_32 wwl_0_3 rwl_1_3 rwl_0_3
+ cell_2r1w
Xcell_2r1w_1343 vdd_uq0 gnd read_bl_0_43 read_bl_1_43 write_bl_0_43 wwl_0_0 rwl_1_0
+ rwl_0_0 cell_2r1w
Xcell_2r1w_1332 vdd_uq4 gnd read_bl_0_43 read_bl_1_43 write_bl_0_43 wwl_0_11 rwl_1_11
+ rwl_0_11 cell_2r1w
Xcell_2r1w_2033 vdd_uq6 gnd read_bl_0_32 read_bl_1_32 write_bl_0_32 wwl_0_14 rwl_1_14
+ rwl_0_14 cell_2r1w
Xcell_2r1w_1321 vdd_uq10 gnd read_bl_0_43 read_bl_1_43 write_bl_0_43 wwl_0_22 rwl_1_22
+ rwl_0_22 cell_2r1w
Xcell_2r1w_2088 vdd_uq10 gnd read_bl_0_31 read_bl_1_31 write_bl_0_31 wwl_0_23 rwl_1_23
+ rwl_0_23 cell_2r1w
Xcell_2r1w_581 vdd_uq28 gnd read_bl_0_54 read_bl_1_54 write_bl_0_54 wwl_0_58 rwl_1_58
+ rwl_0_58 cell_2r1w
Xcell_2r1w_592 vdd_uq22 gnd read_bl_0_54 read_bl_1_54 write_bl_0_54 wwl_0_47 rwl_1_47
+ rwl_0_47 cell_2r1w
Xcell_2r1w_1365 vdd_uq20 gnd read_bl_0_42 read_bl_1_42 write_bl_0_42 wwl_0_42 rwl_1_42
+ rwl_0_42 cell_2r1w
Xcell_2r1w_1376 vdd_uq14 gnd read_bl_0_42 read_bl_1_42 write_bl_0_42 wwl_0_31 rwl_1_31
+ rwl_0_31 cell_2r1w
Xcell_2r1w_570 vdd_uq1 gnd read_bl_0_55 read_bl_1_55 write_bl_0_55 wwl_0_5 rwl_1_5
+ rwl_0_5 cell_2r1w
Xcell_2r1w_1398 vdd_uq3 gnd read_bl_0_42 read_bl_1_42 write_bl_0_42 wwl_0_9 rwl_1_9
+ rwl_0_9 cell_2r1w
Xcell_2r1w_2099 vdd_uq5 gnd read_bl_0_31 read_bl_1_31 write_bl_0_31 wwl_0_12 rwl_1_12
+ rwl_0_12 cell_2r1w
Xcell_2r1w_1387 vdd_uq9 gnd read_bl_0_42 read_bl_1_42 write_bl_0_42 wwl_0_20 rwl_1_20
+ rwl_0_20 cell_2r1w
Xcell_2r1w_3290 vdd_uq17 gnd read_bl_0_12 read_bl_1_12 write_bl_0_12 wwl_0_37 rwl_1_37
+ rwl_0_37 cell_2r1w
Xcell_2r1w_1162 vdd_uq25 gnd read_bl_0_45 read_bl_1_45 write_bl_0_45 wwl_0_53 rwl_1_53
+ rwl_0_53 cell_2r1w
Xcell_2r1w_1173 vdd_uq20 gnd read_bl_0_45 read_bl_1_45 write_bl_0_45 wwl_0_42 rwl_1_42
+ rwl_0_42 cell_2r1w
Xcell_2r1w_1184 vdd_uq14 gnd read_bl_0_45 read_bl_1_45 write_bl_0_45 wwl_0_31 rwl_1_31
+ rwl_0_31 cell_2r1w
Xcell_2r1w_1151 vdd_uq0 gnd read_bl_0_46 read_bl_1_46 write_bl_0_46 wwl_0_0 rwl_1_0
+ rwl_0_0 cell_2r1w
Xcell_2r1w_1140 vdd_uq4 gnd read_bl_0_46 read_bl_1_46 write_bl_0_46 wwl_0_11 rwl_1_11
+ rwl_0_11 cell_2r1w
Xcell_2r1w_1195 vdd_uq9 gnd read_bl_0_45 read_bl_1_45 write_bl_0_45 wwl_0_20 rwl_1_20
+ rwl_0_20 cell_2r1w
Xcell_2r1w_1909 vdd_uq4 gnd read_bl_0_34 read_bl_1_34 write_bl_0_34 wwl_0_10 rwl_1_10
+ rwl_0_10 cell_2r1w
Xcell_2r1w_3845 vdd_uq28 gnd read_bl_0_3 read_bl_1_3 write_bl_0_3 wwl_0_58 rwl_1_58
+ rwl_0_58 cell_2r1w
Xcell_2r1w_3856 vdd_uq22 gnd read_bl_0_3 read_bl_1_3 write_bl_0_3 wwl_0_47 rwl_1_47
+ rwl_0_47 cell_2r1w
Xcell_2r1w_3801 vdd_uq18 gnd read_bl_0_4 read_bl_1_4 write_bl_0_4 wwl_0_38 rwl_1_38
+ rwl_0_38 cell_2r1w
Xcell_2r1w_3867 vdd_uq17 gnd read_bl_0_3 read_bl_1_3 write_bl_0_3 wwl_0_36 rwl_1_36
+ rwl_0_36 cell_2r1w
Xcell_2r1w_3812 vdd_uq12 gnd read_bl_0_4 read_bl_1_4 write_bl_0_4 wwl_0_27 rwl_1_27
+ rwl_0_27 cell_2r1w
Xcell_2r1w_3878 vdd_uq11 gnd read_bl_0_3 read_bl_1_3 write_bl_0_3 wwl_0_25 rwl_1_25
+ rwl_0_25 cell_2r1w
Xcell_2r1w_3834 vdd_uq1 gnd read_bl_0_4 read_bl_1_4 write_bl_0_4 wwl_0_5 rwl_1_5 rwl_0_5
+ cell_2r1w
Xcell_2r1w_3823 vdd_uq7 gnd read_bl_0_4 read_bl_1_4 write_bl_0_4 wwl_0_16 rwl_1_16
+ rwl_0_16 cell_2r1w
Xcell_2r1w_3889 vdd_uq6 gnd read_bl_0_3 read_bl_1_3 write_bl_0_3 wwl_0_14 rwl_1_14
+ rwl_0_14 cell_2r1w
Xcell_2r1w_3108 vdd_uq12 gnd read_bl_0_15 read_bl_1_15 write_bl_0_15 wwl_0_27 rwl_1_27
+ rwl_0_27 cell_2r1w
Xcell_2r1w_2407 vdd_uq11 gnd read_bl_0_26 read_bl_1_26 write_bl_0_26 wwl_0_24 rwl_1_24
+ rwl_0_24 cell_2r1w
Xcell_2r1w_2429 vdd gnd read_bl_0_26 read_bl_1_26 write_bl_0_26 wwl_0_2 rwl_1_2 rwl_0_2
+ cell_2r1w
Xcell_2r1w_2418 vdd_uq5 gnd read_bl_0_26 read_bl_1_26 write_bl_0_26 wwl_0_13 rwl_1_13
+ rwl_0_13 cell_2r1w
Xcell_2r1w_3119 vdd_uq7 gnd read_bl_0_15 read_bl_1_15 write_bl_0_15 wwl_0_16 rwl_1_16
+ rwl_0_16 cell_2r1w
Xcell_2r1w_1728 vdd_uq30 gnd read_bl_0_36 read_bl_1_36 write_bl_0_36 wwl_0_63 rwl_1_63
+ rwl_0_63 cell_2r1w
Xcell_2r1w_900 vdd_uq28 gnd read_bl_0_49 read_bl_1_49 write_bl_0_49 wwl_0_59 rwl_1_59
+ rwl_0_59 cell_2r1w
Xcell_2r1w_966 vdd_uq27 gnd read_bl_0_48 read_bl_1_48 write_bl_0_48 wwl_0_57 rwl_1_57
+ rwl_0_57 cell_2r1w
Xcell_2r1w_1739 vdd_uq25 gnd read_bl_0_36 read_bl_1_36 write_bl_0_36 wwl_0_52 rwl_1_52
+ rwl_0_52 cell_2r1w
Xcell_2r1w_911 vdd_uq23 gnd read_bl_0_49 read_bl_1_49 write_bl_0_49 wwl_0_48 rwl_1_48
+ rwl_0_48 cell_2r1w
Xcell_2r1w_977 vdd_uq22 gnd read_bl_0_48 read_bl_1_48 write_bl_0_48 wwl_0_46 rwl_1_46
+ rwl_0_46 cell_2r1w
Xcell_2r1w_922 vdd_uq17 gnd read_bl_0_49 read_bl_1_49 write_bl_0_49 wwl_0_37 rwl_1_37
+ rwl_0_37 cell_2r1w
Xcell_2r1w_988 vdd_uq16 gnd read_bl_0_48 read_bl_1_48 write_bl_0_48 wwl_0_35 rwl_1_35
+ rwl_0_35 cell_2r1w
Xcell_2r1w_933 vdd_uq12 gnd read_bl_0_49 read_bl_1_49 write_bl_0_49 wwl_0_26 rwl_1_26
+ rwl_0_26 cell_2r1w
Xcell_2r1w_955 vdd_uq1 gnd read_bl_0_49 read_bl_1_49 write_bl_0_49 wwl_0_4 rwl_1_4
+ rwl_0_4 cell_2r1w
Xcell_2r1w_1717 vdd_uq4 gnd read_bl_0_37 read_bl_1_37 write_bl_0_37 wwl_0_10 rwl_1_10
+ rwl_0_10 cell_2r1w
Xcell_2r1w_944 vdd_uq6 gnd read_bl_0_49 read_bl_1_49 write_bl_0_49 wwl_0_15 rwl_1_15
+ rwl_0_15 cell_2r1w
Xcell_2r1w_1706 vdd_uq9 gnd read_bl_0_37 read_bl_1_37 write_bl_0_37 wwl_0_21 rwl_1_21
+ rwl_0_21 cell_2r1w
Xcell_2r1w_999 vdd_uq11 gnd read_bl_0_48 read_bl_1_48 write_bl_0_48 wwl_0_24 rwl_1_24
+ rwl_0_24 cell_2r1w
Xcell_2r1w_3653 vdd_uq28 gnd read_bl_0_6 read_bl_1_6 write_bl_0_6 wwl_0_58 rwl_1_58
+ rwl_0_58 cell_2r1w
Xcell_2r1w_2952 vdd_uq26 gnd read_bl_0_17 read_bl_1_17 write_bl_0_17 wwl_0_55 rwl_1_55
+ rwl_0_55 cell_2r1w
Xcell_2r1w_3664 vdd_uq22 gnd read_bl_0_6 read_bl_1_6 write_bl_0_6 wwl_0_47 rwl_1_47
+ rwl_0_47 cell_2r1w
Xcell_2r1w_2963 vdd_uq21 gnd read_bl_0_17 read_bl_1_17 write_bl_0_17 wwl_0_44 rwl_1_44
+ rwl_0_44 cell_2r1w
Xcell_2r1w_3675 vdd_uq17 gnd read_bl_0_6 read_bl_1_6 write_bl_0_6 wwl_0_36 rwl_1_36
+ rwl_0_36 cell_2r1w
Xcell_2r1w_2974 vdd_uq15 gnd read_bl_0_17 read_bl_1_17 write_bl_0_17 wwl_0_33 rwl_1_33
+ rwl_0_33 cell_2r1w
Xcell_2r1w_3620 vdd_uq12 gnd read_bl_0_7 read_bl_1_7 write_bl_0_7 wwl_0_27 rwl_1_27
+ rwl_0_27 cell_2r1w
Xcell_2r1w_3686 vdd_uq11 gnd read_bl_0_6 read_bl_1_6 write_bl_0_6 wwl_0_25 rwl_1_25
+ rwl_0_25 cell_2r1w
Xcell_2r1w_3642 vdd_uq1 gnd read_bl_0_7 read_bl_1_7 write_bl_0_7 wwl_0_5 rwl_1_5 rwl_0_5
+ cell_2r1w
Xcell_2r1w_2941 vdd gnd read_bl_0_18 read_bl_1_18 write_bl_0_18 wwl_0_2 rwl_1_2 rwl_0_2
+ cell_2r1w
Xcell_2r1w_3697 vdd_uq6 gnd read_bl_0_6 read_bl_1_6 write_bl_0_6 wwl_0_14 rwl_1_14
+ rwl_0_14 cell_2r1w
Xcell_2r1w_2930 vdd_uq5 gnd read_bl_0_18 read_bl_1_18 write_bl_0_18 wwl_0_13 rwl_1_13
+ rwl_0_13 cell_2r1w
Xcell_2r1w_3631 vdd_uq7 gnd read_bl_0_7 read_bl_1_7 write_bl_0_7 wwl_0_16 rwl_1_16
+ rwl_0_16 cell_2r1w
Xcell_2r1w_2985 vdd_uq10 gnd read_bl_0_17 read_bl_1_17 write_bl_0_17 wwl_0_22 rwl_1_22
+ rwl_0_22 cell_2r1w
Xcell_2r1w_12 vdd_uq24 gnd read_bl_0_63 read_bl_1_63 write_bl_0_63 wwl_0_51 rwl_1_51
+ rwl_0_51 cell_2r1w
Xcell_2r1w_2996 vdd_uq4 gnd read_bl_0_17 read_bl_1_17 write_bl_0_17 wwl_0_11 rwl_1_11
+ rwl_0_11 cell_2r1w
Xcell_2r1w_67 vdd_uq29 gnd read_bl_0_62 read_bl_1_62 write_bl_0_62 wwl_0_60 rwl_1_60
+ rwl_0_60 cell_2r1w
Xcell_2r1w_78 vdd_uq23 gnd read_bl_0_62 read_bl_1_62 write_bl_0_62 wwl_0_49 rwl_1_49
+ rwl_0_49 cell_2r1w
Xcell_2r1w_23 vdd_uq19 gnd read_bl_0_63 read_bl_1_63 write_bl_0_63 wwl_0_40 rwl_1_40
+ rwl_0_40 cell_2r1w
Xcell_2r1w_89 vdd_uq18 gnd read_bl_0_62 read_bl_1_62 write_bl_0_62 wwl_0_38 rwl_1_38
+ rwl_0_38 cell_2r1w
Xcell_2r1w_34 vdd_uq13 gnd read_bl_0_63 read_bl_1_63 write_bl_0_63 wwl_0_29 rwl_1_29
+ rwl_0_29 cell_2r1w
Xcell_2r1w_56 vdd_uq2 gnd read_bl_0_63 read_bl_1_63 write_bl_0_63 wwl_0_7 rwl_1_7
+ rwl_0_7 cell_2r1w
Xcell_2r1w_45 vdd_uq8 gnd read_bl_0_63 read_bl_1_63 write_bl_0_63 wwl_0_18 rwl_1_18
+ rwl_0_18 cell_2r1w
Xcell_2r1w_207 vdd_uq23 gnd read_bl_0_60 read_bl_1_60 write_bl_0_60 wwl_0_48 rwl_1_48
+ rwl_0_48 cell_2r1w
Xcell_2r1w_218 vdd_uq17 gnd read_bl_0_60 read_bl_1_60 write_bl_0_60 wwl_0_37 rwl_1_37
+ rwl_0_37 cell_2r1w
Xcell_2r1w_229 vdd_uq12 gnd read_bl_0_60 read_bl_1_60 write_bl_0_60 wwl_0_26 rwl_1_26
+ rwl_0_26 cell_2r1w
Xcell_2r1w_1536 vdd_uq30 gnd read_bl_0_39 read_bl_1_39 write_bl_0_39 wwl_0_63 rwl_1_63
+ rwl_0_63 cell_2r1w
Xcell_2r1w_2248 vdd_uq26 gnd read_bl_0_28 read_bl_1_28 write_bl_0_28 wwl_0_55 rwl_1_55
+ rwl_0_55 cell_2r1w
Xcell_2r1w_2259 vdd_uq21 gnd read_bl_0_28 read_bl_1_28 write_bl_0_28 wwl_0_44 rwl_1_44
+ rwl_0_44 cell_2r1w
Xcell_2r1w_2204 vdd_uq16 gnd read_bl_0_29 read_bl_1_29 write_bl_0_29 wwl_0_35 rwl_1_35
+ rwl_0_35 cell_2r1w
Xcell_2r1w_1503 vdd_uq15 gnd read_bl_0_40 read_bl_1_40 write_bl_0_40 wwl_0_32 rwl_1_32
+ rwl_0_32 cell_2r1w
Xcell_2r1w_2215 vdd_uq11 gnd read_bl_0_29 read_bl_1_29 write_bl_0_29 wwl_0_24 rwl_1_24
+ rwl_0_24 cell_2r1w
Xcell_2r1w_2237 vdd gnd read_bl_0_29 read_bl_1_29 write_bl_0_29 wwl_0_2 rwl_1_2 rwl_0_2
+ cell_2r1w
Xcell_2r1w_1525 vdd_uq4 gnd read_bl_0_40 read_bl_1_40 write_bl_0_40 wwl_0_10 rwl_1_10
+ rwl_0_10 cell_2r1w
Xcell_2r1w_2226 vdd_uq5 gnd read_bl_0_29 read_bl_1_29 write_bl_0_29 wwl_0_13 rwl_1_13
+ rwl_0_13 cell_2r1w
Xcell_2r1w_1514 vdd_uq9 gnd read_bl_0_40 read_bl_1_40 write_bl_0_40 wwl_0_21 rwl_1_21
+ rwl_0_21 cell_2r1w
Xcell_2r1w_774 vdd_uq27 gnd read_bl_0_51 read_bl_1_51 write_bl_0_51 wwl_0_57 rwl_1_57
+ rwl_0_57 cell_2r1w
Xcell_2r1w_1547 vdd_uq25 gnd read_bl_0_39 read_bl_1_39 write_bl_0_39 wwl_0_52 rwl_1_52
+ rwl_0_52 cell_2r1w
Xcell_2r1w_785 vdd_uq22 gnd read_bl_0_51 read_bl_1_51 write_bl_0_51 wwl_0_46 rwl_1_46
+ rwl_0_46 cell_2r1w
Xcell_2r1w_1558 vdd_uq19 gnd read_bl_0_39 read_bl_1_39 write_bl_0_39 wwl_0_41 rwl_1_41
+ rwl_0_41 cell_2r1w
Xcell_2r1w_730 vdd_uq17 gnd read_bl_0_52 read_bl_1_52 write_bl_0_52 wwl_0_37 rwl_1_37
+ rwl_0_37 cell_2r1w
Xcell_2r1w_796 vdd_uq16 gnd read_bl_0_51 read_bl_1_51 write_bl_0_51 wwl_0_35 rwl_1_35
+ rwl_0_35 cell_2r1w
Xcell_2r1w_1569 vdd_uq14 gnd read_bl_0_39 read_bl_1_39 write_bl_0_39 wwl_0_30 rwl_1_30
+ rwl_0_30 cell_2r1w
Xcell_2r1w_741 vdd_uq12 gnd read_bl_0_52 read_bl_1_52 write_bl_0_52 wwl_0_26 rwl_1_26
+ rwl_0_26 cell_2r1w
Xcell_2r1w_763 vdd_uq1 gnd read_bl_0_52 read_bl_1_52 write_bl_0_52 wwl_0_4 rwl_1_4
+ rwl_0_4 cell_2r1w
Xcell_2r1w_752 vdd_uq6 gnd read_bl_0_52 read_bl_1_52 write_bl_0_52 wwl_0_15 rwl_1_15
+ rwl_0_15 cell_2r1w
Xcell_2r1w_2 vdd_uq29 gnd read_bl_0_63 read_bl_1_63 write_bl_0_63 wwl_0_61 rwl_1_61
+ rwl_0_61 cell_2r1w
Xcell_2r1w_3461 vdd_uq28 gnd read_bl_0_9 read_bl_1_9 write_bl_0_9 wwl_0_58 rwl_1_58
+ rwl_0_58 cell_2r1w
Xcell_2r1w_2760 vdd_uq26 gnd read_bl_0_20 read_bl_1_20 write_bl_0_20 wwl_0_55 rwl_1_55
+ rwl_0_55 cell_2r1w
Xcell_2r1w_3472 vdd_uq22 gnd read_bl_0_9 read_bl_1_9 write_bl_0_9 wwl_0_47 rwl_1_47
+ rwl_0_47 cell_2r1w
Xcell_2r1w_2771 vdd_uq21 gnd read_bl_0_20 read_bl_1_20 write_bl_0_20 wwl_0_44 rwl_1_44
+ rwl_0_44 cell_2r1w
Xcell_2r1w_3483 vdd_uq17 gnd read_bl_0_9 read_bl_1_9 write_bl_0_9 wwl_0_36 rwl_1_36
+ rwl_0_36 cell_2r1w
Xcell_2r1w_2782 vdd_uq15 gnd read_bl_0_20 read_bl_1_20 write_bl_0_20 wwl_0_33 rwl_1_33
+ rwl_0_33 cell_2r1w
Xcell_2r1w_3494 vdd_uq11 gnd read_bl_0_9 read_bl_1_9 write_bl_0_9 wwl_0_25 rwl_1_25
+ rwl_0_25 cell_2r1w
Xcell_2r1w_3450 vdd_uq1 gnd read_bl_0_10 read_bl_1_10 write_bl_0_10 wwl_0_5 rwl_1_5
+ rwl_0_5 cell_2r1w
Xcell_2r1w_2793 vdd_uq10 gnd read_bl_0_20 read_bl_1_20 write_bl_0_20 wwl_0_22 rwl_1_22
+ rwl_0_22 cell_2r1w
Xcell_2r1w_1344 vdd_uq30 gnd read_bl_0_42 read_bl_1_42 write_bl_0_42 wwl_0_63 rwl_1_63
+ rwl_0_63 cell_2r1w
Xcell_2r1w_2056 vdd_uq26 gnd read_bl_0_31 read_bl_1_31 write_bl_0_31 wwl_0_55 rwl_1_55
+ rwl_0_55 cell_2r1w
Xcell_2r1w_1355 vdd_uq25 gnd read_bl_0_42 read_bl_1_42 write_bl_0_42 wwl_0_52 rwl_1_52
+ rwl_0_52 cell_2r1w
Xcell_2r1w_2001 vdd_uq22 gnd read_bl_0_32 read_bl_1_32 write_bl_0_32 wwl_0_46 rwl_1_46
+ rwl_0_46 cell_2r1w
Xcell_2r1w_2067 vdd_uq21 gnd read_bl_0_31 read_bl_1_31 write_bl_0_31 wwl_0_44 rwl_1_44
+ rwl_0_44 cell_2r1w
Xcell_2r1w_1300 vdd_uq20 gnd read_bl_0_43 read_bl_1_43 write_bl_0_43 wwl_0_43 rwl_1_43
+ rwl_0_43 cell_2r1w
Xcell_2r1w_1366 vdd_uq19 gnd read_bl_0_42 read_bl_1_42 write_bl_0_42 wwl_0_41 rwl_1_41
+ rwl_0_41 cell_2r1w
Xcell_2r1w_2012 vdd_uq16 gnd read_bl_0_32 read_bl_1_32 write_bl_0_32 wwl_0_35 rwl_1_35
+ rwl_0_35 cell_2r1w
Xcell_2r1w_2078 vdd_uq15 gnd read_bl_0_31 read_bl_1_31 write_bl_0_31 wwl_0_33 rwl_1_33
+ rwl_0_33 cell_2r1w
Xcell_2r1w_1311 vdd_uq15 gnd read_bl_0_43 read_bl_1_43 write_bl_0_43 wwl_0_32 rwl_1_32
+ rwl_0_32 cell_2r1w
Xcell_2r1w_1377 vdd_uq14 gnd read_bl_0_42 read_bl_1_42 write_bl_0_42 wwl_0_30 rwl_1_30
+ rwl_0_30 cell_2r1w
Xcell_2r1w_2023 vdd_uq11 gnd read_bl_0_32 read_bl_1_32 write_bl_0_32 wwl_0_24 rwl_1_24
+ rwl_0_24 cell_2r1w
Xcell_2r1w_2045 vdd gnd read_bl_0_32 read_bl_1_32 write_bl_0_32 wwl_0_2 rwl_1_2 rwl_0_2
+ cell_2r1w
Xcell_2r1w_1333 vdd_uq4 gnd read_bl_0_43 read_bl_1_43 write_bl_0_43 wwl_0_10 rwl_1_10
+ rwl_0_10 cell_2r1w
Xcell_2r1w_2034 vdd_uq5 gnd read_bl_0_32 read_bl_1_32 write_bl_0_32 wwl_0_13 rwl_1_13
+ rwl_0_13 cell_2r1w
Xcell_2r1w_1322 vdd_uq9 gnd read_bl_0_43 read_bl_1_43 write_bl_0_43 wwl_0_21 rwl_1_21
+ rwl_0_21 cell_2r1w
Xcell_2r1w_2089 vdd_uq10 gnd read_bl_0_31 read_bl_1_31 write_bl_0_31 wwl_0_22 rwl_1_22
+ rwl_0_22 cell_2r1w
Xcell_2r1w_582 vdd_uq27 gnd read_bl_0_54 read_bl_1_54 write_bl_0_54 wwl_0_57 rwl_1_57
+ rwl_0_57 cell_2r1w
Xcell_2r1w_593 vdd_uq22 gnd read_bl_0_54 read_bl_1_54 write_bl_0_54 wwl_0_46 rwl_1_46
+ rwl_0_46 cell_2r1w
Xcell_2r1w_571 vdd_uq1 gnd read_bl_0_55 read_bl_1_55 write_bl_0_55 wwl_0_4 rwl_1_4
+ rwl_0_4 cell_2r1w
Xcell_2r1w_1399 vdd_uq3 gnd read_bl_0_42 read_bl_1_42 write_bl_0_42 wwl_0_8 rwl_1_8
+ rwl_0_8 cell_2r1w
Xcell_2r1w_560 vdd_uq6 gnd read_bl_0_55 read_bl_1_55 write_bl_0_55 wwl_0_15 rwl_1_15
+ rwl_0_15 cell_2r1w
Xcell_2r1w_1388 vdd_uq8 gnd read_bl_0_42 read_bl_1_42 write_bl_0_42 wwl_0_19 rwl_1_19
+ rwl_0_19 cell_2r1w
Xcell_2r1w_3280 vdd_uq22 gnd read_bl_0_12 read_bl_1_12 write_bl_0_12 wwl_0_47 rwl_1_47
+ rwl_0_47 cell_2r1w
Xcell_2r1w_3291 vdd_uq17 gnd read_bl_0_12 read_bl_1_12 write_bl_0_12 wwl_0_36 rwl_1_36
+ rwl_0_36 cell_2r1w
Xcell_2r1w_2590 vdd_uq15 gnd read_bl_0_23 read_bl_1_23 write_bl_0_23 wwl_0_33 rwl_1_33
+ rwl_0_33 cell_2r1w
Xcell_2r1w_1152 vdd_uq30 gnd read_bl_0_45 read_bl_1_45 write_bl_0_45 wwl_0_63 rwl_1_63
+ rwl_0_63 cell_2r1w
Xcell_2r1w_390 vdd_uq27 gnd read_bl_0_57 read_bl_1_57 write_bl_0_57 wwl_0_57 rwl_1_57
+ rwl_0_57 cell_2r1w
Xcell_2r1w_1163 vdd_uq25 gnd read_bl_0_45 read_bl_1_45 write_bl_0_45 wwl_0_52 rwl_1_52
+ rwl_0_52 cell_2r1w
Xcell_2r1w_1174 vdd_uq19 gnd read_bl_0_45 read_bl_1_45 write_bl_0_45 wwl_0_41 rwl_1_41
+ rwl_0_41 cell_2r1w
Xcell_2r1w_1185 vdd_uq14 gnd read_bl_0_45 read_bl_1_45 write_bl_0_45 wwl_0_30 rwl_1_30
+ rwl_0_30 cell_2r1w
Xcell_2r1w_1141 vdd_uq4 gnd read_bl_0_46 read_bl_1_46 write_bl_0_46 wwl_0_10 rwl_1_10
+ rwl_0_10 cell_2r1w
Xcell_2r1w_1196 vdd_uq8 gnd read_bl_0_45 read_bl_1_45 write_bl_0_45 wwl_0_19 rwl_1_19
+ rwl_0_19 cell_2r1w
Xcell_2r1w_1130 vdd_uq9 gnd read_bl_0_46 read_bl_1_46 write_bl_0_46 wwl_0_21 rwl_1_21
+ rwl_0_21 cell_2r1w
Xcell_2r1w_3846 vdd_uq27 gnd read_bl_0_3 read_bl_1_3 write_bl_0_3 wwl_0_57 rwl_1_57
+ rwl_0_57 cell_2r1w
Xcell_2r1w_3857 vdd_uq22 gnd read_bl_0_3 read_bl_1_3 write_bl_0_3 wwl_0_46 rwl_1_46
+ rwl_0_46 cell_2r1w
Xcell_2r1w_3802 vdd_uq17 gnd read_bl_0_4 read_bl_1_4 write_bl_0_4 wwl_0_37 rwl_1_37
+ rwl_0_37 cell_2r1w
Xcell_2r1w_3868 vdd_uq16 gnd read_bl_0_3 read_bl_1_3 write_bl_0_3 wwl_0_35 rwl_1_35
+ rwl_0_35 cell_2r1w
Xcell_2r1w_3813 vdd_uq12 gnd read_bl_0_4 read_bl_1_4 write_bl_0_4 wwl_0_26 rwl_1_26
+ rwl_0_26 cell_2r1w
Xcell_2r1w_3879 vdd_uq11 gnd read_bl_0_3 read_bl_1_3 write_bl_0_3 wwl_0_24 rwl_1_24
+ rwl_0_24 cell_2r1w
Xcell_2r1w_3835 vdd_uq1 gnd read_bl_0_4 read_bl_1_4 write_bl_0_4 wwl_0_4 rwl_1_4 rwl_0_4
+ cell_2r1w
Xcell_2r1w_3824 vdd_uq6 gnd read_bl_0_4 read_bl_1_4 write_bl_0_4 wwl_0_15 rwl_1_15
+ rwl_0_15 cell_2r1w
Xcell_2r1w_3109 vdd_uq12 gnd read_bl_0_15 read_bl_1_15 write_bl_0_15 wwl_0_26 rwl_1_26
+ rwl_0_26 cell_2r1w
Xcell_2r1w_1718 vdd_uq3 gnd read_bl_0_37 read_bl_1_37 write_bl_0_37 wwl_0_9 rwl_1_9
+ rwl_0_9 cell_2r1w
Xcell_2r1w_2419 vdd_uq5 gnd read_bl_0_26 read_bl_1_26 write_bl_0_26 wwl_0_12 rwl_1_12
+ rwl_0_12 cell_2r1w
Xcell_2r1w_1707 vdd_uq9 gnd read_bl_0_37 read_bl_1_37 write_bl_0_37 wwl_0_20 rwl_1_20
+ rwl_0_20 cell_2r1w
Xcell_2r1w_2408 vdd_uq10 gnd read_bl_0_26 read_bl_1_26 write_bl_0_26 wwl_0_23 rwl_1_23
+ rwl_0_23 cell_2r1w
Xcell_2r1w_1729 vdd_uq30 gnd read_bl_0_36 read_bl_1_36 write_bl_0_36 wwl_0_62 rwl_1_62
+ rwl_0_62 cell_2r1w
Xcell_2r1w_901 vdd_uq28 gnd read_bl_0_49 read_bl_1_49 write_bl_0_49 wwl_0_58 rwl_1_58
+ rwl_0_58 cell_2r1w
Xcell_2r1w_967 vdd_uq27 gnd read_bl_0_48 read_bl_1_48 write_bl_0_48 wwl_0_56 rwl_1_56
+ rwl_0_56 cell_2r1w
Xcell_2r1w_912 vdd_uq22 gnd read_bl_0_49 read_bl_1_49 write_bl_0_49 wwl_0_47 rwl_1_47
+ rwl_0_47 cell_2r1w
Xcell_2r1w_978 vdd_uq21 gnd read_bl_0_48 read_bl_1_48 write_bl_0_48 wwl_0_45 rwl_1_45
+ rwl_0_45 cell_2r1w
Xcell_2r1w_923 vdd_uq17 gnd read_bl_0_49 read_bl_1_49 write_bl_0_49 wwl_0_36 rwl_1_36
+ rwl_0_36 cell_2r1w
Xcell_2r1w_989 vdd_uq16 gnd read_bl_0_48 read_bl_1_48 write_bl_0_48 wwl_0_34 rwl_1_34
+ rwl_0_34 cell_2r1w
Xcell_2r1w_934 vdd_uq11 gnd read_bl_0_49 read_bl_1_49 write_bl_0_49 wwl_0_25 rwl_1_25
+ rwl_0_25 cell_2r1w
Xcell_2r1w_956 vdd gnd read_bl_0_49 read_bl_1_49 write_bl_0_49 wwl_0_3 rwl_1_3 rwl_0_3
+ cell_2r1w
Xcell_2r1w_945 vdd_uq6 gnd read_bl_0_49 read_bl_1_49 write_bl_0_49 wwl_0_14 rwl_1_14
+ rwl_0_14 cell_2r1w
Xcell_2r1w_3610 vdd_uq17 gnd read_bl_0_7 read_bl_1_7 write_bl_0_7 wwl_0_37 rwl_1_37
+ rwl_0_37 cell_2r1w
Xcell_2r1w_3654 vdd_uq27 gnd read_bl_0_6 read_bl_1_6 write_bl_0_6 wwl_0_57 rwl_1_57
+ rwl_0_57 cell_2r1w
Xcell_2r1w_2953 vdd_uq26 gnd read_bl_0_17 read_bl_1_17 write_bl_0_17 wwl_0_54 rwl_1_54
+ rwl_0_54 cell_2r1w
Xcell_2r1w_3665 vdd_uq22 gnd read_bl_0_6 read_bl_1_6 write_bl_0_6 wwl_0_46 rwl_1_46
+ rwl_0_46 cell_2r1w
Xcell_2r1w_2964 vdd_uq20 gnd read_bl_0_17 read_bl_1_17 write_bl_0_17 wwl_0_43 rwl_1_43
+ rwl_0_43 cell_2r1w
Xcell_2r1w_3676 vdd_uq16 gnd read_bl_0_6 read_bl_1_6 write_bl_0_6 wwl_0_35 rwl_1_35
+ rwl_0_35 cell_2r1w
Xcell_2r1w_2975 vdd_uq15 gnd read_bl_0_17 read_bl_1_17 write_bl_0_17 wwl_0_32 rwl_1_32
+ rwl_0_32 cell_2r1w
Xcell_2r1w_3621 vdd_uq12 gnd read_bl_0_7 read_bl_1_7 write_bl_0_7 wwl_0_26 rwl_1_26
+ rwl_0_26 cell_2r1w
Xcell_2r1w_3687 vdd_uq11 gnd read_bl_0_6 read_bl_1_6 write_bl_0_6 wwl_0_24 rwl_1_24
+ rwl_0_24 cell_2r1w
Xcell_2r1w_3643 vdd_uq1 gnd read_bl_0_7 read_bl_1_7 write_bl_0_7 wwl_0_4 rwl_1_4 rwl_0_4
+ cell_2r1w
Xcell_2r1w_2942 vdd_uq0 gnd read_bl_0_18 read_bl_1_18 write_bl_0_18 wwl_0_1 rwl_1_1
+ rwl_0_1 cell_2r1w
Xcell_2r1w_2997 vdd_uq4 gnd read_bl_0_17 read_bl_1_17 write_bl_0_17 wwl_0_10 rwl_1_10
+ rwl_0_10 cell_2r1w
Xcell_2r1w_2931 vdd_uq5 gnd read_bl_0_18 read_bl_1_18 write_bl_0_18 wwl_0_12 rwl_1_12
+ rwl_0_12 cell_2r1w
Xcell_2r1w_3698 vdd_uq5 gnd read_bl_0_6 read_bl_1_6 write_bl_0_6 wwl_0_13 rwl_1_13
+ rwl_0_13 cell_2r1w
Xcell_2r1w_3632 vdd_uq6 gnd read_bl_0_7 read_bl_1_7 write_bl_0_7 wwl_0_15 rwl_1_15
+ rwl_0_15 cell_2r1w
Xcell_2r1w_2986 vdd_uq9 gnd read_bl_0_17 read_bl_1_17 write_bl_0_17 wwl_0_21 rwl_1_21
+ rwl_0_21 cell_2r1w
Xcell_2r1w_2920 vdd_uq10 gnd read_bl_0_18 read_bl_1_18 write_bl_0_18 wwl_0_23 rwl_1_23
+ rwl_0_23 cell_2r1w
Xcell_2r1w_13 vdd_uq24 gnd read_bl_0_63 read_bl_1_63 write_bl_0_63 wwl_0_50 rwl_1_50
+ rwl_0_50 cell_2r1w
Xcell_2r1w_24 vdd_uq18 gnd read_bl_0_63 read_bl_1_63 write_bl_0_63 wwl_0_39 rwl_1_39
+ rwl_0_39 cell_2r1w
Xcell_2r1w_35 vdd_uq13 gnd read_bl_0_63 read_bl_1_63 write_bl_0_63 wwl_0_28 rwl_1_28
+ rwl_0_28 cell_2r1w
Xcell_2r1w_46 vdd_uq7 gnd read_bl_0_63 read_bl_1_63 write_bl_0_63 wwl_0_17 rwl_1_17
+ rwl_0_17 cell_2r1w
Xcell_2r1w_68 vdd_uq28 gnd read_bl_0_62 read_bl_1_62 write_bl_0_62 wwl_0_59 rwl_1_59
+ rwl_0_59 cell_2r1w
Xcell_2r1w_79 vdd_uq23 gnd read_bl_0_62 read_bl_1_62 write_bl_0_62 wwl_0_48 rwl_1_48
+ rwl_0_48 cell_2r1w
Xcell_2r1w_57 vdd_uq2 gnd read_bl_0_63 read_bl_1_63 write_bl_0_63 wwl_0_6 rwl_1_6
+ rwl_0_6 cell_2r1w
Xcell_2r1w_208 vdd_uq22 gnd read_bl_0_60 read_bl_1_60 write_bl_0_60 wwl_0_47 rwl_1_47
+ rwl_0_47 cell_2r1w
Xcell_2r1w_219 vdd_uq17 gnd read_bl_0_60 read_bl_1_60 write_bl_0_60 wwl_0_36 rwl_1_36
+ rwl_0_36 cell_2r1w
Xcell_2r1w_1537 vdd_uq30 gnd read_bl_0_39 read_bl_1_39 write_bl_0_39 wwl_0_62 rwl_1_62
+ rwl_0_62 cell_2r1w
Xcell_2r1w_2249 vdd_uq26 gnd read_bl_0_28 read_bl_1_28 write_bl_0_28 wwl_0_54 rwl_1_54
+ rwl_0_54 cell_2r1w
Xcell_2r1w_1548 vdd_uq24 gnd read_bl_0_39 read_bl_1_39 write_bl_0_39 wwl_0_51 rwl_1_51
+ rwl_0_51 cell_2r1w
Xcell_2r1w_720 vdd_uq22 gnd read_bl_0_52 read_bl_1_52 write_bl_0_52 wwl_0_47 rwl_1_47
+ rwl_0_47 cell_2r1w
Xcell_2r1w_1559 vdd_uq19 gnd read_bl_0_39 read_bl_1_39 write_bl_0_39 wwl_0_40 rwl_1_40
+ rwl_0_40 cell_2r1w
Xcell_2r1w_731 vdd_uq17 gnd read_bl_0_52 read_bl_1_52 write_bl_0_52 wwl_0_36 rwl_1_36
+ rwl_0_36 cell_2r1w
Xcell_2r1w_2205 vdd_uq16 gnd read_bl_0_29 read_bl_1_29 write_bl_0_29 wwl_0_34 rwl_1_34
+ rwl_0_34 cell_2r1w
Xcell_2r1w_1504 vdd_uq14 gnd read_bl_0_40 read_bl_1_40 write_bl_0_40 wwl_0_31 rwl_1_31
+ rwl_0_31 cell_2r1w
Xcell_2r1w_2238 vdd_uq0 gnd read_bl_0_29 read_bl_1_29 write_bl_0_29 wwl_0_1 rwl_1_1
+ rwl_0_1 cell_2r1w
Xcell_2r1w_1526 vdd_uq3 gnd read_bl_0_40 read_bl_1_40 write_bl_0_40 wwl_0_9 rwl_1_9
+ rwl_0_9 cell_2r1w
Xcell_2r1w_2227 vdd_uq5 gnd read_bl_0_29 read_bl_1_29 write_bl_0_29 wwl_0_12 rwl_1_12
+ rwl_0_12 cell_2r1w
Xcell_2r1w_1515 vdd_uq9 gnd read_bl_0_40 read_bl_1_40 write_bl_0_40 wwl_0_20 rwl_1_20
+ rwl_0_20 cell_2r1w
Xcell_2r1w_2216 vdd_uq10 gnd read_bl_0_29 read_bl_1_29 write_bl_0_29 wwl_0_23 rwl_1_23
+ rwl_0_23 cell_2r1w
Xcell_2r1w_775 vdd_uq27 gnd read_bl_0_51 read_bl_1_51 write_bl_0_51 wwl_0_56 rwl_1_56
+ rwl_0_56 cell_2r1w
Xcell_2r1w_786 vdd_uq21 gnd read_bl_0_51 read_bl_1_51 write_bl_0_51 wwl_0_45 rwl_1_45
+ rwl_0_45 cell_2r1w
Xcell_2r1w_797 vdd_uq16 gnd read_bl_0_51 read_bl_1_51 write_bl_0_51 wwl_0_34 rwl_1_34
+ rwl_0_34 cell_2r1w
Xcell_2r1w_742 vdd_uq11 gnd read_bl_0_52 read_bl_1_52 write_bl_0_52 wwl_0_25 rwl_1_25
+ rwl_0_25 cell_2r1w
Xcell_2r1w_764 vdd gnd read_bl_0_52 read_bl_1_52 write_bl_0_52 wwl_0_3 rwl_1_3 rwl_0_3
+ cell_2r1w
Xcell_2r1w_753 vdd_uq6 gnd read_bl_0_52 read_bl_1_52 write_bl_0_52 wwl_0_14 rwl_1_14
+ rwl_0_14 cell_2r1w
Xcell_2r1w_3 vdd_uq29 gnd read_bl_0_63 read_bl_1_63 write_bl_0_63 wwl_0_60 rwl_1_60
+ rwl_0_60 cell_2r1w
Xcell_2r1w_3462 vdd_uq27 gnd read_bl_0_9 read_bl_1_9 write_bl_0_9 wwl_0_57 rwl_1_57
+ rwl_0_57 cell_2r1w
Xcell_2r1w_3451 vdd_uq1 gnd read_bl_0_10 read_bl_1_10 write_bl_0_10 wwl_0_4 rwl_1_4
+ rwl_0_4 cell_2r1w
Xcell_2r1w_3440 vdd_uq6 gnd read_bl_0_10 read_bl_1_10 write_bl_0_10 wwl_0_15 rwl_1_15
+ rwl_0_15 cell_2r1w
Xcell_2r1w_2761 vdd_uq26 gnd read_bl_0_20 read_bl_1_20 write_bl_0_20 wwl_0_54 rwl_1_54
+ rwl_0_54 cell_2r1w
Xcell_2r1w_3473 vdd_uq22 gnd read_bl_0_9 read_bl_1_9 write_bl_0_9 wwl_0_46 rwl_1_46
+ rwl_0_46 cell_2r1w
Xcell_2r1w_2772 vdd_uq20 gnd read_bl_0_20 read_bl_1_20 write_bl_0_20 wwl_0_43 rwl_1_43
+ rwl_0_43 cell_2r1w
Xcell_2r1w_3484 vdd_uq16 gnd read_bl_0_9 read_bl_1_9 write_bl_0_9 wwl_0_35 rwl_1_35
+ rwl_0_35 cell_2r1w
Xcell_2r1w_2783 vdd_uq15 gnd read_bl_0_20 read_bl_1_20 write_bl_0_20 wwl_0_32 rwl_1_32
+ rwl_0_32 cell_2r1w
Xcell_2r1w_3495 vdd_uq11 gnd read_bl_0_9 read_bl_1_9 write_bl_0_9 wwl_0_24 rwl_1_24
+ rwl_0_24 cell_2r1w
Xcell_2r1w_2750 vdd_uq0 gnd read_bl_0_21 read_bl_1_21 write_bl_0_21 wwl_0_1 rwl_1_1
+ rwl_0_1 cell_2r1w
Xcell_2r1w_2794 vdd_uq9 gnd read_bl_0_20 read_bl_1_20 write_bl_0_20 wwl_0_21 rwl_1_21
+ rwl_0_21 cell_2r1w
Xcell_2r1w_2002 vdd_uq21 gnd read_bl_0_32 read_bl_1_32 write_bl_0_32 wwl_0_45 rwl_1_45
+ rwl_0_45 cell_2r1w
Xcell_2r1w_2013 vdd_uq16 gnd read_bl_0_32 read_bl_1_32 write_bl_0_32 wwl_0_34 rwl_1_34
+ rwl_0_34 cell_2r1w
Xcell_2r1w_1345 vdd_uq30 gnd read_bl_0_42 read_bl_1_42 write_bl_0_42 wwl_0_62 rwl_1_62
+ rwl_0_62 cell_2r1w
Xcell_2r1w_2057 vdd_uq26 gnd read_bl_0_31 read_bl_1_31 write_bl_0_31 wwl_0_54 rwl_1_54
+ rwl_0_54 cell_2r1w
Xcell_2r1w_1356 vdd_uq24 gnd read_bl_0_42 read_bl_1_42 write_bl_0_42 wwl_0_51 rwl_1_51
+ rwl_0_51 cell_2r1w
Xcell_2r1w_2068 vdd_uq20 gnd read_bl_0_31 read_bl_1_31 write_bl_0_31 wwl_0_43 rwl_1_43
+ rwl_0_43 cell_2r1w
Xcell_2r1w_1301 vdd_uq20 gnd read_bl_0_43 read_bl_1_43 write_bl_0_43 wwl_0_42 rwl_1_42
+ rwl_0_42 cell_2r1w
Xcell_2r1w_1367 vdd_uq19 gnd read_bl_0_42 read_bl_1_42 write_bl_0_42 wwl_0_40 rwl_1_40
+ rwl_0_40 cell_2r1w
Xcell_2r1w_2079 vdd_uq15 gnd read_bl_0_31 read_bl_1_31 write_bl_0_31 wwl_0_32 rwl_1_32
+ rwl_0_32 cell_2r1w
Xcell_2r1w_1312 vdd_uq14 gnd read_bl_0_43 read_bl_1_43 write_bl_0_43 wwl_0_31 rwl_1_31
+ rwl_0_31 cell_2r1w
Xcell_2r1w_1378 vdd_uq13 gnd read_bl_0_42 read_bl_1_42 write_bl_0_42 wwl_0_29 rwl_1_29
+ rwl_0_29 cell_2r1w
Xcell_2r1w_550 vdd_uq11 gnd read_bl_0_55 read_bl_1_55 write_bl_0_55 wwl_0_25 rwl_1_25
+ rwl_0_25 cell_2r1w
Xcell_2r1w_572 vdd gnd read_bl_0_55 read_bl_1_55 write_bl_0_55 wwl_0_3 rwl_1_3 rwl_0_3
+ cell_2r1w
Xcell_2r1w_2046 vdd_uq0 gnd read_bl_0_32 read_bl_1_32 write_bl_0_32 wwl_0_1 rwl_1_1
+ rwl_0_1 cell_2r1w
Xcell_2r1w_1334 vdd_uq3 gnd read_bl_0_43 read_bl_1_43 write_bl_0_43 wwl_0_9 rwl_1_9
+ rwl_0_9 cell_2r1w
Xcell_2r1w_2035 vdd_uq5 gnd read_bl_0_32 read_bl_1_32 write_bl_0_32 wwl_0_12 rwl_1_12
+ rwl_0_12 cell_2r1w
Xcell_2r1w_561 vdd_uq6 gnd read_bl_0_55 read_bl_1_55 write_bl_0_55 wwl_0_14 rwl_1_14
+ rwl_0_14 cell_2r1w
Xcell_2r1w_1389 vdd_uq8 gnd read_bl_0_42 read_bl_1_42 write_bl_0_42 wwl_0_18 rwl_1_18
+ rwl_0_18 cell_2r1w
Xcell_2r1w_1323 vdd_uq9 gnd read_bl_0_43 read_bl_1_43 write_bl_0_43 wwl_0_20 rwl_1_20
+ rwl_0_20 cell_2r1w
Xcell_2r1w_2024 vdd_uq10 gnd read_bl_0_32 read_bl_1_32 write_bl_0_32 wwl_0_23 rwl_1_23
+ rwl_0_23 cell_2r1w
Xcell_2r1w_583 vdd_uq27 gnd read_bl_0_54 read_bl_1_54 write_bl_0_54 wwl_0_56 rwl_1_56
+ rwl_0_56 cell_2r1w
Xcell_2r1w_594 vdd_uq21 gnd read_bl_0_54 read_bl_1_54 write_bl_0_54 wwl_0_45 rwl_1_45
+ rwl_0_45 cell_2r1w
Xcell_2r1w_3270 vdd_uq27 gnd read_bl_0_12 read_bl_1_12 write_bl_0_12 wwl_0_57 rwl_1_57
+ rwl_0_57 cell_2r1w
Xcell_2r1w_3281 vdd_uq22 gnd read_bl_0_12 read_bl_1_12 write_bl_0_12 wwl_0_46 rwl_1_46
+ rwl_0_46 cell_2r1w
Xcell_2r1w_3292 vdd_uq16 gnd read_bl_0_12 read_bl_1_12 write_bl_0_12 wwl_0_35 rwl_1_35
+ rwl_0_35 cell_2r1w
Xcell_2r1w_2580 vdd_uq20 gnd read_bl_0_23 read_bl_1_23 write_bl_0_23 wwl_0_43 rwl_1_43
+ rwl_0_43 cell_2r1w
Xcell_2r1w_2591 vdd_uq15 gnd read_bl_0_23 read_bl_1_23 write_bl_0_23 wwl_0_32 rwl_1_32
+ rwl_0_32 cell_2r1w
Xcell_2r1w_1890 vdd_uq13 gnd read_bl_0_34 read_bl_1_34 write_bl_0_34 wwl_0_29 rwl_1_29
+ rwl_0_29 cell_2r1w
Xcell_2r1w_1153 vdd_uq30 gnd read_bl_0_45 read_bl_1_45 write_bl_0_45 wwl_0_62 rwl_1_62
+ rwl_0_62 cell_2r1w
Xcell_2r1w_391 vdd_uq27 gnd read_bl_0_57 read_bl_1_57 write_bl_0_57 wwl_0_56 rwl_1_56
+ rwl_0_56 cell_2r1w
Xcell_2r1w_1164 vdd_uq24 gnd read_bl_0_45 read_bl_1_45 write_bl_0_45 wwl_0_51 rwl_1_51
+ rwl_0_51 cell_2r1w
Xcell_2r1w_1175 vdd_uq19 gnd read_bl_0_45 read_bl_1_45 write_bl_0_45 wwl_0_40 rwl_1_40
+ rwl_0_40 cell_2r1w
Xcell_2r1w_1120 vdd_uq14 gnd read_bl_0_46 read_bl_1_46 write_bl_0_46 wwl_0_31 rwl_1_31
+ rwl_0_31 cell_2r1w
Xcell_2r1w_1186 vdd_uq13 gnd read_bl_0_45 read_bl_1_45 write_bl_0_45 wwl_0_29 rwl_1_29
+ rwl_0_29 cell_2r1w
Xcell_2r1w_380 vdd gnd read_bl_0_58 read_bl_1_58 write_bl_0_58 wwl_0_3 rwl_1_3 rwl_0_3
+ cell_2r1w
Xcell_2r1w_1142 vdd_uq3 gnd read_bl_0_46 read_bl_1_46 write_bl_0_46 wwl_0_9 rwl_1_9
+ rwl_0_9 cell_2r1w
Xcell_2r1w_1197 vdd_uq8 gnd read_bl_0_45 read_bl_1_45 write_bl_0_45 wwl_0_18 rwl_1_18
+ rwl_0_18 cell_2r1w
Xcell_2r1w_1131 vdd_uq9 gnd read_bl_0_46 read_bl_1_46 write_bl_0_46 wwl_0_20 rwl_1_20
+ rwl_0_20 cell_2r1w
Xcell_2r1w_3803 vdd_uq17 gnd read_bl_0_4 read_bl_1_4 write_bl_0_4 wwl_0_36 rwl_1_36
+ rwl_0_36 cell_2r1w
Xcell_2r1w_3847 vdd_uq27 gnd read_bl_0_3 read_bl_1_3 write_bl_0_3 wwl_0_56 rwl_1_56
+ rwl_0_56 cell_2r1w
Xcell_2r1w_3858 vdd_uq21 gnd read_bl_0_3 read_bl_1_3 write_bl_0_3 wwl_0_45 rwl_1_45
+ rwl_0_45 cell_2r1w
Xcell_2r1w_3869 vdd_uq16 gnd read_bl_0_3 read_bl_1_3 write_bl_0_3 wwl_0_34 rwl_1_34
+ rwl_0_34 cell_2r1w
Xcell_2r1w_3814 vdd_uq11 gnd read_bl_0_4 read_bl_1_4 write_bl_0_4 wwl_0_25 rwl_1_25
+ rwl_0_25 cell_2r1w
Xcell_2r1w_3836 vdd gnd read_bl_0_4 read_bl_1_4 write_bl_0_4 wwl_0_3 rwl_1_3 rwl_0_3
+ cell_2r1w
Xcell_2r1w_3825 vdd_uq6 gnd read_bl_0_4 read_bl_1_4 write_bl_0_4 wwl_0_14 rwl_1_14
+ rwl_0_14 cell_2r1w
Xcell_2r1w_902 vdd_uq27 gnd read_bl_0_49 read_bl_1_49 write_bl_0_49 wwl_0_57 rwl_1_57
+ rwl_0_57 cell_2r1w
Xcell_2r1w_913 vdd_uq22 gnd read_bl_0_49 read_bl_1_49 write_bl_0_49 wwl_0_46 rwl_1_46
+ rwl_0_46 cell_2r1w
Xcell_2r1w_1719 vdd_uq3 gnd read_bl_0_37 read_bl_1_37 write_bl_0_37 wwl_0_8 rwl_1_8
+ rwl_0_8 cell_2r1w
Xcell_2r1w_1708 vdd_uq8 gnd read_bl_0_37 read_bl_1_37 write_bl_0_37 wwl_0_19 rwl_1_19
+ rwl_0_19 cell_2r1w
Xcell_2r1w_2409 vdd_uq10 gnd read_bl_0_26 read_bl_1_26 write_bl_0_26 wwl_0_22 rwl_1_22
+ rwl_0_22 cell_2r1w
Xcell_2r1w_968 vdd_uq26 gnd read_bl_0_48 read_bl_1_48 write_bl_0_48 wwl_0_55 rwl_1_55
+ rwl_0_55 cell_2r1w
Xcell_2r1w_979 vdd_uq21 gnd read_bl_0_48 read_bl_1_48 write_bl_0_48 wwl_0_44 rwl_1_44
+ rwl_0_44 cell_2r1w
Xcell_2r1w_924 vdd_uq16 gnd read_bl_0_49 read_bl_1_49 write_bl_0_49 wwl_0_35 rwl_1_35
+ rwl_0_35 cell_2r1w
Xcell_2r1w_935 vdd_uq11 gnd read_bl_0_49 read_bl_1_49 write_bl_0_49 wwl_0_24 rwl_1_24
+ rwl_0_24 cell_2r1w
Xcell_2r1w_957 vdd gnd read_bl_0_49 read_bl_1_49 write_bl_0_49 wwl_0_2 rwl_1_2 rwl_0_2
+ cell_2r1w
Xcell_2r1w_946 vdd_uq5 gnd read_bl_0_49 read_bl_1_49 write_bl_0_49 wwl_0_13 rwl_1_13
+ rwl_0_13 cell_2r1w
Xcell_2r1w_3600 vdd_uq22 gnd read_bl_0_7 read_bl_1_7 write_bl_0_7 wwl_0_47 rwl_1_47
+ rwl_0_47 cell_2r1w
Xcell_2r1w_3611 vdd_uq17 gnd read_bl_0_7 read_bl_1_7 write_bl_0_7 wwl_0_36 rwl_1_36
+ rwl_0_36 cell_2r1w
Xcell_2r1w_3622 vdd_uq11 gnd read_bl_0_7 read_bl_1_7 write_bl_0_7 wwl_0_25 rwl_1_25
+ rwl_0_25 cell_2r1w
Xcell_2r1w_3644 vdd gnd read_bl_0_7 read_bl_1_7 write_bl_0_7 wwl_0_3 rwl_1_3 rwl_0_3
+ cell_2r1w
Xcell_2r1w_3633 vdd_uq6 gnd read_bl_0_7 read_bl_1_7 write_bl_0_7 wwl_0_14 rwl_1_14
+ rwl_0_14 cell_2r1w
Xcell_2r1w_3655 vdd_uq27 gnd read_bl_0_6 read_bl_1_6 write_bl_0_6 wwl_0_56 rwl_1_56
+ rwl_0_56 cell_2r1w
Xcell_2r1w_2954 vdd_uq25 gnd read_bl_0_17 read_bl_1_17 write_bl_0_17 wwl_0_53 rwl_1_53
+ rwl_0_53 cell_2r1w
Xcell_2r1w_3666 vdd_uq21 gnd read_bl_0_6 read_bl_1_6 write_bl_0_6 wwl_0_45 rwl_1_45
+ rwl_0_45 cell_2r1w
Xcell_2r1w_2965 vdd_uq20 gnd read_bl_0_17 read_bl_1_17 write_bl_0_17 wwl_0_42 rwl_1_42
+ rwl_0_42 cell_2r1w
Xcell_2r1w_3677 vdd_uq16 gnd read_bl_0_6 read_bl_1_6 write_bl_0_6 wwl_0_34 rwl_1_34
+ rwl_0_34 cell_2r1w
Xcell_2r1w_2910 vdd_uq15 gnd read_bl_0_18 read_bl_1_18 write_bl_0_18 wwl_0_33 rwl_1_33
+ rwl_0_33 cell_2r1w
Xcell_2r1w_2976 vdd_uq14 gnd read_bl_0_17 read_bl_1_17 write_bl_0_17 wwl_0_31 rwl_1_31
+ rwl_0_31 cell_2r1w
Xcell_2r1w_2943 vdd_uq0 gnd read_bl_0_18 read_bl_1_18 write_bl_0_18 wwl_0_0 rwl_1_0
+ rwl_0_0 cell_2r1w
Xcell_2r1w_2998 vdd_uq3 gnd read_bl_0_17 read_bl_1_17 write_bl_0_17 wwl_0_9 rwl_1_9
+ rwl_0_9 cell_2r1w
Xcell_2r1w_2932 vdd_uq4 gnd read_bl_0_18 read_bl_1_18 write_bl_0_18 wwl_0_11 rwl_1_11
+ rwl_0_11 cell_2r1w
Xcell_2r1w_3699 vdd_uq5 gnd read_bl_0_6 read_bl_1_6 write_bl_0_6 wwl_0_12 rwl_1_12
+ rwl_0_12 cell_2r1w
Xcell_2r1w_2987 vdd_uq9 gnd read_bl_0_17 read_bl_1_17 write_bl_0_17 wwl_0_20 rwl_1_20
+ rwl_0_20 cell_2r1w
Xcell_2r1w_2921 vdd_uq10 gnd read_bl_0_18 read_bl_1_18 write_bl_0_18 wwl_0_22 rwl_1_22
+ rwl_0_22 cell_2r1w
Xcell_2r1w_3688 vdd_uq10 gnd read_bl_0_6 read_bl_1_6 write_bl_0_6 wwl_0_23 rwl_1_23
+ rwl_0_23 cell_2r1w
Xcell_2r1w_69 vdd_uq28 gnd read_bl_0_62 read_bl_1_62 write_bl_0_62 wwl_0_58 rwl_1_58
+ rwl_0_58 cell_2r1w
Xcell_2r1w_14 vdd_uq23 gnd read_bl_0_63 read_bl_1_63 write_bl_0_63 wwl_0_49 rwl_1_49
+ rwl_0_49 cell_2r1w
Xcell_2r1w_25 vdd_uq18 gnd read_bl_0_63 read_bl_1_63 write_bl_0_63 wwl_0_38 rwl_1_38
+ rwl_0_38 cell_2r1w
Xcell_2r1w_36 vdd_uq12 gnd read_bl_0_63 read_bl_1_63 write_bl_0_63 wwl_0_27 rwl_1_27
+ rwl_0_27 cell_2r1w
Xcell_2r1w_58 vdd_uq1 gnd read_bl_0_63 read_bl_1_63 write_bl_0_63 wwl_0_5 rwl_1_5
+ rwl_0_5 cell_2r1w
Xcell_2r1w_47 vdd_uq7 gnd read_bl_0_63 read_bl_1_63 write_bl_0_63 wwl_0_16 rwl_1_16
+ rwl_0_16 cell_2r1w
Xcell_2r1w_209 vdd_uq22 gnd read_bl_0_60 read_bl_1_60 write_bl_0_60 wwl_0_46 rwl_1_46
+ rwl_0_46 cell_2r1w
Xcell_2r1w_1538 vdd_uq29 gnd read_bl_0_39 read_bl_1_39 write_bl_0_39 wwl_0_61 rwl_1_61
+ rwl_0_61 cell_2r1w
Xcell_2r1w_710 vdd_uq27 gnd read_bl_0_52 read_bl_1_52 write_bl_0_52 wwl_0_57 rwl_1_57
+ rwl_0_57 cell_2r1w
Xcell_2r1w_1549 vdd_uq24 gnd read_bl_0_39 read_bl_1_39 write_bl_0_39 wwl_0_50 rwl_1_50
+ rwl_0_50 cell_2r1w
Xcell_2r1w_721 vdd_uq22 gnd read_bl_0_52 read_bl_1_52 write_bl_0_52 wwl_0_46 rwl_1_46
+ rwl_0_46 cell_2r1w
Xcell_2r1w_732 vdd_uq16 gnd read_bl_0_52 read_bl_1_52 write_bl_0_52 wwl_0_35 rwl_1_35
+ rwl_0_35 cell_2r1w
Xcell_2r1w_2206 vdd_uq15 gnd read_bl_0_29 read_bl_1_29 write_bl_0_29 wwl_0_33 rwl_1_33
+ rwl_0_33 cell_2r1w
Xcell_2r1w_1505 vdd_uq14 gnd read_bl_0_40 read_bl_1_40 write_bl_0_40 wwl_0_30 rwl_1_30
+ rwl_0_30 cell_2r1w
Xcell_2r1w_743 vdd_uq11 gnd read_bl_0_52 read_bl_1_52 write_bl_0_52 wwl_0_24 rwl_1_24
+ rwl_0_24 cell_2r1w
Xcell_2r1w_2239 vdd_uq0 gnd read_bl_0_29 read_bl_1_29 write_bl_0_29 wwl_0_0 rwl_1_0
+ rwl_0_0 cell_2r1w
Xcell_2r1w_1527 vdd_uq3 gnd read_bl_0_40 read_bl_1_40 write_bl_0_40 wwl_0_8 rwl_1_8
+ rwl_0_8 cell_2r1w
Xcell_2r1w_2228 vdd_uq4 gnd read_bl_0_29 read_bl_1_29 write_bl_0_29 wwl_0_11 rwl_1_11
+ rwl_0_11 cell_2r1w
Xcell_2r1w_754 vdd_uq5 gnd read_bl_0_52 read_bl_1_52 write_bl_0_52 wwl_0_13 rwl_1_13
+ rwl_0_13 cell_2r1w
Xcell_2r1w_1516 vdd_uq8 gnd read_bl_0_40 read_bl_1_40 write_bl_0_40 wwl_0_19 rwl_1_19
+ rwl_0_19 cell_2r1w
Xcell_2r1w_2217 vdd_uq10 gnd read_bl_0_29 read_bl_1_29 write_bl_0_29 wwl_0_22 rwl_1_22
+ rwl_0_22 cell_2r1w
Xcell_2r1w_776 vdd_uq26 gnd read_bl_0_51 read_bl_1_51 write_bl_0_51 wwl_0_55 rwl_1_55
+ rwl_0_55 cell_2r1w
Xcell_2r1w_787 vdd_uq21 gnd read_bl_0_51 read_bl_1_51 write_bl_0_51 wwl_0_44 rwl_1_44
+ rwl_0_44 cell_2r1w
Xcell_2r1w_798 vdd_uq15 gnd read_bl_0_51 read_bl_1_51 write_bl_0_51 wwl_0_33 rwl_1_33
+ rwl_0_33 cell_2r1w
Xcell_2r1w_765 vdd gnd read_bl_0_52 read_bl_1_52 write_bl_0_52 wwl_0_2 rwl_1_2 rwl_0_2
+ cell_2r1w
Xcell_2r1w_4 vdd_uq28 gnd read_bl_0_63 read_bl_1_63 write_bl_0_63 wwl_0_59 rwl_1_59
+ rwl_0_59 cell_2r1w
Xcell_2r1w_3463 vdd_uq27 gnd read_bl_0_9 read_bl_1_9 write_bl_0_9 wwl_0_56 rwl_1_56
+ rwl_0_56 cell_2r1w
Xcell_2r1w_3474 vdd_uq21 gnd read_bl_0_9 read_bl_1_9 write_bl_0_9 wwl_0_45 rwl_1_45
+ rwl_0_45 cell_2r1w
Xcell_2r1w_3485 vdd_uq16 gnd read_bl_0_9 read_bl_1_9 write_bl_0_9 wwl_0_34 rwl_1_34
+ rwl_0_34 cell_2r1w
Xcell_2r1w_3430 vdd_uq11 gnd read_bl_0_10 read_bl_1_10 write_bl_0_10 wwl_0_25 rwl_1_25
+ rwl_0_25 cell_2r1w
Xcell_2r1w_3452 vdd gnd read_bl_0_10 read_bl_1_10 write_bl_0_10 wwl_0_3 rwl_1_3 rwl_0_3
+ cell_2r1w
Xcell_2r1w_2751 vdd_uq0 gnd read_bl_0_21 read_bl_1_21 write_bl_0_21 wwl_0_0 rwl_1_0
+ rwl_0_0 cell_2r1w
Xcell_2r1w_2740 vdd_uq4 gnd read_bl_0_21 read_bl_1_21 write_bl_0_21 wwl_0_11 rwl_1_11
+ rwl_0_11 cell_2r1w
Xcell_2r1w_3441 vdd_uq6 gnd read_bl_0_10 read_bl_1_10 write_bl_0_10 wwl_0_14 rwl_1_14
+ rwl_0_14 cell_2r1w
Xcell_2r1w_3496 vdd_uq10 gnd read_bl_0_9 read_bl_1_9 write_bl_0_9 wwl_0_23 rwl_1_23
+ rwl_0_23 cell_2r1w
Xcell_2r1w_2762 vdd_uq25 gnd read_bl_0_20 read_bl_1_20 write_bl_0_20 wwl_0_53 rwl_1_53
+ rwl_0_53 cell_2r1w
Xcell_2r1w_2773 vdd_uq20 gnd read_bl_0_20 read_bl_1_20 write_bl_0_20 wwl_0_42 rwl_1_42
+ rwl_0_42 cell_2r1w
Xcell_2r1w_2784 vdd_uq14 gnd read_bl_0_20 read_bl_1_20 write_bl_0_20 wwl_0_31 rwl_1_31
+ rwl_0_31 cell_2r1w
Xcell_2r1w_2795 vdd_uq9 gnd read_bl_0_20 read_bl_1_20 write_bl_0_20 wwl_0_20 rwl_1_20
+ rwl_0_20 cell_2r1w
Xcell_2r1w_2003 vdd_uq21 gnd read_bl_0_32 read_bl_1_32 write_bl_0_32 wwl_0_44 rwl_1_44
+ rwl_0_44 cell_2r1w
Xcell_2r1w_1302 vdd_uq19 gnd read_bl_0_43 read_bl_1_43 write_bl_0_43 wwl_0_41 rwl_1_41
+ rwl_0_41 cell_2r1w
Xcell_2r1w_2014 vdd_uq15 gnd read_bl_0_32 read_bl_1_32 write_bl_0_32 wwl_0_33 rwl_1_33
+ rwl_0_33 cell_2r1w
Xcell_2r1w_2047 vdd_uq0 gnd read_bl_0_32 read_bl_1_32 write_bl_0_32 wwl_0_0 rwl_1_0
+ rwl_0_0 cell_2r1w
Xcell_2r1w_2036 vdd_uq4 gnd read_bl_0_32 read_bl_1_32 write_bl_0_32 wwl_0_11 rwl_1_11
+ rwl_0_11 cell_2r1w
Xcell_2r1w_2025 vdd_uq10 gnd read_bl_0_32 read_bl_1_32 write_bl_0_32 wwl_0_22 rwl_1_22
+ rwl_0_22 cell_2r1w
Xcell_2r1w_1346 vdd_uq29 gnd read_bl_0_42 read_bl_1_42 write_bl_0_42 wwl_0_61 rwl_1_61
+ rwl_0_61 cell_2r1w
Xcell_2r1w_584 vdd_uq26 gnd read_bl_0_54 read_bl_1_54 write_bl_0_54 wwl_0_55 rwl_1_55
+ rwl_0_55 cell_2r1w
Xcell_2r1w_2058 vdd_uq25 gnd read_bl_0_31 read_bl_1_31 write_bl_0_31 wwl_0_53 rwl_1_53
+ rwl_0_53 cell_2r1w
Xcell_2r1w_1357 vdd_uq24 gnd read_bl_0_42 read_bl_1_42 write_bl_0_42 wwl_0_50 rwl_1_50
+ rwl_0_50 cell_2r1w
Xcell_2r1w_595 vdd_uq21 gnd read_bl_0_54 read_bl_1_54 write_bl_0_54 wwl_0_44 rwl_1_44
+ rwl_0_44 cell_2r1w
Xcell_2r1w_2069 vdd_uq20 gnd read_bl_0_31 read_bl_1_31 write_bl_0_31 wwl_0_42 rwl_1_42
+ rwl_0_42 cell_2r1w
Xcell_2r1w_1368 vdd_uq18 gnd read_bl_0_42 read_bl_1_42 write_bl_0_42 wwl_0_39 rwl_1_39
+ rwl_0_39 cell_2r1w
Xcell_2r1w_540 vdd_uq16 gnd read_bl_0_55 read_bl_1_55 write_bl_0_55 wwl_0_35 rwl_1_35
+ rwl_0_35 cell_2r1w
Xcell_2r1w_1313 vdd_uq14 gnd read_bl_0_43 read_bl_1_43 write_bl_0_43 wwl_0_30 rwl_1_30
+ rwl_0_30 cell_2r1w
Xcell_2r1w_1379 vdd_uq13 gnd read_bl_0_42 read_bl_1_42 write_bl_0_42 wwl_0_28 rwl_1_28
+ rwl_0_28 cell_2r1w
Xcell_2r1w_551 vdd_uq11 gnd read_bl_0_55 read_bl_1_55 write_bl_0_55 wwl_0_24 rwl_1_24
+ rwl_0_24 cell_2r1w
Xcell_2r1w_573 vdd gnd read_bl_0_55 read_bl_1_55 write_bl_0_55 wwl_0_2 rwl_1_2 rwl_0_2
+ cell_2r1w
Xcell_2r1w_1335 vdd_uq3 gnd read_bl_0_43 read_bl_1_43 write_bl_0_43 wwl_0_8 rwl_1_8
+ rwl_0_8 cell_2r1w
Xcell_2r1w_562 vdd_uq5 gnd read_bl_0_55 read_bl_1_55 write_bl_0_55 wwl_0_13 rwl_1_13
+ rwl_0_13 cell_2r1w
Xcell_2r1w_1324 vdd_uq8 gnd read_bl_0_43 read_bl_1_43 write_bl_0_43 wwl_0_19 rwl_1_19
+ rwl_0_19 cell_2r1w
Xcell_2r1w_3271 vdd_uq27 gnd read_bl_0_12 read_bl_1_12 write_bl_0_12 wwl_0_56 rwl_1_56
+ rwl_0_56 cell_2r1w
Xcell_2r1w_2570 vdd_uq25 gnd read_bl_0_23 read_bl_1_23 write_bl_0_23 wwl_0_53 rwl_1_53
+ rwl_0_53 cell_2r1w
Xcell_2r1w_3282 vdd_uq21 gnd read_bl_0_12 read_bl_1_12 write_bl_0_12 wwl_0_45 rwl_1_45
+ rwl_0_45 cell_2r1w
Xcell_2r1w_2581 vdd_uq20 gnd read_bl_0_23 read_bl_1_23 write_bl_0_23 wwl_0_42 rwl_1_42
+ rwl_0_42 cell_2r1w
Xcell_2r1w_3293 vdd_uq16 gnd read_bl_0_12 read_bl_1_12 write_bl_0_12 wwl_0_34 rwl_1_34
+ rwl_0_34 cell_2r1w
Xcell_2r1w_2592 vdd_uq14 gnd read_bl_0_23 read_bl_1_23 write_bl_0_23 wwl_0_31 rwl_1_31
+ rwl_0_31 cell_2r1w
Xcell_2r1w_3260 vdd gnd read_bl_0_13 read_bl_1_13 write_bl_0_13 wwl_0_3 rwl_1_3 rwl_0_3
+ cell_2r1w
Xcell_2r1w_1880 vdd_uq18 gnd read_bl_0_34 read_bl_1_34 write_bl_0_34 wwl_0_39 rwl_1_39
+ rwl_0_39 cell_2r1w
Xcell_2r1w_1891 vdd_uq13 gnd read_bl_0_34 read_bl_1_34 write_bl_0_34 wwl_0_28 rwl_1_28
+ rwl_0_28 cell_2r1w
Xcell_2r1w_1110 vdd_uq19 gnd read_bl_0_46 read_bl_1_46 write_bl_0_46 wwl_0_41 rwl_1_41
+ rwl_0_41 cell_2r1w
Xcell_2r1w_1121 vdd_uq14 gnd read_bl_0_46 read_bl_1_46 write_bl_0_46 wwl_0_30 rwl_1_30
+ rwl_0_30 cell_2r1w
Xcell_2r1w_1143 vdd_uq3 gnd read_bl_0_46 read_bl_1_46 write_bl_0_46 wwl_0_8 rwl_1_8
+ rwl_0_8 cell_2r1w
Xcell_2r1w_1132 vdd_uq8 gnd read_bl_0_46 read_bl_1_46 write_bl_0_46 wwl_0_19 rwl_1_19
+ rwl_0_19 cell_2r1w
Xcell_2r1w_1154 vdd_uq29 gnd read_bl_0_45 read_bl_1_45 write_bl_0_45 wwl_0_61 rwl_1_61
+ rwl_0_61 cell_2r1w
Xcell_2r1w_392 vdd_uq26 gnd read_bl_0_57 read_bl_1_57 write_bl_0_57 wwl_0_55 rwl_1_55
+ rwl_0_55 cell_2r1w
Xcell_2r1w_1165 vdd_uq24 gnd read_bl_0_45 read_bl_1_45 write_bl_0_45 wwl_0_50 rwl_1_50
+ rwl_0_50 cell_2r1w
Xcell_2r1w_1176 vdd_uq18 gnd read_bl_0_45 read_bl_1_45 write_bl_0_45 wwl_0_39 rwl_1_39
+ rwl_0_39 cell_2r1w
Xcell_2r1w_1187 vdd_uq13 gnd read_bl_0_45 read_bl_1_45 write_bl_0_45 wwl_0_28 rwl_1_28
+ rwl_0_28 cell_2r1w
Xcell_2r1w_381 vdd gnd read_bl_0_58 read_bl_1_58 write_bl_0_58 wwl_0_2 rwl_1_2 rwl_0_2
+ cell_2r1w
Xcell_2r1w_370 vdd_uq5 gnd read_bl_0_58 read_bl_1_58 write_bl_0_58 wwl_0_13 rwl_1_13
+ rwl_0_13 cell_2r1w
Xcell_2r1w_1198 vdd_uq7 gnd read_bl_0_45 read_bl_1_45 write_bl_0_45 wwl_0_17 rwl_1_17
+ rwl_0_17 cell_2r1w
Xcell_2r1w_3090 vdd_uq21 gnd read_bl_0_15 read_bl_1_15 write_bl_0_15 wwl_0_45 rwl_1_45
+ rwl_0_45 cell_2r1w
Xcell_2r1w_3804 vdd_uq16 gnd read_bl_0_4 read_bl_1_4 write_bl_0_4 wwl_0_35 rwl_1_35
+ rwl_0_35 cell_2r1w
Xcell_2r1w_3815 vdd_uq11 gnd read_bl_0_4 read_bl_1_4 write_bl_0_4 wwl_0_24 rwl_1_24
+ rwl_0_24 cell_2r1w
Xcell_2r1w_3837 vdd gnd read_bl_0_4 read_bl_1_4 write_bl_0_4 wwl_0_2 rwl_1_2 rwl_0_2
+ cell_2r1w
Xcell_2r1w_3826 vdd_uq5 gnd read_bl_0_4 read_bl_1_4 write_bl_0_4 wwl_0_13 rwl_1_13
+ rwl_0_13 cell_2r1w
Xcell_2r1w_3848 vdd_uq26 gnd read_bl_0_3 read_bl_1_3 write_bl_0_3 wwl_0_55 rwl_1_55
+ rwl_0_55 cell_2r1w
Xcell_2r1w_3859 vdd_uq21 gnd read_bl_0_3 read_bl_1_3 write_bl_0_3 wwl_0_44 rwl_1_44
+ rwl_0_44 cell_2r1w
Xcell_2r1w_903 vdd_uq27 gnd read_bl_0_49 read_bl_1_49 write_bl_0_49 wwl_0_56 rwl_1_56
+ rwl_0_56 cell_2r1w
Xcell_2r1w_914 vdd_uq21 gnd read_bl_0_49 read_bl_1_49 write_bl_0_49 wwl_0_45 rwl_1_45
+ rwl_0_45 cell_2r1w
Xcell_2r1w_925 vdd_uq16 gnd read_bl_0_49 read_bl_1_49 write_bl_0_49 wwl_0_34 rwl_1_34
+ rwl_0_34 cell_2r1w
Xcell_2r1w_947 vdd_uq5 gnd read_bl_0_49 read_bl_1_49 write_bl_0_49 wwl_0_12 rwl_1_12
+ rwl_0_12 cell_2r1w
Xcell_2r1w_1709 vdd_uq8 gnd read_bl_0_37 read_bl_1_37 write_bl_0_37 wwl_0_18 rwl_1_18
+ rwl_0_18 cell_2r1w
Xcell_2r1w_936 vdd_uq10 gnd read_bl_0_49 read_bl_1_49 write_bl_0_49 wwl_0_23 rwl_1_23
+ rwl_0_23 cell_2r1w
Xcell_2r1w_969 vdd_uq26 gnd read_bl_0_48 read_bl_1_48 write_bl_0_48 wwl_0_54 rwl_1_54
+ rwl_0_54 cell_2r1w
Xcell_2r1w_958 vdd_uq0 gnd read_bl_0_49 read_bl_1_49 write_bl_0_49 wwl_0_1 rwl_1_1
+ rwl_0_1 cell_2r1w
Xcell_2r1w_3656 vdd_uq26 gnd read_bl_0_6 read_bl_1_6 write_bl_0_6 wwl_0_55 rwl_1_55
+ rwl_0_55 cell_2r1w
Xcell_2r1w_3601 vdd_uq22 gnd read_bl_0_7 read_bl_1_7 write_bl_0_7 wwl_0_46 rwl_1_46
+ rwl_0_46 cell_2r1w
Xcell_2r1w_3667 vdd_uq21 gnd read_bl_0_6 read_bl_1_6 write_bl_0_6 wwl_0_44 rwl_1_44
+ rwl_0_44 cell_2r1w
Xcell_2r1w_2900 vdd_uq20 gnd read_bl_0_18 read_bl_1_18 write_bl_0_18 wwl_0_43 rwl_1_43
+ rwl_0_43 cell_2r1w
Xcell_2r1w_3612 vdd_uq16 gnd read_bl_0_7 read_bl_1_7 write_bl_0_7 wwl_0_35 rwl_1_35
+ rwl_0_35 cell_2r1w
Xcell_2r1w_3678 vdd_uq15 gnd read_bl_0_6 read_bl_1_6 write_bl_0_6 wwl_0_33 rwl_1_33
+ rwl_0_33 cell_2r1w
Xcell_2r1w_2911 vdd_uq15 gnd read_bl_0_18 read_bl_1_18 write_bl_0_18 wwl_0_32 rwl_1_32
+ rwl_0_32 cell_2r1w
Xcell_2r1w_3623 vdd_uq11 gnd read_bl_0_7 read_bl_1_7 write_bl_0_7 wwl_0_24 rwl_1_24
+ rwl_0_24 cell_2r1w
Xcell_2r1w_3645 vdd gnd read_bl_0_7 read_bl_1_7 write_bl_0_7 wwl_0_2 rwl_1_2 rwl_0_2
+ cell_2r1w
Xcell_2r1w_2933 vdd_uq4 gnd read_bl_0_18 read_bl_1_18 write_bl_0_18 wwl_0_10 rwl_1_10
+ rwl_0_10 cell_2r1w
Xcell_2r1w_3634 vdd_uq5 gnd read_bl_0_7 read_bl_1_7 write_bl_0_7 wwl_0_13 rwl_1_13
+ rwl_0_13 cell_2r1w
Xcell_2r1w_2922 vdd_uq9 gnd read_bl_0_18 read_bl_1_18 write_bl_0_18 wwl_0_21 rwl_1_21
+ rwl_0_21 cell_2r1w
Xcell_2r1w_2944 vdd_uq30 gnd read_bl_0_17 read_bl_1_17 write_bl_0_17 wwl_0_63 rwl_1_63
+ rwl_0_63 cell_2r1w
Xcell_2r1w_2955 vdd_uq25 gnd read_bl_0_17 read_bl_1_17 write_bl_0_17 wwl_0_52 rwl_1_52
+ rwl_0_52 cell_2r1w
Xcell_2r1w_2966 vdd_uq19 gnd read_bl_0_17 read_bl_1_17 write_bl_0_17 wwl_0_41 rwl_1_41
+ rwl_0_41 cell_2r1w
Xcell_2r1w_2977 vdd_uq14 gnd read_bl_0_17 read_bl_1_17 write_bl_0_17 wwl_0_30 rwl_1_30
+ rwl_0_30 cell_2r1w
Xcell_2r1w_2999 vdd_uq3 gnd read_bl_0_17 read_bl_1_17 write_bl_0_17 wwl_0_8 rwl_1_8
+ rwl_0_8 cell_2r1w
Xcell_2r1w_2988 vdd_uq8 gnd read_bl_0_17 read_bl_1_17 write_bl_0_17 wwl_0_19 rwl_1_19
+ rwl_0_19 cell_2r1w
Xcell_2r1w_3689 vdd_uq10 gnd read_bl_0_6 read_bl_1_6 write_bl_0_6 wwl_0_22 rwl_1_22
+ rwl_0_22 cell_2r1w
Xcell_2r1w_15 vdd_uq23 gnd read_bl_0_63 read_bl_1_63 write_bl_0_63 wwl_0_48 rwl_1_48
+ rwl_0_48 cell_2r1w
Xcell_2r1w_26 vdd_uq17 gnd read_bl_0_63 read_bl_1_63 write_bl_0_63 wwl_0_37 rwl_1_37
+ rwl_0_37 cell_2r1w
Xcell_2r1w_37 vdd_uq12 gnd read_bl_0_63 read_bl_1_63 write_bl_0_63 wwl_0_26 rwl_1_26
+ rwl_0_26 cell_2r1w
Xcell_2r1w_59 vdd_uq1 gnd read_bl_0_63 read_bl_1_63 write_bl_0_63 wwl_0_4 rwl_1_4
+ rwl_0_4 cell_2r1w
Xcell_2r1w_48 vdd_uq6 gnd read_bl_0_63 read_bl_1_63 write_bl_0_63 wwl_0_15 rwl_1_15
+ rwl_0_15 cell_2r1w
Xcell_2r1w_2207 vdd_uq15 gnd read_bl_0_29 read_bl_1_29 write_bl_0_29 wwl_0_32 rwl_1_32
+ rwl_0_32 cell_2r1w
Xcell_2r1w_2229 vdd_uq4 gnd read_bl_0_29 read_bl_1_29 write_bl_0_29 wwl_0_10 rwl_1_10
+ rwl_0_10 cell_2r1w
Xcell_2r1w_2218 vdd_uq9 gnd read_bl_0_29 read_bl_1_29 write_bl_0_29 wwl_0_21 rwl_1_21
+ rwl_0_21 cell_2r1w
Xcell_2r1w_1539 vdd_uq29 gnd read_bl_0_39 read_bl_1_39 write_bl_0_39 wwl_0_60 rwl_1_60
+ rwl_0_60 cell_2r1w
Xcell_2r1w_711 vdd_uq27 gnd read_bl_0_52 read_bl_1_52 write_bl_0_52 wwl_0_56 rwl_1_56
+ rwl_0_56 cell_2r1w
Xcell_2r1w_777 vdd_uq26 gnd read_bl_0_51 read_bl_1_51 write_bl_0_51 wwl_0_54 rwl_1_54
+ rwl_0_54 cell_2r1w
Xcell_2r1w_722 vdd_uq21 gnd read_bl_0_52 read_bl_1_52 write_bl_0_52 wwl_0_45 rwl_1_45
+ rwl_0_45 cell_2r1w
Xcell_2r1w_788 vdd_uq20 gnd read_bl_0_51 read_bl_1_51 write_bl_0_51 wwl_0_43 rwl_1_43
+ rwl_0_43 cell_2r1w
Xcell_2r1w_733 vdd_uq16 gnd read_bl_0_52 read_bl_1_52 write_bl_0_52 wwl_0_34 rwl_1_34
+ rwl_0_34 cell_2r1w
Xcell_2r1w_1506 vdd_uq13 gnd read_bl_0_40 read_bl_1_40 write_bl_0_40 wwl_0_29 rwl_1_29
+ rwl_0_29 cell_2r1w
Xcell_2r1w_700 vdd gnd read_bl_0_53 read_bl_1_53 write_bl_0_53 wwl_0_3 rwl_1_3 rwl_0_3
+ cell_2r1w
Xcell_2r1w_766 vdd_uq0 gnd read_bl_0_52 read_bl_1_52 write_bl_0_52 wwl_0_1 rwl_1_1
+ rwl_0_1 cell_2r1w
Xcell_2r1w_1528 vdd_uq2 gnd read_bl_0_40 read_bl_1_40 write_bl_0_40 wwl_0_7 rwl_1_7
+ rwl_0_7 cell_2r1w
Xcell_2r1w_755 vdd_uq5 gnd read_bl_0_52 read_bl_1_52 write_bl_0_52 wwl_0_12 rwl_1_12
+ rwl_0_12 cell_2r1w
Xcell_2r1w_1517 vdd_uq8 gnd read_bl_0_40 read_bl_1_40 write_bl_0_40 wwl_0_18 rwl_1_18
+ rwl_0_18 cell_2r1w
Xcell_2r1w_744 vdd_uq10 gnd read_bl_0_52 read_bl_1_52 write_bl_0_52 wwl_0_23 rwl_1_23
+ rwl_0_23 cell_2r1w
Xcell_2r1w_799 vdd_uq15 gnd read_bl_0_51 read_bl_1_51 write_bl_0_51 wwl_0_32 rwl_1_32
+ rwl_0_32 cell_2r1w
Xcell_2r1w_5 vdd_uq28 gnd read_bl_0_63 read_bl_1_63 write_bl_0_63 wwl_0_58 rwl_1_58
+ rwl_0_58 cell_2r1w
Xcell_2r1w_2752 vdd_uq30 gnd read_bl_0_20 read_bl_1_20 write_bl_0_20 wwl_0_63 rwl_1_63
+ rwl_0_63 cell_2r1w
Xcell_2r1w_3464 vdd_uq26 gnd read_bl_0_9 read_bl_1_9 write_bl_0_9 wwl_0_55 rwl_1_55
+ rwl_0_55 cell_2r1w
Xcell_2r1w_2763 vdd_uq25 gnd read_bl_0_20 read_bl_1_20 write_bl_0_20 wwl_0_52 rwl_1_52
+ rwl_0_52 cell_2r1w
Xcell_2r1w_3475 vdd_uq21 gnd read_bl_0_9 read_bl_1_9 write_bl_0_9 wwl_0_44 rwl_1_44
+ rwl_0_44 cell_2r1w
Xcell_2r1w_2774 vdd_uq19 gnd read_bl_0_20 read_bl_1_20 write_bl_0_20 wwl_0_41 rwl_1_41
+ rwl_0_41 cell_2r1w
Xcell_2r1w_3420 vdd_uq16 gnd read_bl_0_10 read_bl_1_10 write_bl_0_10 wwl_0_35 rwl_1_35
+ rwl_0_35 cell_2r1w
Xcell_2r1w_3486 vdd_uq15 gnd read_bl_0_9 read_bl_1_9 write_bl_0_9 wwl_0_33 rwl_1_33
+ rwl_0_33 cell_2r1w
Xcell_2r1w_2785 vdd_uq14 gnd read_bl_0_20 read_bl_1_20 write_bl_0_20 wwl_0_30 rwl_1_30
+ rwl_0_30 cell_2r1w
Xcell_2r1w_3431 vdd_uq11 gnd read_bl_0_10 read_bl_1_10 write_bl_0_10 wwl_0_24 rwl_1_24
+ rwl_0_24 cell_2r1w
Xcell_2r1w_3453 vdd gnd read_bl_0_10 read_bl_1_10 write_bl_0_10 wwl_0_2 rwl_1_2 rwl_0_2
+ cell_2r1w
Xcell_2r1w_2741 vdd_uq4 gnd read_bl_0_21 read_bl_1_21 write_bl_0_21 wwl_0_10 rwl_1_10
+ rwl_0_10 cell_2r1w
Xcell_2r1w_3442 vdd_uq5 gnd read_bl_0_10 read_bl_1_10 write_bl_0_10 wwl_0_13 rwl_1_13
+ rwl_0_13 cell_2r1w
Xcell_2r1w_2730 vdd_uq9 gnd read_bl_0_21 read_bl_1_21 write_bl_0_21 wwl_0_21 rwl_1_21
+ rwl_0_21 cell_2r1w
Xcell_2r1w_3497 vdd_uq10 gnd read_bl_0_9 read_bl_1_9 write_bl_0_9 wwl_0_22 rwl_1_22
+ rwl_0_22 cell_2r1w
Xcell_2r1w_2796 vdd_uq8 gnd read_bl_0_20 read_bl_1_20 write_bl_0_20 wwl_0_19 rwl_1_19
+ rwl_0_19 cell_2r1w
Xcell_2r1w_2048 vdd_uq30 gnd read_bl_0_31 read_bl_1_31 write_bl_0_31 wwl_0_63 rwl_1_63
+ rwl_0_63 cell_2r1w
Xcell_2r1w_2059 vdd_uq25 gnd read_bl_0_31 read_bl_1_31 write_bl_0_31 wwl_0_52 rwl_1_52
+ rwl_0_52 cell_2r1w
Xcell_2r1w_2004 vdd_uq20 gnd read_bl_0_32 read_bl_1_32 write_bl_0_32 wwl_0_43 rwl_1_43
+ rwl_0_43 cell_2r1w
Xcell_2r1w_1303 vdd_uq19 gnd read_bl_0_43 read_bl_1_43 write_bl_0_43 wwl_0_40 rwl_1_40
+ rwl_0_40 cell_2r1w
Xcell_2r1w_2015 vdd_uq15 gnd read_bl_0_32 read_bl_1_32 write_bl_0_32 wwl_0_32 rwl_1_32
+ rwl_0_32 cell_2r1w
Xcell_2r1w_1314 vdd_uq13 gnd read_bl_0_43 read_bl_1_43 write_bl_0_43 wwl_0_29 rwl_1_29
+ rwl_0_29 cell_2r1w
Xcell_2r1w_2037 vdd_uq4 gnd read_bl_0_32 read_bl_1_32 write_bl_0_32 wwl_0_10 rwl_1_10
+ rwl_0_10 cell_2r1w
Xcell_2r1w_1325 vdd_uq8 gnd read_bl_0_43 read_bl_1_43 write_bl_0_43 wwl_0_18 rwl_1_18
+ rwl_0_18 cell_2r1w
Xcell_2r1w_2026 vdd_uq9 gnd read_bl_0_32 read_bl_1_32 write_bl_0_32 wwl_0_21 rwl_1_21
+ rwl_0_21 cell_2r1w
Xcell_2r1w_1347 vdd_uq29 gnd read_bl_0_42 read_bl_1_42 write_bl_0_42 wwl_0_60 rwl_1_60
+ rwl_0_60 cell_2r1w
Xcell_2r1w_585 vdd_uq26 gnd read_bl_0_54 read_bl_1_54 write_bl_0_54 wwl_0_54 rwl_1_54
+ rwl_0_54 cell_2r1w
Xcell_2r1w_1358 vdd_uq23 gnd read_bl_0_42 read_bl_1_42 write_bl_0_42 wwl_0_49 rwl_1_49
+ rwl_0_49 cell_2r1w
Xcell_2r1w_530 vdd_uq21 gnd read_bl_0_55 read_bl_1_55 write_bl_0_55 wwl_0_45 rwl_1_45
+ rwl_0_45 cell_2r1w
Xcell_2r1w_596 vdd_uq20 gnd read_bl_0_54 read_bl_1_54 write_bl_0_54 wwl_0_43 rwl_1_43
+ rwl_0_43 cell_2r1w
Xcell_2r1w_1369 vdd_uq18 gnd read_bl_0_42 read_bl_1_42 write_bl_0_42 wwl_0_38 rwl_1_38
+ rwl_0_38 cell_2r1w
Xcell_2r1w_541 vdd_uq16 gnd read_bl_0_55 read_bl_1_55 write_bl_0_55 wwl_0_34 rwl_1_34
+ rwl_0_34 cell_2r1w
Xcell_2r1w_574 vdd_uq0 gnd read_bl_0_55 read_bl_1_55 write_bl_0_55 wwl_0_1 rwl_1_1
+ rwl_0_1 cell_2r1w
Xcell_2r1w_1336 vdd_uq2 gnd read_bl_0_43 read_bl_1_43 write_bl_0_43 wwl_0_7 rwl_1_7
+ rwl_0_7 cell_2r1w
Xcell_2r1w_563 vdd_uq5 gnd read_bl_0_55 read_bl_1_55 write_bl_0_55 wwl_0_12 rwl_1_12
+ rwl_0_12 cell_2r1w
Xcell_2r1w_552 vdd_uq10 gnd read_bl_0_55 read_bl_1_55 write_bl_0_55 wwl_0_23 rwl_1_23
+ rwl_0_23 cell_2r1w
Xcell_2r1w_2560 vdd_uq30 gnd read_bl_0_23 read_bl_1_23 write_bl_0_23 wwl_0_63 rwl_1_63
+ rwl_0_63 cell_2r1w
Xcell_2r1w_3272 vdd_uq26 gnd read_bl_0_12 read_bl_1_12 write_bl_0_12 wwl_0_55 rwl_1_55
+ rwl_0_55 cell_2r1w
Xcell_2r1w_2571 vdd_uq25 gnd read_bl_0_23 read_bl_1_23 write_bl_0_23 wwl_0_52 rwl_1_52
+ rwl_0_52 cell_2r1w
Xcell_2r1w_1870 vdd_uq23 gnd read_bl_0_34 read_bl_1_34 write_bl_0_34 wwl_0_49 rwl_1_49
+ rwl_0_49 cell_2r1w
Xcell_2r1w_3283 vdd_uq21 gnd read_bl_0_12 read_bl_1_12 write_bl_0_12 wwl_0_44 rwl_1_44
+ rwl_0_44 cell_2r1w
Xcell_2r1w_2582 vdd_uq19 gnd read_bl_0_23 read_bl_1_23 write_bl_0_23 wwl_0_41 rwl_1_41
+ rwl_0_41 cell_2r1w
Xcell_2r1w_1881 vdd_uq18 gnd read_bl_0_34 read_bl_1_34 write_bl_0_34 wwl_0_38 rwl_1_38
+ rwl_0_38 cell_2r1w
Xcell_2r1w_3294 vdd_uq15 gnd read_bl_0_12 read_bl_1_12 write_bl_0_12 wwl_0_33 rwl_1_33
+ rwl_0_33 cell_2r1w
Xcell_2r1w_2593 vdd_uq14 gnd read_bl_0_23 read_bl_1_23 write_bl_0_23 wwl_0_30 rwl_1_30
+ rwl_0_30 cell_2r1w
Xcell_2r1w_3261 vdd gnd read_bl_0_13 read_bl_1_13 write_bl_0_13 wwl_0_2 rwl_1_2 rwl_0_2
+ cell_2r1w
Xcell_2r1w_3250 vdd_uq5 gnd read_bl_0_13 read_bl_1_13 write_bl_0_13 wwl_0_13 rwl_1_13
+ rwl_0_13 cell_2r1w
Xcell_2r1w_1892 vdd_uq12 gnd read_bl_0_34 read_bl_1_34 write_bl_0_34 wwl_0_27 rwl_1_27
+ rwl_0_27 cell_2r1w
Xcell_2r1w_1155 vdd_uq29 gnd read_bl_0_45 read_bl_1_45 write_bl_0_45 wwl_0_60 rwl_1_60
+ rwl_0_60 cell_2r1w
Xcell_2r1w_1100 vdd_uq24 gnd read_bl_0_46 read_bl_1_46 write_bl_0_46 wwl_0_51 rwl_1_51
+ rwl_0_51 cell_2r1w
Xcell_2r1w_1166 vdd_uq23 gnd read_bl_0_45 read_bl_1_45 write_bl_0_45 wwl_0_49 rwl_1_49
+ rwl_0_49 cell_2r1w
Xcell_2r1w_1111 vdd_uq19 gnd read_bl_0_46 read_bl_1_46 write_bl_0_46 wwl_0_40 rwl_1_40
+ rwl_0_40 cell_2r1w
Xcell_2r1w_1177 vdd_uq18 gnd read_bl_0_45 read_bl_1_45 write_bl_0_45 wwl_0_38 rwl_1_38
+ rwl_0_38 cell_2r1w
Xcell_2r1w_1122 vdd_uq13 gnd read_bl_0_46 read_bl_1_46 write_bl_0_46 wwl_0_29 rwl_1_29
+ rwl_0_29 cell_2r1w
Xcell_2r1w_1144 vdd_uq2 gnd read_bl_0_46 read_bl_1_46 write_bl_0_46 wwl_0_7 rwl_1_7
+ rwl_0_7 cell_2r1w
Xcell_2r1w_1133 vdd_uq8 gnd read_bl_0_46 read_bl_1_46 write_bl_0_46 wwl_0_18 rwl_1_18
+ rwl_0_18 cell_2r1w
Xcell_2r1w_393 vdd_uq26 gnd read_bl_0_57 read_bl_1_57 write_bl_0_57 wwl_0_54 rwl_1_54
+ rwl_0_54 cell_2r1w
Xcell_2r1w_1188 vdd_uq12 gnd read_bl_0_45 read_bl_1_45 write_bl_0_45 wwl_0_27 rwl_1_27
+ rwl_0_27 cell_2r1w
Xcell_2r1w_382 vdd_uq0 gnd read_bl_0_58 read_bl_1_58 write_bl_0_58 wwl_0_1 rwl_1_1
+ rwl_0_1 cell_2r1w
Xcell_2r1w_371 vdd_uq5 gnd read_bl_0_58 read_bl_1_58 write_bl_0_58 wwl_0_12 rwl_1_12
+ rwl_0_12 cell_2r1w
Xcell_2r1w_1199 vdd_uq7 gnd read_bl_0_45 read_bl_1_45 write_bl_0_45 wwl_0_16 rwl_1_16
+ rwl_0_16 cell_2r1w
Xcell_2r1w_360 vdd_uq10 gnd read_bl_0_58 read_bl_1_58 write_bl_0_58 wwl_0_23 rwl_1_23
+ rwl_0_23 cell_2r1w
Xcell_2r1w_3080 vdd_uq26 gnd read_bl_0_15 read_bl_1_15 write_bl_0_15 wwl_0_55 rwl_1_55
+ rwl_0_55 cell_2r1w
Xcell_2r1w_3091 vdd_uq21 gnd read_bl_0_15 read_bl_1_15 write_bl_0_15 wwl_0_44 rwl_1_44
+ rwl_0_44 cell_2r1w
Xcell_2r1w_2390 vdd_uq19 gnd read_bl_0_26 read_bl_1_26 write_bl_0_26 wwl_0_41 rwl_1_41
+ rwl_0_41 cell_2r1w
Xcell_2r1w_190 vdd_uq0 gnd read_bl_0_61 read_bl_1_61 write_bl_0_61 wwl_0_1 rwl_1_1
+ rwl_0_1 cell_2r1w
Xcell_2r1w_3849 vdd_uq26 gnd read_bl_0_3 read_bl_1_3 write_bl_0_3 wwl_0_54 rwl_1_54
+ rwl_0_54 cell_2r1w
Xcell_2r1w_3805 vdd_uq16 gnd read_bl_0_4 read_bl_1_4 write_bl_0_4 wwl_0_34 rwl_1_34
+ rwl_0_34 cell_2r1w
Xcell_2r1w_3838 vdd_uq0 gnd read_bl_0_4 read_bl_1_4 write_bl_0_4 wwl_0_1 rwl_1_1 rwl_0_1
+ cell_2r1w
Xcell_2r1w_3827 vdd_uq5 gnd read_bl_0_4 read_bl_1_4 write_bl_0_4 wwl_0_12 rwl_1_12
+ rwl_0_12 cell_2r1w
Xcell_2r1w_3816 vdd_uq10 gnd read_bl_0_4 read_bl_1_4 write_bl_0_4 wwl_0_23 rwl_1_23
+ rwl_0_23 cell_2r1w
Xcell_2r1w_904 vdd_uq26 gnd read_bl_0_49 read_bl_1_49 write_bl_0_49 wwl_0_55 rwl_1_55
+ rwl_0_55 cell_2r1w
Xcell_2r1w_915 vdd_uq21 gnd read_bl_0_49 read_bl_1_49 write_bl_0_49 wwl_0_44 rwl_1_44
+ rwl_0_44 cell_2r1w
Xcell_2r1w_926 vdd_uq15 gnd read_bl_0_49 read_bl_1_49 write_bl_0_49 wwl_0_33 rwl_1_33
+ rwl_0_33 cell_2r1w
Xcell_2r1w_959 vdd_uq0 gnd read_bl_0_49 read_bl_1_49 write_bl_0_49 wwl_0_0 rwl_1_0
+ rwl_0_0 cell_2r1w
Xcell_2r1w_948 vdd_uq4 gnd read_bl_0_49 read_bl_1_49 write_bl_0_49 wwl_0_11 rwl_1_11
+ rwl_0_11 cell_2r1w
Xcell_2r1w_937 vdd_uq10 gnd read_bl_0_49 read_bl_1_49 write_bl_0_49 wwl_0_22 rwl_1_22
+ rwl_0_22 cell_2r1w
Xcell_2r1w_2945 vdd_uq30 gnd read_bl_0_17 read_bl_1_17 write_bl_0_17 wwl_0_62 rwl_1_62
+ rwl_0_62 cell_2r1w
Xcell_2r1w_3657 vdd_uq26 gnd read_bl_0_6 read_bl_1_6 write_bl_0_6 wwl_0_54 rwl_1_54
+ rwl_0_54 cell_2r1w
Xcell_2r1w_2956 vdd_uq24 gnd read_bl_0_17 read_bl_1_17 write_bl_0_17 wwl_0_51 rwl_1_51
+ rwl_0_51 cell_2r1w
Xcell_2r1w_3602 vdd_uq21 gnd read_bl_0_7 read_bl_1_7 write_bl_0_7 wwl_0_45 rwl_1_45
+ rwl_0_45 cell_2r1w
Xcell_2r1w_3668 vdd_uq20 gnd read_bl_0_6 read_bl_1_6 write_bl_0_6 wwl_0_43 rwl_1_43
+ rwl_0_43 cell_2r1w
Xcell_2r1w_2901 vdd_uq20 gnd read_bl_0_18 read_bl_1_18 write_bl_0_18 wwl_0_42 rwl_1_42
+ rwl_0_42 cell_2r1w
Xcell_2r1w_2967 vdd_uq19 gnd read_bl_0_17 read_bl_1_17 write_bl_0_17 wwl_0_40 rwl_1_40
+ rwl_0_40 cell_2r1w
Xcell_2r1w_3613 vdd_uq16 gnd read_bl_0_7 read_bl_1_7 write_bl_0_7 wwl_0_34 rwl_1_34
+ rwl_0_34 cell_2r1w
Xcell_2r1w_3679 vdd_uq15 gnd read_bl_0_6 read_bl_1_6 write_bl_0_6 wwl_0_32 rwl_1_32
+ rwl_0_32 cell_2r1w
Xcell_2r1w_2912 vdd_uq14 gnd read_bl_0_18 read_bl_1_18 write_bl_0_18 wwl_0_31 rwl_1_31
+ rwl_0_31 cell_2r1w
Xcell_2r1w_3646 vdd_uq0 gnd read_bl_0_7 read_bl_1_7 write_bl_0_7 wwl_0_1 rwl_1_1 rwl_0_1
+ cell_2r1w
Xcell_2r1w_2934 vdd_uq3 gnd read_bl_0_18 read_bl_1_18 write_bl_0_18 wwl_0_9 rwl_1_9
+ rwl_0_9 cell_2r1w
Xcell_2r1w_3635 vdd_uq5 gnd read_bl_0_7 read_bl_1_7 write_bl_0_7 wwl_0_12 rwl_1_12
+ rwl_0_12 cell_2r1w
Xcell_2r1w_2923 vdd_uq9 gnd read_bl_0_18 read_bl_1_18 write_bl_0_18 wwl_0_20 rwl_1_20
+ rwl_0_20 cell_2r1w
Xcell_2r1w_3624 vdd_uq10 gnd read_bl_0_7 read_bl_1_7 write_bl_0_7 wwl_0_23 rwl_1_23
+ rwl_0_23 cell_2r1w
Xcell_2r1w_2978 vdd_uq13 gnd read_bl_0_17 read_bl_1_17 write_bl_0_17 wwl_0_29 rwl_1_29
+ rwl_0_29 cell_2r1w
Xcell_2r1w_2989 vdd_uq8 gnd read_bl_0_17 read_bl_1_17 write_bl_0_17 wwl_0_18 rwl_1_18
+ rwl_0_18 cell_2r1w
Xcell_2r1w_16 vdd_uq22 gnd read_bl_0_63 read_bl_1_63 write_bl_0_63 wwl_0_47 rwl_1_47
+ rwl_0_47 cell_2r1w
Xcell_2r1w_27 vdd_uq17 gnd read_bl_0_63 read_bl_1_63 write_bl_0_63 wwl_0_36 rwl_1_36
+ rwl_0_36 cell_2r1w
Xcell_2r1w_38 vdd_uq11 gnd read_bl_0_63 read_bl_1_63 write_bl_0_63 wwl_0_25 rwl_1_25
+ rwl_0_25 cell_2r1w
Xcell_2r1w_49 vdd_uq6 gnd read_bl_0_63 read_bl_1_63 write_bl_0_63 wwl_0_14 rwl_1_14
+ rwl_0_14 cell_2r1w
Xcell_2r1w_2208 vdd_uq14 gnd read_bl_0_29 read_bl_1_29 write_bl_0_29 wwl_0_31 rwl_1_31
+ rwl_0_31 cell_2r1w
Xcell_2r1w_1507 vdd_uq13 gnd read_bl_0_40 read_bl_1_40 write_bl_0_40 wwl_0_28 rwl_1_28
+ rwl_0_28 cell_2r1w
Xcell_2r1w_1518 vdd_uq7 gnd read_bl_0_40 read_bl_1_40 write_bl_0_40 wwl_0_17 rwl_1_17
+ rwl_0_17 cell_2r1w
Xcell_2r1w_2219 vdd_uq9 gnd read_bl_0_29 read_bl_1_29 write_bl_0_29 wwl_0_20 rwl_1_20
+ rwl_0_20 cell_2r1w
Xcell_2r1w_712 vdd_uq26 gnd read_bl_0_52 read_bl_1_52 write_bl_0_52 wwl_0_55 rwl_1_55
+ rwl_0_55 cell_2r1w
Xcell_2r1w_778 vdd_uq25 gnd read_bl_0_51 read_bl_1_51 write_bl_0_51 wwl_0_53 rwl_1_53
+ rwl_0_53 cell_2r1w
Xcell_2r1w_723 vdd_uq21 gnd read_bl_0_52 read_bl_1_52 write_bl_0_52 wwl_0_44 rwl_1_44
+ rwl_0_44 cell_2r1w
Xcell_2r1w_789 vdd_uq20 gnd read_bl_0_51 read_bl_1_51 write_bl_0_51 wwl_0_42 rwl_1_42
+ rwl_0_42 cell_2r1w
Xcell_2r1w_734 vdd_uq15 gnd read_bl_0_52 read_bl_1_52 write_bl_0_52 wwl_0_33 rwl_1_33
+ rwl_0_33 cell_2r1w
Xcell_2r1w_701 vdd gnd read_bl_0_53 read_bl_1_53 write_bl_0_53 wwl_0_2 rwl_1_2 rwl_0_2
+ cell_2r1w
Xcell_2r1w_767 vdd_uq0 gnd read_bl_0_52 read_bl_1_52 write_bl_0_52 wwl_0_0 rwl_1_0
+ rwl_0_0 cell_2r1w
Xcell_2r1w_1529 vdd_uq2 gnd read_bl_0_40 read_bl_1_40 write_bl_0_40 wwl_0_6 rwl_1_6
+ rwl_0_6 cell_2r1w
Xcell_2r1w_756 vdd_uq4 gnd read_bl_0_52 read_bl_1_52 write_bl_0_52 wwl_0_11 rwl_1_11
+ rwl_0_11 cell_2r1w
Xcell_2r1w_745 vdd_uq10 gnd read_bl_0_52 read_bl_1_52 write_bl_0_52 wwl_0_22 rwl_1_22
+ rwl_0_22 cell_2r1w
Xcell_2r1w_6 vdd_uq27 gnd read_bl_0_63 read_bl_1_63 write_bl_0_63 wwl_0_57 rwl_1_57
+ rwl_0_57 cell_2r1w
Xcell_2r1w_3410 vdd_uq21 gnd read_bl_0_10 read_bl_1_10 write_bl_0_10 wwl_0_45 rwl_1_45
+ rwl_0_45 cell_2r1w
Xcell_2r1w_2753 vdd_uq30 gnd read_bl_0_20 read_bl_1_20 write_bl_0_20 wwl_0_62 rwl_1_62
+ rwl_0_62 cell_2r1w
Xcell_2r1w_3465 vdd_uq26 gnd read_bl_0_9 read_bl_1_9 write_bl_0_9 wwl_0_54 rwl_1_54
+ rwl_0_54 cell_2r1w
Xcell_2r1w_2764 vdd_uq24 gnd read_bl_0_20 read_bl_1_20 write_bl_0_20 wwl_0_51 rwl_1_51
+ rwl_0_51 cell_2r1w
Xcell_2r1w_3476 vdd_uq20 gnd read_bl_0_9 read_bl_1_9 write_bl_0_9 wwl_0_43 rwl_1_43
+ rwl_0_43 cell_2r1w
Xcell_2r1w_2775 vdd_uq19 gnd read_bl_0_20 read_bl_1_20 write_bl_0_20 wwl_0_40 rwl_1_40
+ rwl_0_40 cell_2r1w
Xcell_2r1w_3421 vdd_uq16 gnd read_bl_0_10 read_bl_1_10 write_bl_0_10 wwl_0_34 rwl_1_34
+ rwl_0_34 cell_2r1w
Xcell_2r1w_3487 vdd_uq15 gnd read_bl_0_9 read_bl_1_9 write_bl_0_9 wwl_0_32 rwl_1_32
+ rwl_0_32 cell_2r1w
Xcell_2r1w_2720 vdd_uq14 gnd read_bl_0_21 read_bl_1_21 write_bl_0_21 wwl_0_31 rwl_1_31
+ rwl_0_31 cell_2r1w
Xcell_2r1w_2786 vdd_uq13 gnd read_bl_0_20 read_bl_1_20 write_bl_0_20 wwl_0_29 rwl_1_29
+ rwl_0_29 cell_2r1w
Xcell_2r1w_3454 vdd_uq0 gnd read_bl_0_10 read_bl_1_10 write_bl_0_10 wwl_0_1 rwl_1_1
+ rwl_0_1 cell_2r1w
Xcell_2r1w_2742 vdd_uq3 gnd read_bl_0_21 read_bl_1_21 write_bl_0_21 wwl_0_9 rwl_1_9
+ rwl_0_9 cell_2r1w
Xcell_2r1w_3443 vdd_uq5 gnd read_bl_0_10 read_bl_1_10 write_bl_0_10 wwl_0_12 rwl_1_12
+ rwl_0_12 cell_2r1w
Xcell_2r1w_2797 vdd_uq8 gnd read_bl_0_20 read_bl_1_20 write_bl_0_20 wwl_0_18 rwl_1_18
+ rwl_0_18 cell_2r1w
Xcell_2r1w_2731 vdd_uq9 gnd read_bl_0_21 read_bl_1_21 write_bl_0_21 wwl_0_20 rwl_1_20
+ rwl_0_20 cell_2r1w
Xcell_2r1w_3498 vdd_uq9 gnd read_bl_0_9 read_bl_1_9 write_bl_0_9 wwl_0_21 rwl_1_21
+ rwl_0_21 cell_2r1w
Xcell_2r1w_3432 vdd_uq10 gnd read_bl_0_10 read_bl_1_10 write_bl_0_10 wwl_0_23 rwl_1_23
+ rwl_0_23 cell_2r1w
Xcell_2r1w_2049 vdd_uq30 gnd read_bl_0_31 read_bl_1_31 write_bl_0_31 wwl_0_62 rwl_1_62
+ rwl_0_62 cell_2r1w
Xcell_2r1w_1348 vdd_uq28 gnd read_bl_0_42 read_bl_1_42 write_bl_0_42 wwl_0_59 rwl_1_59
+ rwl_0_59 cell_2r1w
Xcell_2r1w_520 vdd_uq26 gnd read_bl_0_55 read_bl_1_55 write_bl_0_55 wwl_0_55 rwl_1_55
+ rwl_0_55 cell_2r1w
Xcell_2r1w_1359 vdd_uq23 gnd read_bl_0_42 read_bl_1_42 write_bl_0_42 wwl_0_48 rwl_1_48
+ rwl_0_48 cell_2r1w
Xcell_2r1w_2005 vdd_uq20 gnd read_bl_0_32 read_bl_1_32 write_bl_0_32 wwl_0_42 rwl_1_42
+ rwl_0_42 cell_2r1w
Xcell_2r1w_1304 vdd_uq18 gnd read_bl_0_43 read_bl_1_43 write_bl_0_43 wwl_0_39 rwl_1_39
+ rwl_0_39 cell_2r1w
Xcell_2r1w_2016 vdd_uq14 gnd read_bl_0_32 read_bl_1_32 write_bl_0_32 wwl_0_31 rwl_1_31
+ rwl_0_31 cell_2r1w
Xcell_2r1w_1315 vdd_uq13 gnd read_bl_0_43 read_bl_1_43 write_bl_0_43 wwl_0_28 rwl_1_28
+ rwl_0_28 cell_2r1w
Xcell_2r1w_1337 vdd_uq2 gnd read_bl_0_43 read_bl_1_43 write_bl_0_43 wwl_0_6 rwl_1_6
+ rwl_0_6 cell_2r1w
Xcell_2r1w_2038 vdd_uq3 gnd read_bl_0_32 read_bl_1_32 write_bl_0_32 wwl_0_9 rwl_1_9
+ rwl_0_9 cell_2r1w
Xcell_2r1w_1326 vdd_uq7 gnd read_bl_0_43 read_bl_1_43 write_bl_0_43 wwl_0_17 rwl_1_17
+ rwl_0_17 cell_2r1w
Xcell_2r1w_2027 vdd_uq9 gnd read_bl_0_32 read_bl_1_32 write_bl_0_32 wwl_0_20 rwl_1_20
+ rwl_0_20 cell_2r1w
Xcell_2r1w_586 vdd_uq25 gnd read_bl_0_54 read_bl_1_54 write_bl_0_54 wwl_0_53 rwl_1_53
+ rwl_0_53 cell_2r1w
Xcell_2r1w_531 vdd_uq21 gnd read_bl_0_55 read_bl_1_55 write_bl_0_55 wwl_0_44 rwl_1_44
+ rwl_0_44 cell_2r1w
Xcell_2r1w_597 vdd_uq20 gnd read_bl_0_54 read_bl_1_54 write_bl_0_54 wwl_0_42 rwl_1_42
+ rwl_0_42 cell_2r1w
Xcell_2r1w_542 vdd_uq15 gnd read_bl_0_55 read_bl_1_55 write_bl_0_55 wwl_0_33 rwl_1_33
+ rwl_0_33 cell_2r1w
Xcell_2r1w_575 vdd_uq0 gnd read_bl_0_55 read_bl_1_55 write_bl_0_55 wwl_0_0 rwl_1_0
+ rwl_0_0 cell_2r1w
Xcell_2r1w_564 vdd_uq4 gnd read_bl_0_55 read_bl_1_55 write_bl_0_55 wwl_0_11 rwl_1_11
+ rwl_0_11 cell_2r1w
Xcell_2r1w_553 vdd_uq10 gnd read_bl_0_55 read_bl_1_55 write_bl_0_55 wwl_0_22 rwl_1_22
+ rwl_0_22 cell_2r1w
Xcell_2r1w_3262 vdd_uq0 gnd read_bl_0_13 read_bl_1_13 write_bl_0_13 wwl_0_1 rwl_1_1
+ rwl_0_1 cell_2r1w
Xcell_2r1w_3251 vdd_uq5 gnd read_bl_0_13 read_bl_1_13 write_bl_0_13 wwl_0_12 rwl_1_12
+ rwl_0_12 cell_2r1w
Xcell_2r1w_3240 vdd_uq10 gnd read_bl_0_13 read_bl_1_13 write_bl_0_13 wwl_0_23 rwl_1_23
+ rwl_0_23 cell_2r1w
Xcell_2r1w_2561 vdd_uq30 gnd read_bl_0_23 read_bl_1_23 write_bl_0_23 wwl_0_62 rwl_1_62
+ rwl_0_62 cell_2r1w
Xcell_2r1w_1860 vdd_uq28 gnd read_bl_0_34 read_bl_1_34 write_bl_0_34 wwl_0_59 rwl_1_59
+ rwl_0_59 cell_2r1w
Xcell_2r1w_3273 vdd_uq26 gnd read_bl_0_12 read_bl_1_12 write_bl_0_12 wwl_0_54 rwl_1_54
+ rwl_0_54 cell_2r1w
Xcell_2r1w_2572 vdd_uq24 gnd read_bl_0_23 read_bl_1_23 write_bl_0_23 wwl_0_51 rwl_1_51
+ rwl_0_51 cell_2r1w
Xcell_2r1w_1871 vdd_uq23 gnd read_bl_0_34 read_bl_1_34 write_bl_0_34 wwl_0_48 rwl_1_48
+ rwl_0_48 cell_2r1w
Xcell_2r1w_3284 vdd_uq20 gnd read_bl_0_12 read_bl_1_12 write_bl_0_12 wwl_0_43 rwl_1_43
+ rwl_0_43 cell_2r1w
Xcell_2r1w_2583 vdd_uq19 gnd read_bl_0_23 read_bl_1_23 write_bl_0_23 wwl_0_40 rwl_1_40
+ rwl_0_40 cell_2r1w
Xcell_2r1w_1882 vdd_uq17 gnd read_bl_0_34 read_bl_1_34 write_bl_0_34 wwl_0_37 rwl_1_37
+ rwl_0_37 cell_2r1w
Xcell_2r1w_3295 vdd_uq15 gnd read_bl_0_12 read_bl_1_12 write_bl_0_12 wwl_0_32 rwl_1_32
+ rwl_0_32 cell_2r1w
Xcell_2r1w_2594 vdd_uq13 gnd read_bl_0_23 read_bl_1_23 write_bl_0_23 wwl_0_29 rwl_1_29
+ rwl_0_29 cell_2r1w
Xcell_2r1w_1893 vdd_uq12 gnd read_bl_0_34 read_bl_1_34 write_bl_0_34 wwl_0_26 rwl_1_26
+ rwl_0_26 cell_2r1w
Xcell_2r1w_2550 vdd_uq3 gnd read_bl_0_24 read_bl_1_24 write_bl_0_24 wwl_0_9 rwl_1_9
+ rwl_0_9 cell_2r1w
Xcell_2r1w_1156 vdd_uq28 gnd read_bl_0_45 read_bl_1_45 write_bl_0_45 wwl_0_59 rwl_1_59
+ rwl_0_59 cell_2r1w
Xcell_2r1w_1101 vdd_uq24 gnd read_bl_0_46 read_bl_1_46 write_bl_0_46 wwl_0_50 rwl_1_50
+ rwl_0_50 cell_2r1w
Xcell_2r1w_1167 vdd_uq23 gnd read_bl_0_45 read_bl_1_45 write_bl_0_45 wwl_0_48 rwl_1_48
+ rwl_0_48 cell_2r1w
Xcell_2r1w_1112 vdd_uq18 gnd read_bl_0_46 read_bl_1_46 write_bl_0_46 wwl_0_39 rwl_1_39
+ rwl_0_39 cell_2r1w
Xcell_2r1w_1178 vdd_uq17 gnd read_bl_0_45 read_bl_1_45 write_bl_0_45 wwl_0_37 rwl_1_37
+ rwl_0_37 cell_2r1w
Xcell_2r1w_350 vdd_uq15 gnd read_bl_0_58 read_bl_1_58 write_bl_0_58 wwl_0_33 rwl_1_33
+ rwl_0_33 cell_2r1w
Xcell_2r1w_1123 vdd_uq13 gnd read_bl_0_46 read_bl_1_46 write_bl_0_46 wwl_0_28 rwl_1_28
+ rwl_0_28 cell_2r1w
Xcell_2r1w_1189 vdd_uq12 gnd read_bl_0_45 read_bl_1_45 write_bl_0_45 wwl_0_26 rwl_1_26
+ rwl_0_26 cell_2r1w
Xcell_2r1w_1145 vdd_uq2 gnd read_bl_0_46 read_bl_1_46 write_bl_0_46 wwl_0_6 rwl_1_6
+ rwl_0_6 cell_2r1w
Xcell_2r1w_372 vdd_uq4 gnd read_bl_0_58 read_bl_1_58 write_bl_0_58 wwl_0_11 rwl_1_11
+ rwl_0_11 cell_2r1w
Xcell_2r1w_1134 vdd_uq7 gnd read_bl_0_46 read_bl_1_46 write_bl_0_46 wwl_0_17 rwl_1_17
+ rwl_0_17 cell_2r1w
Xcell_2r1w_361 vdd_uq10 gnd read_bl_0_58 read_bl_1_58 write_bl_0_58 wwl_0_22 rwl_1_22
+ rwl_0_22 cell_2r1w
Xcell_2r1w_394 vdd_uq25 gnd read_bl_0_57 read_bl_1_57 write_bl_0_57 wwl_0_53 rwl_1_53
+ rwl_0_53 cell_2r1w
Xcell_2r1w_383 vdd_uq0 gnd read_bl_0_58 read_bl_1_58 write_bl_0_58 wwl_0_0 rwl_1_0
+ rwl_0_0 cell_2r1w
Xcell_2r1w_3081 vdd_uq26 gnd read_bl_0_15 read_bl_1_15 write_bl_0_15 wwl_0_54 rwl_1_54
+ rwl_0_54 cell_2r1w
Xcell_2r1w_3092 vdd_uq20 gnd read_bl_0_15 read_bl_1_15 write_bl_0_15 wwl_0_43 rwl_1_43
+ rwl_0_43 cell_2r1w
Xcell_2r1w_3070 vdd_uq0 gnd read_bl_0_16 read_bl_1_16 write_bl_0_16 wwl_0_1 rwl_1_1
+ rwl_0_1 cell_2r1w
Xcell_2r1w_2380 vdd_uq24 gnd read_bl_0_26 read_bl_1_26 write_bl_0_26 wwl_0_51 rwl_1_51
+ rwl_0_51 cell_2r1w
Xcell_2r1w_2391 vdd_uq19 gnd read_bl_0_26 read_bl_1_26 write_bl_0_26 wwl_0_40 rwl_1_40
+ rwl_0_40 cell_2r1w
Xcell_2r1w_1690 vdd_uq17 gnd read_bl_0_37 read_bl_1_37 write_bl_0_37 wwl_0_37 rwl_1_37
+ rwl_0_37 cell_2r1w
Xcell_2r1w_191 vdd_uq0 gnd read_bl_0_61 read_bl_1_61 write_bl_0_61 wwl_0_0 rwl_1_0
+ rwl_0_0 cell_2r1w
Xcell_2r1w_180 vdd_uq4 gnd read_bl_0_61 read_bl_1_61 write_bl_0_61 wwl_0_11 rwl_1_11
+ rwl_0_11 cell_2r1w
Xcell_2r1w_3806 vdd_uq15 gnd read_bl_0_4 read_bl_1_4 write_bl_0_4 wwl_0_33 rwl_1_33
+ rwl_0_33 cell_2r1w
Xcell_2r1w_3839 vdd_uq0 gnd read_bl_0_4 read_bl_1_4 write_bl_0_4 wwl_0_0 rwl_1_0 rwl_0_0
+ cell_2r1w
Xcell_2r1w_3828 vdd_uq4 gnd read_bl_0_4 read_bl_1_4 write_bl_0_4 wwl_0_11 rwl_1_11
+ rwl_0_11 cell_2r1w
Xcell_2r1w_3817 vdd_uq10 gnd read_bl_0_4 read_bl_1_4 write_bl_0_4 wwl_0_22 rwl_1_22
+ rwl_0_22 cell_2r1w
Xcell_2r1w_905 vdd_uq26 gnd read_bl_0_49 read_bl_1_49 write_bl_0_49 wwl_0_54 rwl_1_54
+ rwl_0_54 cell_2r1w
Xcell_2r1w_916 vdd_uq20 gnd read_bl_0_49 read_bl_1_49 write_bl_0_49 wwl_0_43 rwl_1_43
+ rwl_0_43 cell_2r1w
Xcell_2r1w_927 vdd_uq15 gnd read_bl_0_49 read_bl_1_49 write_bl_0_49 wwl_0_32 rwl_1_32
+ rwl_0_32 cell_2r1w
Xcell_2r1w_949 vdd_uq4 gnd read_bl_0_49 read_bl_1_49 write_bl_0_49 wwl_0_10 rwl_1_10
+ rwl_0_10 cell_2r1w
Xcell_2r1w_938 vdd_uq9 gnd read_bl_0_49 read_bl_1_49 write_bl_0_49 wwl_0_21 rwl_1_21
+ rwl_0_21 cell_2r1w
Xcell_2r1w_2946 vdd_uq29 gnd read_bl_0_17 read_bl_1_17 write_bl_0_17 wwl_0_61 rwl_1_61
+ rwl_0_61 cell_2r1w
Xcell_2r1w_3658 vdd_uq25 gnd read_bl_0_6 read_bl_1_6 write_bl_0_6 wwl_0_53 rwl_1_53
+ rwl_0_53 cell_2r1w
Xcell_2r1w_2957 vdd_uq24 gnd read_bl_0_17 read_bl_1_17 write_bl_0_17 wwl_0_50 rwl_1_50
+ rwl_0_50 cell_2r1w
Xcell_2r1w_3603 vdd_uq21 gnd read_bl_0_7 read_bl_1_7 write_bl_0_7 wwl_0_44 rwl_1_44
+ rwl_0_44 cell_2r1w
Xcell_2r1w_2902 vdd_uq19 gnd read_bl_0_18 read_bl_1_18 write_bl_0_18 wwl_0_41 rwl_1_41
+ rwl_0_41 cell_2r1w
Xcell_2r1w_3669 vdd_uq20 gnd read_bl_0_6 read_bl_1_6 write_bl_0_6 wwl_0_42 rwl_1_42
+ rwl_0_42 cell_2r1w
Xcell_2r1w_2968 vdd_uq18 gnd read_bl_0_17 read_bl_1_17 write_bl_0_17 wwl_0_39 rwl_1_39
+ rwl_0_39 cell_2r1w
Xcell_2r1w_3614 vdd_uq15 gnd read_bl_0_7 read_bl_1_7 write_bl_0_7 wwl_0_33 rwl_1_33
+ rwl_0_33 cell_2r1w
Xcell_2r1w_2913 vdd_uq14 gnd read_bl_0_18 read_bl_1_18 write_bl_0_18 wwl_0_30 rwl_1_30
+ rwl_0_30 cell_2r1w
Xcell_2r1w_2979 vdd_uq13 gnd read_bl_0_17 read_bl_1_17 write_bl_0_17 wwl_0_28 rwl_1_28
+ rwl_0_28 cell_2r1w
Xcell_2r1w_3647 vdd_uq0 gnd read_bl_0_7 read_bl_1_7 write_bl_0_7 wwl_0_0 rwl_1_0 rwl_0_0
+ cell_2r1w
Xcell_2r1w_2935 vdd_uq3 gnd read_bl_0_18 read_bl_1_18 write_bl_0_18 wwl_0_8 rwl_1_8
+ rwl_0_8 cell_2r1w
Xcell_2r1w_3636 vdd_uq4 gnd read_bl_0_7 read_bl_1_7 write_bl_0_7 wwl_0_11 rwl_1_11
+ rwl_0_11 cell_2r1w
Xcell_2r1w_2924 vdd_uq8 gnd read_bl_0_18 read_bl_1_18 write_bl_0_18 wwl_0_19 rwl_1_19
+ rwl_0_19 cell_2r1w
Xcell_2r1w_3625 vdd_uq10 gnd read_bl_0_7 read_bl_1_7 write_bl_0_7 wwl_0_22 rwl_1_22
+ rwl_0_22 cell_2r1w
Xcell_2r1w_17 vdd_uq22 gnd read_bl_0_63 read_bl_1_63 write_bl_0_63 wwl_0_46 rwl_1_46
+ rwl_0_46 cell_2r1w
Xcell_2r1w_28 vdd_uq16 gnd read_bl_0_63 read_bl_1_63 write_bl_0_63 wwl_0_35 rwl_1_35
+ rwl_0_35 cell_2r1w
Xcell_2r1w_39 vdd_uq11 gnd read_bl_0_63 read_bl_1_63 write_bl_0_63 wwl_0_24 rwl_1_24
+ rwl_0_24 cell_2r1w
Xcell_2r1w_2209 vdd_uq14 gnd read_bl_0_29 read_bl_1_29 write_bl_0_29 wwl_0_30 rwl_1_30
+ rwl_0_30 cell_2r1w
Xcell_2r1w_1508 vdd_uq12 gnd read_bl_0_40 read_bl_1_40 write_bl_0_40 wwl_0_27 rwl_1_27
+ rwl_0_27 cell_2r1w
Xcell_2r1w_702 vdd_uq0 gnd read_bl_0_53 read_bl_1_53 write_bl_0_53 wwl_0_1 rwl_1_1
+ rwl_0_1 cell_2r1w
Xcell_2r1w_1519 vdd_uq7 gnd read_bl_0_40 read_bl_1_40 write_bl_0_40 wwl_0_16 rwl_1_16
+ rwl_0_16 cell_2r1w
Xcell_2r1w_768 vdd_uq30 gnd read_bl_0_51 read_bl_1_51 write_bl_0_51 wwl_0_63 rwl_1_63
+ rwl_0_63 cell_2r1w
Xcell_2r1w_713 vdd_uq26 gnd read_bl_0_52 read_bl_1_52 write_bl_0_52 wwl_0_54 rwl_1_54
+ rwl_0_54 cell_2r1w
Xcell_2r1w_779 vdd_uq25 gnd read_bl_0_51 read_bl_1_51 write_bl_0_51 wwl_0_52 rwl_1_52
+ rwl_0_52 cell_2r1w
Xcell_2r1w_724 vdd_uq20 gnd read_bl_0_52 read_bl_1_52 write_bl_0_52 wwl_0_43 rwl_1_43
+ rwl_0_43 cell_2r1w
Xcell_2r1w_735 vdd_uq15 gnd read_bl_0_52 read_bl_1_52 write_bl_0_52 wwl_0_32 rwl_1_32
+ rwl_0_32 cell_2r1w
Xcell_2r1w_757 vdd_uq4 gnd read_bl_0_52 read_bl_1_52 write_bl_0_52 wwl_0_10 rwl_1_10
+ rwl_0_10 cell_2r1w
Xcell_2r1w_746 vdd_uq9 gnd read_bl_0_52 read_bl_1_52 write_bl_0_52 wwl_0_21 rwl_1_21
+ rwl_0_21 cell_2r1w
Xcell_2r1w_7 vdd_uq27 gnd read_bl_0_63 read_bl_1_63 write_bl_0_63 wwl_0_56 rwl_1_56
+ rwl_0_56 cell_2r1w
Xcell_2r1w_3400 vdd_uq26 gnd read_bl_0_10 read_bl_1_10 write_bl_0_10 wwl_0_55 rwl_1_55
+ rwl_0_55 cell_2r1w
Xcell_2r1w_3411 vdd_uq21 gnd read_bl_0_10 read_bl_1_10 write_bl_0_10 wwl_0_44 rwl_1_44
+ rwl_0_44 cell_2r1w
Xcell_2r1w_3422 vdd_uq15 gnd read_bl_0_10 read_bl_1_10 write_bl_0_10 wwl_0_33 rwl_1_33
+ rwl_0_33 cell_2r1w
Xcell_2r1w_3444 vdd_uq4 gnd read_bl_0_10 read_bl_1_10 write_bl_0_10 wwl_0_11 rwl_1_11
+ rwl_0_11 cell_2r1w
Xcell_2r1w_3433 vdd_uq10 gnd read_bl_0_10 read_bl_1_10 write_bl_0_10 wwl_0_22 rwl_1_22
+ rwl_0_22 cell_2r1w
Xcell_2r1w_2754 vdd_uq29 gnd read_bl_0_20 read_bl_1_20 write_bl_0_20 wwl_0_61 rwl_1_61
+ rwl_0_61 cell_2r1w
Xcell_2r1w_3466 vdd_uq25 gnd read_bl_0_9 read_bl_1_9 write_bl_0_9 wwl_0_53 rwl_1_53
+ rwl_0_53 cell_2r1w
Xcell_2r1w_2765 vdd_uq24 gnd read_bl_0_20 read_bl_1_20 write_bl_0_20 wwl_0_50 rwl_1_50
+ rwl_0_50 cell_2r1w
Xcell_2r1w_2710 vdd_uq19 gnd read_bl_0_21 read_bl_1_21 write_bl_0_21 wwl_0_41 rwl_1_41
+ rwl_0_41 cell_2r1w
Xcell_2r1w_3477 vdd_uq20 gnd read_bl_0_9 read_bl_1_9 write_bl_0_9 wwl_0_42 rwl_1_42
+ rwl_0_42 cell_2r1w
Xcell_2r1w_2776 vdd_uq18 gnd read_bl_0_20 read_bl_1_20 write_bl_0_20 wwl_0_39 rwl_1_39
+ rwl_0_39 cell_2r1w
Xcell_2r1w_3488 vdd_uq14 gnd read_bl_0_9 read_bl_1_9 write_bl_0_9 wwl_0_31 rwl_1_31
+ rwl_0_31 cell_2r1w
Xcell_2r1w_2721 vdd_uq14 gnd read_bl_0_21 read_bl_1_21 write_bl_0_21 wwl_0_30 rwl_1_30
+ rwl_0_30 cell_2r1w
Xcell_2r1w_2787 vdd_uq13 gnd read_bl_0_20 read_bl_1_20 write_bl_0_20 wwl_0_28 rwl_1_28
+ rwl_0_28 cell_2r1w
Xcell_2r1w_3455 vdd_uq0 gnd read_bl_0_10 read_bl_1_10 write_bl_0_10 wwl_0_0 rwl_1_0
+ rwl_0_0 cell_2r1w
Xcell_2r1w_2743 vdd_uq3 gnd read_bl_0_21 read_bl_1_21 write_bl_0_21 wwl_0_8 rwl_1_8
+ rwl_0_8 cell_2r1w
Xcell_2r1w_2798 vdd_uq7 gnd read_bl_0_20 read_bl_1_20 write_bl_0_20 wwl_0_17 rwl_1_17
+ rwl_0_17 cell_2r1w
Xcell_2r1w_2732 vdd_uq8 gnd read_bl_0_21 read_bl_1_21 write_bl_0_21 wwl_0_19 rwl_1_19
+ rwl_0_19 cell_2r1w
Xcell_2r1w_3499 vdd_uq9 gnd read_bl_0_9 read_bl_1_9 write_bl_0_9 wwl_0_20 rwl_1_20
+ rwl_0_20 cell_2r1w
Xcell_2r1w_1349 vdd_uq28 gnd read_bl_0_42 read_bl_1_42 write_bl_0_42 wwl_0_58 rwl_1_58
+ rwl_0_58 cell_2r1w
Xcell_2r1w_521 vdd_uq26 gnd read_bl_0_55 read_bl_1_55 write_bl_0_55 wwl_0_54 rwl_1_54
+ rwl_0_54 cell_2r1w
Xcell_2r1w_532 vdd_uq20 gnd read_bl_0_55 read_bl_1_55 write_bl_0_55 wwl_0_43 rwl_1_43
+ rwl_0_43 cell_2r1w
Xcell_2r1w_2006 vdd_uq19 gnd read_bl_0_32 read_bl_1_32 write_bl_0_32 wwl_0_41 rwl_1_41
+ rwl_0_41 cell_2r1w
Xcell_2r1w_1305 vdd_uq18 gnd read_bl_0_43 read_bl_1_43 write_bl_0_43 wwl_0_38 rwl_1_38
+ rwl_0_38 cell_2r1w
Xcell_2r1w_543 vdd_uq15 gnd read_bl_0_55 read_bl_1_55 write_bl_0_55 wwl_0_32 rwl_1_32
+ rwl_0_32 cell_2r1w
Xcell_2r1w_2017 vdd_uq14 gnd read_bl_0_32 read_bl_1_32 write_bl_0_32 wwl_0_30 rwl_1_30
+ rwl_0_30 cell_2r1w
Xcell_2r1w_1316 vdd_uq12 gnd read_bl_0_43 read_bl_1_43 write_bl_0_43 wwl_0_27 rwl_1_27
+ rwl_0_27 cell_2r1w
Xcell_2r1w_1338 vdd_uq1 gnd read_bl_0_43 read_bl_1_43 write_bl_0_43 wwl_0_5 rwl_1_5
+ rwl_0_5 cell_2r1w
Xcell_2r1w_510 vdd_uq0 gnd read_bl_0_56 read_bl_1_56 write_bl_0_56 wwl_0_1 rwl_1_1
+ rwl_0_1 cell_2r1w
Xcell_2r1w_2039 vdd_uq3 gnd read_bl_0_32 read_bl_1_32 write_bl_0_32 wwl_0_8 rwl_1_8
+ rwl_0_8 cell_2r1w
Xcell_2r1w_1327 vdd_uq7 gnd read_bl_0_43 read_bl_1_43 write_bl_0_43 wwl_0_16 rwl_1_16
+ rwl_0_16 cell_2r1w
Xcell_2r1w_2028 vdd_uq8 gnd read_bl_0_32 read_bl_1_32 write_bl_0_32 wwl_0_19 rwl_1_19
+ rwl_0_19 cell_2r1w
Xcell_2r1w_554 vdd_uq9 gnd read_bl_0_55 read_bl_1_55 write_bl_0_55 wwl_0_21 rwl_1_21
+ rwl_0_21 cell_2r1w
Xcell_2r1w_576 vdd_uq30 gnd read_bl_0_54 read_bl_1_54 write_bl_0_54 wwl_0_63 rwl_1_63
+ rwl_0_63 cell_2r1w
Xcell_2r1w_587 vdd_uq25 gnd read_bl_0_54 read_bl_1_54 write_bl_0_54 wwl_0_52 rwl_1_52
+ rwl_0_52 cell_2r1w
Xcell_2r1w_598 vdd_uq19 gnd read_bl_0_54 read_bl_1_54 write_bl_0_54 wwl_0_41 rwl_1_41
+ rwl_0_41 cell_2r1w
Xcell_2r1w_565 vdd_uq4 gnd read_bl_0_55 read_bl_1_55 write_bl_0_55 wwl_0_10 rwl_1_10
+ rwl_0_10 cell_2r1w
Xcell_2r1w_3274 vdd_uq25 gnd read_bl_0_12 read_bl_1_12 write_bl_0_12 wwl_0_53 rwl_1_53
+ rwl_0_53 cell_2r1w
Xcell_2r1w_3285 vdd_uq20 gnd read_bl_0_12 read_bl_1_12 write_bl_0_12 wwl_0_42 rwl_1_42
+ rwl_0_42 cell_2r1w
Xcell_2r1w_3230 vdd_uq15 gnd read_bl_0_13 read_bl_1_13 write_bl_0_13 wwl_0_33 rwl_1_33
+ rwl_0_33 cell_2r1w
Xcell_2r1w_3263 vdd_uq0 gnd read_bl_0_13 read_bl_1_13 write_bl_0_13 wwl_0_0 rwl_1_0
+ rwl_0_0 cell_2r1w
Xcell_2r1w_2551 vdd_uq3 gnd read_bl_0_24 read_bl_1_24 write_bl_0_24 wwl_0_8 rwl_1_8
+ rwl_0_8 cell_2r1w
Xcell_2r1w_3252 vdd_uq4 gnd read_bl_0_13 read_bl_1_13 write_bl_0_13 wwl_0_11 rwl_1_11
+ rwl_0_11 cell_2r1w
Xcell_2r1w_2540 vdd_uq8 gnd read_bl_0_24 read_bl_1_24 write_bl_0_24 wwl_0_19 rwl_1_19
+ rwl_0_19 cell_2r1w
Xcell_2r1w_3241 vdd_uq10 gnd read_bl_0_13 read_bl_1_13 write_bl_0_13 wwl_0_22 rwl_1_22
+ rwl_0_22 cell_2r1w
Xcell_2r1w_2562 vdd_uq29 gnd read_bl_0_23 read_bl_1_23 write_bl_0_23 wwl_0_61 rwl_1_61
+ rwl_0_61 cell_2r1w
Xcell_2r1w_1861 vdd_uq28 gnd read_bl_0_34 read_bl_1_34 write_bl_0_34 wwl_0_58 rwl_1_58
+ rwl_0_58 cell_2r1w
Xcell_2r1w_2573 vdd_uq24 gnd read_bl_0_23 read_bl_1_23 write_bl_0_23 wwl_0_50 rwl_1_50
+ rwl_0_50 cell_2r1w
Xcell_2r1w_1872 vdd_uq22 gnd read_bl_0_34 read_bl_1_34 write_bl_0_34 wwl_0_47 rwl_1_47
+ rwl_0_47 cell_2r1w
Xcell_2r1w_2584 vdd_uq18 gnd read_bl_0_23 read_bl_1_23 write_bl_0_23 wwl_0_39 rwl_1_39
+ rwl_0_39 cell_2r1w
Xcell_2r1w_1883 vdd_uq17 gnd read_bl_0_34 read_bl_1_34 write_bl_0_34 wwl_0_36 rwl_1_36
+ rwl_0_36 cell_2r1w
Xcell_2r1w_3296 vdd_uq14 gnd read_bl_0_12 read_bl_1_12 write_bl_0_12 wwl_0_31 rwl_1_31
+ rwl_0_31 cell_2r1w
Xcell_2r1w_2595 vdd_uq13 gnd read_bl_0_23 read_bl_1_23 write_bl_0_23 wwl_0_28 rwl_1_28
+ rwl_0_28 cell_2r1w
Xcell_2r1w_1894 vdd_uq11 gnd read_bl_0_34 read_bl_1_34 write_bl_0_34 wwl_0_25 rwl_1_25
+ rwl_0_25 cell_2r1w
Xcell_2r1w_1850 vdd_uq1 gnd read_bl_0_35 read_bl_1_35 write_bl_0_35 wwl_0_5 rwl_1_5
+ rwl_0_5 cell_2r1w
Xcell_2r1w_384 vdd_uq30 gnd read_bl_0_57 read_bl_1_57 write_bl_0_57 wwl_0_63 rwl_1_63
+ rwl_0_63 cell_2r1w
Xcell_2r1w_1157 vdd_uq28 gnd read_bl_0_45 read_bl_1_45 write_bl_0_45 wwl_0_58 rwl_1_58
+ rwl_0_58 cell_2r1w
Xcell_2r1w_395 vdd_uq25 gnd read_bl_0_57 read_bl_1_57 write_bl_0_57 wwl_0_52 rwl_1_52
+ rwl_0_52 cell_2r1w
Xcell_2r1w_1102 vdd_uq23 gnd read_bl_0_46 read_bl_1_46 write_bl_0_46 wwl_0_49 rwl_1_49
+ rwl_0_49 cell_2r1w
Xcell_2r1w_1168 vdd_uq22 gnd read_bl_0_45 read_bl_1_45 write_bl_0_45 wwl_0_47 rwl_1_47
+ rwl_0_47 cell_2r1w
Xcell_2r1w_340 vdd_uq20 gnd read_bl_0_58 read_bl_1_58 write_bl_0_58 wwl_0_43 rwl_1_43
+ rwl_0_43 cell_2r1w
Xcell_2r1w_1113 vdd_uq18 gnd read_bl_0_46 read_bl_1_46 write_bl_0_46 wwl_0_38 rwl_1_38
+ rwl_0_38 cell_2r1w
Xcell_2r1w_1179 vdd_uq17 gnd read_bl_0_45 read_bl_1_45 write_bl_0_45 wwl_0_36 rwl_1_36
+ rwl_0_36 cell_2r1w
Xcell_2r1w_351 vdd_uq15 gnd read_bl_0_58 read_bl_1_58 write_bl_0_58 wwl_0_32 rwl_1_32
+ rwl_0_32 cell_2r1w
Xcell_2r1w_1124 vdd_uq12 gnd read_bl_0_46 read_bl_1_46 write_bl_0_46 wwl_0_27 rwl_1_27
+ rwl_0_27 cell_2r1w
Xcell_2r1w_1146 vdd_uq1 gnd read_bl_0_46 read_bl_1_46 write_bl_0_46 wwl_0_5 rwl_1_5
+ rwl_0_5 cell_2r1w
Xcell_2r1w_373 vdd_uq4 gnd read_bl_0_58 read_bl_1_58 write_bl_0_58 wwl_0_10 rwl_1_10
+ rwl_0_10 cell_2r1w
Xcell_2r1w_1135 vdd_uq7 gnd read_bl_0_46 read_bl_1_46 write_bl_0_46 wwl_0_16 rwl_1_16
+ rwl_0_16 cell_2r1w
Xcell_2r1w_362 vdd_uq9 gnd read_bl_0_58 read_bl_1_58 write_bl_0_58 wwl_0_21 rwl_1_21
+ rwl_0_21 cell_2r1w
Xcell_2r1w_2370 vdd_uq29 gnd read_bl_0_26 read_bl_1_26 write_bl_0_26 wwl_0_61 rwl_1_61
+ rwl_0_61 cell_2r1w
Xcell_2r1w_3082 vdd_uq25 gnd read_bl_0_15 read_bl_1_15 write_bl_0_15 wwl_0_53 rwl_1_53
+ rwl_0_53 cell_2r1w
Xcell_2r1w_2381 vdd_uq24 gnd read_bl_0_26 read_bl_1_26 write_bl_0_26 wwl_0_50 rwl_1_50
+ rwl_0_50 cell_2r1w
Xcell_2r1w_3093 vdd_uq20 gnd read_bl_0_15 read_bl_1_15 write_bl_0_15 wwl_0_42 rwl_1_42
+ rwl_0_42 cell_2r1w
Xcell_2r1w_2392 vdd_uq18 gnd read_bl_0_26 read_bl_1_26 write_bl_0_26 wwl_0_39 rwl_1_39
+ rwl_0_39 cell_2r1w
Xcell_2r1w_3071 vdd_uq0 gnd read_bl_0_16 read_bl_1_16 write_bl_0_16 wwl_0_0 rwl_1_0
+ rwl_0_0 cell_2r1w
Xcell_2r1w_3060 vdd_uq4 gnd read_bl_0_16 read_bl_1_16 write_bl_0_16 wwl_0_11 rwl_1_11
+ rwl_0_11 cell_2r1w
Xcell_2r1w_1680 vdd_uq22 gnd read_bl_0_37 read_bl_1_37 write_bl_0_37 wwl_0_47 rwl_1_47
+ rwl_0_47 cell_2r1w
Xcell_2r1w_1691 vdd_uq17 gnd read_bl_0_37 read_bl_1_37 write_bl_0_37 wwl_0_36 rwl_1_36
+ rwl_0_36 cell_2r1w
Xcell_2r1w_192 vdd_uq30 gnd read_bl_0_60 read_bl_1_60 write_bl_0_60 wwl_0_63 rwl_1_63
+ rwl_0_63 cell_2r1w
Xcell_2r1w_181 vdd_uq4 gnd read_bl_0_61 read_bl_1_61 write_bl_0_61 wwl_0_10 rwl_1_10
+ rwl_0_10 cell_2r1w
Xcell_2r1w_170 vdd_uq9 gnd read_bl_0_61 read_bl_1_61 write_bl_0_61 wwl_0_21 rwl_1_21
+ rwl_0_21 cell_2r1w
Xcell_2r1w_3807 vdd_uq15 gnd read_bl_0_4 read_bl_1_4 write_bl_0_4 wwl_0_32 rwl_1_32
+ rwl_0_32 cell_2r1w
Xcell_2r1w_3829 vdd_uq4 gnd read_bl_0_4 read_bl_1_4 write_bl_0_4 wwl_0_10 rwl_1_10
+ rwl_0_10 cell_2r1w
Xcell_2r1w_3818 vdd_uq9 gnd read_bl_0_4 read_bl_1_4 write_bl_0_4 wwl_0_21 rwl_1_21
+ rwl_0_21 cell_2r1w
Xcell_2r1w_906 vdd_uq25 gnd read_bl_0_49 read_bl_1_49 write_bl_0_49 wwl_0_53 rwl_1_53
+ rwl_0_53 cell_2r1w
Xcell_2r1w_917 vdd_uq20 gnd read_bl_0_49 read_bl_1_49 write_bl_0_49 wwl_0_42 rwl_1_42
+ rwl_0_42 cell_2r1w
Xcell_2r1w_928 vdd_uq14 gnd read_bl_0_49 read_bl_1_49 write_bl_0_49 wwl_0_31 rwl_1_31
+ rwl_0_31 cell_2r1w
Xcell_2r1w_939 vdd_uq9 gnd read_bl_0_49 read_bl_1_49 write_bl_0_49 wwl_0_20 rwl_1_20
+ rwl_0_20 cell_2r1w
Xcell_2r1w_3604 vdd_uq20 gnd read_bl_0_7 read_bl_1_7 write_bl_0_7 wwl_0_43 rwl_1_43
+ rwl_0_43 cell_2r1w
Xcell_2r1w_3615 vdd_uq15 gnd read_bl_0_7 read_bl_1_7 write_bl_0_7 wwl_0_32 rwl_1_32
+ rwl_0_32 cell_2r1w
Xcell_2r1w_3626 vdd_uq9 gnd read_bl_0_7 read_bl_1_7 write_bl_0_7 wwl_0_21 rwl_1_21
+ rwl_0_21 cell_2r1w
Xcell_2r1w_3648 vdd_uq30 gnd read_bl_0_6 read_bl_1_6 write_bl_0_6 wwl_0_63 rwl_1_63
+ rwl_0_63 cell_2r1w
Xcell_2r1w_2947 vdd_uq29 gnd read_bl_0_17 read_bl_1_17 write_bl_0_17 wwl_0_60 rwl_1_60
+ rwl_0_60 cell_2r1w
Xcell_2r1w_3659 vdd_uq25 gnd read_bl_0_6 read_bl_1_6 write_bl_0_6 wwl_0_52 rwl_1_52
+ rwl_0_52 cell_2r1w
Xcell_2r1w_2958 vdd_uq23 gnd read_bl_0_17 read_bl_1_17 write_bl_0_17 wwl_0_49 rwl_1_49
+ rwl_0_49 cell_2r1w
Xcell_2r1w_2903 vdd_uq19 gnd read_bl_0_18 read_bl_1_18 write_bl_0_18 wwl_0_40 rwl_1_40
+ rwl_0_40 cell_2r1w
Xcell_2r1w_2969 vdd_uq18 gnd read_bl_0_17 read_bl_1_17 write_bl_0_17 wwl_0_38 rwl_1_38
+ rwl_0_38 cell_2r1w
Xcell_2r1w_2914 vdd_uq13 gnd read_bl_0_18 read_bl_1_18 write_bl_0_18 wwl_0_29 rwl_1_29
+ rwl_0_29 cell_2r1w
Xcell_2r1w_2936 vdd_uq2 gnd read_bl_0_18 read_bl_1_18 write_bl_0_18 wwl_0_7 rwl_1_7
+ rwl_0_7 cell_2r1w
Xcell_2r1w_3637 vdd_uq4 gnd read_bl_0_7 read_bl_1_7 write_bl_0_7 wwl_0_10 rwl_1_10
+ rwl_0_10 cell_2r1w
Xcell_2r1w_2925 vdd_uq8 gnd read_bl_0_18 read_bl_1_18 write_bl_0_18 wwl_0_18 rwl_1_18
+ rwl_0_18 cell_2r1w
Xcell_2r1w_18 vdd_uq21 gnd read_bl_0_63 read_bl_1_63 write_bl_0_63 wwl_0_45 rwl_1_45
+ rwl_0_45 cell_2r1w
Xcell_2r1w_29 vdd_uq16 gnd read_bl_0_63 read_bl_1_63 write_bl_0_63 wwl_0_34 rwl_1_34
+ rwl_0_34 cell_2r1w
Xcell_2r1w_714 vdd_uq25 gnd read_bl_0_52 read_bl_1_52 write_bl_0_52 wwl_0_53 rwl_1_53
+ rwl_0_53 cell_2r1w
Xcell_2r1w_725 vdd_uq20 gnd read_bl_0_52 read_bl_1_52 write_bl_0_52 wwl_0_42 rwl_1_42
+ rwl_0_42 cell_2r1w
Xcell_2r1w_736 vdd_uq14 gnd read_bl_0_52 read_bl_1_52 write_bl_0_52 wwl_0_31 rwl_1_31
+ rwl_0_31 cell_2r1w
Xcell_2r1w_1509 vdd_uq12 gnd read_bl_0_40 read_bl_1_40 write_bl_0_40 wwl_0_26 rwl_1_26
+ rwl_0_26 cell_2r1w
Xcell_2r1w_703 vdd_uq0 gnd read_bl_0_53 read_bl_1_53 write_bl_0_53 wwl_0_0 rwl_1_0
+ rwl_0_0 cell_2r1w
Xcell_2r1w_769 vdd_uq30 gnd read_bl_0_51 read_bl_1_51 write_bl_0_51 wwl_0_62 rwl_1_62
+ rwl_0_62 cell_2r1w
Xcell_2r1w_758 vdd_uq3 gnd read_bl_0_52 read_bl_1_52 write_bl_0_52 wwl_0_9 rwl_1_9
+ rwl_0_9 cell_2r1w
Xcell_2r1w_747 vdd_uq9 gnd read_bl_0_52 read_bl_1_52 write_bl_0_52 wwl_0_20 rwl_1_20
+ rwl_0_20 cell_2r1w
Xcell_2r1w_8 vdd_uq26 gnd read_bl_0_63 read_bl_1_63 write_bl_0_63 wwl_0_55 rwl_1_55
+ rwl_0_55 cell_2r1w
Xcell_2r1w_3456 vdd_uq30 gnd read_bl_0_9 read_bl_1_9 write_bl_0_9 wwl_0_63 rwl_1_63
+ rwl_0_63 cell_2r1w
Xcell_2r1w_3401 vdd_uq26 gnd read_bl_0_10 read_bl_1_10 write_bl_0_10 wwl_0_54 rwl_1_54
+ rwl_0_54 cell_2r1w
Xcell_2r1w_3467 vdd_uq25 gnd read_bl_0_9 read_bl_1_9 write_bl_0_9 wwl_0_52 rwl_1_52
+ rwl_0_52 cell_2r1w
Xcell_2r1w_2700 vdd_uq24 gnd read_bl_0_21 read_bl_1_21 write_bl_0_21 wwl_0_51 rwl_1_51
+ rwl_0_51 cell_2r1w
Xcell_2r1w_3412 vdd_uq20 gnd read_bl_0_10 read_bl_1_10 write_bl_0_10 wwl_0_43 rwl_1_43
+ rwl_0_43 cell_2r1w
Xcell_2r1w_3478 vdd_uq19 gnd read_bl_0_9 read_bl_1_9 write_bl_0_9 wwl_0_41 rwl_1_41
+ rwl_0_41 cell_2r1w
Xcell_2r1w_2711 vdd_uq19 gnd read_bl_0_21 read_bl_1_21 write_bl_0_21 wwl_0_40 rwl_1_40
+ rwl_0_40 cell_2r1w
Xcell_2r1w_3423 vdd_uq15 gnd read_bl_0_10 read_bl_1_10 write_bl_0_10 wwl_0_32 rwl_1_32
+ rwl_0_32 cell_2r1w
Xcell_2r1w_2722 vdd_uq13 gnd read_bl_0_21 read_bl_1_21 write_bl_0_21 wwl_0_29 rwl_1_29
+ rwl_0_29 cell_2r1w
Xcell_2r1w_3445 vdd_uq4 gnd read_bl_0_10 read_bl_1_10 write_bl_0_10 wwl_0_10 rwl_1_10
+ rwl_0_10 cell_2r1w
Xcell_2r1w_2733 vdd_uq8 gnd read_bl_0_21 read_bl_1_21 write_bl_0_21 wwl_0_18 rwl_1_18
+ rwl_0_18 cell_2r1w
Xcell_2r1w_3434 vdd_uq9 gnd read_bl_0_10 read_bl_1_10 write_bl_0_10 wwl_0_21 rwl_1_21
+ rwl_0_21 cell_2r1w
Xcell_2r1w_2755 vdd_uq29 gnd read_bl_0_20 read_bl_1_20 write_bl_0_20 wwl_0_60 rwl_1_60
+ rwl_0_60 cell_2r1w
Xcell_2r1w_2766 vdd_uq23 gnd read_bl_0_20 read_bl_1_20 write_bl_0_20 wwl_0_49 rwl_1_49
+ rwl_0_49 cell_2r1w
Xcell_2r1w_2777 vdd_uq18 gnd read_bl_0_20 read_bl_1_20 write_bl_0_20 wwl_0_38 rwl_1_38
+ rwl_0_38 cell_2r1w
Xcell_2r1w_3489 vdd_uq14 gnd read_bl_0_9 read_bl_1_9 write_bl_0_9 wwl_0_30 rwl_1_30
+ rwl_0_30 cell_2r1w
Xcell_2r1w_2788 vdd_uq12 gnd read_bl_0_20 read_bl_1_20 write_bl_0_20 wwl_0_27 rwl_1_27
+ rwl_0_27 cell_2r1w
Xcell_2r1w_2744 vdd_uq2 gnd read_bl_0_21 read_bl_1_21 write_bl_0_21 wwl_0_7 rwl_1_7
+ rwl_0_7 cell_2r1w
Xcell_2r1w_2799 vdd_uq7 gnd read_bl_0_20 read_bl_1_20 write_bl_0_20 wwl_0_16 rwl_1_16
+ rwl_0_16 cell_2r1w
Xcell_2r1w_3990 vdd_uq19 gnd read_bl_0_1 read_bl_1_1 write_bl_0_1 wwl_0_41 rwl_1_41
+ rwl_0_41 cell_2r1w
Xcell_2r1w_2007 vdd_uq19 gnd read_bl_0_32 read_bl_1_32 write_bl_0_32 wwl_0_40 rwl_1_40
+ rwl_0_40 cell_2r1w
Xcell_2r1w_2018 vdd_uq13 gnd read_bl_0_32 read_bl_1_32 write_bl_0_32 wwl_0_29 rwl_1_29
+ rwl_0_29 cell_2r1w
Xcell_2r1w_2029 vdd_uq8 gnd read_bl_0_32 read_bl_1_32 write_bl_0_32 wwl_0_18 rwl_1_18
+ rwl_0_18 cell_2r1w
Xcell_2r1w_577 vdd_uq30 gnd read_bl_0_54 read_bl_1_54 write_bl_0_54 wwl_0_62 rwl_1_62
+ rwl_0_62 cell_2r1w
Xcell_2r1w_522 vdd_uq25 gnd read_bl_0_55 read_bl_1_55 write_bl_0_55 wwl_0_53 rwl_1_53
+ rwl_0_53 cell_2r1w
Xcell_2r1w_588 vdd_uq24 gnd read_bl_0_54 read_bl_1_54 write_bl_0_54 wwl_0_51 rwl_1_51
+ rwl_0_51 cell_2r1w
Xcell_2r1w_533 vdd_uq20 gnd read_bl_0_55 read_bl_1_55 write_bl_0_55 wwl_0_42 rwl_1_42
+ rwl_0_42 cell_2r1w
Xcell_2r1w_1306 vdd_uq17 gnd read_bl_0_43 read_bl_1_43 write_bl_0_43 wwl_0_37 rwl_1_37
+ rwl_0_37 cell_2r1w
Xcell_2r1w_544 vdd_uq14 gnd read_bl_0_55 read_bl_1_55 write_bl_0_55 wwl_0_31 rwl_1_31
+ rwl_0_31 cell_2r1w
Xcell_2r1w_1317 vdd_uq12 gnd read_bl_0_43 read_bl_1_43 write_bl_0_43 wwl_0_26 rwl_1_26
+ rwl_0_26 cell_2r1w
Xcell_2r1w_1339 vdd_uq1 gnd read_bl_0_43 read_bl_1_43 write_bl_0_43 wwl_0_4 rwl_1_4
+ rwl_0_4 cell_2r1w
Xcell_2r1w_511 vdd_uq0 gnd read_bl_0_56 read_bl_1_56 write_bl_0_56 wwl_0_0 rwl_1_0
+ rwl_0_0 cell_2r1w
Xcell_2r1w_566 vdd_uq3 gnd read_bl_0_55 read_bl_1_55 write_bl_0_55 wwl_0_9 rwl_1_9
+ rwl_0_9 cell_2r1w
Xcell_2r1w_500 vdd_uq4 gnd read_bl_0_56 read_bl_1_56 write_bl_0_56 wwl_0_11 rwl_1_11
+ rwl_0_11 cell_2r1w
Xcell_2r1w_1328 vdd_uq6 gnd read_bl_0_43 read_bl_1_43 write_bl_0_43 wwl_0_15 rwl_1_15
+ rwl_0_15 cell_2r1w
Xcell_2r1w_555 vdd_uq9 gnd read_bl_0_55 read_bl_1_55 write_bl_0_55 wwl_0_20 rwl_1_20
+ rwl_0_20 cell_2r1w
Xcell_2r1w_599 vdd_uq19 gnd read_bl_0_54 read_bl_1_54 write_bl_0_54 wwl_0_40 rwl_1_40
+ rwl_0_40 cell_2r1w
Xcell_2r1w_3264 vdd_uq30 gnd read_bl_0_12 read_bl_1_12 write_bl_0_12 wwl_0_63 rwl_1_63
+ rwl_0_63 cell_2r1w
Xcell_2r1w_2563 vdd_uq29 gnd read_bl_0_23 read_bl_1_23 write_bl_0_23 wwl_0_60 rwl_1_60
+ rwl_0_60 cell_2r1w
Xcell_2r1w_3275 vdd_uq25 gnd read_bl_0_12 read_bl_1_12 write_bl_0_12 wwl_0_52 rwl_1_52
+ rwl_0_52 cell_2r1w
Xcell_2r1w_2574 vdd_uq23 gnd read_bl_0_23 read_bl_1_23 write_bl_0_23 wwl_0_49 rwl_1_49
+ rwl_0_49 cell_2r1w
Xcell_2r1w_3220 vdd_uq20 gnd read_bl_0_13 read_bl_1_13 write_bl_0_13 wwl_0_43 rwl_1_43
+ rwl_0_43 cell_2r1w
Xcell_2r1w_3286 vdd_uq19 gnd read_bl_0_12 read_bl_1_12 write_bl_0_12 wwl_0_41 rwl_1_41
+ rwl_0_41 cell_2r1w
Xcell_2r1w_3231 vdd_uq15 gnd read_bl_0_13 read_bl_1_13 write_bl_0_13 wwl_0_32 rwl_1_32
+ rwl_0_32 cell_2r1w
Xcell_2r1w_3297 vdd_uq14 gnd read_bl_0_12 read_bl_1_12 write_bl_0_12 wwl_0_30 rwl_1_30
+ rwl_0_30 cell_2r1w
Xcell_2r1w_2530 vdd_uq13 gnd read_bl_0_24 read_bl_1_24 write_bl_0_24 wwl_0_29 rwl_1_29
+ rwl_0_29 cell_2r1w
Xcell_2r1w_2552 vdd_uq2 gnd read_bl_0_24 read_bl_1_24 write_bl_0_24 wwl_0_7 rwl_1_7
+ rwl_0_7 cell_2r1w
Xcell_2r1w_3253 vdd_uq4 gnd read_bl_0_13 read_bl_1_13 write_bl_0_13 wwl_0_10 rwl_1_10
+ rwl_0_10 cell_2r1w
Xcell_2r1w_2541 vdd_uq8 gnd read_bl_0_24 read_bl_1_24 write_bl_0_24 wwl_0_18 rwl_1_18
+ rwl_0_18 cell_2r1w
Xcell_2r1w_3242 vdd_uq9 gnd read_bl_0_13 read_bl_1_13 write_bl_0_13 wwl_0_21 rwl_1_21
+ rwl_0_21 cell_2r1w
Xcell_2r1w_1862 vdd_uq27 gnd read_bl_0_34 read_bl_1_34 write_bl_0_34 wwl_0_57 rwl_1_57
+ rwl_0_57 cell_2r1w
Xcell_2r1w_1873 vdd_uq22 gnd read_bl_0_34 read_bl_1_34 write_bl_0_34 wwl_0_46 rwl_1_46
+ rwl_0_46 cell_2r1w
Xcell_2r1w_2585 vdd_uq18 gnd read_bl_0_23 read_bl_1_23 write_bl_0_23 wwl_0_38 rwl_1_38
+ rwl_0_38 cell_2r1w
Xcell_2r1w_1884 vdd_uq16 gnd read_bl_0_34 read_bl_1_34 write_bl_0_34 wwl_0_35 rwl_1_35
+ rwl_0_35 cell_2r1w
Xcell_2r1w_2596 vdd_uq12 gnd read_bl_0_23 read_bl_1_23 write_bl_0_23 wwl_0_27 rwl_1_27
+ rwl_0_27 cell_2r1w
Xcell_2r1w_1895 vdd_uq11 gnd read_bl_0_34 read_bl_1_34 write_bl_0_34 wwl_0_24 rwl_1_24
+ rwl_0_24 cell_2r1w
Xcell_2r1w_1851 vdd_uq1 gnd read_bl_0_35 read_bl_1_35 write_bl_0_35 wwl_0_4 rwl_1_4
+ rwl_0_4 cell_2r1w
Xcell_2r1w_1840 vdd_uq6 gnd read_bl_0_35 read_bl_1_35 write_bl_0_35 wwl_0_15 rwl_1_15
+ rwl_0_15 cell_2r1w
Xcell_2r1w_1103 vdd_uq23 gnd read_bl_0_46 read_bl_1_46 write_bl_0_46 wwl_0_48 rwl_1_48
+ rwl_0_48 cell_2r1w
Xcell_2r1w_1114 vdd_uq17 gnd read_bl_0_46 read_bl_1_46 write_bl_0_46 wwl_0_37 rwl_1_37
+ rwl_0_37 cell_2r1w
Xcell_2r1w_1125 vdd_uq12 gnd read_bl_0_46 read_bl_1_46 write_bl_0_46 wwl_0_26 rwl_1_26
+ rwl_0_26 cell_2r1w
Xcell_2r1w_385 vdd_uq30 gnd read_bl_0_57 read_bl_1_57 write_bl_0_57 wwl_0_62 rwl_1_62
+ rwl_0_62 cell_2r1w
Xcell_2r1w_1158 vdd_uq27 gnd read_bl_0_45 read_bl_1_45 write_bl_0_45 wwl_0_57 rwl_1_57
+ rwl_0_57 cell_2r1w
Xcell_2r1w_330 vdd_uq25 gnd read_bl_0_58 read_bl_1_58 write_bl_0_58 wwl_0_53 rwl_1_53
+ rwl_0_53 cell_2r1w
Xcell_2r1w_396 vdd_uq24 gnd read_bl_0_57 read_bl_1_57 write_bl_0_57 wwl_0_51 rwl_1_51
+ rwl_0_51 cell_2r1w
Xcell_2r1w_1169 vdd_uq22 gnd read_bl_0_45 read_bl_1_45 write_bl_0_45 wwl_0_46 rwl_1_46
+ rwl_0_46 cell_2r1w
Xcell_2r1w_341 vdd_uq20 gnd read_bl_0_58 read_bl_1_58 write_bl_0_58 wwl_0_42 rwl_1_42
+ rwl_0_42 cell_2r1w
Xcell_2r1w_352 vdd_uq14 gnd read_bl_0_58 read_bl_1_58 write_bl_0_58 wwl_0_31 rwl_1_31
+ rwl_0_31 cell_2r1w
Xcell_2r1w_1147 vdd_uq1 gnd read_bl_0_46 read_bl_1_46 write_bl_0_46 wwl_0_4 rwl_1_4
+ rwl_0_4 cell_2r1w
Xcell_2r1w_374 vdd_uq3 gnd read_bl_0_58 read_bl_1_58 write_bl_0_58 wwl_0_9 rwl_1_9
+ rwl_0_9 cell_2r1w
Xcell_2r1w_1136 vdd_uq6 gnd read_bl_0_46 read_bl_1_46 write_bl_0_46 wwl_0_15 rwl_1_15
+ rwl_0_15 cell_2r1w
Xcell_2r1w_363 vdd_uq9 gnd read_bl_0_58 read_bl_1_58 write_bl_0_58 wwl_0_20 rwl_1_20
+ rwl_0_20 cell_2r1w
Xcell_2r1w_3072 vdd_uq30 gnd read_bl_0_15 read_bl_1_15 write_bl_0_15 wwl_0_63 rwl_1_63
+ rwl_0_63 cell_2r1w
Xcell_2r1w_2371 vdd_uq29 gnd read_bl_0_26 read_bl_1_26 write_bl_0_26 wwl_0_60 rwl_1_60
+ rwl_0_60 cell_2r1w
Xcell_2r1w_1670 vdd_uq27 gnd read_bl_0_37 read_bl_1_37 write_bl_0_37 wwl_0_57 rwl_1_57
+ rwl_0_57 cell_2r1w
Xcell_2r1w_3083 vdd_uq25 gnd read_bl_0_15 read_bl_1_15 write_bl_0_15 wwl_0_52 rwl_1_52
+ rwl_0_52 cell_2r1w
Xcell_2r1w_2382 vdd_uq23 gnd read_bl_0_26 read_bl_1_26 write_bl_0_26 wwl_0_49 rwl_1_49
+ rwl_0_49 cell_2r1w
Xcell_2r1w_1681 vdd_uq22 gnd read_bl_0_37 read_bl_1_37 write_bl_0_37 wwl_0_46 rwl_1_46
+ rwl_0_46 cell_2r1w
Xcell_2r1w_3094 vdd_uq19 gnd read_bl_0_15 read_bl_1_15 write_bl_0_15 wwl_0_41 rwl_1_41
+ rwl_0_41 cell_2r1w
Xcell_2r1w_2393 vdd_uq18 gnd read_bl_0_26 read_bl_1_26 write_bl_0_26 wwl_0_38 rwl_1_38
+ rwl_0_38 cell_2r1w
Xcell_2r1w_2360 vdd_uq2 gnd read_bl_0_27 read_bl_1_27 write_bl_0_27 wwl_0_7 rwl_1_7
+ rwl_0_7 cell_2r1w
Xcell_2r1w_3061 vdd_uq4 gnd read_bl_0_16 read_bl_1_16 write_bl_0_16 wwl_0_10 rwl_1_10
+ rwl_0_10 cell_2r1w
Xcell_2r1w_3050 vdd_uq9 gnd read_bl_0_16 read_bl_1_16 write_bl_0_16 wwl_0_21 rwl_1_21
+ rwl_0_21 cell_2r1w
Xcell_2r1w_1692 vdd_uq16 gnd read_bl_0_37 read_bl_1_37 write_bl_0_37 wwl_0_35 rwl_1_35
+ rwl_0_35 cell_2r1w
Xcell_2r1w_193 vdd_uq30 gnd read_bl_0_60 read_bl_1_60 write_bl_0_60 wwl_0_62 rwl_1_62
+ rwl_0_62 cell_2r1w
Xcell_2r1w_160 vdd_uq14 gnd read_bl_0_61 read_bl_1_61 write_bl_0_61 wwl_0_31 rwl_1_31
+ rwl_0_31 cell_2r1w
Xcell_2r1w_182 vdd_uq3 gnd read_bl_0_61 read_bl_1_61 write_bl_0_61 wwl_0_9 rwl_1_9
+ rwl_0_9 cell_2r1w
Xcell_2r1w_171 vdd_uq9 gnd read_bl_0_61 read_bl_1_61 write_bl_0_61 wwl_0_20 rwl_1_20
+ rwl_0_20 cell_2r1w
Xcell_2r1w_2190 vdd_uq23 gnd read_bl_0_29 read_bl_1_29 write_bl_0_29 wwl_0_49 rwl_1_49
+ rwl_0_49 cell_2r1w
Xcell_2r1w_3808 vdd_uq14 gnd read_bl_0_4 read_bl_1_4 write_bl_0_4 wwl_0_31 rwl_1_31
+ rwl_0_31 cell_2r1w
Xcell_2r1w_3819 vdd_uq9 gnd read_bl_0_4 read_bl_1_4 write_bl_0_4 wwl_0_20 rwl_1_20
+ rwl_0_20 cell_2r1w
Xcell_2r1w_907 vdd_uq25 gnd read_bl_0_49 read_bl_1_49 write_bl_0_49 wwl_0_52 rwl_1_52
+ rwl_0_52 cell_2r1w
Xcell_2r1w_918 vdd_uq19 gnd read_bl_0_49 read_bl_1_49 write_bl_0_49 wwl_0_41 rwl_1_41
+ rwl_0_41 cell_2r1w
Xcell_2r1w_929 vdd_uq14 gnd read_bl_0_49 read_bl_1_49 write_bl_0_49 wwl_0_30 rwl_1_30
+ rwl_0_30 cell_2r1w
Xcell_2r1w_3649 vdd_uq30 gnd read_bl_0_6 read_bl_1_6 write_bl_0_6 wwl_0_62 rwl_1_62
+ rwl_0_62 cell_2r1w
Xcell_2r1w_3605 vdd_uq20 gnd read_bl_0_7 read_bl_1_7 write_bl_0_7 wwl_0_42 rwl_1_42
+ rwl_0_42 cell_2r1w
Xcell_2r1w_2904 vdd_uq18 gnd read_bl_0_18 read_bl_1_18 write_bl_0_18 wwl_0_39 rwl_1_39
+ rwl_0_39 cell_2r1w
Xcell_2r1w_3616 vdd_uq14 gnd read_bl_0_7 read_bl_1_7 write_bl_0_7 wwl_0_31 rwl_1_31
+ rwl_0_31 cell_2r1w
Xcell_2r1w_2915 vdd_uq13 gnd read_bl_0_18 read_bl_1_18 write_bl_0_18 wwl_0_28 rwl_1_28
+ rwl_0_28 cell_2r1w
Xcell_2r1w_3638 vdd_uq3 gnd read_bl_0_7 read_bl_1_7 write_bl_0_7 wwl_0_9 rwl_1_9 rwl_0_9
+ cell_2r1w
Xcell_2r1w_3627 vdd_uq9 gnd read_bl_0_7 read_bl_1_7 write_bl_0_7 wwl_0_20 rwl_1_20
+ rwl_0_20 cell_2r1w
Xcell_2r1w_2948 vdd_uq28 gnd read_bl_0_17 read_bl_1_17 write_bl_0_17 wwl_0_59 rwl_1_59
+ rwl_0_59 cell_2r1w
Xcell_2r1w_2959 vdd_uq23 gnd read_bl_0_17 read_bl_1_17 write_bl_0_17 wwl_0_48 rwl_1_48
+ rwl_0_48 cell_2r1w
Xcell_2r1w_2937 vdd_uq2 gnd read_bl_0_18 read_bl_1_18 write_bl_0_18 wwl_0_6 rwl_1_6
+ rwl_0_6 cell_2r1w
Xcell_2r1w_2926 vdd_uq7 gnd read_bl_0_18 read_bl_1_18 write_bl_0_18 wwl_0_17 rwl_1_17
+ rwl_0_17 cell_2r1w
Xcell_2r1w_19 vdd_uq21 gnd read_bl_0_63 read_bl_1_63 write_bl_0_63 wwl_0_44 rwl_1_44
+ rwl_0_44 cell_2r1w
Xcell_2r1w_704 vdd_uq30 gnd read_bl_0_52 read_bl_1_52 write_bl_0_52 wwl_0_63 rwl_1_63
+ rwl_0_63 cell_2r1w
Xcell_2r1w_715 vdd_uq25 gnd read_bl_0_52 read_bl_1_52 write_bl_0_52 wwl_0_52 rwl_1_52
+ rwl_0_52 cell_2r1w
Xcell_2r1w_726 vdd_uq19 gnd read_bl_0_52 read_bl_1_52 write_bl_0_52 wwl_0_41 rwl_1_41
+ rwl_0_41 cell_2r1w
Xcell_2r1w_737 vdd_uq14 gnd read_bl_0_52 read_bl_1_52 write_bl_0_52 wwl_0_30 rwl_1_30
+ rwl_0_30 cell_2r1w
Xcell_2r1w_759 vdd_uq3 gnd read_bl_0_52 read_bl_1_52 write_bl_0_52 wwl_0_8 rwl_1_8
+ rwl_0_8 cell_2r1w
Xcell_2r1w_748 vdd_uq8 gnd read_bl_0_52 read_bl_1_52 write_bl_0_52 wwl_0_19 rwl_1_19
+ rwl_0_19 cell_2r1w
Xcell_2r1w_9 vdd_uq26 gnd read_bl_0_63 read_bl_1_63 write_bl_0_63 wwl_0_54 rwl_1_54
+ rwl_0_54 cell_2r1w
Xcell_2r1w_3457 vdd_uq30 gnd read_bl_0_9 read_bl_1_9 write_bl_0_9 wwl_0_62 rwl_1_62
+ rwl_0_62 cell_2r1w
Xcell_2r1w_2756 vdd_uq28 gnd read_bl_0_20 read_bl_1_20 write_bl_0_20 wwl_0_59 rwl_1_59
+ rwl_0_59 cell_2r1w
Xcell_2r1w_3402 vdd_uq25 gnd read_bl_0_10 read_bl_1_10 write_bl_0_10 wwl_0_53 rwl_1_53
+ rwl_0_53 cell_2r1w
Xcell_2r1w_3468 vdd_uq24 gnd read_bl_0_9 read_bl_1_9 write_bl_0_9 wwl_0_51 rwl_1_51
+ rwl_0_51 cell_2r1w
Xcell_2r1w_2701 vdd_uq24 gnd read_bl_0_21 read_bl_1_21 write_bl_0_21 wwl_0_50 rwl_1_50
+ rwl_0_50 cell_2r1w
Xcell_2r1w_2767 vdd_uq23 gnd read_bl_0_20 read_bl_1_20 write_bl_0_20 wwl_0_48 rwl_1_48
+ rwl_0_48 cell_2r1w
Xcell_2r1w_3413 vdd_uq20 gnd read_bl_0_10 read_bl_1_10 write_bl_0_10 wwl_0_42 rwl_1_42
+ rwl_0_42 cell_2r1w
Xcell_2r1w_3479 vdd_uq19 gnd read_bl_0_9 read_bl_1_9 write_bl_0_9 wwl_0_40 rwl_1_40
+ rwl_0_40 cell_2r1w
Xcell_2r1w_2712 vdd_uq18 gnd read_bl_0_21 read_bl_1_21 write_bl_0_21 wwl_0_39 rwl_1_39
+ rwl_0_39 cell_2r1w
Xcell_2r1w_3424 vdd_uq14 gnd read_bl_0_10 read_bl_1_10 write_bl_0_10 wwl_0_31 rwl_1_31
+ rwl_0_31 cell_2r1w
Xcell_2r1w_2723 vdd_uq13 gnd read_bl_0_21 read_bl_1_21 write_bl_0_21 wwl_0_28 rwl_1_28
+ rwl_0_28 cell_2r1w
Xcell_2r1w_2745 vdd_uq2 gnd read_bl_0_21 read_bl_1_21 write_bl_0_21 wwl_0_6 rwl_1_6
+ rwl_0_6 cell_2r1w
Xcell_2r1w_3446 vdd_uq3 gnd read_bl_0_10 read_bl_1_10 write_bl_0_10 wwl_0_9 rwl_1_9
+ rwl_0_9 cell_2r1w
Xcell_2r1w_2734 vdd_uq7 gnd read_bl_0_21 read_bl_1_21 write_bl_0_21 wwl_0_17 rwl_1_17
+ rwl_0_17 cell_2r1w
Xcell_2r1w_3435 vdd_uq9 gnd read_bl_0_10 read_bl_1_10 write_bl_0_10 wwl_0_20 rwl_1_20
+ rwl_0_20 cell_2r1w
Xcell_2r1w_2778 vdd_uq17 gnd read_bl_0_20 read_bl_1_20 write_bl_0_20 wwl_0_37 rwl_1_37
+ rwl_0_37 cell_2r1w
Xcell_2r1w_2789 vdd_uq12 gnd read_bl_0_20 read_bl_1_20 write_bl_0_20 wwl_0_26 rwl_1_26
+ rwl_0_26 cell_2r1w
Xcell_2r1w_3980 vdd_uq24 gnd read_bl_0_1 read_bl_1_1 write_bl_0_1 wwl_0_51 rwl_1_51
+ rwl_0_51 cell_2r1w
Xcell_2r1w_3991 vdd_uq19 gnd read_bl_0_1 read_bl_1_1 write_bl_0_1 wwl_0_40 rwl_1_40
+ rwl_0_40 cell_2r1w
Xcell_2r1w_2008 vdd_uq18 gnd read_bl_0_32 read_bl_1_32 write_bl_0_32 wwl_0_39 rwl_1_39
+ rwl_0_39 cell_2r1w
Xcell_2r1w_1307 vdd_uq17 gnd read_bl_0_43 read_bl_1_43 write_bl_0_43 wwl_0_36 rwl_1_36
+ rwl_0_36 cell_2r1w
Xcell_2r1w_2019 vdd_uq13 gnd read_bl_0_32 read_bl_1_32 write_bl_0_32 wwl_0_28 rwl_1_28
+ rwl_0_28 cell_2r1w
Xcell_2r1w_512 vdd_uq30 gnd read_bl_0_55 read_bl_1_55 write_bl_0_55 wwl_0_63 rwl_1_63
+ rwl_0_63 cell_2r1w
Xcell_2r1w_578 vdd_uq29 gnd read_bl_0_54 read_bl_1_54 write_bl_0_54 wwl_0_61 rwl_1_61
+ rwl_0_61 cell_2r1w
Xcell_2r1w_523 vdd_uq25 gnd read_bl_0_55 read_bl_1_55 write_bl_0_55 wwl_0_52 rwl_1_52
+ rwl_0_52 cell_2r1w
Xcell_2r1w_589 vdd_uq24 gnd read_bl_0_54 read_bl_1_54 write_bl_0_54 wwl_0_50 rwl_1_50
+ rwl_0_50 cell_2r1w
Xcell_2r1w_534 vdd_uq19 gnd read_bl_0_55 read_bl_1_55 write_bl_0_55 wwl_0_41 rwl_1_41
+ rwl_0_41 cell_2r1w
Xcell_2r1w_545 vdd_uq14 gnd read_bl_0_55 read_bl_1_55 write_bl_0_55 wwl_0_30 rwl_1_30
+ rwl_0_30 cell_2r1w
Xcell_2r1w_1318 vdd_uq11 gnd read_bl_0_43 read_bl_1_43 write_bl_0_43 wwl_0_25 rwl_1_25
+ rwl_0_25 cell_2r1w
Xcell_2r1w_567 vdd_uq3 gnd read_bl_0_55 read_bl_1_55 write_bl_0_55 wwl_0_8 rwl_1_8
+ rwl_0_8 cell_2r1w
Xcell_2r1w_501 vdd_uq4 gnd read_bl_0_56 read_bl_1_56 write_bl_0_56 wwl_0_10 rwl_1_10
+ rwl_0_10 cell_2r1w
Xcell_2r1w_1329 vdd_uq6 gnd read_bl_0_43 read_bl_1_43 write_bl_0_43 wwl_0_14 rwl_1_14
+ rwl_0_14 cell_2r1w
Xcell_2r1w_556 vdd_uq8 gnd read_bl_0_55 read_bl_1_55 write_bl_0_55 wwl_0_19 rwl_1_19
+ rwl_0_19 cell_2r1w
Xcell_2r1w_3210 vdd_uq25 gnd read_bl_0_13 read_bl_1_13 write_bl_0_13 wwl_0_53 rwl_1_53
+ rwl_0_53 cell_2r1w
Xcell_2r1w_3265 vdd_uq30 gnd read_bl_0_12 read_bl_1_12 write_bl_0_12 wwl_0_62 rwl_1_62
+ rwl_0_62 cell_2r1w
Xcell_2r1w_2564 vdd_uq28 gnd read_bl_0_23 read_bl_1_23 write_bl_0_23 wwl_0_59 rwl_1_59
+ rwl_0_59 cell_2r1w
Xcell_2r1w_1863 vdd_uq27 gnd read_bl_0_34 read_bl_1_34 write_bl_0_34 wwl_0_56 rwl_1_56
+ rwl_0_56 cell_2r1w
Xcell_2r1w_3276 vdd_uq24 gnd read_bl_0_12 read_bl_1_12 write_bl_0_12 wwl_0_51 rwl_1_51
+ rwl_0_51 cell_2r1w
Xcell_2r1w_2575 vdd_uq23 gnd read_bl_0_23 read_bl_1_23 write_bl_0_23 wwl_0_48 rwl_1_48
+ rwl_0_48 cell_2r1w
Xcell_2r1w_3221 vdd_uq20 gnd read_bl_0_13 read_bl_1_13 write_bl_0_13 wwl_0_42 rwl_1_42
+ rwl_0_42 cell_2r1w
Xcell_2r1w_3287 vdd_uq19 gnd read_bl_0_12 read_bl_1_12 write_bl_0_12 wwl_0_40 rwl_1_40
+ rwl_0_40 cell_2r1w
Xcell_2r1w_2520 vdd_uq18 gnd read_bl_0_24 read_bl_1_24 write_bl_0_24 wwl_0_39 rwl_1_39
+ rwl_0_39 cell_2r1w
Xcell_2r1w_2586 vdd_uq17 gnd read_bl_0_23 read_bl_1_23 write_bl_0_23 wwl_0_37 rwl_1_37
+ rwl_0_37 cell_2r1w
Xcell_2r1w_3232 vdd_uq14 gnd read_bl_0_13 read_bl_1_13 write_bl_0_13 wwl_0_31 rwl_1_31
+ rwl_0_31 cell_2r1w
Xcell_2r1w_3298 vdd_uq13 gnd read_bl_0_12 read_bl_1_12 write_bl_0_12 wwl_0_29 rwl_1_29
+ rwl_0_29 cell_2r1w
Xcell_2r1w_2531 vdd_uq13 gnd read_bl_0_24 read_bl_1_24 write_bl_0_24 wwl_0_28 rwl_1_28
+ rwl_0_28 cell_2r1w
Xcell_2r1w_2597 vdd_uq12 gnd read_bl_0_23 read_bl_1_23 write_bl_0_23 wwl_0_26 rwl_1_26
+ rwl_0_26 cell_2r1w
Xcell_2r1w_1830 vdd_uq11 gnd read_bl_0_35 read_bl_1_35 write_bl_0_35 wwl_0_25 rwl_1_25
+ rwl_0_25 cell_2r1w
Xcell_2r1w_1852 vdd gnd read_bl_0_35 read_bl_1_35 write_bl_0_35 wwl_0_3 rwl_1_3 rwl_0_3
+ cell_2r1w
Xcell_2r1w_2553 vdd_uq2 gnd read_bl_0_24 read_bl_1_24 write_bl_0_24 wwl_0_6 rwl_1_6
+ rwl_0_6 cell_2r1w
Xcell_2r1w_3254 vdd_uq3 gnd read_bl_0_13 read_bl_1_13 write_bl_0_13 wwl_0_9 rwl_1_9
+ rwl_0_9 cell_2r1w
Xcell_2r1w_1841 vdd_uq6 gnd read_bl_0_35 read_bl_1_35 write_bl_0_35 wwl_0_14 rwl_1_14
+ rwl_0_14 cell_2r1w
Xcell_2r1w_2542 vdd_uq7 gnd read_bl_0_24 read_bl_1_24 write_bl_0_24 wwl_0_17 rwl_1_17
+ rwl_0_17 cell_2r1w
Xcell_2r1w_3243 vdd_uq9 gnd read_bl_0_13 read_bl_1_13 write_bl_0_13 wwl_0_20 rwl_1_20
+ rwl_0_20 cell_2r1w
Xcell_2r1w_1874 vdd_uq21 gnd read_bl_0_34 read_bl_1_34 write_bl_0_34 wwl_0_45 rwl_1_45
+ rwl_0_45 cell_2r1w
Xcell_2r1w_1885 vdd_uq16 gnd read_bl_0_34 read_bl_1_34 write_bl_0_34 wwl_0_34 rwl_1_34
+ rwl_0_34 cell_2r1w
Xcell_2r1w_1896 vdd_uq10 gnd read_bl_0_34 read_bl_1_34 write_bl_0_34 wwl_0_23 rwl_1_23
+ rwl_0_23 cell_2r1w
Xcell_2r1w_320 vdd_uq30 gnd read_bl_0_58 read_bl_1_58 write_bl_0_58 wwl_0_63 rwl_1_63
+ rwl_0_63 cell_2r1w
Xcell_2r1w_1159 vdd_uq27 gnd read_bl_0_45 read_bl_1_45 write_bl_0_45 wwl_0_56 rwl_1_56
+ rwl_0_56 cell_2r1w
Xcell_2r1w_1104 vdd_uq22 gnd read_bl_0_46 read_bl_1_46 write_bl_0_46 wwl_0_47 rwl_1_47
+ rwl_0_47 cell_2r1w
Xcell_2r1w_1115 vdd_uq17 gnd read_bl_0_46 read_bl_1_46 write_bl_0_46 wwl_0_36 rwl_1_36
+ rwl_0_36 cell_2r1w
Xcell_2r1w_1126 vdd_uq11 gnd read_bl_0_46 read_bl_1_46 write_bl_0_46 wwl_0_25 rwl_1_25
+ rwl_0_25 cell_2r1w
Xcell_2r1w_1148 vdd gnd read_bl_0_46 read_bl_1_46 write_bl_0_46 wwl_0_3 rwl_1_3 rwl_0_3
+ cell_2r1w
Xcell_2r1w_1137 vdd_uq6 gnd read_bl_0_46 read_bl_1_46 write_bl_0_46 wwl_0_14 rwl_1_14
+ rwl_0_14 cell_2r1w
Xcell_2r1w_386 vdd_uq29 gnd read_bl_0_57 read_bl_1_57 write_bl_0_57 wwl_0_61 rwl_1_61
+ rwl_0_61 cell_2r1w
Xcell_2r1w_331 vdd_uq25 gnd read_bl_0_58 read_bl_1_58 write_bl_0_58 wwl_0_52 rwl_1_52
+ rwl_0_52 cell_2r1w
Xcell_2r1w_397 vdd_uq24 gnd read_bl_0_57 read_bl_1_57 write_bl_0_57 wwl_0_50 rwl_1_50
+ rwl_0_50 cell_2r1w
Xcell_2r1w_342 vdd_uq19 gnd read_bl_0_58 read_bl_1_58 write_bl_0_58 wwl_0_41 rwl_1_41
+ rwl_0_41 cell_2r1w
Xcell_2r1w_353 vdd_uq14 gnd read_bl_0_58 read_bl_1_58 write_bl_0_58 wwl_0_30 rwl_1_30
+ rwl_0_30 cell_2r1w
Xcell_2r1w_375 vdd_uq3 gnd read_bl_0_58 read_bl_1_58 write_bl_0_58 wwl_0_8 rwl_1_8
+ rwl_0_8 cell_2r1w
Xcell_2r1w_364 vdd_uq8 gnd read_bl_0_58 read_bl_1_58 write_bl_0_58 wwl_0_19 rwl_1_19
+ rwl_0_19 cell_2r1w
Xcell_2r1w_3040 vdd_uq14 gnd read_bl_0_16 read_bl_1_16 write_bl_0_16 wwl_0_31 rwl_1_31
+ rwl_0_31 cell_2r1w
Xcell_2r1w_3051 vdd_uq9 gnd read_bl_0_16 read_bl_1_16 write_bl_0_16 wwl_0_20 rwl_1_20
+ rwl_0_20 cell_2r1w
Xcell_2r1w_3073 vdd_uq30 gnd read_bl_0_15 read_bl_1_15 write_bl_0_15 wwl_0_62 rwl_1_62
+ rwl_0_62 cell_2r1w
Xcell_2r1w_2372 vdd_uq28 gnd read_bl_0_26 read_bl_1_26 write_bl_0_26 wwl_0_59 rwl_1_59
+ rwl_0_59 cell_2r1w
Xcell_2r1w_1671 vdd_uq27 gnd read_bl_0_37 read_bl_1_37 write_bl_0_37 wwl_0_56 rwl_1_56
+ rwl_0_56 cell_2r1w
Xcell_2r1w_3084 vdd_uq24 gnd read_bl_0_15 read_bl_1_15 write_bl_0_15 wwl_0_51 rwl_1_51
+ rwl_0_51 cell_2r1w
Xcell_2r1w_2383 vdd_uq23 gnd read_bl_0_26 read_bl_1_26 write_bl_0_26 wwl_0_48 rwl_1_48
+ rwl_0_48 cell_2r1w
Xcell_2r1w_1682 vdd_uq21 gnd read_bl_0_37 read_bl_1_37 write_bl_0_37 wwl_0_45 rwl_1_45
+ rwl_0_45 cell_2r1w
Xcell_2r1w_3095 vdd_uq19 gnd read_bl_0_15 read_bl_1_15 write_bl_0_15 wwl_0_40 rwl_1_40
+ rwl_0_40 cell_2r1w
Xcell_2r1w_2394 vdd_uq17 gnd read_bl_0_26 read_bl_1_26 write_bl_0_26 wwl_0_37 rwl_1_37
+ rwl_0_37 cell_2r1w
Xcell_2r1w_1693 vdd_uq16 gnd read_bl_0_37 read_bl_1_37 write_bl_0_37 wwl_0_34 rwl_1_34
+ rwl_0_34 cell_2r1w
Xcell_2r1w_1660 vdd gnd read_bl_0_38 read_bl_1_38 write_bl_0_38 wwl_0_3 rwl_1_3 rwl_0_3
+ cell_2r1w
Xcell_2r1w_2361 vdd_uq2 gnd read_bl_0_27 read_bl_1_27 write_bl_0_27 wwl_0_6 rwl_1_6
+ rwl_0_6 cell_2r1w
Xcell_2r1w_3062 vdd_uq3 gnd read_bl_0_16 read_bl_1_16 write_bl_0_16 wwl_0_9 rwl_1_9
+ rwl_0_9 cell_2r1w
Xcell_2r1w_2350 vdd_uq7 gnd read_bl_0_27 read_bl_1_27 write_bl_0_27 wwl_0_17 rwl_1_17
+ rwl_0_17 cell_2r1w
Xcell_2r1w_150 vdd_uq19 gnd read_bl_0_61 read_bl_1_61 write_bl_0_61 wwl_0_41 rwl_1_41
+ rwl_0_41 cell_2r1w
Xcell_2r1w_161 vdd_uq14 gnd read_bl_0_61 read_bl_1_61 write_bl_0_61 wwl_0_30 rwl_1_30
+ rwl_0_30 cell_2r1w
Xcell_2r1w_194 vdd_uq29 gnd read_bl_0_60 read_bl_1_60 write_bl_0_60 wwl_0_61 rwl_1_61
+ rwl_0_61 cell_2r1w
Xcell_2r1w_183 vdd_uq3 gnd read_bl_0_61 read_bl_1_61 write_bl_0_61 wwl_0_8 rwl_1_8
+ rwl_0_8 cell_2r1w
Xcell_2r1w_172 vdd_uq8 gnd read_bl_0_61 read_bl_1_61 write_bl_0_61 wwl_0_19 rwl_1_19
+ rwl_0_19 cell_2r1w
Xcell_2r1w_2180 vdd_uq28 gnd read_bl_0_29 read_bl_1_29 write_bl_0_29 wwl_0_59 rwl_1_59
+ rwl_0_59 cell_2r1w
Xcell_2r1w_2191 vdd_uq23 gnd read_bl_0_29 read_bl_1_29 write_bl_0_29 wwl_0_48 rwl_1_48
+ rwl_0_48 cell_2r1w
Xcell_2r1w_1490 vdd_uq21 gnd read_bl_0_40 read_bl_1_40 write_bl_0_40 wwl_0_45 rwl_1_45
+ rwl_0_45 cell_2r1w
Xcell_2r1w_3809 vdd_uq14 gnd read_bl_0_4 read_bl_1_4 write_bl_0_4 wwl_0_30 rwl_1_30
+ rwl_0_30 cell_2r1w
Xcell_2r1w_908 vdd_uq24 gnd read_bl_0_49 read_bl_1_49 write_bl_0_49 wwl_0_51 rwl_1_51
+ rwl_0_51 cell_2r1w
Xcell_2r1w_919 vdd_uq19 gnd read_bl_0_49 read_bl_1_49 write_bl_0_49 wwl_0_40 rwl_1_40
+ rwl_0_40 cell_2r1w
Xcell_2r1w_2949 vdd_uq28 gnd read_bl_0_17 read_bl_1_17 write_bl_0_17 wwl_0_58 rwl_1_58
+ rwl_0_58 cell_2r1w
Xcell_2r1w_3606 vdd_uq19 gnd read_bl_0_7 read_bl_1_7 write_bl_0_7 wwl_0_41 rwl_1_41
+ rwl_0_41 cell_2r1w
Xcell_2r1w_2905 vdd_uq18 gnd read_bl_0_18 read_bl_1_18 write_bl_0_18 wwl_0_38 rwl_1_38
+ rwl_0_38 cell_2r1w
Xcell_2r1w_3617 vdd_uq14 gnd read_bl_0_7 read_bl_1_7 write_bl_0_7 wwl_0_30 rwl_1_30
+ rwl_0_30 cell_2r1w
Xcell_2r1w_2916 vdd_uq12 gnd read_bl_0_18 read_bl_1_18 write_bl_0_18 wwl_0_27 rwl_1_27
+ rwl_0_27 cell_2r1w
Xcell_2r1w_2938 vdd_uq1 gnd read_bl_0_18 read_bl_1_18 write_bl_0_18 wwl_0_5 rwl_1_5
+ rwl_0_5 cell_2r1w
Xcell_2r1w_3639 vdd_uq3 gnd read_bl_0_7 read_bl_1_7 write_bl_0_7 wwl_0_8 rwl_1_8 rwl_0_8
+ cell_2r1w
Xcell_2r1w_2927 vdd_uq7 gnd read_bl_0_18 read_bl_1_18 write_bl_0_18 wwl_0_16 rwl_1_16
+ rwl_0_16 cell_2r1w
Xcell_2r1w_3628 vdd_uq8 gnd read_bl_0_7 read_bl_1_7 write_bl_0_7 wwl_0_19 rwl_1_19
+ rwl_0_19 cell_2r1w
Xcell_2r1w_705 vdd_uq30 gnd read_bl_0_52 read_bl_1_52 write_bl_0_52 wwl_0_62 rwl_1_62
+ rwl_0_62 cell_2r1w
Xcell_2r1w_716 vdd_uq24 gnd read_bl_0_52 read_bl_1_52 write_bl_0_52 wwl_0_51 rwl_1_51
+ rwl_0_51 cell_2r1w
Xcell_2r1w_727 vdd_uq19 gnd read_bl_0_52 read_bl_1_52 write_bl_0_52 wwl_0_40 rwl_1_40
+ rwl_0_40 cell_2r1w
Xcell_2r1w_738 vdd_uq13 gnd read_bl_0_52 read_bl_1_52 write_bl_0_52 wwl_0_29 rwl_1_29
+ rwl_0_29 cell_2r1w
Xcell_2r1w_749 vdd_uq8 gnd read_bl_0_52 read_bl_1_52 write_bl_0_52 wwl_0_18 rwl_1_18
+ rwl_0_18 cell_2r1w
Xcell_2r1w_3458 vdd_uq29 gnd read_bl_0_9 read_bl_1_9 write_bl_0_9 wwl_0_61 rwl_1_61
+ rwl_0_61 cell_2r1w
Xcell_2r1w_2757 vdd_uq28 gnd read_bl_0_20 read_bl_1_20 write_bl_0_20 wwl_0_58 rwl_1_58
+ rwl_0_58 cell_2r1w
Xcell_2r1w_3403 vdd_uq25 gnd read_bl_0_10 read_bl_1_10 write_bl_0_10 wwl_0_52 rwl_1_52
+ rwl_0_52 cell_2r1w
Xcell_2r1w_3469 vdd_uq24 gnd read_bl_0_9 read_bl_1_9 write_bl_0_9 wwl_0_50 rwl_1_50
+ rwl_0_50 cell_2r1w
Xcell_2r1w_2702 vdd_uq23 gnd read_bl_0_21 read_bl_1_21 write_bl_0_21 wwl_0_49 rwl_1_49
+ rwl_0_49 cell_2r1w
Xcell_2r1w_2768 vdd_uq22 gnd read_bl_0_20 read_bl_1_20 write_bl_0_20 wwl_0_47 rwl_1_47
+ rwl_0_47 cell_2r1w
Xcell_2r1w_3414 vdd_uq19 gnd read_bl_0_10 read_bl_1_10 write_bl_0_10 wwl_0_41 rwl_1_41
+ rwl_0_41 cell_2r1w
Xcell_2r1w_2713 vdd_uq18 gnd read_bl_0_21 read_bl_1_21 write_bl_0_21 wwl_0_38 rwl_1_38
+ rwl_0_38 cell_2r1w
Xcell_2r1w_2779 vdd_uq17 gnd read_bl_0_20 read_bl_1_20 write_bl_0_20 wwl_0_36 rwl_1_36
+ rwl_0_36 cell_2r1w
Xcell_2r1w_3425 vdd_uq14 gnd read_bl_0_10 read_bl_1_10 write_bl_0_10 wwl_0_30 rwl_1_30
+ rwl_0_30 cell_2r1w
Xcell_2r1w_2724 vdd_uq12 gnd read_bl_0_21 read_bl_1_21 write_bl_0_21 wwl_0_27 rwl_1_27
+ rwl_0_27 cell_2r1w
Xcell_2r1w_2746 vdd_uq1 gnd read_bl_0_21 read_bl_1_21 write_bl_0_21 wwl_0_5 rwl_1_5
+ rwl_0_5 cell_2r1w
Xcell_2r1w_3447 vdd_uq3 gnd read_bl_0_10 read_bl_1_10 write_bl_0_10 wwl_0_8 rwl_1_8
+ rwl_0_8 cell_2r1w
Xcell_2r1w_2735 vdd_uq7 gnd read_bl_0_21 read_bl_1_21 write_bl_0_21 wwl_0_16 rwl_1_16
+ rwl_0_16 cell_2r1w
Xcell_2r1w_3436 vdd_uq8 gnd read_bl_0_10 read_bl_1_10 write_bl_0_10 wwl_0_19 rwl_1_19
+ rwl_0_19 cell_2r1w
Xcell_2r1w_3970 vdd_uq29 gnd read_bl_0_1 read_bl_1_1 write_bl_0_1 wwl_0_61 rwl_1_61
+ rwl_0_61 cell_2r1w
Xcell_2r1w_3981 vdd_uq24 gnd read_bl_0_1 read_bl_1_1 write_bl_0_1 wwl_0_50 rwl_1_50
+ rwl_0_50 cell_2r1w
Xcell_2r1w_3992 vdd_uq18 gnd read_bl_0_1 read_bl_1_1 write_bl_0_1 wwl_0_39 rwl_1_39
+ rwl_0_39 cell_2r1w
Xcell_2r1w_2009 vdd_uq18 gnd read_bl_0_32 read_bl_1_32 write_bl_0_32 wwl_0_38 rwl_1_38
+ rwl_0_38 cell_2r1w
Xcell_2r1w_1308 vdd_uq16 gnd read_bl_0_43 read_bl_1_43 write_bl_0_43 wwl_0_35 rwl_1_35
+ rwl_0_35 cell_2r1w
Xcell_2r1w_1319 vdd_uq11 gnd read_bl_0_43 read_bl_1_43 write_bl_0_43 wwl_0_24 rwl_1_24
+ rwl_0_24 cell_2r1w
Xcell_2r1w_502 vdd_uq3 gnd read_bl_0_56 read_bl_1_56 write_bl_0_56 wwl_0_9 rwl_1_9
+ rwl_0_9 cell_2r1w
Xcell_2r1w_513 vdd_uq30 gnd read_bl_0_55 read_bl_1_55 write_bl_0_55 wwl_0_62 rwl_1_62
+ rwl_0_62 cell_2r1w
Xcell_2r1w_579 vdd_uq29 gnd read_bl_0_54 read_bl_1_54 write_bl_0_54 wwl_0_60 rwl_1_60
+ rwl_0_60 cell_2r1w
Xcell_2r1w_524 vdd_uq24 gnd read_bl_0_55 read_bl_1_55 write_bl_0_55 wwl_0_51 rwl_1_51
+ rwl_0_51 cell_2r1w
Xcell_2r1w_535 vdd_uq19 gnd read_bl_0_55 read_bl_1_55 write_bl_0_55 wwl_0_40 rwl_1_40
+ rwl_0_40 cell_2r1w
Xcell_2r1w_546 vdd_uq13 gnd read_bl_0_55 read_bl_1_55 write_bl_0_55 wwl_0_29 rwl_1_29
+ rwl_0_29 cell_2r1w
Xcell_2r1w_568 vdd_uq2 gnd read_bl_0_55 read_bl_1_55 write_bl_0_55 wwl_0_7 rwl_1_7
+ rwl_0_7 cell_2r1w
Xcell_2r1w_557 vdd_uq8 gnd read_bl_0_55 read_bl_1_55 write_bl_0_55 wwl_0_18 rwl_1_18
+ rwl_0_18 cell_2r1w
Xcell_2r1w_3200 vdd_uq30 gnd read_bl_0_13 read_bl_1_13 write_bl_0_13 wwl_0_63 rwl_1_63
+ rwl_0_63 cell_2r1w
Xcell_2r1w_3211 vdd_uq25 gnd read_bl_0_13 read_bl_1_13 write_bl_0_13 wwl_0_52 rwl_1_52
+ rwl_0_52 cell_2r1w
Xcell_2r1w_3222 vdd_uq19 gnd read_bl_0_13 read_bl_1_13 write_bl_0_13 wwl_0_41 rwl_1_41
+ rwl_0_41 cell_2r1w
Xcell_2r1w_3233 vdd_uq14 gnd read_bl_0_13 read_bl_1_13 write_bl_0_13 wwl_0_30 rwl_1_30
+ rwl_0_30 cell_2r1w
Xcell_2r1w_3244 vdd_uq8 gnd read_bl_0_13 read_bl_1_13 write_bl_0_13 wwl_0_19 rwl_1_19
+ rwl_0_19 cell_2r1w
Xcell_2r1w_3266 vdd_uq29 gnd read_bl_0_12 read_bl_1_12 write_bl_0_12 wwl_0_61 rwl_1_61
+ rwl_0_61 cell_2r1w
Xcell_2r1w_2565 vdd_uq28 gnd read_bl_0_23 read_bl_1_23 write_bl_0_23 wwl_0_58 rwl_1_58
+ rwl_0_58 cell_2r1w
Xcell_2r1w_1864 vdd_uq26 gnd read_bl_0_34 read_bl_1_34 write_bl_0_34 wwl_0_55 rwl_1_55
+ rwl_0_55 cell_2r1w
Xcell_2r1w_3277 vdd_uq24 gnd read_bl_0_12 read_bl_1_12 write_bl_0_12 wwl_0_50 rwl_1_50
+ rwl_0_50 cell_2r1w
Xcell_2r1w_2510 vdd_uq23 gnd read_bl_0_24 read_bl_1_24 write_bl_0_24 wwl_0_49 rwl_1_49
+ rwl_0_49 cell_2r1w
Xcell_2r1w_2576 vdd_uq22 gnd read_bl_0_23 read_bl_1_23 write_bl_0_23 wwl_0_47 rwl_1_47
+ rwl_0_47 cell_2r1w
Xcell_2r1w_1875 vdd_uq21 gnd read_bl_0_34 read_bl_1_34 write_bl_0_34 wwl_0_44 rwl_1_44
+ rwl_0_44 cell_2r1w
Xcell_2r1w_3288 vdd_uq18 gnd read_bl_0_12 read_bl_1_12 write_bl_0_12 wwl_0_39 rwl_1_39
+ rwl_0_39 cell_2r1w
Xcell_2r1w_2521 vdd_uq18 gnd read_bl_0_24 read_bl_1_24 write_bl_0_24 wwl_0_38 rwl_1_38
+ rwl_0_38 cell_2r1w
Xcell_2r1w_2587 vdd_uq17 gnd read_bl_0_23 read_bl_1_23 write_bl_0_23 wwl_0_36 rwl_1_36
+ rwl_0_36 cell_2r1w
Xcell_2r1w_1820 vdd_uq16 gnd read_bl_0_35 read_bl_1_35 write_bl_0_35 wwl_0_35 rwl_1_35
+ rwl_0_35 cell_2r1w
Xcell_2r1w_1886 vdd_uq15 gnd read_bl_0_34 read_bl_1_34 write_bl_0_34 wwl_0_33 rwl_1_33
+ rwl_0_33 cell_2r1w
Xcell_2r1w_2532 vdd_uq12 gnd read_bl_0_24 read_bl_1_24 write_bl_0_24 wwl_0_27 rwl_1_27
+ rwl_0_27 cell_2r1w
Xcell_2r1w_3299 vdd_uq13 gnd read_bl_0_12 read_bl_1_12 write_bl_0_12 wwl_0_28 rwl_1_28
+ rwl_0_28 cell_2r1w
Xcell_2r1w_2598 vdd_uq11 gnd read_bl_0_23 read_bl_1_23 write_bl_0_23 wwl_0_25 rwl_1_25
+ rwl_0_25 cell_2r1w
Xcell_2r1w_1831 vdd_uq11 gnd read_bl_0_35 read_bl_1_35 write_bl_0_35 wwl_0_24 rwl_1_24
+ rwl_0_24 cell_2r1w
Xcell_2r1w_2554 vdd_uq1 gnd read_bl_0_24 read_bl_1_24 write_bl_0_24 wwl_0_5 rwl_1_5
+ rwl_0_5 cell_2r1w
Xcell_2r1w_1853 vdd gnd read_bl_0_35 read_bl_1_35 write_bl_0_35 wwl_0_2 rwl_1_2 rwl_0_2
+ cell_2r1w
Xcell_2r1w_3255 vdd_uq3 gnd read_bl_0_13 read_bl_1_13 write_bl_0_13 wwl_0_8 rwl_1_8
+ rwl_0_8 cell_2r1w
Xcell_2r1w_1842 vdd_uq5 gnd read_bl_0_35 read_bl_1_35 write_bl_0_35 wwl_0_13 rwl_1_13
+ rwl_0_13 cell_2r1w
Xcell_2r1w_2543 vdd_uq7 gnd read_bl_0_24 read_bl_1_24 write_bl_0_24 wwl_0_16 rwl_1_16
+ rwl_0_16 cell_2r1w
Xcell_2r1w_1897 vdd_uq10 gnd read_bl_0_34 read_bl_1_34 write_bl_0_34 wwl_0_22 rwl_1_22
+ rwl_0_22 cell_2r1w
Xcell_2r1w_321 vdd_uq30 gnd read_bl_0_58 read_bl_1_58 write_bl_0_58 wwl_0_62 rwl_1_62
+ rwl_0_62 cell_2r1w
Xcell_2r1w_332 vdd_uq24 gnd read_bl_0_58 read_bl_1_58 write_bl_0_58 wwl_0_51 rwl_1_51
+ rwl_0_51 cell_2r1w
Xcell_2r1w_1105 vdd_uq22 gnd read_bl_0_46 read_bl_1_46 write_bl_0_46 wwl_0_46 rwl_1_46
+ rwl_0_46 cell_2r1w
Xcell_2r1w_343 vdd_uq19 gnd read_bl_0_58 read_bl_1_58 write_bl_0_58 wwl_0_40 rwl_1_40
+ rwl_0_40 cell_2r1w
Xcell_2r1w_1116 vdd_uq16 gnd read_bl_0_46 read_bl_1_46 write_bl_0_46 wwl_0_35 rwl_1_35
+ rwl_0_35 cell_2r1w
Xcell_2r1w_354 vdd_uq13 gnd read_bl_0_58 read_bl_1_58 write_bl_0_58 wwl_0_29 rwl_1_29
+ rwl_0_29 cell_2r1w
Xcell_2r1w_1127 vdd_uq11 gnd read_bl_0_46 read_bl_1_46 write_bl_0_46 wwl_0_24 rwl_1_24
+ rwl_0_24 cell_2r1w
Xcell_2r1w_1149 vdd gnd read_bl_0_46 read_bl_1_46 write_bl_0_46 wwl_0_2 rwl_1_2 rwl_0_2
+ cell_2r1w
Xcell_2r1w_310 vdd_uq3 gnd read_bl_0_59 read_bl_1_59 write_bl_0_59 wwl_0_9 rwl_1_9
+ rwl_0_9 cell_2r1w
Xcell_2r1w_1138 vdd_uq5 gnd read_bl_0_46 read_bl_1_46 write_bl_0_46 wwl_0_13 rwl_1_13
+ rwl_0_13 cell_2r1w
Xcell_2r1w_387 vdd_uq29 gnd read_bl_0_57 read_bl_1_57 write_bl_0_57 wwl_0_60 rwl_1_60
+ rwl_0_60 cell_2r1w
Xcell_2r1w_398 vdd_uq23 gnd read_bl_0_57 read_bl_1_57 write_bl_0_57 wwl_0_49 rwl_1_49
+ rwl_0_49 cell_2r1w
Xcell_2r1w_376 vdd_uq2 gnd read_bl_0_58 read_bl_1_58 write_bl_0_58 wwl_0_7 rwl_1_7
+ rwl_0_7 cell_2r1w
Xcell_2r1w_365 vdd_uq8 gnd read_bl_0_58 read_bl_1_58 write_bl_0_58 wwl_0_18 rwl_1_18
+ rwl_0_18 cell_2r1w
Xcell_2r1w_3074 vdd_uq29 gnd read_bl_0_15 read_bl_1_15 write_bl_0_15 wwl_0_61 rwl_1_61
+ rwl_0_61 cell_2r1w
Xcell_2r1w_3085 vdd_uq24 gnd read_bl_0_15 read_bl_1_15 write_bl_0_15 wwl_0_50 rwl_1_50
+ rwl_0_50 cell_2r1w
Xcell_2r1w_3030 vdd_uq19 gnd read_bl_0_16 read_bl_1_16 write_bl_0_16 wwl_0_41 rwl_1_41
+ rwl_0_41 cell_2r1w
Xcell_2r1w_3041 vdd_uq14 gnd read_bl_0_16 read_bl_1_16 write_bl_0_16 wwl_0_30 rwl_1_30
+ rwl_0_30 cell_2r1w
Xcell_2r1w_2340 vdd_uq12 gnd read_bl_0_27 read_bl_1_27 write_bl_0_27 wwl_0_27 rwl_1_27
+ rwl_0_27 cell_2r1w
Xcell_2r1w_3063 vdd_uq3 gnd read_bl_0_16 read_bl_1_16 write_bl_0_16 wwl_0_8 rwl_1_8
+ rwl_0_8 cell_2r1w
Xcell_2r1w_3052 vdd_uq8 gnd read_bl_0_16 read_bl_1_16 write_bl_0_16 wwl_0_19 rwl_1_19
+ rwl_0_19 cell_2r1w
Xcell_2r1w_2373 vdd_uq28 gnd read_bl_0_26 read_bl_1_26 write_bl_0_26 wwl_0_58 rwl_1_58
+ rwl_0_58 cell_2r1w
Xcell_2r1w_1672 vdd_uq26 gnd read_bl_0_37 read_bl_1_37 write_bl_0_37 wwl_0_55 rwl_1_55
+ rwl_0_55 cell_2r1w
Xcell_2r1w_2384 vdd_uq22 gnd read_bl_0_26 read_bl_1_26 write_bl_0_26 wwl_0_47 rwl_1_47
+ rwl_0_47 cell_2r1w
Xcell_2r1w_1683 vdd_uq21 gnd read_bl_0_37 read_bl_1_37 write_bl_0_37 wwl_0_44 rwl_1_44
+ rwl_0_44 cell_2r1w
Xcell_2r1w_3096 vdd_uq18 gnd read_bl_0_15 read_bl_1_15 write_bl_0_15 wwl_0_39 rwl_1_39
+ rwl_0_39 cell_2r1w
Xcell_2r1w_2395 vdd_uq17 gnd read_bl_0_26 read_bl_1_26 write_bl_0_26 wwl_0_36 rwl_1_36
+ rwl_0_36 cell_2r1w
Xcell_2r1w_1694 vdd_uq15 gnd read_bl_0_37 read_bl_1_37 write_bl_0_37 wwl_0_33 rwl_1_33
+ rwl_0_33 cell_2r1w
Xcell_2r1w_2362 vdd_uq1 gnd read_bl_0_27 read_bl_1_27 write_bl_0_27 wwl_0_5 rwl_1_5
+ rwl_0_5 cell_2r1w
Xcell_2r1w_1661 vdd gnd read_bl_0_38 read_bl_1_38 write_bl_0_38 wwl_0_2 rwl_1_2 rwl_0_2
+ cell_2r1w
Xcell_2r1w_1650 vdd_uq5 gnd read_bl_0_38 read_bl_1_38 write_bl_0_38 wwl_0_13 rwl_1_13
+ rwl_0_13 cell_2r1w
Xcell_2r1w_2351 vdd_uq7 gnd read_bl_0_27 read_bl_1_27 write_bl_0_27 wwl_0_16 rwl_1_16
+ rwl_0_16 cell_2r1w
Xcell_2r1w_195 vdd_uq29 gnd read_bl_0_60 read_bl_1_60 write_bl_0_60 wwl_0_60 rwl_1_60
+ rwl_0_60 cell_2r1w
Xcell_2r1w_140 vdd_uq24 gnd read_bl_0_61 read_bl_1_61 write_bl_0_61 wwl_0_51 rwl_1_51
+ rwl_0_51 cell_2r1w
Xcell_2r1w_151 vdd_uq19 gnd read_bl_0_61 read_bl_1_61 write_bl_0_61 wwl_0_40 rwl_1_40
+ rwl_0_40 cell_2r1w
Xcell_2r1w_162 vdd_uq13 gnd read_bl_0_61 read_bl_1_61 write_bl_0_61 wwl_0_29 rwl_1_29
+ rwl_0_29 cell_2r1w
Xcell_2r1w_184 vdd_uq2 gnd read_bl_0_61 read_bl_1_61 write_bl_0_61 wwl_0_7 rwl_1_7
+ rwl_0_7 cell_2r1w
Xcell_2r1w_173 vdd_uq8 gnd read_bl_0_61 read_bl_1_61 write_bl_0_61 wwl_0_18 rwl_1_18
+ rwl_0_18 cell_2r1w
Xcell_2r1w_2181 vdd_uq28 gnd read_bl_0_29 read_bl_1_29 write_bl_0_29 wwl_0_58 rwl_1_58
+ rwl_0_58 cell_2r1w
Xcell_2r1w_2192 vdd_uq22 gnd read_bl_0_29 read_bl_1_29 write_bl_0_29 wwl_0_47 rwl_1_47
+ rwl_0_47 cell_2r1w
Xcell_2r1w_2170 vdd_uq1 gnd read_bl_0_30 read_bl_1_30 write_bl_0_30 wwl_0_5 rwl_1_5
+ rwl_0_5 cell_2r1w
Xcell_2r1w_1480 vdd_uq26 gnd read_bl_0_40 read_bl_1_40 write_bl_0_40 wwl_0_55 rwl_1_55
+ rwl_0_55 cell_2r1w
Xcell_2r1w_1491 vdd_uq21 gnd read_bl_0_40 read_bl_1_40 write_bl_0_40 wwl_0_44 rwl_1_44
+ rwl_0_44 cell_2r1w
Xcell_2r1w_909 vdd_uq24 gnd read_bl_0_49 read_bl_1_49 write_bl_0_49 wwl_0_50 rwl_1_50
+ rwl_0_50 cell_2r1w
Xcell_2r1w_3607 vdd_uq19 gnd read_bl_0_7 read_bl_1_7 write_bl_0_7 wwl_0_40 rwl_1_40
+ rwl_0_40 cell_2r1w
Xcell_2r1w_2906 vdd_uq17 gnd read_bl_0_18 read_bl_1_18 write_bl_0_18 wwl_0_37 rwl_1_37
+ rwl_0_37 cell_2r1w
Xcell_2r1w_3618 vdd_uq13 gnd read_bl_0_7 read_bl_1_7 write_bl_0_7 wwl_0_29 rwl_1_29
+ rwl_0_29 cell_2r1w
Xcell_2r1w_2917 vdd_uq12 gnd read_bl_0_18 read_bl_1_18 write_bl_0_18 wwl_0_26 rwl_1_26
+ rwl_0_26 cell_2r1w
Xcell_2r1w_2939 vdd_uq1 gnd read_bl_0_18 read_bl_1_18 write_bl_0_18 wwl_0_4 rwl_1_4
+ rwl_0_4 cell_2r1w
Xcell_2r1w_2928 vdd_uq6 gnd read_bl_0_18 read_bl_1_18 write_bl_0_18 wwl_0_15 rwl_1_15
+ rwl_0_15 cell_2r1w
Xcell_2r1w_3629 vdd_uq8 gnd read_bl_0_7 read_bl_1_7 write_bl_0_7 wwl_0_18 rwl_1_18
+ rwl_0_18 cell_2r1w
Xcell_2r1w_706 vdd_uq29 gnd read_bl_0_52 read_bl_1_52 write_bl_0_52 wwl_0_61 rwl_1_61
+ rwl_0_61 cell_2r1w
Xcell_2r1w_717 vdd_uq24 gnd read_bl_0_52 read_bl_1_52 write_bl_0_52 wwl_0_50 rwl_1_50
+ rwl_0_50 cell_2r1w
Xcell_2r1w_728 vdd_uq18 gnd read_bl_0_52 read_bl_1_52 write_bl_0_52 wwl_0_39 rwl_1_39
+ rwl_0_39 cell_2r1w
Xcell_2r1w_739 vdd_uq13 gnd read_bl_0_52 read_bl_1_52 write_bl_0_52 wwl_0_28 rwl_1_28
+ rwl_0_28 cell_2r1w
Xcell_2r1w_3404 vdd_uq24 gnd read_bl_0_10 read_bl_1_10 write_bl_0_10 wwl_0_51 rwl_1_51
+ rwl_0_51 cell_2r1w
Xcell_2r1w_3415 vdd_uq19 gnd read_bl_0_10 read_bl_1_10 write_bl_0_10 wwl_0_40 rwl_1_40
+ rwl_0_40 cell_2r1w
Xcell_2r1w_3426 vdd_uq13 gnd read_bl_0_10 read_bl_1_10 write_bl_0_10 wwl_0_29 rwl_1_29
+ rwl_0_29 cell_2r1w
Xcell_2r1w_3459 vdd_uq29 gnd read_bl_0_9 read_bl_1_9 write_bl_0_9 wwl_0_60 rwl_1_60
+ rwl_0_60 cell_2r1w
Xcell_2r1w_2758 vdd_uq27 gnd read_bl_0_20 read_bl_1_20 write_bl_0_20 wwl_0_57 rwl_1_57
+ rwl_0_57 cell_2r1w
Xcell_2r1w_2703 vdd_uq23 gnd read_bl_0_21 read_bl_1_21 write_bl_0_21 wwl_0_48 rwl_1_48
+ rwl_0_48 cell_2r1w
Xcell_2r1w_2769 vdd_uq22 gnd read_bl_0_20 read_bl_1_20 write_bl_0_20 wwl_0_46 rwl_1_46
+ rwl_0_46 cell_2r1w
Xcell_2r1w_2714 vdd_uq17 gnd read_bl_0_21 read_bl_1_21 write_bl_0_21 wwl_0_37 rwl_1_37
+ rwl_0_37 cell_2r1w
Xcell_2r1w_2725 vdd_uq12 gnd read_bl_0_21 read_bl_1_21 write_bl_0_21 wwl_0_26 rwl_1_26
+ rwl_0_26 cell_2r1w
Xcell_2r1w_2747 vdd_uq1 gnd read_bl_0_21 read_bl_1_21 write_bl_0_21 wwl_0_4 rwl_1_4
+ rwl_0_4 cell_2r1w
Xcell_2r1w_3448 vdd_uq2 gnd read_bl_0_10 read_bl_1_10 write_bl_0_10 wwl_0_7 rwl_1_7
+ rwl_0_7 cell_2r1w
Xcell_2r1w_2736 vdd_uq6 gnd read_bl_0_21 read_bl_1_21 write_bl_0_21 wwl_0_15 rwl_1_15
+ rwl_0_15 cell_2r1w
Xcell_2r1w_3437 vdd_uq8 gnd read_bl_0_10 read_bl_1_10 write_bl_0_10 wwl_0_18 rwl_1_18
+ rwl_0_18 cell_2r1w
Xcell_2r1w_3971 vdd_uq29 gnd read_bl_0_1 read_bl_1_1 write_bl_0_1 wwl_0_60 rwl_1_60
+ rwl_0_60 cell_2r1w
Xcell_2r1w_3982 vdd_uq23 gnd read_bl_0_1 read_bl_1_1 write_bl_0_1 wwl_0_49 rwl_1_49
+ rwl_0_49 cell_2r1w
Xcell_2r1w_3960 vdd_uq2 gnd read_bl_0_2 read_bl_1_2 write_bl_0_2 wwl_0_7 rwl_1_7 rwl_0_7
+ cell_2r1w
Xcell_2r1w_3993 vdd_uq18 gnd read_bl_0_1 read_bl_1_1 write_bl_0_1 wwl_0_38 rwl_1_38
+ rwl_0_38 cell_2r1w
Xcell_2r1w_514 vdd_uq29 gnd read_bl_0_55 read_bl_1_55 write_bl_0_55 wwl_0_61 rwl_1_61
+ rwl_0_61 cell_2r1w
Xcell_2r1w_525 vdd_uq24 gnd read_bl_0_55 read_bl_1_55 write_bl_0_55 wwl_0_50 rwl_1_50
+ rwl_0_50 cell_2r1w
Xcell_2r1w_536 vdd_uq18 gnd read_bl_0_55 read_bl_1_55 write_bl_0_55 wwl_0_39 rwl_1_39
+ rwl_0_39 cell_2r1w
Xcell_2r1w_1309 vdd_uq16 gnd read_bl_0_43 read_bl_1_43 write_bl_0_43 wwl_0_34 rwl_1_34
+ rwl_0_34 cell_2r1w
Xcell_2r1w_503 vdd_uq3 gnd read_bl_0_56 read_bl_1_56 write_bl_0_56 wwl_0_8 rwl_1_8
+ rwl_0_8 cell_2r1w
Xcell_2r1w_547 vdd_uq13 gnd read_bl_0_55 read_bl_1_55 write_bl_0_55 wwl_0_28 rwl_1_28
+ rwl_0_28 cell_2r1w
Xcell_2r1w_569 vdd_uq2 gnd read_bl_0_55 read_bl_1_55 write_bl_0_55 wwl_0_6 rwl_1_6
+ rwl_0_6 cell_2r1w
Xcell_2r1w_558 vdd_uq7 gnd read_bl_0_55 read_bl_1_55 write_bl_0_55 wwl_0_17 rwl_1_17
+ rwl_0_17 cell_2r1w
Xcell_2r1w_3201 vdd_uq30 gnd read_bl_0_13 read_bl_1_13 write_bl_0_13 wwl_0_62 rwl_1_62
+ rwl_0_62 cell_2r1w
Xcell_2r1w_3267 vdd_uq29 gnd read_bl_0_12 read_bl_1_12 write_bl_0_12 wwl_0_60 rwl_1_60
+ rwl_0_60 cell_2r1w
Xcell_2r1w_2500 vdd_uq28 gnd read_bl_0_24 read_bl_1_24 write_bl_0_24 wwl_0_59 rwl_1_59
+ rwl_0_59 cell_2r1w
Xcell_2r1w_3212 vdd_uq24 gnd read_bl_0_13 read_bl_1_13 write_bl_0_13 wwl_0_51 rwl_1_51
+ rwl_0_51 cell_2r1w
Xcell_2r1w_2511 vdd_uq23 gnd read_bl_0_24 read_bl_1_24 write_bl_0_24 wwl_0_48 rwl_1_48
+ rwl_0_48 cell_2r1w
Xcell_2r1w_3223 vdd_uq19 gnd read_bl_0_13 read_bl_1_13 write_bl_0_13 wwl_0_40 rwl_1_40
+ rwl_0_40 cell_2r1w
Xcell_2r1w_2522 vdd_uq17 gnd read_bl_0_24 read_bl_1_24 write_bl_0_24 wwl_0_37 rwl_1_37
+ rwl_0_37 cell_2r1w
Xcell_2r1w_3234 vdd_uq13 gnd read_bl_0_13 read_bl_1_13 write_bl_0_13 wwl_0_29 rwl_1_29
+ rwl_0_29 cell_2r1w
Xcell_2r1w_2533 vdd_uq12 gnd read_bl_0_24 read_bl_1_24 write_bl_0_24 wwl_0_26 rwl_1_26
+ rwl_0_26 cell_2r1w
Xcell_2r1w_3256 vdd_uq2 gnd read_bl_0_13 read_bl_1_13 write_bl_0_13 wwl_0_7 rwl_1_7
+ rwl_0_7 cell_2r1w
Xcell_2r1w_3245 vdd_uq8 gnd read_bl_0_13 read_bl_1_13 write_bl_0_13 wwl_0_18 rwl_1_18
+ rwl_0_18 cell_2r1w
Xcell_2r1w_2566 vdd_uq27 gnd read_bl_0_23 read_bl_1_23 write_bl_0_23 wwl_0_57 rwl_1_57
+ rwl_0_57 cell_2r1w
Xcell_2r1w_1865 vdd_uq26 gnd read_bl_0_34 read_bl_1_34 write_bl_0_34 wwl_0_54 rwl_1_54
+ rwl_0_54 cell_2r1w
Xcell_2r1w_3278 vdd_uq23 gnd read_bl_0_12 read_bl_1_12 write_bl_0_12 wwl_0_49 rwl_1_49
+ rwl_0_49 cell_2r1w
Xcell_2r1w_2577 vdd_uq22 gnd read_bl_0_23 read_bl_1_23 write_bl_0_23 wwl_0_46 rwl_1_46
+ rwl_0_46 cell_2r1w
Xcell_2r1w_1810 vdd_uq21 gnd read_bl_0_35 read_bl_1_35 write_bl_0_35 wwl_0_45 rwl_1_45
+ rwl_0_45 cell_2r1w
Xcell_2r1w_1876 vdd_uq20 gnd read_bl_0_34 read_bl_1_34 write_bl_0_34 wwl_0_43 rwl_1_43
+ rwl_0_43 cell_2r1w
Xcell_2r1w_3289 vdd_uq18 gnd read_bl_0_12 read_bl_1_12 write_bl_0_12 wwl_0_38 rwl_1_38
+ rwl_0_38 cell_2r1w
Xcell_2r1w_2588 vdd_uq16 gnd read_bl_0_23 read_bl_1_23 write_bl_0_23 wwl_0_35 rwl_1_35
+ rwl_0_35 cell_2r1w
Xcell_2r1w_1821 vdd_uq16 gnd read_bl_0_35 read_bl_1_35 write_bl_0_35 wwl_0_34 rwl_1_34
+ rwl_0_34 cell_2r1w
Xcell_2r1w_1887 vdd_uq15 gnd read_bl_0_34 read_bl_1_34 write_bl_0_34 wwl_0_32 rwl_1_32
+ rwl_0_32 cell_2r1w
Xcell_2r1w_2599 vdd_uq11 gnd read_bl_0_23 read_bl_1_23 write_bl_0_23 wwl_0_24 rwl_1_24
+ rwl_0_24 cell_2r1w
Xcell_2r1w_2555 vdd_uq1 gnd read_bl_0_24 read_bl_1_24 write_bl_0_24 wwl_0_4 rwl_1_4
+ rwl_0_4 cell_2r1w
Xcell_2r1w_1854 vdd_uq0 gnd read_bl_0_35 read_bl_1_35 write_bl_0_35 wwl_0_1 rwl_1_1
+ rwl_0_1 cell_2r1w
Xcell_2r1w_1843 vdd_uq5 gnd read_bl_0_35 read_bl_1_35 write_bl_0_35 wwl_0_12 rwl_1_12
+ rwl_0_12 cell_2r1w
Xcell_2r1w_2544 vdd_uq6 gnd read_bl_0_24 read_bl_1_24 write_bl_0_24 wwl_0_15 rwl_1_15
+ rwl_0_15 cell_2r1w
Xcell_2r1w_1898 vdd_uq9 gnd read_bl_0_34 read_bl_1_34 write_bl_0_34 wwl_0_21 rwl_1_21
+ rwl_0_21 cell_2r1w
Xcell_2r1w_1832 vdd_uq10 gnd read_bl_0_35 read_bl_1_35 write_bl_0_35 wwl_0_23 rwl_1_23
+ rwl_0_23 cell_2r1w
Xcell_2r1w_3790 vdd_uq23 gnd read_bl_0_4 read_bl_1_4 write_bl_0_4 wwl_0_49 rwl_1_49
+ rwl_0_49 cell_2r1w
Xcell_2r1w_322 vdd_uq29 gnd read_bl_0_58 read_bl_1_58 write_bl_0_58 wwl_0_61 rwl_1_61
+ rwl_0_61 cell_2r1w
Xcell_2r1w_333 vdd_uq24 gnd read_bl_0_58 read_bl_1_58 write_bl_0_58 wwl_0_50 rwl_1_50
+ rwl_0_50 cell_2r1w
Xcell_2r1w_1106 vdd_uq21 gnd read_bl_0_46 read_bl_1_46 write_bl_0_46 wwl_0_45 rwl_1_45
+ rwl_0_45 cell_2r1w
Xcell_2r1w_344 vdd_uq18 gnd read_bl_0_58 read_bl_1_58 write_bl_0_58 wwl_0_39 rwl_1_39
+ rwl_0_39 cell_2r1w
Xcell_2r1w_1117 vdd_uq16 gnd read_bl_0_46 read_bl_1_46 write_bl_0_46 wwl_0_34 rwl_1_34
+ rwl_0_34 cell_2r1w
Xcell_2r1w_355 vdd_uq13 gnd read_bl_0_58 read_bl_1_58 write_bl_0_58 wwl_0_28 rwl_1_28
+ rwl_0_28 cell_2r1w
Xcell_2r1w_377 vdd_uq2 gnd read_bl_0_58 read_bl_1_58 write_bl_0_58 wwl_0_6 rwl_1_6
+ rwl_0_6 cell_2r1w
Xcell_2r1w_311 vdd_uq3 gnd read_bl_0_59 read_bl_1_59 write_bl_0_59 wwl_0_8 rwl_1_8
+ rwl_0_8 cell_2r1w
Xcell_2r1w_1139 vdd_uq5 gnd read_bl_0_46 read_bl_1_46 write_bl_0_46 wwl_0_12 rwl_1_12
+ rwl_0_12 cell_2r1w
Xcell_2r1w_366 vdd_uq7 gnd read_bl_0_58 read_bl_1_58 write_bl_0_58 wwl_0_17 rwl_1_17
+ rwl_0_17 cell_2r1w
Xcell_2r1w_300 vdd_uq8 gnd read_bl_0_59 read_bl_1_59 write_bl_0_59 wwl_0_19 rwl_1_19
+ rwl_0_19 cell_2r1w
Xcell_2r1w_1128 vdd_uq10 gnd read_bl_0_46 read_bl_1_46 write_bl_0_46 wwl_0_23 rwl_1_23
+ rwl_0_23 cell_2r1w
Xcell_2r1w_388 vdd_uq28 gnd read_bl_0_57 read_bl_1_57 write_bl_0_57 wwl_0_59 rwl_1_59
+ rwl_0_59 cell_2r1w
Xcell_2r1w_399 vdd_uq23 gnd read_bl_0_57 read_bl_1_57 write_bl_0_57 wwl_0_48 rwl_1_48
+ rwl_0_48 cell_2r1w
Xcell_2r1w_3075 vdd_uq29 gnd read_bl_0_15 read_bl_1_15 write_bl_0_15 wwl_0_60 rwl_1_60
+ rwl_0_60 cell_2r1w
Xcell_2r1w_2374 vdd_uq27 gnd read_bl_0_26 read_bl_1_26 write_bl_0_26 wwl_0_57 rwl_1_57
+ rwl_0_57 cell_2r1w
Xcell_2r1w_3020 vdd_uq24 gnd read_bl_0_16 read_bl_1_16 write_bl_0_16 wwl_0_51 rwl_1_51
+ rwl_0_51 cell_2r1w
Xcell_2r1w_3086 vdd_uq23 gnd read_bl_0_15 read_bl_1_15 write_bl_0_15 wwl_0_49 rwl_1_49
+ rwl_0_49 cell_2r1w
Xcell_2r1w_3031 vdd_uq19 gnd read_bl_0_16 read_bl_1_16 write_bl_0_16 wwl_0_40 rwl_1_40
+ rwl_0_40 cell_2r1w
Xcell_2r1w_3097 vdd_uq18 gnd read_bl_0_15 read_bl_1_15 write_bl_0_15 wwl_0_38 rwl_1_38
+ rwl_0_38 cell_2r1w
Xcell_2r1w_2330 vdd_uq17 gnd read_bl_0_27 read_bl_1_27 write_bl_0_27 wwl_0_37 rwl_1_37
+ rwl_0_37 cell_2r1w
Xcell_2r1w_3042 vdd_uq13 gnd read_bl_0_16 read_bl_1_16 write_bl_0_16 wwl_0_29 rwl_1_29
+ rwl_0_29 cell_2r1w
Xcell_2r1w_2341 vdd_uq12 gnd read_bl_0_27 read_bl_1_27 write_bl_0_27 wwl_0_26 rwl_1_26
+ rwl_0_26 cell_2r1w
Xcell_2r1w_2363 vdd_uq1 gnd read_bl_0_27 read_bl_1_27 write_bl_0_27 wwl_0_4 rwl_1_4
+ rwl_0_4 cell_2r1w
Xcell_2r1w_3064 vdd_uq2 gnd read_bl_0_16 read_bl_1_16 write_bl_0_16 wwl_0_7 rwl_1_7
+ rwl_0_7 cell_2r1w
Xcell_2r1w_2352 vdd_uq6 gnd read_bl_0_27 read_bl_1_27 write_bl_0_27 wwl_0_15 rwl_1_15
+ rwl_0_15 cell_2r1w
Xcell_2r1w_3053 vdd_uq8 gnd read_bl_0_16 read_bl_1_16 write_bl_0_16 wwl_0_18 rwl_1_18
+ rwl_0_18 cell_2r1w
Xcell_2r1w_1673 vdd_uq26 gnd read_bl_0_37 read_bl_1_37 write_bl_0_37 wwl_0_54 rwl_1_54
+ rwl_0_54 cell_2r1w
Xcell_2r1w_2385 vdd_uq22 gnd read_bl_0_26 read_bl_1_26 write_bl_0_26 wwl_0_46 rwl_1_46
+ rwl_0_46 cell_2r1w
Xcell_2r1w_1684 vdd_uq20 gnd read_bl_0_37 read_bl_1_37 write_bl_0_37 wwl_0_43 rwl_1_43
+ rwl_0_43 cell_2r1w
Xcell_2r1w_2396 vdd_uq16 gnd read_bl_0_26 read_bl_1_26 write_bl_0_26 wwl_0_35 rwl_1_35
+ rwl_0_35 cell_2r1w
Xcell_2r1w_1695 vdd_uq15 gnd read_bl_0_37 read_bl_1_37 write_bl_0_37 wwl_0_32 rwl_1_32
+ rwl_0_32 cell_2r1w
Xcell_2r1w_1662 vdd_uq0 gnd read_bl_0_38 read_bl_1_38 write_bl_0_38 wwl_0_1 rwl_1_1
+ rwl_0_1 cell_2r1w
Xcell_2r1w_1651 vdd_uq5 gnd read_bl_0_38 read_bl_1_38 write_bl_0_38 wwl_0_12 rwl_1_12
+ rwl_0_12 cell_2r1w
Xcell_2r1w_1640 vdd_uq10 gnd read_bl_0_38 read_bl_1_38 write_bl_0_38 wwl_0_23 rwl_1_23
+ rwl_0_23 cell_2r1w
Xcell_2r1w_130 vdd_uq29 gnd read_bl_0_61 read_bl_1_61 write_bl_0_61 wwl_0_61 rwl_1_61
+ rwl_0_61 cell_2r1w
Xcell_2r1w_196 vdd_uq28 gnd read_bl_0_60 read_bl_1_60 write_bl_0_60 wwl_0_59 rwl_1_59
+ rwl_0_59 cell_2r1w
Xcell_2r1w_141 vdd_uq24 gnd read_bl_0_61 read_bl_1_61 write_bl_0_61 wwl_0_50 rwl_1_50
+ rwl_0_50 cell_2r1w
Xcell_2r1w_152 vdd_uq18 gnd read_bl_0_61 read_bl_1_61 write_bl_0_61 wwl_0_39 rwl_1_39
+ rwl_0_39 cell_2r1w
Xcell_2r1w_163 vdd_uq13 gnd read_bl_0_61 read_bl_1_61 write_bl_0_61 wwl_0_28 rwl_1_28
+ rwl_0_28 cell_2r1w
Xcell_2r1w_185 vdd_uq2 gnd read_bl_0_61 read_bl_1_61 write_bl_0_61 wwl_0_6 rwl_1_6
+ rwl_0_6 cell_2r1w
Xcell_2r1w_174 vdd_uq7 gnd read_bl_0_61 read_bl_1_61 write_bl_0_61 wwl_0_17 rwl_1_17
+ rwl_0_17 cell_2r1w
Xcell_2r1w_2182 vdd_uq27 gnd read_bl_0_29 read_bl_1_29 write_bl_0_29 wwl_0_57 rwl_1_57
+ rwl_0_57 cell_2r1w
Xcell_2r1w_1481 vdd_uq26 gnd read_bl_0_40 read_bl_1_40 write_bl_0_40 wwl_0_54 rwl_1_54
+ rwl_0_54 cell_2r1w
Xcell_2r1w_2193 vdd_uq22 gnd read_bl_0_29 read_bl_1_29 write_bl_0_29 wwl_0_46 rwl_1_46
+ rwl_0_46 cell_2r1w
Xcell_2r1w_2171 vdd_uq1 gnd read_bl_0_30 read_bl_1_30 write_bl_0_30 wwl_0_4 rwl_1_4
+ rwl_0_4 cell_2r1w
Xcell_2r1w_1470 vdd_uq0 gnd read_bl_0_41 read_bl_1_41 write_bl_0_41 wwl_0_1 rwl_1_1
+ rwl_0_1 cell_2r1w
Xcell_2r1w_2160 vdd_uq6 gnd read_bl_0_30 read_bl_1_30 write_bl_0_30 wwl_0_15 rwl_1_15
+ rwl_0_15 cell_2r1w
Xcell_2r1w_1492 vdd_uq20 gnd read_bl_0_40 read_bl_1_40 write_bl_0_40 wwl_0_43 rwl_1_43
+ rwl_0_43 cell_2r1w
Xcell_2r1w_3608 vdd_uq18 gnd read_bl_0_7 read_bl_1_7 write_bl_0_7 wwl_0_39 rwl_1_39
+ rwl_0_39 cell_2r1w
Xcell_2r1w_2907 vdd_uq17 gnd read_bl_0_18 read_bl_1_18 write_bl_0_18 wwl_0_36 rwl_1_36
+ rwl_0_36 cell_2r1w
Xcell_2r1w_3619 vdd_uq13 gnd read_bl_0_7 read_bl_1_7 write_bl_0_7 wwl_0_28 rwl_1_28
+ rwl_0_28 cell_2r1w
Xcell_2r1w_2918 vdd_uq11 gnd read_bl_0_18 read_bl_1_18 write_bl_0_18 wwl_0_25 rwl_1_25
+ rwl_0_25 cell_2r1w
Xcell_2r1w_2929 vdd_uq6 gnd read_bl_0_18 read_bl_1_18 write_bl_0_18 wwl_0_14 rwl_1_14
+ rwl_0_14 cell_2r1w
Xcell_2r1w_707 vdd_uq29 gnd read_bl_0_52 read_bl_1_52 write_bl_0_52 wwl_0_60 rwl_1_60
+ rwl_0_60 cell_2r1w
Xcell_2r1w_718 vdd_uq23 gnd read_bl_0_52 read_bl_1_52 write_bl_0_52 wwl_0_49 rwl_1_49
+ rwl_0_49 cell_2r1w
Xcell_2r1w_729 vdd_uq18 gnd read_bl_0_52 read_bl_1_52 write_bl_0_52 wwl_0_38 rwl_1_38
+ rwl_0_38 cell_2r1w
Xcell_2r1w_3405 vdd_uq24 gnd read_bl_0_10 read_bl_1_10 write_bl_0_10 wwl_0_50 rwl_1_50
+ rwl_0_50 cell_2r1w
Xcell_2r1w_2704 vdd_uq22 gnd read_bl_0_21 read_bl_1_21 write_bl_0_21 wwl_0_47 rwl_1_47
+ rwl_0_47 cell_2r1w
Xcell_2r1w_3416 vdd_uq18 gnd read_bl_0_10 read_bl_1_10 write_bl_0_10 wwl_0_39 rwl_1_39
+ rwl_0_39 cell_2r1w
Xcell_2r1w_2715 vdd_uq17 gnd read_bl_0_21 read_bl_1_21 write_bl_0_21 wwl_0_36 rwl_1_36
+ rwl_0_36 cell_2r1w
Xcell_2r1w_3427 vdd_uq13 gnd read_bl_0_10 read_bl_1_10 write_bl_0_10 wwl_0_28 rwl_1_28
+ rwl_0_28 cell_2r1w
Xcell_2r1w_3449 vdd_uq2 gnd read_bl_0_10 read_bl_1_10 write_bl_0_10 wwl_0_6 rwl_1_6
+ rwl_0_6 cell_2r1w
Xcell_2r1w_3438 vdd_uq7 gnd read_bl_0_10 read_bl_1_10 write_bl_0_10 wwl_0_17 rwl_1_17
+ rwl_0_17 cell_2r1w
Xcell_2r1w_2759 vdd_uq27 gnd read_bl_0_20 read_bl_1_20 write_bl_0_20 wwl_0_56 rwl_1_56
+ rwl_0_56 cell_2r1w
Xcell_2r1w_2726 vdd_uq11 gnd read_bl_0_21 read_bl_1_21 write_bl_0_21 wwl_0_25 rwl_1_25
+ rwl_0_25 cell_2r1w
Xcell_2r1w_2748 vdd gnd read_bl_0_21 read_bl_1_21 write_bl_0_21 wwl_0_3 rwl_1_3 rwl_0_3
+ cell_2r1w
Xcell_2r1w_2737 vdd_uq6 gnd read_bl_0_21 read_bl_1_21 write_bl_0_21 wwl_0_14 rwl_1_14
+ rwl_0_14 cell_2r1w
Xcell_2r1w_3972 vdd_uq28 gnd read_bl_0_1 read_bl_1_1 write_bl_0_1 wwl_0_59 rwl_1_59
+ rwl_0_59 cell_2r1w
Xcell_2r1w_3983 vdd_uq23 gnd read_bl_0_1 read_bl_1_1 write_bl_0_1 wwl_0_48 rwl_1_48
+ rwl_0_48 cell_2r1w
Xcell_2r1w_3994 vdd_uq17 gnd read_bl_0_1 read_bl_1_1 write_bl_0_1 wwl_0_37 rwl_1_37
+ rwl_0_37 cell_2r1w
Xcell_2r1w_3961 vdd_uq2 gnd read_bl_0_2 read_bl_1_2 write_bl_0_2 wwl_0_6 rwl_1_6 rwl_0_6
+ cell_2r1w
Xcell_2r1w_3950 vdd_uq7 gnd read_bl_0_2 read_bl_1_2 write_bl_0_2 wwl_0_17 rwl_1_17
+ rwl_0_17 cell_2r1w
Xcell_2r1w_515 vdd_uq29 gnd read_bl_0_55 read_bl_1_55 write_bl_0_55 wwl_0_60 rwl_1_60
+ rwl_0_60 cell_2r1w
Xcell_2r1w_526 vdd_uq23 gnd read_bl_0_55 read_bl_1_55 write_bl_0_55 wwl_0_49 rwl_1_49
+ rwl_0_49 cell_2r1w
Xcell_2r1w_537 vdd_uq18 gnd read_bl_0_55 read_bl_1_55 write_bl_0_55 wwl_0_38 rwl_1_38
+ rwl_0_38 cell_2r1w
Xcell_2r1w_548 vdd_uq12 gnd read_bl_0_55 read_bl_1_55 write_bl_0_55 wwl_0_27 rwl_1_27
+ rwl_0_27 cell_2r1w
Xcell_2r1w_504 vdd_uq2 gnd read_bl_0_56 read_bl_1_56 write_bl_0_56 wwl_0_7 rwl_1_7
+ rwl_0_7 cell_2r1w
Xcell_2r1w_559 vdd_uq7 gnd read_bl_0_55 read_bl_1_55 write_bl_0_55 wwl_0_16 rwl_1_16
+ rwl_0_16 cell_2r1w
Xcell_2r1w_3202 vdd_uq29 gnd read_bl_0_13 read_bl_1_13 write_bl_0_13 wwl_0_61 rwl_1_61
+ rwl_0_61 cell_2r1w
Xcell_2r1w_3268 vdd_uq28 gnd read_bl_0_12 read_bl_1_12 write_bl_0_12 wwl_0_59 rwl_1_59
+ rwl_0_59 cell_2r1w
Xcell_2r1w_2501 vdd_uq28 gnd read_bl_0_24 read_bl_1_24 write_bl_0_24 wwl_0_58 rwl_1_58
+ rwl_0_58 cell_2r1w
Xcell_2r1w_1800 vdd_uq26 gnd read_bl_0_35 read_bl_1_35 write_bl_0_35 wwl_0_55 rwl_1_55
+ rwl_0_55 cell_2r1w
Xcell_2r1w_3213 vdd_uq24 gnd read_bl_0_13 read_bl_1_13 write_bl_0_13 wwl_0_50 rwl_1_50
+ rwl_0_50 cell_2r1w
Xcell_2r1w_3279 vdd_uq23 gnd read_bl_0_12 read_bl_1_12 write_bl_0_12 wwl_0_48 rwl_1_48
+ rwl_0_48 cell_2r1w
Xcell_2r1w_2512 vdd_uq22 gnd read_bl_0_24 read_bl_1_24 write_bl_0_24 wwl_0_47 rwl_1_47
+ rwl_0_47 cell_2r1w
Xcell_2r1w_1811 vdd_uq21 gnd read_bl_0_35 read_bl_1_35 write_bl_0_35 wwl_0_44 rwl_1_44
+ rwl_0_44 cell_2r1w
Xcell_2r1w_3224 vdd_uq18 gnd read_bl_0_13 read_bl_1_13 write_bl_0_13 wwl_0_39 rwl_1_39
+ rwl_0_39 cell_2r1w
Xcell_2r1w_2523 vdd_uq17 gnd read_bl_0_24 read_bl_1_24 write_bl_0_24 wwl_0_36 rwl_1_36
+ rwl_0_36 cell_2r1w
Xcell_2r1w_3235 vdd_uq13 gnd read_bl_0_13 read_bl_1_13 write_bl_0_13 wwl_0_28 rwl_1_28
+ rwl_0_28 cell_2r1w
Xcell_2r1w_2534 vdd_uq11 gnd read_bl_0_24 read_bl_1_24 write_bl_0_24 wwl_0_25 rwl_1_25
+ rwl_0_25 cell_2r1w
Xcell_2r1w_2556 vdd gnd read_bl_0_24 read_bl_1_24 write_bl_0_24 wwl_0_3 rwl_1_3 rwl_0_3
+ cell_2r1w
Xcell_2r1w_3257 vdd_uq2 gnd read_bl_0_13 read_bl_1_13 write_bl_0_13 wwl_0_6 rwl_1_6
+ rwl_0_6 cell_2r1w
Xcell_2r1w_2545 vdd_uq6 gnd read_bl_0_24 read_bl_1_24 write_bl_0_24 wwl_0_14 rwl_1_14
+ rwl_0_14 cell_2r1w
Xcell_2r1w_3246 vdd_uq7 gnd read_bl_0_13 read_bl_1_13 write_bl_0_13 wwl_0_17 rwl_1_17
+ rwl_0_17 cell_2r1w
Xcell_2r1w_2567 vdd_uq27 gnd read_bl_0_23 read_bl_1_23 write_bl_0_23 wwl_0_56 rwl_1_56
+ rwl_0_56 cell_2r1w
Xcell_2r1w_1866 vdd_uq25 gnd read_bl_0_34 read_bl_1_34 write_bl_0_34 wwl_0_53 rwl_1_53
+ rwl_0_53 cell_2r1w
Xcell_2r1w_2578 vdd_uq21 gnd read_bl_0_23 read_bl_1_23 write_bl_0_23 wwl_0_45 rwl_1_45
+ rwl_0_45 cell_2r1w
Xcell_2r1w_1877 vdd_uq20 gnd read_bl_0_34 read_bl_1_34 write_bl_0_34 wwl_0_42 rwl_1_42
+ rwl_0_42 cell_2r1w
Xcell_2r1w_2589 vdd_uq16 gnd read_bl_0_23 read_bl_1_23 write_bl_0_23 wwl_0_34 rwl_1_34
+ rwl_0_34 cell_2r1w
Xcell_2r1w_1822 vdd_uq15 gnd read_bl_0_35 read_bl_1_35 write_bl_0_35 wwl_0_33 rwl_1_33
+ rwl_0_33 cell_2r1w
Xcell_2r1w_1888 vdd_uq14 gnd read_bl_0_34 read_bl_1_34 write_bl_0_34 wwl_0_31 rwl_1_31
+ rwl_0_31 cell_2r1w
Xcell_2r1w_1855 vdd_uq0 gnd read_bl_0_35 read_bl_1_35 write_bl_0_35 wwl_0_0 rwl_1_0
+ rwl_0_0 cell_2r1w
Xcell_2r1w_1844 vdd_uq4 gnd read_bl_0_35 read_bl_1_35 write_bl_0_35 wwl_0_11 rwl_1_11
+ rwl_0_11 cell_2r1w
Xcell_2r1w_1899 vdd_uq9 gnd read_bl_0_34 read_bl_1_34 write_bl_0_34 wwl_0_20 rwl_1_20
+ rwl_0_20 cell_2r1w
Xcell_2r1w_1833 vdd_uq10 gnd read_bl_0_35 read_bl_1_35 write_bl_0_35 wwl_0_22 rwl_1_22
+ rwl_0_22 cell_2r1w
Xcell_2r1w_3780 vdd_uq28 gnd read_bl_0_4 read_bl_1_4 write_bl_0_4 wwl_0_59 rwl_1_59
+ rwl_0_59 cell_2r1w
Xcell_2r1w_3791 vdd_uq23 gnd read_bl_0_4 read_bl_1_4 write_bl_0_4 wwl_0_48 rwl_1_48
+ rwl_0_48 cell_2r1w
Xcell_2r1w_1107 vdd_uq21 gnd read_bl_0_46 read_bl_1_46 write_bl_0_46 wwl_0_44 rwl_1_44
+ rwl_0_44 cell_2r1w
Xcell_2r1w_323 vdd_uq29 gnd read_bl_0_58 read_bl_1_58 write_bl_0_58 wwl_0_60 rwl_1_60
+ rwl_0_60 cell_2r1w
Xcell_2r1w_389 vdd_uq28 gnd read_bl_0_57 read_bl_1_57 write_bl_0_57 wwl_0_58 rwl_1_58
+ rwl_0_58 cell_2r1w
Xcell_2r1w_334 vdd_uq23 gnd read_bl_0_58 read_bl_1_58 write_bl_0_58 wwl_0_49 rwl_1_49
+ rwl_0_49 cell_2r1w
Xcell_2r1w_345 vdd_uq18 gnd read_bl_0_58 read_bl_1_58 write_bl_0_58 wwl_0_38 rwl_1_38
+ rwl_0_38 cell_2r1w
Xcell_2r1w_1118 vdd_uq15 gnd read_bl_0_46 read_bl_1_46 write_bl_0_46 wwl_0_33 rwl_1_33
+ rwl_0_33 cell_2r1w
Xcell_2r1w_356 vdd_uq12 gnd read_bl_0_58 read_bl_1_58 write_bl_0_58 wwl_0_27 rwl_1_27
+ rwl_0_27 cell_2r1w
Xcell_2r1w_378 vdd_uq1 gnd read_bl_0_58 read_bl_1_58 write_bl_0_58 wwl_0_5 rwl_1_5
+ rwl_0_5 cell_2r1w
Xcell_2r1w_312 vdd_uq2 gnd read_bl_0_59 read_bl_1_59 write_bl_0_59 wwl_0_7 rwl_1_7
+ rwl_0_7 cell_2r1w
Xcell_2r1w_367 vdd_uq7 gnd read_bl_0_58 read_bl_1_58 write_bl_0_58 wwl_0_16 rwl_1_16
+ rwl_0_16 cell_2r1w
Xcell_2r1w_301 vdd_uq8 gnd read_bl_0_59 read_bl_1_59 write_bl_0_59 wwl_0_18 rwl_1_18
+ rwl_0_18 cell_2r1w
Xcell_2r1w_1129 vdd_uq10 gnd read_bl_0_46 read_bl_1_46 write_bl_0_46 wwl_0_22 rwl_1_22
+ rwl_0_22 cell_2r1w
Xcell_2r1w_3010 vdd_uq29 gnd read_bl_0_16 read_bl_1_16 write_bl_0_16 wwl_0_61 rwl_1_61
+ rwl_0_61 cell_2r1w
Xcell_2r1w_3076 vdd_uq28 gnd read_bl_0_15 read_bl_1_15 write_bl_0_15 wwl_0_59 rwl_1_59
+ rwl_0_59 cell_2r1w
Xcell_2r1w_2375 vdd_uq27 gnd read_bl_0_26 read_bl_1_26 write_bl_0_26 wwl_0_56 rwl_1_56
+ rwl_0_56 cell_2r1w
Xcell_2r1w_3021 vdd_uq24 gnd read_bl_0_16 read_bl_1_16 write_bl_0_16 wwl_0_50 rwl_1_50
+ rwl_0_50 cell_2r1w
Xcell_2r1w_3087 vdd_uq23 gnd read_bl_0_15 read_bl_1_15 write_bl_0_15 wwl_0_48 rwl_1_48
+ rwl_0_48 cell_2r1w
Xcell_2r1w_2320 vdd_uq22 gnd read_bl_0_27 read_bl_1_27 write_bl_0_27 wwl_0_47 rwl_1_47
+ rwl_0_47 cell_2r1w
Xcell_2r1w_2386 vdd_uq21 gnd read_bl_0_26 read_bl_1_26 write_bl_0_26 wwl_0_45 rwl_1_45
+ rwl_0_45 cell_2r1w
Xcell_2r1w_3032 vdd_uq18 gnd read_bl_0_16 read_bl_1_16 write_bl_0_16 wwl_0_39 rwl_1_39
+ rwl_0_39 cell_2r1w
Xcell_2r1w_3098 vdd_uq17 gnd read_bl_0_15 read_bl_1_15 write_bl_0_15 wwl_0_37 rwl_1_37
+ rwl_0_37 cell_2r1w
Xcell_2r1w_2331 vdd_uq17 gnd read_bl_0_27 read_bl_1_27 write_bl_0_27 wwl_0_36 rwl_1_36
+ rwl_0_36 cell_2r1w
Xcell_2r1w_2397 vdd_uq16 gnd read_bl_0_26 read_bl_1_26 write_bl_0_26 wwl_0_34 rwl_1_34
+ rwl_0_34 cell_2r1w
Xcell_2r1w_1630 vdd_uq15 gnd read_bl_0_38 read_bl_1_38 write_bl_0_38 wwl_0_33 rwl_1_33
+ rwl_0_33 cell_2r1w
Xcell_2r1w_3043 vdd_uq13 gnd read_bl_0_16 read_bl_1_16 write_bl_0_16 wwl_0_28 rwl_1_28
+ rwl_0_28 cell_2r1w
Xcell_2r1w_2342 vdd_uq11 gnd read_bl_0_27 read_bl_1_27 write_bl_0_27 wwl_0_25 rwl_1_25
+ rwl_0_25 cell_2r1w
Xcell_2r1w_2364 vdd gnd read_bl_0_27 read_bl_1_27 write_bl_0_27 wwl_0_3 rwl_1_3 rwl_0_3
+ cell_2r1w
Xcell_2r1w_1663 vdd_uq0 gnd read_bl_0_38 read_bl_1_38 write_bl_0_38 wwl_0_0 rwl_1_0
+ rwl_0_0 cell_2r1w
Xcell_2r1w_3065 vdd_uq2 gnd read_bl_0_16 read_bl_1_16 write_bl_0_16 wwl_0_6 rwl_1_6
+ rwl_0_6 cell_2r1w
Xcell_2r1w_1652 vdd_uq4 gnd read_bl_0_38 read_bl_1_38 write_bl_0_38 wwl_0_11 rwl_1_11
+ rwl_0_11 cell_2r1w
Xcell_2r1w_2353 vdd_uq6 gnd read_bl_0_27 read_bl_1_27 write_bl_0_27 wwl_0_14 rwl_1_14
+ rwl_0_14 cell_2r1w
Xcell_2r1w_3054 vdd_uq7 gnd read_bl_0_16 read_bl_1_16 write_bl_0_16 wwl_0_17 rwl_1_17
+ rwl_0_17 cell_2r1w
Xcell_2r1w_1641 vdd_uq10 gnd read_bl_0_38 read_bl_1_38 write_bl_0_38 wwl_0_22 rwl_1_22
+ rwl_0_22 cell_2r1w
Xcell_2r1w_1674 vdd_uq25 gnd read_bl_0_37 read_bl_1_37 write_bl_0_37 wwl_0_53 rwl_1_53
+ rwl_0_53 cell_2r1w
Xcell_2r1w_1685 vdd_uq20 gnd read_bl_0_37 read_bl_1_37 write_bl_0_37 wwl_0_42 rwl_1_42
+ rwl_0_42 cell_2r1w
Xcell_2r1w_1696 vdd_uq14 gnd read_bl_0_37 read_bl_1_37 write_bl_0_37 wwl_0_31 rwl_1_31
+ rwl_0_31 cell_2r1w
Xcell_2r1w_890 vdd_uq1 gnd read_bl_0_50 read_bl_1_50 write_bl_0_50 wwl_0_5 rwl_1_5
+ rwl_0_5 cell_2r1w
Xcell_2r1w_120 vdd_uq2 gnd read_bl_0_62 read_bl_1_62 write_bl_0_62 wwl_0_7 rwl_1_7
+ rwl_0_7 cell_2r1w
Xcell_2r1w_131 vdd_uq29 gnd read_bl_0_61 read_bl_1_61 write_bl_0_61 wwl_0_60 rwl_1_60
+ rwl_0_60 cell_2r1w
Xcell_2r1w_197 vdd_uq28 gnd read_bl_0_60 read_bl_1_60 write_bl_0_60 wwl_0_58 rwl_1_58
+ rwl_0_58 cell_2r1w
Xcell_2r1w_142 vdd_uq23 gnd read_bl_0_61 read_bl_1_61 write_bl_0_61 wwl_0_49 rwl_1_49
+ rwl_0_49 cell_2r1w
Xcell_2r1w_153 vdd_uq18 gnd read_bl_0_61 read_bl_1_61 write_bl_0_61 wwl_0_38 rwl_1_38
+ rwl_0_38 cell_2r1w
Xcell_2r1w_164 vdd_uq12 gnd read_bl_0_61 read_bl_1_61 write_bl_0_61 wwl_0_27 rwl_1_27
+ rwl_0_27 cell_2r1w
Xcell_2r1w_186 vdd_uq1 gnd read_bl_0_61 read_bl_1_61 write_bl_0_61 wwl_0_5 rwl_1_5
+ rwl_0_5 cell_2r1w
Xcell_2r1w_175 vdd_uq7 gnd read_bl_0_61 read_bl_1_61 write_bl_0_61 wwl_0_16 rwl_1_16
+ rwl_0_16 cell_2r1w
Xcell_2r1w_2183 vdd_uq27 gnd read_bl_0_29 read_bl_1_29 write_bl_0_29 wwl_0_56 rwl_1_56
+ rwl_0_56 cell_2r1w
Xcell_2r1w_1482 vdd_uq25 gnd read_bl_0_40 read_bl_1_40 write_bl_0_40 wwl_0_53 rwl_1_53
+ rwl_0_53 cell_2r1w
Xcell_2r1w_2194 vdd_uq21 gnd read_bl_0_29 read_bl_1_29 write_bl_0_29 wwl_0_45 rwl_1_45
+ rwl_0_45 cell_2r1w
Xcell_2r1w_1493 vdd_uq20 gnd read_bl_0_40 read_bl_1_40 write_bl_0_40 wwl_0_42 rwl_1_42
+ rwl_0_42 cell_2r1w
Xcell_2r1w_2150 vdd_uq11 gnd read_bl_0_30 read_bl_1_30 write_bl_0_30 wwl_0_25 rwl_1_25
+ rwl_0_25 cell_2r1w
Xcell_2r1w_2172 vdd gnd read_bl_0_30 read_bl_1_30 write_bl_0_30 wwl_0_3 rwl_1_3 rwl_0_3
+ cell_2r1w
Xcell_2r1w_1471 vdd_uq0 gnd read_bl_0_41 read_bl_1_41 write_bl_0_41 wwl_0_0 rwl_1_0
+ rwl_0_0 cell_2r1w
Xcell_2r1w_1460 vdd_uq4 gnd read_bl_0_41 read_bl_1_41 write_bl_0_41 wwl_0_11 rwl_1_11
+ rwl_0_11 cell_2r1w
Xcell_2r1w_2161 vdd_uq6 gnd read_bl_0_30 read_bl_1_30 write_bl_0_30 wwl_0_14 rwl_1_14
+ rwl_0_14 cell_2r1w
Xcell_2r1w_1290 vdd_uq25 gnd read_bl_0_43 read_bl_1_43 write_bl_0_43 wwl_0_53 rwl_1_53
+ rwl_0_53 cell_2r1w
Xcell_2r1w_3609 vdd_uq18 gnd read_bl_0_7 read_bl_1_7 write_bl_0_7 wwl_0_38 rwl_1_38
+ rwl_0_38 cell_2r1w
Xcell_2r1w_2908 vdd_uq16 gnd read_bl_0_18 read_bl_1_18 write_bl_0_18 wwl_0_35 rwl_1_35
+ rwl_0_35 cell_2r1w
Xcell_2r1w_2919 vdd_uq11 gnd read_bl_0_18 read_bl_1_18 write_bl_0_18 wwl_0_24 rwl_1_24
+ rwl_0_24 cell_2r1w
Xcell_2r1w_708 vdd_uq28 gnd read_bl_0_52 read_bl_1_52 write_bl_0_52 wwl_0_59 rwl_1_59
+ rwl_0_59 cell_2r1w
Xcell_2r1w_719 vdd_uq23 gnd read_bl_0_52 read_bl_1_52 write_bl_0_52 wwl_0_48 rwl_1_48
+ rwl_0_48 cell_2r1w
Xcell_2r1w_3406 vdd_uq23 gnd read_bl_0_10 read_bl_1_10 write_bl_0_10 wwl_0_49 rwl_1_49
+ rwl_0_49 cell_2r1w
Xcell_2r1w_2705 vdd_uq22 gnd read_bl_0_21 read_bl_1_21 write_bl_0_21 wwl_0_46 rwl_1_46
+ rwl_0_46 cell_2r1w
Xcell_2r1w_3417 vdd_uq18 gnd read_bl_0_10 read_bl_1_10 write_bl_0_10 wwl_0_38 rwl_1_38
+ rwl_0_38 cell_2r1w
Xcell_2r1w_2716 vdd_uq16 gnd read_bl_0_21 read_bl_1_21 write_bl_0_21 wwl_0_35 rwl_1_35
+ rwl_0_35 cell_2r1w
Xcell_2r1w_3428 vdd_uq12 gnd read_bl_0_10 read_bl_1_10 write_bl_0_10 wwl_0_27 rwl_1_27
+ rwl_0_27 cell_2r1w
Xcell_2r1w_2727 vdd_uq11 gnd read_bl_0_21 read_bl_1_21 write_bl_0_21 wwl_0_24 rwl_1_24
+ rwl_0_24 cell_2r1w
Xcell_2r1w_2749 vdd gnd read_bl_0_21 read_bl_1_21 write_bl_0_21 wwl_0_2 rwl_1_2 rwl_0_2
+ cell_2r1w
Xcell_2r1w_2738 vdd_uq5 gnd read_bl_0_21 read_bl_1_21 write_bl_0_21 wwl_0_13 rwl_1_13
+ rwl_0_13 cell_2r1w
Xcell_2r1w_3439 vdd_uq7 gnd read_bl_0_10 read_bl_1_10 write_bl_0_10 wwl_0_16 rwl_1_16
+ rwl_0_16 cell_2r1w
Xcell_2r1w_3973 vdd_uq28 gnd read_bl_0_1 read_bl_1_1 write_bl_0_1 wwl_0_58 rwl_1_58
+ rwl_0_58 cell_2r1w
Xcell_2r1w_3984 vdd_uq22 gnd read_bl_0_1 read_bl_1_1 write_bl_0_1 wwl_0_47 rwl_1_47
+ rwl_0_47 cell_2r1w
Xcell_2r1w_3995 vdd_uq17 gnd read_bl_0_1 read_bl_1_1 write_bl_0_1 wwl_0_36 rwl_1_36
+ rwl_0_36 cell_2r1w
Xcell_2r1w_3940 vdd_uq12 gnd read_bl_0_2 read_bl_1_2 write_bl_0_2 wwl_0_27 rwl_1_27
+ rwl_0_27 cell_2r1w
Xcell_2r1w_3962 vdd_uq1 gnd read_bl_0_2 read_bl_1_2 write_bl_0_2 wwl_0_5 rwl_1_5 rwl_0_5
+ cell_2r1w
Xcell_2r1w_3951 vdd_uq7 gnd read_bl_0_2 read_bl_1_2 write_bl_0_2 wwl_0_16 rwl_1_16
+ rwl_0_16 cell_2r1w
Xcell_2r1w_516 vdd_uq28 gnd read_bl_0_55 read_bl_1_55 write_bl_0_55 wwl_0_59 rwl_1_59
+ rwl_0_59 cell_2r1w
Xcell_2r1w_527 vdd_uq23 gnd read_bl_0_55 read_bl_1_55 write_bl_0_55 wwl_0_48 rwl_1_48
+ rwl_0_48 cell_2r1w
Xcell_2r1w_538 vdd_uq17 gnd read_bl_0_55 read_bl_1_55 write_bl_0_55 wwl_0_37 rwl_1_37
+ rwl_0_37 cell_2r1w
Xcell_2r1w_549 vdd_uq12 gnd read_bl_0_55 read_bl_1_55 write_bl_0_55 wwl_0_26 rwl_1_26
+ rwl_0_26 cell_2r1w
Xcell_2r1w_505 vdd_uq2 gnd read_bl_0_56 read_bl_1_56 write_bl_0_56 wwl_0_6 rwl_1_6
+ rwl_0_6 cell_2r1w
Xcell_2r1w_3203 vdd_uq29 gnd read_bl_0_13 read_bl_1_13 write_bl_0_13 wwl_0_60 rwl_1_60
+ rwl_0_60 cell_2r1w
Xcell_2r1w_3269 vdd_uq28 gnd read_bl_0_12 read_bl_1_12 write_bl_0_12 wwl_0_58 rwl_1_58
+ rwl_0_58 cell_2r1w
Xcell_2r1w_2502 vdd_uq27 gnd read_bl_0_24 read_bl_1_24 write_bl_0_24 wwl_0_57 rwl_1_57
+ rwl_0_57 cell_2r1w
Xcell_2r1w_2568 vdd_uq26 gnd read_bl_0_23 read_bl_1_23 write_bl_0_23 wwl_0_55 rwl_1_55
+ rwl_0_55 cell_2r1w
Xcell_2r1w_1801 vdd_uq26 gnd read_bl_0_35 read_bl_1_35 write_bl_0_35 wwl_0_54 rwl_1_54
+ rwl_0_54 cell_2r1w
Xcell_2r1w_3214 vdd_uq23 gnd read_bl_0_13 read_bl_1_13 write_bl_0_13 wwl_0_49 rwl_1_49
+ rwl_0_49 cell_2r1w
Xcell_2r1w_2513 vdd_uq22 gnd read_bl_0_24 read_bl_1_24 write_bl_0_24 wwl_0_46 rwl_1_46
+ rwl_0_46 cell_2r1w
Xcell_2r1w_2579 vdd_uq21 gnd read_bl_0_23 read_bl_1_23 write_bl_0_23 wwl_0_44 rwl_1_44
+ rwl_0_44 cell_2r1w
Xcell_2r1w_1812 vdd_uq20 gnd read_bl_0_35 read_bl_1_35 write_bl_0_35 wwl_0_43 rwl_1_43
+ rwl_0_43 cell_2r1w
Xcell_2r1w_3225 vdd_uq18 gnd read_bl_0_13 read_bl_1_13 write_bl_0_13 wwl_0_38 rwl_1_38
+ rwl_0_38 cell_2r1w
Xcell_2r1w_2524 vdd_uq16 gnd read_bl_0_24 read_bl_1_24 write_bl_0_24 wwl_0_35 rwl_1_35
+ rwl_0_35 cell_2r1w
Xcell_2r1w_1823 vdd_uq15 gnd read_bl_0_35 read_bl_1_35 write_bl_0_35 wwl_0_32 rwl_1_32
+ rwl_0_32 cell_2r1w
Xcell_2r1w_3236 vdd_uq12 gnd read_bl_0_13 read_bl_1_13 write_bl_0_13 wwl_0_27 rwl_1_27
+ rwl_0_27 cell_2r1w
Xcell_2r1w_2535 vdd_uq11 gnd read_bl_0_24 read_bl_1_24 write_bl_0_24 wwl_0_24 rwl_1_24
+ rwl_0_24 cell_2r1w
Xcell_2r1w_3258 vdd_uq1 gnd read_bl_0_13 read_bl_1_13 write_bl_0_13 wwl_0_5 rwl_1_5
+ rwl_0_5 cell_2r1w
Xcell_2r1w_2557 vdd gnd read_bl_0_24 read_bl_1_24 write_bl_0_24 wwl_0_2 rwl_1_2 rwl_0_2
+ cell_2r1w
Xcell_2r1w_1845 vdd_uq4 gnd read_bl_0_35 read_bl_1_35 write_bl_0_35 wwl_0_10 rwl_1_10
+ rwl_0_10 cell_2r1w
Xcell_2r1w_2546 vdd_uq5 gnd read_bl_0_24 read_bl_1_24 write_bl_0_24 wwl_0_13 rwl_1_13
+ rwl_0_13 cell_2r1w
Xcell_2r1w_3247 vdd_uq7 gnd read_bl_0_13 read_bl_1_13 write_bl_0_13 wwl_0_16 rwl_1_16
+ rwl_0_16 cell_2r1w
Xcell_2r1w_1834 vdd_uq9 gnd read_bl_0_35 read_bl_1_35 write_bl_0_35 wwl_0_21 rwl_1_21
+ rwl_0_21 cell_2r1w
Xcell_2r1w_1856 vdd_uq30 gnd read_bl_0_34 read_bl_1_34 write_bl_0_34 wwl_0_63 rwl_1_63
+ rwl_0_63 cell_2r1w
Xcell_2r1w_1867 vdd_uq25 gnd read_bl_0_34 read_bl_1_34 write_bl_0_34 wwl_0_52 rwl_1_52
+ rwl_0_52 cell_2r1w
Xcell_2r1w_1878 vdd_uq19 gnd read_bl_0_34 read_bl_1_34 write_bl_0_34 wwl_0_41 rwl_1_41
+ rwl_0_41 cell_2r1w
Xcell_2r1w_1889 vdd_uq14 gnd read_bl_0_34 read_bl_1_34 write_bl_0_34 wwl_0_30 rwl_1_30
+ rwl_0_30 cell_2r1w
Xcell_2r1w_3781 vdd_uq28 gnd read_bl_0_4 read_bl_1_4 write_bl_0_4 wwl_0_58 rwl_1_58
+ rwl_0_58 cell_2r1w
Xcell_2r1w_3792 vdd_uq22 gnd read_bl_0_4 read_bl_1_4 write_bl_0_4 wwl_0_47 rwl_1_47
+ rwl_0_47 cell_2r1w
Xcell_2r1w_3770 vdd_uq1 gnd read_bl_0_5 read_bl_1_5 write_bl_0_5 wwl_0_5 rwl_1_5 rwl_0_5
+ cell_2r1w
Xcell_2r1w_1108 vdd_uq20 gnd read_bl_0_46 read_bl_1_46 write_bl_0_46 wwl_0_43 rwl_1_43
+ rwl_0_43 cell_2r1w
Xcell_2r1w_1119 vdd_uq15 gnd read_bl_0_46 read_bl_1_46 write_bl_0_46 wwl_0_32 rwl_1_32
+ rwl_0_32 cell_2r1w
Xcell_2r1w_302 vdd_uq7 gnd read_bl_0_59 read_bl_1_59 write_bl_0_59 wwl_0_17 rwl_1_17
+ rwl_0_17 cell_2r1w
Xcell_2r1w_324 vdd_uq28 gnd read_bl_0_58 read_bl_1_58 write_bl_0_58 wwl_0_59 rwl_1_59
+ rwl_0_59 cell_2r1w
Xcell_2r1w_335 vdd_uq23 gnd read_bl_0_58 read_bl_1_58 write_bl_0_58 wwl_0_48 rwl_1_48
+ rwl_0_48 cell_2r1w
Xcell_2r1w_346 vdd_uq17 gnd read_bl_0_58 read_bl_1_58 write_bl_0_58 wwl_0_37 rwl_1_37
+ rwl_0_37 cell_2r1w
Xcell_2r1w_357 vdd_uq12 gnd read_bl_0_58 read_bl_1_58 write_bl_0_58 wwl_0_26 rwl_1_26
+ rwl_0_26 cell_2r1w
Xcell_2r1w_379 vdd_uq1 gnd read_bl_0_58 read_bl_1_58 write_bl_0_58 wwl_0_4 rwl_1_4
+ rwl_0_4 cell_2r1w
Xcell_2r1w_313 vdd_uq2 gnd read_bl_0_59 read_bl_1_59 write_bl_0_59 wwl_0_6 rwl_1_6
+ rwl_0_6 cell_2r1w
Xcell_2r1w_368 vdd_uq6 gnd read_bl_0_58 read_bl_1_58 write_bl_0_58 wwl_0_15 rwl_1_15
+ rwl_0_15 cell_2r1w
Xcell_2r1w_3011 vdd_uq29 gnd read_bl_0_16 read_bl_1_16 write_bl_0_16 wwl_0_60 rwl_1_60
+ rwl_0_60 cell_2r1w
Xcell_2r1w_3022 vdd_uq23 gnd read_bl_0_16 read_bl_1_16 write_bl_0_16 wwl_0_49 rwl_1_49
+ rwl_0_49 cell_2r1w
Xcell_2r1w_3033 vdd_uq18 gnd read_bl_0_16 read_bl_1_16 write_bl_0_16 wwl_0_38 rwl_1_38
+ rwl_0_38 cell_2r1w
Xcell_2r1w_3000 vdd_uq2 gnd read_bl_0_17 read_bl_1_17 write_bl_0_17 wwl_0_7 rwl_1_7
+ rwl_0_7 cell_2r1w
Xcell_2r1w_1664 vdd_uq30 gnd read_bl_0_37 read_bl_1_37 write_bl_0_37 wwl_0_63 rwl_1_63
+ rwl_0_63 cell_2r1w
Xcell_2r1w_3077 vdd_uq28 gnd read_bl_0_15 read_bl_1_15 write_bl_0_15 wwl_0_58 rwl_1_58
+ rwl_0_58 cell_2r1w
Xcell_2r1w_2310 vdd_uq27 gnd read_bl_0_27 read_bl_1_27 write_bl_0_27 wwl_0_57 rwl_1_57
+ rwl_0_57 cell_2r1w
Xcell_2r1w_2376 vdd_uq26 gnd read_bl_0_26 read_bl_1_26 write_bl_0_26 wwl_0_55 rwl_1_55
+ rwl_0_55 cell_2r1w
Xcell_2r1w_1675 vdd_uq25 gnd read_bl_0_37 read_bl_1_37 write_bl_0_37 wwl_0_52 rwl_1_52
+ rwl_0_52 cell_2r1w
Xcell_2r1w_3088 vdd_uq22 gnd read_bl_0_15 read_bl_1_15 write_bl_0_15 wwl_0_47 rwl_1_47
+ rwl_0_47 cell_2r1w
Xcell_2r1w_2321 vdd_uq22 gnd read_bl_0_27 read_bl_1_27 write_bl_0_27 wwl_0_46 rwl_1_46
+ rwl_0_46 cell_2r1w
Xcell_2r1w_2387 vdd_uq21 gnd read_bl_0_26 read_bl_1_26 write_bl_0_26 wwl_0_44 rwl_1_44
+ rwl_0_44 cell_2r1w
Xcell_2r1w_1620 vdd_uq20 gnd read_bl_0_38 read_bl_1_38 write_bl_0_38 wwl_0_43 rwl_1_43
+ rwl_0_43 cell_2r1w
Xcell_2r1w_1686 vdd_uq19 gnd read_bl_0_37 read_bl_1_37 write_bl_0_37 wwl_0_41 rwl_1_41
+ rwl_0_41 cell_2r1w
Xcell_2r1w_3099 vdd_uq17 gnd read_bl_0_15 read_bl_1_15 write_bl_0_15 wwl_0_36 rwl_1_36
+ rwl_0_36 cell_2r1w
Xcell_2r1w_2332 vdd_uq16 gnd read_bl_0_27 read_bl_1_27 write_bl_0_27 wwl_0_35 rwl_1_35
+ rwl_0_35 cell_2r1w
Xcell_2r1w_2398 vdd_uq15 gnd read_bl_0_26 read_bl_1_26 write_bl_0_26 wwl_0_33 rwl_1_33
+ rwl_0_33 cell_2r1w
Xcell_2r1w_1631 vdd_uq15 gnd read_bl_0_38 read_bl_1_38 write_bl_0_38 wwl_0_32 rwl_1_32
+ rwl_0_32 cell_2r1w
Xcell_2r1w_1697 vdd_uq14 gnd read_bl_0_37 read_bl_1_37 write_bl_0_37 wwl_0_30 rwl_1_30
+ rwl_0_30 cell_2r1w
Xcell_2r1w_3044 vdd_uq12 gnd read_bl_0_16 read_bl_1_16 write_bl_0_16 wwl_0_27 rwl_1_27
+ rwl_0_27 cell_2r1w
Xcell_2r1w_2343 vdd_uq11 gnd read_bl_0_27 read_bl_1_27 write_bl_0_27 wwl_0_24 rwl_1_24
+ rwl_0_24 cell_2r1w
Xcell_2r1w_3066 vdd_uq1 gnd read_bl_0_16 read_bl_1_16 write_bl_0_16 wwl_0_5 rwl_1_5
+ rwl_0_5 cell_2r1w
Xcell_2r1w_2365 vdd gnd read_bl_0_27 read_bl_1_27 write_bl_0_27 wwl_0_2 rwl_1_2 rwl_0_2
+ cell_2r1w
Xcell_2r1w_1653 vdd_uq4 gnd read_bl_0_38 read_bl_1_38 write_bl_0_38 wwl_0_10 rwl_1_10
+ rwl_0_10 cell_2r1w
Xcell_2r1w_2354 vdd_uq5 gnd read_bl_0_27 read_bl_1_27 write_bl_0_27 wwl_0_13 rwl_1_13
+ rwl_0_13 cell_2r1w
Xcell_2r1w_3055 vdd_uq7 gnd read_bl_0_16 read_bl_1_16 write_bl_0_16 wwl_0_16 rwl_1_16
+ rwl_0_16 cell_2r1w
Xcell_2r1w_1642 vdd_uq9 gnd read_bl_0_38 read_bl_1_38 write_bl_0_38 wwl_0_21 rwl_1_21
+ rwl_0_21 cell_2r1w
Xcell_2r1w_891 vdd_uq1 gnd read_bl_0_50 read_bl_1_50 write_bl_0_50 wwl_0_4 rwl_1_4
+ rwl_0_4 cell_2r1w
Xcell_2r1w_880 vdd_uq6 gnd read_bl_0_50 read_bl_1_50 write_bl_0_50 wwl_0_15 rwl_1_15
+ rwl_0_15 cell_2r1w
Xcell_2r1w_132 vdd_uq28 gnd read_bl_0_61 read_bl_1_61 write_bl_0_61 wwl_0_59 rwl_1_59
+ rwl_0_59 cell_2r1w
Xcell_2r1w_143 vdd_uq23 gnd read_bl_0_61 read_bl_1_61 write_bl_0_61 wwl_0_48 rwl_1_48
+ rwl_0_48 cell_2r1w
Xcell_2r1w_121 vdd_uq2 gnd read_bl_0_62 read_bl_1_62 write_bl_0_62 wwl_0_6 rwl_1_6
+ rwl_0_6 cell_2r1w
Xcell_2r1w_110 vdd_uq7 gnd read_bl_0_62 read_bl_1_62 write_bl_0_62 wwl_0_17 rwl_1_17
+ rwl_0_17 cell_2r1w
Xcell_2r1w_198 vdd_uq27 gnd read_bl_0_60 read_bl_1_60 write_bl_0_60 wwl_0_57 rwl_1_57
+ rwl_0_57 cell_2r1w
Xcell_2r1w_154 vdd_uq17 gnd read_bl_0_61 read_bl_1_61 write_bl_0_61 wwl_0_37 rwl_1_37
+ rwl_0_37 cell_2r1w
Xcell_2r1w_165 vdd_uq12 gnd read_bl_0_61 read_bl_1_61 write_bl_0_61 wwl_0_26 rwl_1_26
+ rwl_0_26 cell_2r1w
Xcell_2r1w_187 vdd_uq1 gnd read_bl_0_61 read_bl_1_61 write_bl_0_61 wwl_0_4 rwl_1_4
+ rwl_0_4 cell_2r1w
Xcell_2r1w_176 vdd_uq6 gnd read_bl_0_61 read_bl_1_61 write_bl_0_61 wwl_0_15 rwl_1_15
+ rwl_0_15 cell_2r1w
Xcell_2r1w_2140 vdd_uq16 gnd read_bl_0_30 read_bl_1_30 write_bl_0_30 wwl_0_35 rwl_1_35
+ rwl_0_35 cell_2r1w
Xcell_2r1w_1472 vdd_uq30 gnd read_bl_0_40 read_bl_1_40 write_bl_0_40 wwl_0_63 rwl_1_63
+ rwl_0_63 cell_2r1w
Xcell_2r1w_2184 vdd_uq26 gnd read_bl_0_29 read_bl_1_29 write_bl_0_29 wwl_0_55 rwl_1_55
+ rwl_0_55 cell_2r1w
Xcell_2r1w_1483 vdd_uq25 gnd read_bl_0_40 read_bl_1_40 write_bl_0_40 wwl_0_52 rwl_1_52
+ rwl_0_52 cell_2r1w
Xcell_2r1w_2195 vdd_uq21 gnd read_bl_0_29 read_bl_1_29 write_bl_0_29 wwl_0_44 rwl_1_44
+ rwl_0_44 cell_2r1w
Xcell_2r1w_1494 vdd_uq19 gnd read_bl_0_40 read_bl_1_40 write_bl_0_40 wwl_0_41 rwl_1_41
+ rwl_0_41 cell_2r1w
Xcell_2r1w_2151 vdd_uq11 gnd read_bl_0_30 read_bl_1_30 write_bl_0_30 wwl_0_24 rwl_1_24
+ rwl_0_24 cell_2r1w
Xcell_2r1w_2173 vdd gnd read_bl_0_30 read_bl_1_30 write_bl_0_30 wwl_0_2 rwl_1_2 rwl_0_2
+ cell_2r1w
Xcell_2r1w_1461 vdd_uq4 gnd read_bl_0_41 read_bl_1_41 write_bl_0_41 wwl_0_10 rwl_1_10
+ rwl_0_10 cell_2r1w
Xcell_2r1w_2162 vdd_uq5 gnd read_bl_0_30 read_bl_1_30 write_bl_0_30 wwl_0_13 rwl_1_13
+ rwl_0_13 cell_2r1w
Xcell_2r1w_1450 vdd_uq9 gnd read_bl_0_41 read_bl_1_41 write_bl_0_41 wwl_0_21 rwl_1_21
+ rwl_0_21 cell_2r1w
Xcell_2r1w_1280 vdd_uq30 gnd read_bl_0_43 read_bl_1_43 write_bl_0_43 wwl_0_63 rwl_1_63
+ rwl_0_63 cell_2r1w
Xcell_2r1w_1291 vdd_uq25 gnd read_bl_0_43 read_bl_1_43 write_bl_0_43 wwl_0_52 rwl_1_52
+ rwl_0_52 cell_2r1w
Xcell_2r1w_2909 vdd_uq16 gnd read_bl_0_18 read_bl_1_18 write_bl_0_18 wwl_0_34 rwl_1_34
+ rwl_0_34 cell_2r1w
Xcell_2r1w_709 vdd_uq28 gnd read_bl_0_52 read_bl_1_52 write_bl_0_52 wwl_0_58 rwl_1_58
+ rwl_0_58 cell_2r1w
Xcell_2r1w_3407 vdd_uq23 gnd read_bl_0_10 read_bl_1_10 write_bl_0_10 wwl_0_48 rwl_1_48
+ rwl_0_48 cell_2r1w
Xcell_2r1w_2706 vdd_uq21 gnd read_bl_0_21 read_bl_1_21 write_bl_0_21 wwl_0_45 rwl_1_45
+ rwl_0_45 cell_2r1w
Xcell_2r1w_3418 vdd_uq17 gnd read_bl_0_10 read_bl_1_10 write_bl_0_10 wwl_0_37 rwl_1_37
+ rwl_0_37 cell_2r1w
Xcell_2r1w_2717 vdd_uq16 gnd read_bl_0_21 read_bl_1_21 write_bl_0_21 wwl_0_34 rwl_1_34
+ rwl_0_34 cell_2r1w
Xcell_2r1w_3429 vdd_uq12 gnd read_bl_0_10 read_bl_1_10 write_bl_0_10 wwl_0_26 rwl_1_26
+ rwl_0_26 cell_2r1w
Xcell_2r1w_2739 vdd_uq5 gnd read_bl_0_21 read_bl_1_21 write_bl_0_21 wwl_0_12 rwl_1_12
+ rwl_0_12 cell_2r1w
Xcell_2r1w_2728 vdd_uq10 gnd read_bl_0_21 read_bl_1_21 write_bl_0_21 wwl_0_23 rwl_1_23
+ rwl_0_23 cell_2r1w
Xcell_2r1w_3930 vdd_uq17 gnd read_bl_0_2 read_bl_1_2 write_bl_0_2 wwl_0_37 rwl_1_37
+ rwl_0_37 cell_2r1w
Xcell_2r1w_3974 vdd_uq27 gnd read_bl_0_1 read_bl_1_1 write_bl_0_1 wwl_0_57 rwl_1_57
+ rwl_0_57 cell_2r1w
Xcell_2r1w_3985 vdd_uq22 gnd read_bl_0_1 read_bl_1_1 write_bl_0_1 wwl_0_46 rwl_1_46
+ rwl_0_46 cell_2r1w
Xcell_2r1w_3996 vdd_uq16 gnd read_bl_0_1 read_bl_1_1 write_bl_0_1 wwl_0_35 rwl_1_35
+ rwl_0_35 cell_2r1w
Xcell_2r1w_3941 vdd_uq12 gnd read_bl_0_2 read_bl_1_2 write_bl_0_2 wwl_0_26 rwl_1_26
+ rwl_0_26 cell_2r1w
Xcell_2r1w_3963 vdd_uq1 gnd read_bl_0_2 read_bl_1_2 write_bl_0_2 wwl_0_4 rwl_1_4 rwl_0_4
+ cell_2r1w
Xcell_2r1w_3952 vdd_uq6 gnd read_bl_0_2 read_bl_1_2 write_bl_0_2 wwl_0_15 rwl_1_15
+ rwl_0_15 cell_2r1w
Xcell_2r1w_517 vdd_uq28 gnd read_bl_0_55 read_bl_1_55 write_bl_0_55 wwl_0_58 rwl_1_58
+ rwl_0_58 cell_2r1w
Xcell_2r1w_528 vdd_uq22 gnd read_bl_0_55 read_bl_1_55 write_bl_0_55 wwl_0_47 rwl_1_47
+ rwl_0_47 cell_2r1w
Xcell_2r1w_539 vdd_uq17 gnd read_bl_0_55 read_bl_1_55 write_bl_0_55 wwl_0_36 rwl_1_36
+ rwl_0_36 cell_2r1w
Xcell_2r1w_506 vdd_uq1 gnd read_bl_0_56 read_bl_1_56 write_bl_0_56 wwl_0_5 rwl_1_5
+ rwl_0_5 cell_2r1w
Xcell_2r1w_3204 vdd_uq28 gnd read_bl_0_13 read_bl_1_13 write_bl_0_13 wwl_0_59 rwl_1_59
+ rwl_0_59 cell_2r1w
Xcell_2r1w_3215 vdd_uq23 gnd read_bl_0_13 read_bl_1_13 write_bl_0_13 wwl_0_48 rwl_1_48
+ rwl_0_48 cell_2r1w
Xcell_2r1w_3226 vdd_uq17 gnd read_bl_0_13 read_bl_1_13 write_bl_0_13 wwl_0_37 rwl_1_37
+ rwl_0_37 cell_2r1w
Xcell_2r1w_1857 vdd_uq30 gnd read_bl_0_34 read_bl_1_34 write_bl_0_34 wwl_0_62 rwl_1_62
+ rwl_0_62 cell_2r1w
Xcell_2r1w_2503 vdd_uq27 gnd read_bl_0_24 read_bl_1_24 write_bl_0_24 wwl_0_56 rwl_1_56
+ rwl_0_56 cell_2r1w
Xcell_2r1w_2569 vdd_uq26 gnd read_bl_0_23 read_bl_1_23 write_bl_0_23 wwl_0_54 rwl_1_54
+ rwl_0_54 cell_2r1w
Xcell_2r1w_1802 vdd_uq25 gnd read_bl_0_35 read_bl_1_35 write_bl_0_35 wwl_0_53 rwl_1_53
+ rwl_0_53 cell_2r1w
Xcell_2r1w_1868 vdd_uq24 gnd read_bl_0_34 read_bl_1_34 write_bl_0_34 wwl_0_51 rwl_1_51
+ rwl_0_51 cell_2r1w
Xcell_2r1w_2514 vdd_uq21 gnd read_bl_0_24 read_bl_1_24 write_bl_0_24 wwl_0_45 rwl_1_45
+ rwl_0_45 cell_2r1w
Xcell_2r1w_1813 vdd_uq20 gnd read_bl_0_35 read_bl_1_35 write_bl_0_35 wwl_0_42 rwl_1_42
+ rwl_0_42 cell_2r1w
Xcell_2r1w_1879 vdd_uq19 gnd read_bl_0_34 read_bl_1_34 write_bl_0_34 wwl_0_40 rwl_1_40
+ rwl_0_40 cell_2r1w
Xcell_2r1w_2525 vdd_uq16 gnd read_bl_0_24 read_bl_1_24 write_bl_0_24 wwl_0_34 rwl_1_34
+ rwl_0_34 cell_2r1w
Xcell_2r1w_1824 vdd_uq14 gnd read_bl_0_35 read_bl_1_35 write_bl_0_35 wwl_0_31 rwl_1_31
+ rwl_0_31 cell_2r1w
Xcell_2r1w_3237 vdd_uq12 gnd read_bl_0_13 read_bl_1_13 write_bl_0_13 wwl_0_26 rwl_1_26
+ rwl_0_26 cell_2r1w
Xcell_2r1w_3259 vdd_uq1 gnd read_bl_0_13 read_bl_1_13 write_bl_0_13 wwl_0_4 rwl_1_4
+ rwl_0_4 cell_2r1w
Xcell_2r1w_2558 vdd_uq0 gnd read_bl_0_24 read_bl_1_24 write_bl_0_24 wwl_0_1 rwl_1_1
+ rwl_0_1 cell_2r1w
Xcell_2r1w_1846 vdd_uq3 gnd read_bl_0_35 read_bl_1_35 write_bl_0_35 wwl_0_9 rwl_1_9
+ rwl_0_9 cell_2r1w
Xcell_2r1w_2547 vdd_uq5 gnd read_bl_0_24 read_bl_1_24 write_bl_0_24 wwl_0_12 rwl_1_12
+ rwl_0_12 cell_2r1w
Xcell_2r1w_3248 vdd_uq6 gnd read_bl_0_13 read_bl_1_13 write_bl_0_13 wwl_0_15 rwl_1_15
+ rwl_0_15 cell_2r1w
Xcell_2r1w_1835 vdd_uq9 gnd read_bl_0_35 read_bl_1_35 write_bl_0_35 wwl_0_20 rwl_1_20
+ rwl_0_20 cell_2r1w
Xcell_2r1w_2536 vdd_uq10 gnd read_bl_0_24 read_bl_1_24 write_bl_0_24 wwl_0_23 rwl_1_23
+ rwl_0_23 cell_2r1w
Xcell_2r1w_3771 vdd_uq1 gnd read_bl_0_5 read_bl_1_5 write_bl_0_5 wwl_0_4 rwl_1_4 rwl_0_4
+ cell_2r1w
Xcell_2r1w_3760 vdd_uq6 gnd read_bl_0_5 read_bl_1_5 write_bl_0_5 wwl_0_15 rwl_1_15
+ rwl_0_15 cell_2r1w
Xcell_2r1w_3782 vdd_uq27 gnd read_bl_0_4 read_bl_1_4 write_bl_0_4 wwl_0_57 rwl_1_57
+ rwl_0_57 cell_2r1w
Xcell_2r1w_3793 vdd_uq22 gnd read_bl_0_4 read_bl_1_4 write_bl_0_4 wwl_0_46 rwl_1_46
+ rwl_0_46 cell_2r1w
Xcell_2r1w_325 vdd_uq28 gnd read_bl_0_58 read_bl_1_58 write_bl_0_58 wwl_0_58 rwl_1_58
+ rwl_0_58 cell_2r1w
Xcell_2r1w_336 vdd_uq22 gnd read_bl_0_58 read_bl_1_58 write_bl_0_58 wwl_0_47 rwl_1_47
+ rwl_0_47 cell_2r1w
Xcell_2r1w_1109 vdd_uq20 gnd read_bl_0_46 read_bl_1_46 write_bl_0_46 wwl_0_42 rwl_1_42
+ rwl_0_42 cell_2r1w
Xcell_2r1w_314 vdd_uq1 gnd read_bl_0_59 read_bl_1_59 write_bl_0_59 wwl_0_5 rwl_1_5
+ rwl_0_5 cell_2r1w
Xcell_2r1w_303 vdd_uq7 gnd read_bl_0_59 read_bl_1_59 write_bl_0_59 wwl_0_16 rwl_1_16
+ rwl_0_16 cell_2r1w
Xcell_2r1w_347 vdd_uq17 gnd read_bl_0_58 read_bl_1_58 write_bl_0_58 wwl_0_36 rwl_1_36
+ rwl_0_36 cell_2r1w
Xcell_2r1w_358 vdd_uq11 gnd read_bl_0_58 read_bl_1_58 write_bl_0_58 wwl_0_25 rwl_1_25
+ rwl_0_25 cell_2r1w
Xcell_2r1w_369 vdd_uq6 gnd read_bl_0_58 read_bl_1_58 write_bl_0_58 wwl_0_14 rwl_1_14
+ rwl_0_14 cell_2r1w
Xcell_2r1w_3012 vdd_uq28 gnd read_bl_0_16 read_bl_1_16 write_bl_0_16 wwl_0_59 rwl_1_59
+ rwl_0_59 cell_2r1w
Xcell_2r1w_2311 vdd_uq27 gnd read_bl_0_27 read_bl_1_27 write_bl_0_27 wwl_0_56 rwl_1_56
+ rwl_0_56 cell_2r1w
Xcell_2r1w_3023 vdd_uq23 gnd read_bl_0_16 read_bl_1_16 write_bl_0_16 wwl_0_48 rwl_1_48
+ rwl_0_48 cell_2r1w
Xcell_2r1w_2322 vdd_uq21 gnd read_bl_0_27 read_bl_1_27 write_bl_0_27 wwl_0_45 rwl_1_45
+ rwl_0_45 cell_2r1w
Xcell_2r1w_3034 vdd_uq17 gnd read_bl_0_16 read_bl_1_16 write_bl_0_16 wwl_0_37 rwl_1_37
+ rwl_0_37 cell_2r1w
Xcell_2r1w_3045 vdd_uq12 gnd read_bl_0_16 read_bl_1_16 write_bl_0_16 wwl_0_26 rwl_1_26
+ rwl_0_26 cell_2r1w
Xcell_2r1w_3067 vdd_uq1 gnd read_bl_0_16 read_bl_1_16 write_bl_0_16 wwl_0_4 rwl_1_4
+ rwl_0_4 cell_2r1w
Xcell_2r1w_2300 vdd gnd read_bl_0_28 read_bl_1_28 write_bl_0_28 wwl_0_3 rwl_1_3 rwl_0_3
+ cell_2r1w
Xcell_2r1w_3001 vdd_uq2 gnd read_bl_0_17 read_bl_1_17 write_bl_0_17 wwl_0_6 rwl_1_6
+ rwl_0_6 cell_2r1w
Xcell_2r1w_3056 vdd_uq6 gnd read_bl_0_16 read_bl_1_16 write_bl_0_16 wwl_0_15 rwl_1_15
+ rwl_0_15 cell_2r1w
Xcell_2r1w_1665 vdd_uq30 gnd read_bl_0_37 read_bl_1_37 write_bl_0_37 wwl_0_62 rwl_1_62
+ rwl_0_62 cell_2r1w
Xcell_2r1w_3078 vdd_uq27 gnd read_bl_0_15 read_bl_1_15 write_bl_0_15 wwl_0_57 rwl_1_57
+ rwl_0_57 cell_2r1w
Xcell_2r1w_2377 vdd_uq26 gnd read_bl_0_26 read_bl_1_26 write_bl_0_26 wwl_0_54 rwl_1_54
+ rwl_0_54 cell_2r1w
Xcell_2r1w_1610 vdd_uq25 gnd read_bl_0_38 read_bl_1_38 write_bl_0_38 wwl_0_53 rwl_1_53
+ rwl_0_53 cell_2r1w
Xcell_2r1w_1676 vdd_uq24 gnd read_bl_0_37 read_bl_1_37 write_bl_0_37 wwl_0_51 rwl_1_51
+ rwl_0_51 cell_2r1w
Xcell_2r1w_3089 vdd_uq22 gnd read_bl_0_15 read_bl_1_15 write_bl_0_15 wwl_0_46 rwl_1_46
+ rwl_0_46 cell_2r1w
Xcell_2r1w_2388 vdd_uq20 gnd read_bl_0_26 read_bl_1_26 write_bl_0_26 wwl_0_43 rwl_1_43
+ rwl_0_43 cell_2r1w
Xcell_2r1w_1621 vdd_uq20 gnd read_bl_0_38 read_bl_1_38 write_bl_0_38 wwl_0_42 rwl_1_42
+ rwl_0_42 cell_2r1w
Xcell_2r1w_1687 vdd_uq19 gnd read_bl_0_37 read_bl_1_37 write_bl_0_37 wwl_0_40 rwl_1_40
+ rwl_0_40 cell_2r1w
Xcell_2r1w_2333 vdd_uq16 gnd read_bl_0_27 read_bl_1_27 write_bl_0_27 wwl_0_34 rwl_1_34
+ rwl_0_34 cell_2r1w
Xcell_2r1w_2399 vdd_uq15 gnd read_bl_0_26 read_bl_1_26 write_bl_0_26 wwl_0_32 rwl_1_32
+ rwl_0_32 cell_2r1w
Xcell_2r1w_1632 vdd_uq14 gnd read_bl_0_38 read_bl_1_38 write_bl_0_38 wwl_0_31 rwl_1_31
+ rwl_0_31 cell_2r1w
Xcell_2r1w_1698 vdd_uq13 gnd read_bl_0_37 read_bl_1_37 write_bl_0_37 wwl_0_29 rwl_1_29
+ rwl_0_29 cell_2r1w
Xcell_2r1w_870 vdd_uq11 gnd read_bl_0_50 read_bl_1_50 write_bl_0_50 wwl_0_25 rwl_1_25
+ rwl_0_25 cell_2r1w
Xcell_2r1w_2366 vdd_uq0 gnd read_bl_0_27 read_bl_1_27 write_bl_0_27 wwl_0_1 rwl_1_1
+ rwl_0_1 cell_2r1w
Xcell_2r1w_1654 vdd_uq3 gnd read_bl_0_38 read_bl_1_38 write_bl_0_38 wwl_0_9 rwl_1_9
+ rwl_0_9 cell_2r1w
Xcell_2r1w_2355 vdd_uq5 gnd read_bl_0_27 read_bl_1_27 write_bl_0_27 wwl_0_12 rwl_1_12
+ rwl_0_12 cell_2r1w
Xcell_2r1w_881 vdd_uq6 gnd read_bl_0_50 read_bl_1_50 write_bl_0_50 wwl_0_14 rwl_1_14
+ rwl_0_14 cell_2r1w
Xcell_2r1w_1643 vdd_uq9 gnd read_bl_0_38 read_bl_1_38 write_bl_0_38 wwl_0_20 rwl_1_20
+ rwl_0_20 cell_2r1w
Xcell_2r1w_2344 vdd_uq10 gnd read_bl_0_27 read_bl_1_27 write_bl_0_27 wwl_0_23 rwl_1_23
+ rwl_0_23 cell_2r1w
Xcell_2r1w_892 vdd gnd read_bl_0_50 read_bl_1_50 write_bl_0_50 wwl_0_3 rwl_1_3 rwl_0_3
+ cell_2r1w
Xcell_2r1w_3590 vdd_uq27 gnd read_bl_0_7 read_bl_1_7 write_bl_0_7 wwl_0_57 rwl_1_57
+ rwl_0_57 cell_2r1w
Xcell_2r1w_133 vdd_uq28 gnd read_bl_0_61 read_bl_1_61 write_bl_0_61 wwl_0_58 rwl_1_58
+ rwl_0_58 cell_2r1w
Xcell_2r1w_144 vdd_uq22 gnd read_bl_0_61 read_bl_1_61 write_bl_0_61 wwl_0_47 rwl_1_47
+ rwl_0_47 cell_2r1w
Xcell_2r1w_155 vdd_uq17 gnd read_bl_0_61 read_bl_1_61 write_bl_0_61 wwl_0_36 rwl_1_36
+ rwl_0_36 cell_2r1w
Xcell_2r1w_100 vdd_uq12 gnd read_bl_0_62 read_bl_1_62 write_bl_0_62 wwl_0_27 rwl_1_27
+ rwl_0_27 cell_2r1w
Xcell_2r1w_166 vdd_uq11 gnd read_bl_0_61 read_bl_1_61 write_bl_0_61 wwl_0_25 rwl_1_25
+ rwl_0_25 cell_2r1w
Xcell_2r1w_122 vdd_uq1 gnd read_bl_0_62 read_bl_1_62 write_bl_0_62 wwl_0_5 rwl_1_5
+ rwl_0_5 cell_2r1w
Xcell_2r1w_177 vdd_uq6 gnd read_bl_0_61 read_bl_1_61 write_bl_0_61 wwl_0_14 rwl_1_14
+ rwl_0_14 cell_2r1w
Xcell_2r1w_111 vdd_uq7 gnd read_bl_0_62 read_bl_1_62 write_bl_0_62 wwl_0_16 rwl_1_16
+ rwl_0_16 cell_2r1w
Xcell_2r1w_199 vdd_uq27 gnd read_bl_0_60 read_bl_1_60 write_bl_0_60 wwl_0_56 rwl_1_56
+ rwl_0_56 cell_2r1w
Xcell_2r1w_188 vdd gnd read_bl_0_61 read_bl_1_61 write_bl_0_61 wwl_0_3 rwl_1_3 rwl_0_3
+ cell_2r1w
Xcell_2r1w_2130 vdd_uq21 gnd read_bl_0_30 read_bl_1_30 write_bl_0_30 wwl_0_45 rwl_1_45
+ rwl_0_45 cell_2r1w
Xcell_2r1w_2141 vdd_uq16 gnd read_bl_0_30 read_bl_1_30 write_bl_0_30 wwl_0_34 rwl_1_34
+ rwl_0_34 cell_2r1w
Xcell_2r1w_2174 vdd_uq0 gnd read_bl_0_30 read_bl_1_30 write_bl_0_30 wwl_0_1 rwl_1_1
+ rwl_0_1 cell_2r1w
Xcell_2r1w_2163 vdd_uq5 gnd read_bl_0_30 read_bl_1_30 write_bl_0_30 wwl_0_12 rwl_1_12
+ rwl_0_12 cell_2r1w
Xcell_2r1w_2152 vdd_uq10 gnd read_bl_0_30 read_bl_1_30 write_bl_0_30 wwl_0_23 rwl_1_23
+ rwl_0_23 cell_2r1w
Xcell_2r1w_1473 vdd_uq30 gnd read_bl_0_40 read_bl_1_40 write_bl_0_40 wwl_0_62 rwl_1_62
+ rwl_0_62 cell_2r1w
Xcell_2r1w_2185 vdd_uq26 gnd read_bl_0_29 read_bl_1_29 write_bl_0_29 wwl_0_54 rwl_1_54
+ rwl_0_54 cell_2r1w
Xcell_2r1w_1484 vdd_uq24 gnd read_bl_0_40 read_bl_1_40 write_bl_0_40 wwl_0_51 rwl_1_51
+ rwl_0_51 cell_2r1w
Xcell_2r1w_2196 vdd_uq20 gnd read_bl_0_29 read_bl_1_29 write_bl_0_29 wwl_0_43 rwl_1_43
+ rwl_0_43 cell_2r1w
Xcell_2r1w_1495 vdd_uq19 gnd read_bl_0_40 read_bl_1_40 write_bl_0_40 wwl_0_40 rwl_1_40
+ rwl_0_40 cell_2r1w
Xcell_2r1w_1440 vdd_uq14 gnd read_bl_0_41 read_bl_1_41 write_bl_0_41 wwl_0_31 rwl_1_31
+ rwl_0_31 cell_2r1w
Xcell_2r1w_1462 vdd_uq3 gnd read_bl_0_41 read_bl_1_41 write_bl_0_41 wwl_0_9 rwl_1_9
+ rwl_0_9 cell_2r1w
Xcell_2r1w_1451 vdd_uq9 gnd read_bl_0_41 read_bl_1_41 write_bl_0_41 wwl_0_20 rwl_1_20
+ rwl_0_20 cell_2r1w
Xcell_2r1w_1270 vdd_uq3 gnd read_bl_0_44 read_bl_1_44 write_bl_0_44 wwl_0_9 rwl_1_9
+ rwl_0_9 cell_2r1w
Xcell_2r1w_1281 vdd_uq30 gnd read_bl_0_43 read_bl_1_43 write_bl_0_43 wwl_0_62 rwl_1_62
+ rwl_0_62 cell_2r1w
Xcell_2r1w_1292 vdd_uq24 gnd read_bl_0_43 read_bl_1_43 write_bl_0_43 wwl_0_51 rwl_1_51
+ rwl_0_51 cell_2r1w
Xcell_2r1w_3408 vdd_uq22 gnd read_bl_0_10 read_bl_1_10 write_bl_0_10 wwl_0_47 rwl_1_47
+ rwl_0_47 cell_2r1w
Xcell_2r1w_2707 vdd_uq21 gnd read_bl_0_21 read_bl_1_21 write_bl_0_21 wwl_0_44 rwl_1_44
+ rwl_0_44 cell_2r1w
Xcell_2r1w_3419 vdd_uq17 gnd read_bl_0_10 read_bl_1_10 write_bl_0_10 wwl_0_36 rwl_1_36
+ rwl_0_36 cell_2r1w
Xcell_2r1w_2718 vdd_uq15 gnd read_bl_0_21 read_bl_1_21 write_bl_0_21 wwl_0_33 rwl_1_33
+ rwl_0_33 cell_2r1w
Xcell_2r1w_2729 vdd_uq10 gnd read_bl_0_21 read_bl_1_21 write_bl_0_21 wwl_0_22 rwl_1_22
+ rwl_0_22 cell_2r1w
Xcell_2r1w_3920 vdd_uq22 gnd read_bl_0_2 read_bl_1_2 write_bl_0_2 wwl_0_47 rwl_1_47
+ rwl_0_47 cell_2r1w
Xcell_2r1w_3931 vdd_uq17 gnd read_bl_0_2 read_bl_1_2 write_bl_0_2 wwl_0_36 rwl_1_36
+ rwl_0_36 cell_2r1w
Xcell_2r1w_3942 vdd_uq11 gnd read_bl_0_2 read_bl_1_2 write_bl_0_2 wwl_0_25 rwl_1_25
+ rwl_0_25 cell_2r1w
Xcell_2r1w_3964 vdd gnd read_bl_0_2 read_bl_1_2 write_bl_0_2 wwl_0_3 rwl_1_3 rwl_0_3
+ cell_2r1w
Xcell_2r1w_3953 vdd_uq6 gnd read_bl_0_2 read_bl_1_2 write_bl_0_2 wwl_0_14 rwl_1_14
+ rwl_0_14 cell_2r1w
Xcell_2r1w_3975 vdd_uq27 gnd read_bl_0_1 read_bl_1_1 write_bl_0_1 wwl_0_56 rwl_1_56
+ rwl_0_56 cell_2r1w
Xcell_2r1w_3986 vdd_uq21 gnd read_bl_0_1 read_bl_1_1 write_bl_0_1 wwl_0_45 rwl_1_45
+ rwl_0_45 cell_2r1w
Xcell_2r1w_3997 vdd_uq16 gnd read_bl_0_1 read_bl_1_1 write_bl_0_1 wwl_0_34 rwl_1_34
+ rwl_0_34 cell_2r1w
Xcell_2r1w_518 vdd_uq27 gnd read_bl_0_55 read_bl_1_55 write_bl_0_55 wwl_0_57 rwl_1_57
+ rwl_0_57 cell_2r1w
Xcell_2r1w_507 vdd_uq1 gnd read_bl_0_56 read_bl_1_56 write_bl_0_56 wwl_0_4 rwl_1_4
+ rwl_0_4 cell_2r1w
Xcell_2r1w_529 vdd_uq22 gnd read_bl_0_55 read_bl_1_55 write_bl_0_55 wwl_0_46 rwl_1_46
+ rwl_0_46 cell_2r1w
Xcell_2r1w_3205 vdd_uq28 gnd read_bl_0_13 read_bl_1_13 write_bl_0_13 wwl_0_58 rwl_1_58
+ rwl_0_58 cell_2r1w
Xcell_2r1w_2504 vdd_uq26 gnd read_bl_0_24 read_bl_1_24 write_bl_0_24 wwl_0_55 rwl_1_55
+ rwl_0_55 cell_2r1w
Xcell_2r1w_3216 vdd_uq22 gnd read_bl_0_13 read_bl_1_13 write_bl_0_13 wwl_0_47 rwl_1_47
+ rwl_0_47 cell_2r1w
Xcell_2r1w_2515 vdd_uq21 gnd read_bl_0_24 read_bl_1_24 write_bl_0_24 wwl_0_44 rwl_1_44
+ rwl_0_44 cell_2r1w
Xcell_2r1w_3227 vdd_uq17 gnd read_bl_0_13 read_bl_1_13 write_bl_0_13 wwl_0_36 rwl_1_36
+ rwl_0_36 cell_2r1w
Xcell_2r1w_3238 vdd_uq11 gnd read_bl_0_13 read_bl_1_13 write_bl_0_13 wwl_0_25 rwl_1_25
+ rwl_0_25 cell_2r1w
Xcell_2r1w_3249 vdd_uq6 gnd read_bl_0_13 read_bl_1_13 write_bl_0_13 wwl_0_14 rwl_1_14
+ rwl_0_14 cell_2r1w
Xcell_2r1w_1858 vdd_uq29 gnd read_bl_0_34 read_bl_1_34 write_bl_0_34 wwl_0_61 rwl_1_61
+ rwl_0_61 cell_2r1w
Xcell_2r1w_1803 vdd_uq25 gnd read_bl_0_35 read_bl_1_35 write_bl_0_35 wwl_0_52 rwl_1_52
+ rwl_0_52 cell_2r1w
Xcell_2r1w_1869 vdd_uq24 gnd read_bl_0_34 read_bl_1_34 write_bl_0_34 wwl_0_50 rwl_1_50
+ rwl_0_50 cell_2r1w
Xcell_2r1w_1814 vdd_uq19 gnd read_bl_0_35 read_bl_1_35 write_bl_0_35 wwl_0_41 rwl_1_41
+ rwl_0_41 cell_2r1w
Xcell_2r1w_2526 vdd_uq15 gnd read_bl_0_24 read_bl_1_24 write_bl_0_24 wwl_0_33 rwl_1_33
+ rwl_0_33 cell_2r1w
Xcell_2r1w_1825 vdd_uq14 gnd read_bl_0_35 read_bl_1_35 write_bl_0_35 wwl_0_30 rwl_1_30
+ rwl_0_30 cell_2r1w
Xcell_2r1w_2559 vdd_uq0 gnd read_bl_0_24 read_bl_1_24 write_bl_0_24 wwl_0_0 rwl_1_0
+ rwl_0_0 cell_2r1w
Xcell_2r1w_1847 vdd_uq3 gnd read_bl_0_35 read_bl_1_35 write_bl_0_35 wwl_0_8 rwl_1_8
+ rwl_0_8 cell_2r1w
Xcell_2r1w_2548 vdd_uq4 gnd read_bl_0_24 read_bl_1_24 write_bl_0_24 wwl_0_11 rwl_1_11
+ rwl_0_11 cell_2r1w
Xcell_2r1w_1836 vdd_uq8 gnd read_bl_0_35 read_bl_1_35 write_bl_0_35 wwl_0_19 rwl_1_19
+ rwl_0_19 cell_2r1w
Xcell_2r1w_2537 vdd_uq10 gnd read_bl_0_24 read_bl_1_24 write_bl_0_24 wwl_0_22 rwl_1_22
+ rwl_0_22 cell_2r1w
Xcell_2r1w_3783 vdd_uq27 gnd read_bl_0_4 read_bl_1_4 write_bl_0_4 wwl_0_56 rwl_1_56
+ rwl_0_56 cell_2r1w
Xcell_2r1w_3794 vdd_uq21 gnd read_bl_0_4 read_bl_1_4 write_bl_0_4 wwl_0_45 rwl_1_45
+ rwl_0_45 cell_2r1w
Xcell_2r1w_3750 vdd_uq11 gnd read_bl_0_5 read_bl_1_5 write_bl_0_5 wwl_0_25 rwl_1_25
+ rwl_0_25 cell_2r1w
Xcell_2r1w_3772 vdd gnd read_bl_0_5 read_bl_1_5 write_bl_0_5 wwl_0_3 rwl_1_3 rwl_0_3
+ cell_2r1w
Xcell_2r1w_3761 vdd_uq6 gnd read_bl_0_5 read_bl_1_5 write_bl_0_5 wwl_0_14 rwl_1_14
+ rwl_0_14 cell_2r1w
Xcell_2r1w_326 vdd_uq27 gnd read_bl_0_58 read_bl_1_58 write_bl_0_58 wwl_0_57 rwl_1_57
+ rwl_0_57 cell_2r1w
Xcell_2r1w_337 vdd_uq22 gnd read_bl_0_58 read_bl_1_58 write_bl_0_58 wwl_0_46 rwl_1_46
+ rwl_0_46 cell_2r1w
Xcell_2r1w_348 vdd_uq16 gnd read_bl_0_58 read_bl_1_58 write_bl_0_58 wwl_0_35 rwl_1_35
+ rwl_0_35 cell_2r1w
Xcell_2r1w_359 vdd_uq11 gnd read_bl_0_58 read_bl_1_58 write_bl_0_58 wwl_0_24 rwl_1_24
+ rwl_0_24 cell_2r1w
Xcell_2r1w_315 vdd_uq1 gnd read_bl_0_59 read_bl_1_59 write_bl_0_59 wwl_0_4 rwl_1_4
+ rwl_0_4 cell_2r1w
Xcell_2r1w_304 vdd_uq6 gnd read_bl_0_59 read_bl_1_59 write_bl_0_59 wwl_0_15 rwl_1_15
+ rwl_0_15 cell_2r1w
Xcell_2r1w_1600 vdd_uq30 gnd read_bl_0_38 read_bl_1_38 write_bl_0_38 wwl_0_63 rwl_1_63
+ rwl_0_63 cell_2r1w
Xcell_2r1w_3013 vdd_uq28 gnd read_bl_0_16 read_bl_1_16 write_bl_0_16 wwl_0_58 rwl_1_58
+ rwl_0_58 cell_2r1w
Xcell_2r1w_2312 vdd_uq26 gnd read_bl_0_27 read_bl_1_27 write_bl_0_27 wwl_0_55 rwl_1_55
+ rwl_0_55 cell_2r1w
Xcell_2r1w_3079 vdd_uq27 gnd read_bl_0_15 read_bl_1_15 write_bl_0_15 wwl_0_56 rwl_1_56
+ rwl_0_56 cell_2r1w
Xcell_2r1w_1611 vdd_uq25 gnd read_bl_0_38 read_bl_1_38 write_bl_0_38 wwl_0_52 rwl_1_52
+ rwl_0_52 cell_2r1w
Xcell_2r1w_3024 vdd_uq22 gnd read_bl_0_16 read_bl_1_16 write_bl_0_16 wwl_0_47 rwl_1_47
+ rwl_0_47 cell_2r1w
Xcell_2r1w_2323 vdd_uq21 gnd read_bl_0_27 read_bl_1_27 write_bl_0_27 wwl_0_44 rwl_1_44
+ rwl_0_44 cell_2r1w
Xcell_2r1w_3035 vdd_uq17 gnd read_bl_0_16 read_bl_1_16 write_bl_0_16 wwl_0_36 rwl_1_36
+ rwl_0_36 cell_2r1w
Xcell_2r1w_2334 vdd_uq15 gnd read_bl_0_27 read_bl_1_27 write_bl_0_27 wwl_0_33 rwl_1_33
+ rwl_0_33 cell_2r1w
Xcell_2r1w_3046 vdd_uq11 gnd read_bl_0_16 read_bl_1_16 write_bl_0_16 wwl_0_25 rwl_1_25
+ rwl_0_25 cell_2r1w
Xcell_2r1w_3002 vdd_uq1 gnd read_bl_0_17 read_bl_1_17 write_bl_0_17 wwl_0_5 rwl_1_5
+ rwl_0_5 cell_2r1w
Xcell_2r1w_3068 vdd gnd read_bl_0_16 read_bl_1_16 write_bl_0_16 wwl_0_3 rwl_1_3 rwl_0_3
+ cell_2r1w
Xcell_2r1w_2301 vdd gnd read_bl_0_28 read_bl_1_28 write_bl_0_28 wwl_0_2 rwl_1_2 rwl_0_2
+ cell_2r1w
Xcell_2r1w_2356 vdd_uq4 gnd read_bl_0_27 read_bl_1_27 write_bl_0_27 wwl_0_11 rwl_1_11
+ rwl_0_11 cell_2r1w
Xcell_2r1w_3057 vdd_uq6 gnd read_bl_0_16 read_bl_1_16 write_bl_0_16 wwl_0_14 rwl_1_14
+ rwl_0_14 cell_2r1w
Xcell_2r1w_2345 vdd_uq10 gnd read_bl_0_27 read_bl_1_27 write_bl_0_27 wwl_0_22 rwl_1_22
+ rwl_0_22 cell_2r1w
Xcell_2r1w_1666 vdd_uq29 gnd read_bl_0_37 read_bl_1_37 write_bl_0_37 wwl_0_61 rwl_1_61
+ rwl_0_61 cell_2r1w
Xcell_2r1w_2378 vdd_uq25 gnd read_bl_0_26 read_bl_1_26 write_bl_0_26 wwl_0_53 rwl_1_53
+ rwl_0_53 cell_2r1w
Xcell_2r1w_1677 vdd_uq24 gnd read_bl_0_37 read_bl_1_37 write_bl_0_37 wwl_0_50 rwl_1_50
+ rwl_0_50 cell_2r1w
Xcell_2r1w_1622 vdd_uq19 gnd read_bl_0_38 read_bl_1_38 write_bl_0_38 wwl_0_41 rwl_1_41
+ rwl_0_41 cell_2r1w
Xcell_2r1w_2389 vdd_uq20 gnd read_bl_0_26 read_bl_1_26 write_bl_0_26 wwl_0_42 rwl_1_42
+ rwl_0_42 cell_2r1w
Xcell_2r1w_1688 vdd_uq18 gnd read_bl_0_37 read_bl_1_37 write_bl_0_37 wwl_0_39 rwl_1_39
+ rwl_0_39 cell_2r1w
Xcell_2r1w_860 vdd_uq16 gnd read_bl_0_50 read_bl_1_50 write_bl_0_50 wwl_0_35 rwl_1_35
+ rwl_0_35 cell_2r1w
Xcell_2r1w_1633 vdd_uq14 gnd read_bl_0_38 read_bl_1_38 write_bl_0_38 wwl_0_30 rwl_1_30
+ rwl_0_30 cell_2r1w
Xcell_2r1w_1699 vdd_uq13 gnd read_bl_0_37 read_bl_1_37 write_bl_0_37 wwl_0_28 rwl_1_28
+ rwl_0_28 cell_2r1w
Xcell_2r1w_871 vdd_uq11 gnd read_bl_0_50 read_bl_1_50 write_bl_0_50 wwl_0_24 rwl_1_24
+ rwl_0_24 cell_2r1w
Xcell_2r1w_893 vdd gnd read_bl_0_50 read_bl_1_50 write_bl_0_50 wwl_0_2 rwl_1_2 rwl_0_2
+ cell_2r1w
Xcell_2r1w_2367 vdd_uq0 gnd read_bl_0_27 read_bl_1_27 write_bl_0_27 wwl_0_0 rwl_1_0
+ rwl_0_0 cell_2r1w
Xcell_2r1w_1655 vdd_uq3 gnd read_bl_0_38 read_bl_1_38 write_bl_0_38 wwl_0_8 rwl_1_8
+ rwl_0_8 cell_2r1w
Xcell_2r1w_882 vdd_uq5 gnd read_bl_0_50 read_bl_1_50 write_bl_0_50 wwl_0_13 rwl_1_13
+ rwl_0_13 cell_2r1w
Xcell_2r1w_1644 vdd_uq8 gnd read_bl_0_38 read_bl_1_38 write_bl_0_38 wwl_0_19 rwl_1_19
+ rwl_0_19 cell_2r1w
Xcell_2r1w_3591 vdd_uq27 gnd read_bl_0_7 read_bl_1_7 write_bl_0_7 wwl_0_56 rwl_1_56
+ rwl_0_56 cell_2r1w
Xcell_2r1w_2890 vdd_uq25 gnd read_bl_0_18 read_bl_1_18 write_bl_0_18 wwl_0_53 rwl_1_53
+ rwl_0_53 cell_2r1w
Xcell_2r1w_3580 vdd gnd read_bl_0_8 read_bl_1_8 write_bl_0_8 wwl_0_3 rwl_1_3 rwl_0_3
+ cell_2r1w
Xcell_2r1w_134 vdd_uq27 gnd read_bl_0_61 read_bl_1_61 write_bl_0_61 wwl_0_57 rwl_1_57
+ rwl_0_57 cell_2r1w
Xcell_2r1w_145 vdd_uq22 gnd read_bl_0_61 read_bl_1_61 write_bl_0_61 wwl_0_46 rwl_1_46
+ rwl_0_46 cell_2r1w
Xcell_2r1w_156 vdd_uq16 gnd read_bl_0_61 read_bl_1_61 write_bl_0_61 wwl_0_35 rwl_1_35
+ rwl_0_35 cell_2r1w
Xcell_2r1w_101 vdd_uq12 gnd read_bl_0_62 read_bl_1_62 write_bl_0_62 wwl_0_26 rwl_1_26
+ rwl_0_26 cell_2r1w
Xcell_2r1w_167 vdd_uq11 gnd read_bl_0_61 read_bl_1_61 write_bl_0_61 wwl_0_24 rwl_1_24
+ rwl_0_24 cell_2r1w
Xcell_2r1w_123 vdd_uq1 gnd read_bl_0_62 read_bl_1_62 write_bl_0_62 wwl_0_4 rwl_1_4
+ rwl_0_4 cell_2r1w
Xcell_2r1w_189 vdd gnd read_bl_0_61 read_bl_1_61 write_bl_0_61 wwl_0_2 rwl_1_2 rwl_0_2
+ cell_2r1w
Xcell_2r1w_178 vdd_uq5 gnd read_bl_0_61 read_bl_1_61 write_bl_0_61 wwl_0_13 rwl_1_13
+ rwl_0_13 cell_2r1w
Xcell_2r1w_112 vdd_uq6 gnd read_bl_0_62 read_bl_1_62 write_bl_0_62 wwl_0_15 rwl_1_15
+ rwl_0_15 cell_2r1w
Xcell_2r1w_2120 vdd_uq26 gnd read_bl_0_30 read_bl_1_30 write_bl_0_30 wwl_0_55 rwl_1_55
+ rwl_0_55 cell_2r1w
Xcell_2r1w_2186 vdd_uq25 gnd read_bl_0_29 read_bl_1_29 write_bl_0_29 wwl_0_53 rwl_1_53
+ rwl_0_53 cell_2r1w
Xcell_2r1w_2131 vdd_uq21 gnd read_bl_0_30 read_bl_1_30 write_bl_0_30 wwl_0_44 rwl_1_44
+ rwl_0_44 cell_2r1w
Xcell_2r1w_1430 vdd_uq19 gnd read_bl_0_41 read_bl_1_41 write_bl_0_41 wwl_0_41 rwl_1_41
+ rwl_0_41 cell_2r1w
Xcell_2r1w_2197 vdd_uq20 gnd read_bl_0_29 read_bl_1_29 write_bl_0_29 wwl_0_42 rwl_1_42
+ rwl_0_42 cell_2r1w
Xcell_2r1w_2142 vdd_uq15 gnd read_bl_0_30 read_bl_1_30 write_bl_0_30 wwl_0_33 rwl_1_33
+ rwl_0_33 cell_2r1w
Xcell_2r1w_1441 vdd_uq14 gnd read_bl_0_41 read_bl_1_41 write_bl_0_41 wwl_0_30 rwl_1_30
+ rwl_0_30 cell_2r1w
Xcell_2r1w_2175 vdd_uq0 gnd read_bl_0_30 read_bl_1_30 write_bl_0_30 wwl_0_0 rwl_1_0
+ rwl_0_0 cell_2r1w
Xcell_2r1w_1463 vdd_uq3 gnd read_bl_0_41 read_bl_1_41 write_bl_0_41 wwl_0_8 rwl_1_8
+ rwl_0_8 cell_2r1w
Xcell_2r1w_2164 vdd_uq4 gnd read_bl_0_30 read_bl_1_30 write_bl_0_30 wwl_0_11 rwl_1_11
+ rwl_0_11 cell_2r1w
Xcell_2r1w_1452 vdd_uq8 gnd read_bl_0_41 read_bl_1_41 write_bl_0_41 wwl_0_19 rwl_1_19
+ rwl_0_19 cell_2r1w
Xcell_2r1w_2153 vdd_uq10 gnd read_bl_0_30 read_bl_1_30 write_bl_0_30 wwl_0_22 rwl_1_22
+ rwl_0_22 cell_2r1w
Xcell_2r1w_1474 vdd_uq29 gnd read_bl_0_40 read_bl_1_40 write_bl_0_40 wwl_0_61 rwl_1_61
+ rwl_0_61 cell_2r1w
Xcell_2r1w_1485 vdd_uq24 gnd read_bl_0_40 read_bl_1_40 write_bl_0_40 wwl_0_50 rwl_1_50
+ rwl_0_50 cell_2r1w
Xcell_2r1w_1496 vdd_uq18 gnd read_bl_0_40 read_bl_1_40 write_bl_0_40 wwl_0_39 rwl_1_39
+ rwl_0_39 cell_2r1w
Xcell_2r1w_690 vdd_uq5 gnd read_bl_0_53 read_bl_1_53 write_bl_0_53 wwl_0_13 rwl_1_13
+ rwl_0_13 cell_2r1w
Xcell_2r1w_1282 vdd_uq29 gnd read_bl_0_43 read_bl_1_43 write_bl_0_43 wwl_0_61 rwl_1_61
+ rwl_0_61 cell_2r1w
Xcell_2r1w_1293 vdd_uq24 gnd read_bl_0_43 read_bl_1_43 write_bl_0_43 wwl_0_50 rwl_1_50
+ rwl_0_50 cell_2r1w
Xcell_2r1w_1271 vdd_uq3 gnd read_bl_0_44 read_bl_1_44 write_bl_0_44 wwl_0_8 rwl_1_8
+ rwl_0_8 cell_2r1w
Xcell_2r1w_1260 vdd_uq8 gnd read_bl_0_44 read_bl_1_44 write_bl_0_44 wwl_0_19 rwl_1_19
+ rwl_0_19 cell_2r1w
Xcell_2r1w_1090 vdd_uq29 gnd read_bl_0_46 read_bl_1_46 write_bl_0_46 wwl_0_61 rwl_1_61
+ rwl_0_61 cell_2r1w
Xcell_2r1w_3409 vdd_uq22 gnd read_bl_0_10 read_bl_1_10 write_bl_0_10 wwl_0_46 rwl_1_46
+ rwl_0_46 cell_2r1w
Xcell_2r1w_2708 vdd_uq20 gnd read_bl_0_21 read_bl_1_21 write_bl_0_21 wwl_0_43 rwl_1_43
+ rwl_0_43 cell_2r1w
Xcell_2r1w_2719 vdd_uq15 gnd read_bl_0_21 read_bl_1_21 write_bl_0_21 wwl_0_32 rwl_1_32
+ rwl_0_32 cell_2r1w
Xcell_2r1w_3910 vdd_uq27 gnd read_bl_0_2 read_bl_1_2 write_bl_0_2 wwl_0_57 rwl_1_57
+ rwl_0_57 cell_2r1w
Xcell_2r1w_3976 vdd_uq26 gnd read_bl_0_1 read_bl_1_1 write_bl_0_1 wwl_0_55 rwl_1_55
+ rwl_0_55 cell_2r1w
Xcell_2r1w_3921 vdd_uq22 gnd read_bl_0_2 read_bl_1_2 write_bl_0_2 wwl_0_46 rwl_1_46
+ rwl_0_46 cell_2r1w
Xcell_2r1w_3987 vdd_uq21 gnd read_bl_0_1 read_bl_1_1 write_bl_0_1 wwl_0_44 rwl_1_44
+ rwl_0_44 cell_2r1w
Xcell_2r1w_3932 vdd_uq16 gnd read_bl_0_2 read_bl_1_2 write_bl_0_2 wwl_0_35 rwl_1_35
+ rwl_0_35 cell_2r1w
Xcell_2r1w_3943 vdd_uq11 gnd read_bl_0_2 read_bl_1_2 write_bl_0_2 wwl_0_24 rwl_1_24
+ rwl_0_24 cell_2r1w
Xcell_2r1w_3965 vdd gnd read_bl_0_2 read_bl_1_2 write_bl_0_2 wwl_0_2 rwl_1_2 rwl_0_2
+ cell_2r1w
Xcell_2r1w_3954 vdd_uq5 gnd read_bl_0_2 read_bl_1_2 write_bl_0_2 wwl_0_13 rwl_1_13
+ rwl_0_13 cell_2r1w
Xcell_2r1w_3998 vdd_uq15 gnd read_bl_0_1 read_bl_1_1 write_bl_0_1 wwl_0_33 rwl_1_33
+ rwl_0_33 cell_2r1w
Xcell_2r1w_519 vdd_uq27 gnd read_bl_0_55 read_bl_1_55 write_bl_0_55 wwl_0_56 rwl_1_56
+ rwl_0_56 cell_2r1w
Xcell_2r1w_508 vdd gnd read_bl_0_56 read_bl_1_56 write_bl_0_56 wwl_0_3 rwl_1_3 rwl_0_3
+ cell_2r1w
Xcell_2r1w_3206 vdd_uq27 gnd read_bl_0_13 read_bl_1_13 write_bl_0_13 wwl_0_57 rwl_1_57
+ rwl_0_57 cell_2r1w
Xcell_2r1w_2505 vdd_uq26 gnd read_bl_0_24 read_bl_1_24 write_bl_0_24 wwl_0_54 rwl_1_54
+ rwl_0_54 cell_2r1w
Xcell_2r1w_3217 vdd_uq22 gnd read_bl_0_13 read_bl_1_13 write_bl_0_13 wwl_0_46 rwl_1_46
+ rwl_0_46 cell_2r1w
Xcell_2r1w_2516 vdd_uq20 gnd read_bl_0_24 read_bl_1_24 write_bl_0_24 wwl_0_43 rwl_1_43
+ rwl_0_43 cell_2r1w
Xcell_2r1w_3228 vdd_uq16 gnd read_bl_0_13 read_bl_1_13 write_bl_0_13 wwl_0_35 rwl_1_35
+ rwl_0_35 cell_2r1w
Xcell_2r1w_2527 vdd_uq15 gnd read_bl_0_24 read_bl_1_24 write_bl_0_24 wwl_0_32 rwl_1_32
+ rwl_0_32 cell_2r1w
Xcell_2r1w_3239 vdd_uq11 gnd read_bl_0_13 read_bl_1_13 write_bl_0_13 wwl_0_24 rwl_1_24
+ rwl_0_24 cell_2r1w
Xcell_2r1w_2538 vdd_uq9 gnd read_bl_0_24 read_bl_1_24 write_bl_0_24 wwl_0_21 rwl_1_21
+ rwl_0_21 cell_2r1w
Xcell_2r1w_1859 vdd_uq29 gnd read_bl_0_34 read_bl_1_34 write_bl_0_34 wwl_0_60 rwl_1_60
+ rwl_0_60 cell_2r1w
Xcell_2r1w_1804 vdd_uq24 gnd read_bl_0_35 read_bl_1_35 write_bl_0_35 wwl_0_51 rwl_1_51
+ rwl_0_51 cell_2r1w
Xcell_2r1w_1815 vdd_uq19 gnd read_bl_0_35 read_bl_1_35 write_bl_0_35 wwl_0_40 rwl_1_40
+ rwl_0_40 cell_2r1w
Xcell_2r1w_1826 vdd_uq13 gnd read_bl_0_35 read_bl_1_35 write_bl_0_35 wwl_0_29 rwl_1_29
+ rwl_0_29 cell_2r1w
Xcell_2r1w_1848 vdd_uq2 gnd read_bl_0_35 read_bl_1_35 write_bl_0_35 wwl_0_7 rwl_1_7
+ rwl_0_7 cell_2r1w
Xcell_2r1w_2549 vdd_uq4 gnd read_bl_0_24 read_bl_1_24 write_bl_0_24 wwl_0_10 rwl_1_10
+ rwl_0_10 cell_2r1w
Xcell_2r1w_1837 vdd_uq8 gnd read_bl_0_35 read_bl_1_35 write_bl_0_35 wwl_0_18 rwl_1_18
+ rwl_0_18 cell_2r1w
Xcell_2r1w_3784 vdd_uq26 gnd read_bl_0_4 read_bl_1_4 write_bl_0_4 wwl_0_55 rwl_1_55
+ rwl_0_55 cell_2r1w
Xcell_2r1w_3795 vdd_uq21 gnd read_bl_0_4 read_bl_1_4 write_bl_0_4 wwl_0_44 rwl_1_44
+ rwl_0_44 cell_2r1w
Xcell_2r1w_3740 vdd_uq16 gnd read_bl_0_5 read_bl_1_5 write_bl_0_5 wwl_0_35 rwl_1_35
+ rwl_0_35 cell_2r1w
Xcell_2r1w_3751 vdd_uq11 gnd read_bl_0_5 read_bl_1_5 write_bl_0_5 wwl_0_24 rwl_1_24
+ rwl_0_24 cell_2r1w
Xcell_2r1w_3773 vdd gnd read_bl_0_5 read_bl_1_5 write_bl_0_5 wwl_0_2 rwl_1_2 rwl_0_2
+ cell_2r1w
Xcell_2r1w_3762 vdd_uq5 gnd read_bl_0_5 read_bl_1_5 write_bl_0_5 wwl_0_13 rwl_1_13
+ rwl_0_13 cell_2r1w
Xcell_2r1w_327 vdd_uq27 gnd read_bl_0_58 read_bl_1_58 write_bl_0_58 wwl_0_56 rwl_1_56
+ rwl_0_56 cell_2r1w
Xcell_2r1w_338 vdd_uq21 gnd read_bl_0_58 read_bl_1_58 write_bl_0_58 wwl_0_45 rwl_1_45
+ rwl_0_45 cell_2r1w
Xcell_2r1w_349 vdd_uq16 gnd read_bl_0_58 read_bl_1_58 write_bl_0_58 wwl_0_34 rwl_1_34
+ rwl_0_34 cell_2r1w
Xcell_2r1w_316 vdd gnd read_bl_0_59 read_bl_1_59 write_bl_0_59 wwl_0_3 rwl_1_3 rwl_0_3
+ cell_2r1w
Xcell_2r1w_305 vdd_uq6 gnd read_bl_0_59 read_bl_1_59 write_bl_0_59 wwl_0_14 rwl_1_14
+ rwl_0_14 cell_2r1w
Xcell_2r1w_2368 vdd_uq30 gnd read_bl_0_26 read_bl_1_26 write_bl_0_26 wwl_0_63 rwl_1_63
+ rwl_0_63 cell_2r1w
Xcell_2r1w_1601 vdd_uq30 gnd read_bl_0_38 read_bl_1_38 write_bl_0_38 wwl_0_62 rwl_1_62
+ rwl_0_62 cell_2r1w
Xcell_2r1w_3014 vdd_uq27 gnd read_bl_0_16 read_bl_1_16 write_bl_0_16 wwl_0_57 rwl_1_57
+ rwl_0_57 cell_2r1w
Xcell_2r1w_2313 vdd_uq26 gnd read_bl_0_27 read_bl_1_27 write_bl_0_27 wwl_0_54 rwl_1_54
+ rwl_0_54 cell_2r1w
Xcell_2r1w_2379 vdd_uq25 gnd read_bl_0_26 read_bl_1_26 write_bl_0_26 wwl_0_52 rwl_1_52
+ rwl_0_52 cell_2r1w
Xcell_2r1w_1612 vdd_uq24 gnd read_bl_0_38 read_bl_1_38 write_bl_0_38 wwl_0_51 rwl_1_51
+ rwl_0_51 cell_2r1w
Xcell_2r1w_3025 vdd_uq22 gnd read_bl_0_16 read_bl_1_16 write_bl_0_16 wwl_0_46 rwl_1_46
+ rwl_0_46 cell_2r1w
Xcell_2r1w_2324 vdd_uq20 gnd read_bl_0_27 read_bl_1_27 write_bl_0_27 wwl_0_43 rwl_1_43
+ rwl_0_43 cell_2r1w
Xcell_2r1w_1623 vdd_uq19 gnd read_bl_0_38 read_bl_1_38 write_bl_0_38 wwl_0_40 rwl_1_40
+ rwl_0_40 cell_2r1w
Xcell_2r1w_3036 vdd_uq16 gnd read_bl_0_16 read_bl_1_16 write_bl_0_16 wwl_0_35 rwl_1_35
+ rwl_0_35 cell_2r1w
Xcell_2r1w_2335 vdd_uq15 gnd read_bl_0_27 read_bl_1_27 write_bl_0_27 wwl_0_32 rwl_1_32
+ rwl_0_32 cell_2r1w
Xcell_2r1w_1634 vdd_uq13 gnd read_bl_0_38 read_bl_1_38 write_bl_0_38 wwl_0_29 rwl_1_29
+ rwl_0_29 cell_2r1w
Xcell_2r1w_3047 vdd_uq11 gnd read_bl_0_16 read_bl_1_16 write_bl_0_16 wwl_0_24 rwl_1_24
+ rwl_0_24 cell_2r1w
Xcell_2r1w_3003 vdd_uq1 gnd read_bl_0_17 read_bl_1_17 write_bl_0_17 wwl_0_4 rwl_1_4
+ rwl_0_4 cell_2r1w
Xcell_2r1w_3069 vdd gnd read_bl_0_16 read_bl_1_16 write_bl_0_16 wwl_0_2 rwl_1_2 rwl_0_2
+ cell_2r1w
Xcell_2r1w_2302 vdd_uq0 gnd read_bl_0_28 read_bl_1_28 write_bl_0_28 wwl_0_1 rwl_1_1
+ rwl_0_1 cell_2r1w
Xcell_2r1w_2357 vdd_uq4 gnd read_bl_0_27 read_bl_1_27 write_bl_0_27 wwl_0_10 rwl_1_10
+ rwl_0_10 cell_2r1w
Xcell_2r1w_3058 vdd_uq5 gnd read_bl_0_16 read_bl_1_16 write_bl_0_16 wwl_0_13 rwl_1_13
+ rwl_0_13 cell_2r1w
Xcell_2r1w_1645 vdd_uq8 gnd read_bl_0_38 read_bl_1_38 write_bl_0_38 wwl_0_18 rwl_1_18
+ rwl_0_18 cell_2r1w
Xcell_2r1w_2346 vdd_uq9 gnd read_bl_0_27 read_bl_1_27 write_bl_0_27 wwl_0_21 rwl_1_21
+ rwl_0_21 cell_2r1w
Xcell_2r1w_1667 vdd_uq29 gnd read_bl_0_37 read_bl_1_37 write_bl_0_37 wwl_0_60 rwl_1_60
+ rwl_0_60 cell_2r1w
Xcell_2r1w_1678 vdd_uq23 gnd read_bl_0_37 read_bl_1_37 write_bl_0_37 wwl_0_49 rwl_1_49
+ rwl_0_49 cell_2r1w
Xcell_2r1w_850 vdd_uq21 gnd read_bl_0_50 read_bl_1_50 write_bl_0_50 wwl_0_45 rwl_1_45
+ rwl_0_45 cell_2r1w
Xcell_2r1w_1689 vdd_uq18 gnd read_bl_0_37 read_bl_1_37 write_bl_0_37 wwl_0_38 rwl_1_38
+ rwl_0_38 cell_2r1w
Xcell_2r1w_861 vdd_uq16 gnd read_bl_0_50 read_bl_1_50 write_bl_0_50 wwl_0_34 rwl_1_34
+ rwl_0_34 cell_2r1w
Xcell_2r1w_894 vdd_uq0 gnd read_bl_0_50 read_bl_1_50 write_bl_0_50 wwl_0_1 rwl_1_1
+ rwl_0_1 cell_2r1w
Xcell_2r1w_1656 vdd_uq2 gnd read_bl_0_38 read_bl_1_38 write_bl_0_38 wwl_0_7 rwl_1_7
+ rwl_0_7 cell_2r1w
Xcell_2r1w_883 vdd_uq5 gnd read_bl_0_50 read_bl_1_50 write_bl_0_50 wwl_0_12 rwl_1_12
+ rwl_0_12 cell_2r1w
Xcell_2r1w_872 vdd_uq10 gnd read_bl_0_50 read_bl_1_50 write_bl_0_50 wwl_0_23 rwl_1_23
+ rwl_0_23 cell_2r1w
Xcell_2r1w_2880 vdd_uq30 gnd read_bl_0_18 read_bl_1_18 write_bl_0_18 wwl_0_63 rwl_1_63
+ rwl_0_63 cell_2r1w
Xcell_2r1w_3592 vdd_uq26 gnd read_bl_0_7 read_bl_1_7 write_bl_0_7 wwl_0_55 rwl_1_55
+ rwl_0_55 cell_2r1w
Xcell_2r1w_2891 vdd_uq25 gnd read_bl_0_18 read_bl_1_18 write_bl_0_18 wwl_0_52 rwl_1_52
+ rwl_0_52 cell_2r1w
Xcell_2r1w_3581 vdd gnd read_bl_0_8 read_bl_1_8 write_bl_0_8 wwl_0_2 rwl_1_2 rwl_0_2
+ cell_2r1w
Xcell_2r1w_3570 vdd_uq5 gnd read_bl_0_8 read_bl_1_8 write_bl_0_8 wwl_0_13 rwl_1_13
+ rwl_0_13 cell_2r1w
Xcell_2r1w_102 vdd_uq11 gnd read_bl_0_62 read_bl_1_62 write_bl_0_62 wwl_0_25 rwl_1_25
+ rwl_0_25 cell_2r1w
Xcell_2r1w_135 vdd_uq27 gnd read_bl_0_61 read_bl_1_61 write_bl_0_61 wwl_0_56 rwl_1_56
+ rwl_0_56 cell_2r1w
Xcell_2r1w_146 vdd_uq21 gnd read_bl_0_61 read_bl_1_61 write_bl_0_61 wwl_0_45 rwl_1_45
+ rwl_0_45 cell_2r1w
Xcell_2r1w_157 vdd_uq16 gnd read_bl_0_61 read_bl_1_61 write_bl_0_61 wwl_0_34 rwl_1_34
+ rwl_0_34 cell_2r1w
Xcell_2r1w_124 vdd gnd read_bl_0_62 read_bl_1_62 write_bl_0_62 wwl_0_3 rwl_1_3 rwl_0_3
+ cell_2r1w
Xcell_2r1w_179 vdd_uq5 gnd read_bl_0_61 read_bl_1_61 write_bl_0_61 wwl_0_12 rwl_1_12
+ rwl_0_12 cell_2r1w
Xcell_2r1w_113 vdd_uq6 gnd read_bl_0_62 read_bl_1_62 write_bl_0_62 wwl_0_14 rwl_1_14
+ rwl_0_14 cell_2r1w
Xcell_2r1w_168 vdd_uq10 gnd read_bl_0_61 read_bl_1_61 write_bl_0_61 wwl_0_23 rwl_1_23
+ rwl_0_23 cell_2r1w
Xcell_2r1w_2176 vdd_uq30 gnd read_bl_0_29 read_bl_1_29 write_bl_0_29 wwl_0_63 rwl_1_63
+ rwl_0_63 cell_2r1w
Xcell_2r1w_1475 vdd_uq29 gnd read_bl_0_40 read_bl_1_40 write_bl_0_40 wwl_0_60 rwl_1_60
+ rwl_0_60 cell_2r1w
Xcell_2r1w_2121 vdd_uq26 gnd read_bl_0_30 read_bl_1_30 write_bl_0_30 wwl_0_54 rwl_1_54
+ rwl_0_54 cell_2r1w
Xcell_2r1w_2187 vdd_uq25 gnd read_bl_0_29 read_bl_1_29 write_bl_0_29 wwl_0_52 rwl_1_52
+ rwl_0_52 cell_2r1w
Xcell_2r1w_1420 vdd_uq24 gnd read_bl_0_41 read_bl_1_41 write_bl_0_41 wwl_0_51 rwl_1_51
+ rwl_0_51 cell_2r1w
Xcell_2r1w_1486 vdd_uq23 gnd read_bl_0_40 read_bl_1_40 write_bl_0_40 wwl_0_49 rwl_1_49
+ rwl_0_49 cell_2r1w
Xcell_2r1w_2132 vdd_uq20 gnd read_bl_0_30 read_bl_1_30 write_bl_0_30 wwl_0_43 rwl_1_43
+ rwl_0_43 cell_2r1w
Xcell_2r1w_2198 vdd_uq19 gnd read_bl_0_29 read_bl_1_29 write_bl_0_29 wwl_0_41 rwl_1_41
+ rwl_0_41 cell_2r1w
Xcell_2r1w_1431 vdd_uq19 gnd read_bl_0_41 read_bl_1_41 write_bl_0_41 wwl_0_40 rwl_1_40
+ rwl_0_40 cell_2r1w
Xcell_2r1w_2143 vdd_uq15 gnd read_bl_0_30 read_bl_1_30 write_bl_0_30 wwl_0_32 rwl_1_32
+ rwl_0_32 cell_2r1w
Xcell_2r1w_1442 vdd_uq13 gnd read_bl_0_41 read_bl_1_41 write_bl_0_41 wwl_0_29 rwl_1_29
+ rwl_0_29 cell_2r1w
Xcell_2r1w_2110 vdd_uq0 gnd read_bl_0_31 read_bl_1_31 write_bl_0_31 wwl_0_1 rwl_1_1
+ rwl_0_1 cell_2r1w
Xcell_2r1w_1464 vdd_uq2 gnd read_bl_0_41 read_bl_1_41 write_bl_0_41 wwl_0_7 rwl_1_7
+ rwl_0_7 cell_2r1w
Xcell_2r1w_2165 vdd_uq4 gnd read_bl_0_30 read_bl_1_30 write_bl_0_30 wwl_0_10 rwl_1_10
+ rwl_0_10 cell_2r1w
Xcell_2r1w_1453 vdd_uq8 gnd read_bl_0_41 read_bl_1_41 write_bl_0_41 wwl_0_18 rwl_1_18
+ rwl_0_18 cell_2r1w
Xcell_2r1w_2154 vdd_uq9 gnd read_bl_0_30 read_bl_1_30 write_bl_0_30 wwl_0_21 rwl_1_21
+ rwl_0_21 cell_2r1w
Xcell_2r1w_1497 vdd_uq18 gnd read_bl_0_40 read_bl_1_40 write_bl_0_40 wwl_0_38 rwl_1_38
+ rwl_0_38 cell_2r1w
Xcell_2r1w_691 vdd_uq5 gnd read_bl_0_53 read_bl_1_53 write_bl_0_53 wwl_0_12 rwl_1_12
+ rwl_0_12 cell_2r1w
Xcell_2r1w_680 vdd_uq10 gnd read_bl_0_53 read_bl_1_53 write_bl_0_53 wwl_0_23 rwl_1_23
+ rwl_0_23 cell_2r1w
Xcell_2r1w_4090 vdd_uq1 gnd read_bl_0_0 read_bl_1_0 write_bl_0_0 wwl_0_5 rwl_1_5 rwl_0_5
+ cell_2r1w
Xcell_2r1w_1283 vdd_uq29 gnd read_bl_0_43 read_bl_1_43 write_bl_0_43 wwl_0_60 rwl_1_60
+ rwl_0_60 cell_2r1w
Xcell_2r1w_1294 vdd_uq23 gnd read_bl_0_43 read_bl_1_43 write_bl_0_43 wwl_0_49 rwl_1_49
+ rwl_0_49 cell_2r1w
Xcell_2r1w_1250 vdd_uq13 gnd read_bl_0_44 read_bl_1_44 write_bl_0_44 wwl_0_29 rwl_1_29
+ rwl_0_29 cell_2r1w
Xcell_2r1w_1272 vdd_uq2 gnd read_bl_0_44 read_bl_1_44 write_bl_0_44 wwl_0_7 rwl_1_7
+ rwl_0_7 cell_2r1w
Xcell_2r1w_1261 vdd_uq8 gnd read_bl_0_44 read_bl_1_44 write_bl_0_44 wwl_0_18 rwl_1_18
+ rwl_0_18 cell_2r1w
Xcell_2r1w_1091 vdd_uq29 gnd read_bl_0_46 read_bl_1_46 write_bl_0_46 wwl_0_60 rwl_1_60
+ rwl_0_60 cell_2r1w
Xcell_2r1w_1080 vdd_uq2 gnd read_bl_0_47 read_bl_1_47 write_bl_0_47 wwl_0_7 rwl_1_7
+ rwl_0_7 cell_2r1w
Xcell_2r1w_2709 vdd_uq20 gnd read_bl_0_21 read_bl_1_21 write_bl_0_21 wwl_0_42 rwl_1_42
+ rwl_0_42 cell_2r1w
Xcell_2r1w_3911 vdd_uq27 gnd read_bl_0_2 read_bl_1_2 write_bl_0_2 wwl_0_56 rwl_1_56
+ rwl_0_56 cell_2r1w
Xcell_2r1w_3977 vdd_uq26 gnd read_bl_0_1 read_bl_1_1 write_bl_0_1 wwl_0_54 rwl_1_54
+ rwl_0_54 cell_2r1w
Xcell_2r1w_3922 vdd_uq21 gnd read_bl_0_2 read_bl_1_2 write_bl_0_2 wwl_0_45 rwl_1_45
+ rwl_0_45 cell_2r1w
Xcell_2r1w_3988 vdd_uq20 gnd read_bl_0_1 read_bl_1_1 write_bl_0_1 wwl_0_43 rwl_1_43
+ rwl_0_43 cell_2r1w
Xcell_2r1w_3933 vdd_uq16 gnd read_bl_0_2 read_bl_1_2 write_bl_0_2 wwl_0_34 rwl_1_34
+ rwl_0_34 cell_2r1w
Xcell_2r1w_3999 vdd_uq15 gnd read_bl_0_1 read_bl_1_1 write_bl_0_1 wwl_0_32 rwl_1_32
+ rwl_0_32 cell_2r1w
Xcell_2r1w_3900 vdd gnd read_bl_0_3 read_bl_1_3 write_bl_0_3 wwl_0_3 rwl_1_3 rwl_0_3
+ cell_2r1w
Xcell_2r1w_3966 vdd_uq0 gnd read_bl_0_2 read_bl_1_2 write_bl_0_2 wwl_0_1 rwl_1_1 rwl_0_1
+ cell_2r1w
Xcell_2r1w_3955 vdd_uq5 gnd read_bl_0_2 read_bl_1_2 write_bl_0_2 wwl_0_12 rwl_1_12
+ rwl_0_12 cell_2r1w
Xcell_2r1w_3944 vdd_uq10 gnd read_bl_0_2 read_bl_1_2 write_bl_0_2 wwl_0_23 rwl_1_23
+ rwl_0_23 cell_2r1w
Xcell_2r1w_509 vdd gnd read_bl_0_56 read_bl_1_56 write_bl_0_56 wwl_0_2 rwl_1_2 rwl_0_2
+ cell_2r1w
Xcell_2r1w_3207 vdd_uq27 gnd read_bl_0_13 read_bl_1_13 write_bl_0_13 wwl_0_56 rwl_1_56
+ rwl_0_56 cell_2r1w
Xcell_2r1w_2506 vdd_uq25 gnd read_bl_0_24 read_bl_1_24 write_bl_0_24 wwl_0_53 rwl_1_53
+ rwl_0_53 cell_2r1w
Xcell_2r1w_1805 vdd_uq24 gnd read_bl_0_35 read_bl_1_35 write_bl_0_35 wwl_0_50 rwl_1_50
+ rwl_0_50 cell_2r1w
Xcell_2r1w_3218 vdd_uq21 gnd read_bl_0_13 read_bl_1_13 write_bl_0_13 wwl_0_45 rwl_1_45
+ rwl_0_45 cell_2r1w
Xcell_2r1w_2517 vdd_uq20 gnd read_bl_0_24 read_bl_1_24 write_bl_0_24 wwl_0_42 rwl_1_42
+ rwl_0_42 cell_2r1w
Xcell_2r1w_1816 vdd_uq18 gnd read_bl_0_35 read_bl_1_35 write_bl_0_35 wwl_0_39 rwl_1_39
+ rwl_0_39 cell_2r1w
Xcell_2r1w_3229 vdd_uq16 gnd read_bl_0_13 read_bl_1_13 write_bl_0_13 wwl_0_34 rwl_1_34
+ rwl_0_34 cell_2r1w
Xcell_2r1w_2528 vdd_uq14 gnd read_bl_0_24 read_bl_1_24 write_bl_0_24 wwl_0_31 rwl_1_31
+ rwl_0_31 cell_2r1w
Xcell_2r1w_1827 vdd_uq13 gnd read_bl_0_35 read_bl_1_35 write_bl_0_35 wwl_0_28 rwl_1_28
+ rwl_0_28 cell_2r1w
Xcell_2r1w_2539 vdd_uq9 gnd read_bl_0_24 read_bl_1_24 write_bl_0_24 wwl_0_20 rwl_1_20
+ rwl_0_20 cell_2r1w
Xcell_2r1w_1849 vdd_uq2 gnd read_bl_0_35 read_bl_1_35 write_bl_0_35 wwl_0_6 rwl_1_6
+ rwl_0_6 cell_2r1w
Xcell_2r1w_1838 vdd_uq7 gnd read_bl_0_35 read_bl_1_35 write_bl_0_35 wwl_0_17 rwl_1_17
+ rwl_0_17 cell_2r1w
Xcell_2r1w_3730 vdd_uq21 gnd read_bl_0_5 read_bl_1_5 write_bl_0_5 wwl_0_45 rwl_1_45
+ rwl_0_45 cell_2r1w
Xcell_2r1w_3785 vdd_uq26 gnd read_bl_0_4 read_bl_1_4 write_bl_0_4 wwl_0_54 rwl_1_54
+ rwl_0_54 cell_2r1w
Xcell_2r1w_3796 vdd_uq20 gnd read_bl_0_4 read_bl_1_4 write_bl_0_4 wwl_0_43 rwl_1_43
+ rwl_0_43 cell_2r1w
Xcell_2r1w_3741 vdd_uq16 gnd read_bl_0_5 read_bl_1_5 write_bl_0_5 wwl_0_34 rwl_1_34
+ rwl_0_34 cell_2r1w
Xcell_2r1w_3774 vdd_uq0 gnd read_bl_0_5 read_bl_1_5 write_bl_0_5 wwl_0_1 rwl_1_1 rwl_0_1
+ cell_2r1w
Xcell_2r1w_3763 vdd_uq5 gnd read_bl_0_5 read_bl_1_5 write_bl_0_5 wwl_0_12 rwl_1_12
+ rwl_0_12 cell_2r1w
Xcell_2r1w_3752 vdd_uq10 gnd read_bl_0_5 read_bl_1_5 write_bl_0_5 wwl_0_23 rwl_1_23
+ rwl_0_23 cell_2r1w
Xcell_2r1w_328 vdd_uq26 gnd read_bl_0_58 read_bl_1_58 write_bl_0_58 wwl_0_55 rwl_1_55
+ rwl_0_55 cell_2r1w
Xcell_2r1w_339 vdd_uq21 gnd read_bl_0_58 read_bl_1_58 write_bl_0_58 wwl_0_44 rwl_1_44
+ rwl_0_44 cell_2r1w
Xcell_2r1w_317 vdd gnd read_bl_0_59 read_bl_1_59 write_bl_0_59 wwl_0_2 rwl_1_2 rwl_0_2
+ cell_2r1w
Xcell_2r1w_306 vdd_uq5 gnd read_bl_0_59 read_bl_1_59 write_bl_0_59 wwl_0_13 rwl_1_13
+ rwl_0_13 cell_2r1w
Xcell_2r1w_3015 vdd_uq27 gnd read_bl_0_16 read_bl_1_16 write_bl_0_16 wwl_0_56 rwl_1_56
+ rwl_0_56 cell_2r1w
Xcell_2r1w_3004 vdd gnd read_bl_0_17 read_bl_1_17 write_bl_0_17 wwl_0_3 rwl_1_3 rwl_0_3
+ cell_2r1w
Xcell_2r1w_2369 vdd_uq30 gnd read_bl_0_26 read_bl_1_26 write_bl_0_26 wwl_0_62 rwl_1_62
+ rwl_0_62 cell_2r1w
Xcell_2r1w_1602 vdd_uq29 gnd read_bl_0_38 read_bl_1_38 write_bl_0_38 wwl_0_61 rwl_1_61
+ rwl_0_61 cell_2r1w
Xcell_2r1w_1668 vdd_uq28 gnd read_bl_0_37 read_bl_1_37 write_bl_0_37 wwl_0_59 rwl_1_59
+ rwl_0_59 cell_2r1w
Xcell_2r1w_840 vdd_uq26 gnd read_bl_0_50 read_bl_1_50 write_bl_0_50 wwl_0_55 rwl_1_55
+ rwl_0_55 cell_2r1w
Xcell_2r1w_2314 vdd_uq25 gnd read_bl_0_27 read_bl_1_27 write_bl_0_27 wwl_0_53 rwl_1_53
+ rwl_0_53 cell_2r1w
Xcell_2r1w_1613 vdd_uq24 gnd read_bl_0_38 read_bl_1_38 write_bl_0_38 wwl_0_50 rwl_1_50
+ rwl_0_50 cell_2r1w
Xcell_2r1w_1679 vdd_uq23 gnd read_bl_0_37 read_bl_1_37 write_bl_0_37 wwl_0_48 rwl_1_48
+ rwl_0_48 cell_2r1w
Xcell_2r1w_3026 vdd_uq21 gnd read_bl_0_16 read_bl_1_16 write_bl_0_16 wwl_0_45 rwl_1_45
+ rwl_0_45 cell_2r1w
Xcell_2r1w_2325 vdd_uq20 gnd read_bl_0_27 read_bl_1_27 write_bl_0_27 wwl_0_42 rwl_1_42
+ rwl_0_42 cell_2r1w
Xcell_2r1w_1624 vdd_uq18 gnd read_bl_0_38 read_bl_1_38 write_bl_0_38 wwl_0_39 rwl_1_39
+ rwl_0_39 cell_2r1w
Xcell_2r1w_3037 vdd_uq16 gnd read_bl_0_16 read_bl_1_16 write_bl_0_16 wwl_0_34 rwl_1_34
+ rwl_0_34 cell_2r1w
Xcell_2r1w_2336 vdd_uq14 gnd read_bl_0_27 read_bl_1_27 write_bl_0_27 wwl_0_31 rwl_1_31
+ rwl_0_31 cell_2r1w
Xcell_2r1w_1635 vdd_uq13 gnd read_bl_0_38 read_bl_1_38 write_bl_0_38 wwl_0_28 rwl_1_28
+ rwl_0_28 cell_2r1w
Xcell_2r1w_2303 vdd_uq0 gnd read_bl_0_28 read_bl_1_28 write_bl_0_28 wwl_0_0 rwl_1_0
+ rwl_0_0 cell_2r1w
Xcell_2r1w_1657 vdd_uq2 gnd read_bl_0_38 read_bl_1_38 write_bl_0_38 wwl_0_6 rwl_1_6
+ rwl_0_6 cell_2r1w
Xcell_2r1w_2358 vdd_uq3 gnd read_bl_0_27 read_bl_1_27 write_bl_0_27 wwl_0_9 rwl_1_9
+ rwl_0_9 cell_2r1w
Xcell_2r1w_3059 vdd_uq5 gnd read_bl_0_16 read_bl_1_16 write_bl_0_16 wwl_0_12 rwl_1_12
+ rwl_0_12 cell_2r1w
Xcell_2r1w_1646 vdd_uq7 gnd read_bl_0_38 read_bl_1_38 write_bl_0_38 wwl_0_17 rwl_1_17
+ rwl_0_17 cell_2r1w
Xcell_2r1w_2347 vdd_uq9 gnd read_bl_0_27 read_bl_1_27 write_bl_0_27 wwl_0_20 rwl_1_20
+ rwl_0_20 cell_2r1w
Xcell_2r1w_3048 vdd_uq10 gnd read_bl_0_16 read_bl_1_16 write_bl_0_16 wwl_0_23 rwl_1_23
+ rwl_0_23 cell_2r1w
Xcell_2r1w_851 vdd_uq21 gnd read_bl_0_50 read_bl_1_50 write_bl_0_50 wwl_0_44 rwl_1_44
+ rwl_0_44 cell_2r1w
Xcell_2r1w_862 vdd_uq15 gnd read_bl_0_50 read_bl_1_50 write_bl_0_50 wwl_0_33 rwl_1_33
+ rwl_0_33 cell_2r1w
Xcell_2r1w_895 vdd_uq0 gnd read_bl_0_50 read_bl_1_50 write_bl_0_50 wwl_0_0 rwl_1_0
+ rwl_0_0 cell_2r1w
Xcell_2r1w_884 vdd_uq4 gnd read_bl_0_50 read_bl_1_50 write_bl_0_50 wwl_0_11 rwl_1_11
+ rwl_0_11 cell_2r1w
Xcell_2r1w_873 vdd_uq10 gnd read_bl_0_50 read_bl_1_50 write_bl_0_50 wwl_0_22 rwl_1_22
+ rwl_0_22 cell_2r1w
Xcell_2r1w_3571 vdd_uq5 gnd read_bl_0_8 read_bl_1_8 write_bl_0_8 wwl_0_12 rwl_1_12
+ rwl_0_12 cell_2r1w
Xcell_2r1w_3560 vdd_uq10 gnd read_bl_0_8 read_bl_1_8 write_bl_0_8 wwl_0_23 rwl_1_23
+ rwl_0_23 cell_2r1w
Xcell_2r1w_2881 vdd_uq30 gnd read_bl_0_18 read_bl_1_18 write_bl_0_18 wwl_0_62 rwl_1_62
+ rwl_0_62 cell_2r1w
Xcell_2r1w_3593 vdd_uq26 gnd read_bl_0_7 read_bl_1_7 write_bl_0_7 wwl_0_54 rwl_1_54
+ rwl_0_54 cell_2r1w
Xcell_2r1w_2892 vdd_uq24 gnd read_bl_0_18 read_bl_1_18 write_bl_0_18 wwl_0_51 rwl_1_51
+ rwl_0_51 cell_2r1w
Xcell_2r1w_3582 vdd_uq0 gnd read_bl_0_8 read_bl_1_8 write_bl_0_8 wwl_0_1 rwl_1_1 rwl_0_1
+ cell_2r1w
Xcell_2r1w_2870 vdd_uq3 gnd read_bl_0_19 read_bl_1_19 write_bl_0_19 wwl_0_9 rwl_1_9
+ rwl_0_9 cell_2r1w
Xcell_2r1w_103 vdd_uq11 gnd read_bl_0_62 read_bl_1_62 write_bl_0_62 wwl_0_24 rwl_1_24
+ rwl_0_24 cell_2r1w
Xcell_2r1w_125 vdd gnd read_bl_0_62 read_bl_1_62 write_bl_0_62 wwl_0_2 rwl_1_2 rwl_0_2
+ cell_2r1w
Xcell_2r1w_114 vdd_uq5 gnd read_bl_0_62 read_bl_1_62 write_bl_0_62 wwl_0_13 rwl_1_13
+ rwl_0_13 cell_2r1w
Xcell_2r1w_136 vdd_uq26 gnd read_bl_0_61 read_bl_1_61 write_bl_0_61 wwl_0_55 rwl_1_55
+ rwl_0_55 cell_2r1w
Xcell_2r1w_147 vdd_uq21 gnd read_bl_0_61 read_bl_1_61 write_bl_0_61 wwl_0_44 rwl_1_44
+ rwl_0_44 cell_2r1w
Xcell_2r1w_158 vdd_uq15 gnd read_bl_0_61 read_bl_1_61 write_bl_0_61 wwl_0_33 rwl_1_33
+ rwl_0_33 cell_2r1w
Xcell_2r1w_169 vdd_uq10 gnd read_bl_0_61 read_bl_1_61 write_bl_0_61 wwl_0_22 rwl_1_22
+ rwl_0_22 cell_2r1w
Xcell_2r1w_2122 vdd_uq25 gnd read_bl_0_30 read_bl_1_30 write_bl_0_30 wwl_0_53 rwl_1_53
+ rwl_0_53 cell_2r1w
Xcell_2r1w_2111 vdd_uq0 gnd read_bl_0_31 read_bl_1_31 write_bl_0_31 wwl_0_0 rwl_1_0
+ rwl_0_0 cell_2r1w
Xcell_2r1w_2100 vdd_uq4 gnd read_bl_0_31 read_bl_1_31 write_bl_0_31 wwl_0_11 rwl_1_11
+ rwl_0_11 cell_2r1w
Xcell_2r1w_2177 vdd_uq30 gnd read_bl_0_29 read_bl_1_29 write_bl_0_29 wwl_0_62 rwl_1_62
+ rwl_0_62 cell_2r1w
Xcell_2r1w_1410 vdd_uq29 gnd read_bl_0_41 read_bl_1_41 write_bl_0_41 wwl_0_61 rwl_1_61
+ rwl_0_61 cell_2r1w
Xcell_2r1w_1476 vdd_uq28 gnd read_bl_0_40 read_bl_1_40 write_bl_0_40 wwl_0_59 rwl_1_59
+ rwl_0_59 cell_2r1w
Xcell_2r1w_2188 vdd_uq24 gnd read_bl_0_29 read_bl_1_29 write_bl_0_29 wwl_0_51 rwl_1_51
+ rwl_0_51 cell_2r1w
Xcell_2r1w_1421 vdd_uq24 gnd read_bl_0_41 read_bl_1_41 write_bl_0_41 wwl_0_50 rwl_1_50
+ rwl_0_50 cell_2r1w
Xcell_2r1w_1487 vdd_uq23 gnd read_bl_0_40 read_bl_1_40 write_bl_0_40 wwl_0_48 rwl_1_48
+ rwl_0_48 cell_2r1w
Xcell_2r1w_2133 vdd_uq20 gnd read_bl_0_30 read_bl_1_30 write_bl_0_30 wwl_0_42 rwl_1_42
+ rwl_0_42 cell_2r1w
Xcell_2r1w_2199 vdd_uq19 gnd read_bl_0_29 read_bl_1_29 write_bl_0_29 wwl_0_40 rwl_1_40
+ rwl_0_40 cell_2r1w
Xcell_2r1w_1432 vdd_uq18 gnd read_bl_0_41 read_bl_1_41 write_bl_0_41 wwl_0_39 rwl_1_39
+ rwl_0_39 cell_2r1w
Xcell_2r1w_1498 vdd_uq17 gnd read_bl_0_40 read_bl_1_40 write_bl_0_40 wwl_0_37 rwl_1_37
+ rwl_0_37 cell_2r1w
Xcell_2r1w_670 vdd_uq15 gnd read_bl_0_53 read_bl_1_53 write_bl_0_53 wwl_0_33 rwl_1_33
+ rwl_0_33 cell_2r1w
Xcell_2r1w_2144 vdd_uq14 gnd read_bl_0_30 read_bl_1_30 write_bl_0_30 wwl_0_31 rwl_1_31
+ rwl_0_31 cell_2r1w
Xcell_2r1w_1443 vdd_uq13 gnd read_bl_0_41 read_bl_1_41 write_bl_0_41 wwl_0_28 rwl_1_28
+ rwl_0_28 cell_2r1w
Xcell_2r1w_1465 vdd_uq2 gnd read_bl_0_41 read_bl_1_41 write_bl_0_41 wwl_0_6 rwl_1_6
+ rwl_0_6 cell_2r1w
Xcell_2r1w_2166 vdd_uq3 gnd read_bl_0_30 read_bl_1_30 write_bl_0_30 wwl_0_9 rwl_1_9
+ rwl_0_9 cell_2r1w
Xcell_2r1w_1454 vdd_uq7 gnd read_bl_0_41 read_bl_1_41 write_bl_0_41 wwl_0_17 rwl_1_17
+ rwl_0_17 cell_2r1w
Xcell_2r1w_2155 vdd_uq9 gnd read_bl_0_30 read_bl_1_30 write_bl_0_30 wwl_0_20 rwl_1_20
+ rwl_0_20 cell_2r1w
Xcell_2r1w_681 vdd_uq10 gnd read_bl_0_53 read_bl_1_53 write_bl_0_53 wwl_0_22 rwl_1_22
+ rwl_0_22 cell_2r1w
Xcell_2r1w_692 vdd_uq4 gnd read_bl_0_53 read_bl_1_53 write_bl_0_53 wwl_0_11 rwl_1_11
+ rwl_0_11 cell_2r1w
Xcell_2r1w_4091 vdd_uq1 gnd read_bl_0_0 read_bl_1_0 write_bl_0_0 wwl_0_4 rwl_1_4 rwl_0_4
+ cell_2r1w
Xcell_2r1w_3390 vdd_uq0 gnd read_bl_0_11 read_bl_1_11 write_bl_0_11 wwl_0_1 rwl_1_1
+ rwl_0_1 cell_2r1w
Xcell_2r1w_4080 vdd_uq6 gnd read_bl_0_0 read_bl_1_0 write_bl_0_0 wwl_0_15 rwl_1_15
+ rwl_0_15 cell_2r1w
Xcell_2r1w_1284 vdd_uq28 gnd read_bl_0_43 read_bl_1_43 write_bl_0_43 wwl_0_59 rwl_1_59
+ rwl_0_59 cell_2r1w
Xcell_2r1w_1295 vdd_uq23 gnd read_bl_0_43 read_bl_1_43 write_bl_0_43 wwl_0_48 rwl_1_48
+ rwl_0_48 cell_2r1w
Xcell_2r1w_1240 vdd_uq18 gnd read_bl_0_44 read_bl_1_44 write_bl_0_44 wwl_0_39 rwl_1_39
+ rwl_0_39 cell_2r1w
Xcell_2r1w_1251 vdd_uq13 gnd read_bl_0_44 read_bl_1_44 write_bl_0_44 wwl_0_28 rwl_1_28
+ rwl_0_28 cell_2r1w
Xcell_2r1w_1273 vdd_uq2 gnd read_bl_0_44 read_bl_1_44 write_bl_0_44 wwl_0_6 rwl_1_6
+ rwl_0_6 cell_2r1w
Xcell_2r1w_1262 vdd_uq7 gnd read_bl_0_44 read_bl_1_44 write_bl_0_44 wwl_0_17 rwl_1_17
+ rwl_0_17 cell_2r1w
Xcell_2r1w_1070 vdd_uq7 gnd read_bl_0_47 read_bl_1_47 write_bl_0_47 wwl_0_17 rwl_1_17
+ rwl_0_17 cell_2r1w
Xcell_2r1w_1092 vdd_uq28 gnd read_bl_0_46 read_bl_1_46 write_bl_0_46 wwl_0_59 rwl_1_59
+ rwl_0_59 cell_2r1w
Xcell_2r1w_1081 vdd_uq2 gnd read_bl_0_47 read_bl_1_47 write_bl_0_47 wwl_0_6 rwl_1_6
+ rwl_0_6 cell_2r1w
Xcell_2r1w_3912 vdd_uq26 gnd read_bl_0_2 read_bl_1_2 write_bl_0_2 wwl_0_55 rwl_1_55
+ rwl_0_55 cell_2r1w
Xcell_2r1w_3901 vdd gnd read_bl_0_3 read_bl_1_3 write_bl_0_3 wwl_0_2 rwl_1_2 rwl_0_2
+ cell_2r1w
Xcell_2r1w_3978 vdd_uq25 gnd read_bl_0_1 read_bl_1_1 write_bl_0_1 wwl_0_53 rwl_1_53
+ rwl_0_53 cell_2r1w
Xcell_2r1w_3923 vdd_uq21 gnd read_bl_0_2 read_bl_1_2 write_bl_0_2 wwl_0_44 rwl_1_44
+ rwl_0_44 cell_2r1w
Xcell_2r1w_3989 vdd_uq20 gnd read_bl_0_1 read_bl_1_1 write_bl_0_1 wwl_0_42 rwl_1_42
+ rwl_0_42 cell_2r1w
Xcell_2r1w_3934 vdd_uq15 gnd read_bl_0_2 read_bl_1_2 write_bl_0_2 wwl_0_33 rwl_1_33
+ rwl_0_33 cell_2r1w
Xcell_2r1w_3967 vdd_uq0 gnd read_bl_0_2 read_bl_1_2 write_bl_0_2 wwl_0_0 rwl_1_0 rwl_0_0
+ cell_2r1w
Xcell_2r1w_3956 vdd_uq4 gnd read_bl_0_2 read_bl_1_2 write_bl_0_2 wwl_0_11 rwl_1_11
+ rwl_0_11 cell_2r1w
Xcell_2r1w_3945 vdd_uq10 gnd read_bl_0_2 read_bl_1_2 write_bl_0_2 wwl_0_22 rwl_1_22
+ rwl_0_22 cell_2r1w
Xcell_2r1w_3208 vdd_uq26 gnd read_bl_0_13 read_bl_1_13 write_bl_0_13 wwl_0_55 rwl_1_55
+ rwl_0_55 cell_2r1w
Xcell_2r1w_2507 vdd_uq25 gnd read_bl_0_24 read_bl_1_24 write_bl_0_24 wwl_0_52 rwl_1_52
+ rwl_0_52 cell_2r1w
Xcell_2r1w_1806 vdd_uq23 gnd read_bl_0_35 read_bl_1_35 write_bl_0_35 wwl_0_49 rwl_1_49
+ rwl_0_49 cell_2r1w
Xcell_2r1w_3219 vdd_uq21 gnd read_bl_0_13 read_bl_1_13 write_bl_0_13 wwl_0_44 rwl_1_44
+ rwl_0_44 cell_2r1w
Xcell_2r1w_2518 vdd_uq19 gnd read_bl_0_24 read_bl_1_24 write_bl_0_24 wwl_0_41 rwl_1_41
+ rwl_0_41 cell_2r1w
Xcell_2r1w_1817 vdd_uq18 gnd read_bl_0_35 read_bl_1_35 write_bl_0_35 wwl_0_38 rwl_1_38
+ rwl_0_38 cell_2r1w
Xcell_2r1w_2529 vdd_uq14 gnd read_bl_0_24 read_bl_1_24 write_bl_0_24 wwl_0_30 rwl_1_30
+ rwl_0_30 cell_2r1w
Xcell_2r1w_1828 vdd_uq12 gnd read_bl_0_35 read_bl_1_35 write_bl_0_35 wwl_0_27 rwl_1_27
+ rwl_0_27 cell_2r1w
Xcell_2r1w_1839 vdd_uq7 gnd read_bl_0_35 read_bl_1_35 write_bl_0_35 wwl_0_16 rwl_1_16
+ rwl_0_16 cell_2r1w
Xcell_2r1w_3720 vdd_uq26 gnd read_bl_0_5 read_bl_1_5 write_bl_0_5 wwl_0_55 rwl_1_55
+ rwl_0_55 cell_2r1w
Xcell_2r1w_3731 vdd_uq21 gnd read_bl_0_5 read_bl_1_5 write_bl_0_5 wwl_0_44 rwl_1_44
+ rwl_0_44 cell_2r1w
Xcell_2r1w_3742 vdd_uq15 gnd read_bl_0_5 read_bl_1_5 write_bl_0_5 wwl_0_33 rwl_1_33
+ rwl_0_33 cell_2r1w
Xcell_2r1w_3753 vdd_uq10 gnd read_bl_0_5 read_bl_1_5 write_bl_0_5 wwl_0_22 rwl_1_22
+ rwl_0_22 cell_2r1w
Xcell_2r1w_3786 vdd_uq25 gnd read_bl_0_4 read_bl_1_4 write_bl_0_4 wwl_0_53 rwl_1_53
+ rwl_0_53 cell_2r1w
Xcell_2r1w_3797 vdd_uq20 gnd read_bl_0_4 read_bl_1_4 write_bl_0_4 wwl_0_42 rwl_1_42
+ rwl_0_42 cell_2r1w
Xcell_2r1w_3775 vdd_uq0 gnd read_bl_0_5 read_bl_1_5 write_bl_0_5 wwl_0_0 rwl_1_0 rwl_0_0
+ cell_2r1w
Xcell_2r1w_3764 vdd_uq4 gnd read_bl_0_5 read_bl_1_5 write_bl_0_5 wwl_0_11 rwl_1_11
+ rwl_0_11 cell_2r1w
Xcell_2r1w_318 vdd_uq0 gnd read_bl_0_59 read_bl_1_59 write_bl_0_59 wwl_0_1 rwl_1_1
+ rwl_0_1 cell_2r1w
Xcell_2r1w_307 vdd_uq5 gnd read_bl_0_59 read_bl_1_59 write_bl_0_59 wwl_0_12 rwl_1_12
+ rwl_0_12 cell_2r1w
Xcell_2r1w_329 vdd_uq26 gnd read_bl_0_58 read_bl_1_58 write_bl_0_58 wwl_0_54 rwl_1_54
+ rwl_0_54 cell_2r1w
Xcell_2r1w_2304 vdd_uq30 gnd read_bl_0_27 read_bl_1_27 write_bl_0_27 wwl_0_63 rwl_1_63
+ rwl_0_63 cell_2r1w
Xcell_2r1w_3016 vdd_uq26 gnd read_bl_0_16 read_bl_1_16 write_bl_0_16 wwl_0_55 rwl_1_55
+ rwl_0_55 cell_2r1w
Xcell_2r1w_3027 vdd_uq21 gnd read_bl_0_16 read_bl_1_16 write_bl_0_16 wwl_0_44 rwl_1_44
+ rwl_0_44 cell_2r1w
Xcell_2r1w_3038 vdd_uq15 gnd read_bl_0_16 read_bl_1_16 write_bl_0_16 wwl_0_33 rwl_1_33
+ rwl_0_33 cell_2r1w
Xcell_2r1w_3005 vdd gnd read_bl_0_17 read_bl_1_17 write_bl_0_17 wwl_0_2 rwl_1_2 rwl_0_2
+ cell_2r1w
Xcell_2r1w_3049 vdd_uq10 gnd read_bl_0_16 read_bl_1_16 write_bl_0_16 wwl_0_22 rwl_1_22
+ rwl_0_22 cell_2r1w
Xcell_2r1w_1603 vdd_uq29 gnd read_bl_0_38 read_bl_1_38 write_bl_0_38 wwl_0_60 rwl_1_60
+ rwl_0_60 cell_2r1w
Xcell_2r1w_1669 vdd_uq28 gnd read_bl_0_37 read_bl_1_37 write_bl_0_37 wwl_0_58 rwl_1_58
+ rwl_0_58 cell_2r1w
Xcell_2r1w_841 vdd_uq26 gnd read_bl_0_50 read_bl_1_50 write_bl_0_50 wwl_0_54 rwl_1_54
+ rwl_0_54 cell_2r1w
Xcell_2r1w_2315 vdd_uq25 gnd read_bl_0_27 read_bl_1_27 write_bl_0_27 wwl_0_52 rwl_1_52
+ rwl_0_52 cell_2r1w
Xcell_2r1w_1614 vdd_uq23 gnd read_bl_0_38 read_bl_1_38 write_bl_0_38 wwl_0_49 rwl_1_49
+ rwl_0_49 cell_2r1w
Xcell_2r1w_852 vdd_uq20 gnd read_bl_0_50 read_bl_1_50 write_bl_0_50 wwl_0_43 rwl_1_43
+ rwl_0_43 cell_2r1w
Xcell_2r1w_2326 vdd_uq19 gnd read_bl_0_27 read_bl_1_27 write_bl_0_27 wwl_0_41 rwl_1_41
+ rwl_0_41 cell_2r1w
Xcell_2r1w_1625 vdd_uq18 gnd read_bl_0_38 read_bl_1_38 write_bl_0_38 wwl_0_38 rwl_1_38
+ rwl_0_38 cell_2r1w
Xcell_2r1w_863 vdd_uq15 gnd read_bl_0_50 read_bl_1_50 write_bl_0_50 wwl_0_32 rwl_1_32
+ rwl_0_32 cell_2r1w
Xcell_2r1w_2337 vdd_uq14 gnd read_bl_0_27 read_bl_1_27 write_bl_0_27 wwl_0_30 rwl_1_30
+ rwl_0_30 cell_2r1w
Xcell_2r1w_1636 vdd_uq12 gnd read_bl_0_38 read_bl_1_38 write_bl_0_38 wwl_0_27 rwl_1_27
+ rwl_0_27 cell_2r1w
Xcell_2r1w_1658 vdd_uq1 gnd read_bl_0_38 read_bl_1_38 write_bl_0_38 wwl_0_5 rwl_1_5
+ rwl_0_5 cell_2r1w
Xcell_2r1w_830 vdd_uq0 gnd read_bl_0_51 read_bl_1_51 write_bl_0_51 wwl_0_1 rwl_1_1
+ rwl_0_1 cell_2r1w
Xcell_2r1w_2359 vdd_uq3 gnd read_bl_0_27 read_bl_1_27 write_bl_0_27 wwl_0_8 rwl_1_8
+ rwl_0_8 cell_2r1w
Xcell_2r1w_1647 vdd_uq7 gnd read_bl_0_38 read_bl_1_38 write_bl_0_38 wwl_0_16 rwl_1_16
+ rwl_0_16 cell_2r1w
Xcell_2r1w_2348 vdd_uq8 gnd read_bl_0_27 read_bl_1_27 write_bl_0_27 wwl_0_19 rwl_1_19
+ rwl_0_19 cell_2r1w
Xcell_2r1w_896 vdd_uq30 gnd read_bl_0_49 read_bl_1_49 write_bl_0_49 wwl_0_63 rwl_1_63
+ rwl_0_63 cell_2r1w
Xcell_2r1w_885 vdd_uq4 gnd read_bl_0_50 read_bl_1_50 write_bl_0_50 wwl_0_10 rwl_1_10
+ rwl_0_10 cell_2r1w
Xcell_2r1w_874 vdd_uq9 gnd read_bl_0_50 read_bl_1_50 write_bl_0_50 wwl_0_21 rwl_1_21
+ rwl_0_21 cell_2r1w
Xcell_2r1w_3594 vdd_uq25 gnd read_bl_0_7 read_bl_1_7 write_bl_0_7 wwl_0_53 rwl_1_53
+ rwl_0_53 cell_2r1w
Xcell_2r1w_3550 vdd_uq15 gnd read_bl_0_8 read_bl_1_8 write_bl_0_8 wwl_0_33 rwl_1_33
+ rwl_0_33 cell_2r1w
Xcell_2r1w_3583 vdd_uq0 gnd read_bl_0_8 read_bl_1_8 write_bl_0_8 wwl_0_0 rwl_1_0 rwl_0_0
+ cell_2r1w
Xcell_2r1w_3572 vdd_uq4 gnd read_bl_0_8 read_bl_1_8 write_bl_0_8 wwl_0_11 rwl_1_11
+ rwl_0_11 cell_2r1w
Xcell_2r1w_2860 vdd_uq8 gnd read_bl_0_19 read_bl_1_19 write_bl_0_19 wwl_0_19 rwl_1_19
+ rwl_0_19 cell_2r1w
Xcell_2r1w_3561 vdd_uq10 gnd read_bl_0_8 read_bl_1_8 write_bl_0_8 wwl_0_22 rwl_1_22
+ rwl_0_22 cell_2r1w
Xcell_2r1w_2882 vdd_uq29 gnd read_bl_0_18 read_bl_1_18 write_bl_0_18 wwl_0_61 rwl_1_61
+ rwl_0_61 cell_2r1w
Xcell_2r1w_2893 vdd_uq24 gnd read_bl_0_18 read_bl_1_18 write_bl_0_18 wwl_0_50 rwl_1_50
+ rwl_0_50 cell_2r1w
Xcell_2r1w_2871 vdd_uq3 gnd read_bl_0_19 read_bl_1_19 write_bl_0_19 wwl_0_8 rwl_1_8
+ rwl_0_8 cell_2r1w
Xcell_2r1w_137 vdd_uq26 gnd read_bl_0_61 read_bl_1_61 write_bl_0_61 wwl_0_54 rwl_1_54
+ rwl_0_54 cell_2r1w
Xcell_2r1w_148 vdd_uq20 gnd read_bl_0_61 read_bl_1_61 write_bl_0_61 wwl_0_43 rwl_1_43
+ rwl_0_43 cell_2r1w
Xcell_2r1w_159 vdd_uq15 gnd read_bl_0_61 read_bl_1_61 write_bl_0_61 wwl_0_32 rwl_1_32
+ rwl_0_32 cell_2r1w
Xcell_2r1w_126 vdd_uq0 gnd read_bl_0_62 read_bl_1_62 write_bl_0_62 wwl_0_1 rwl_1_1
+ rwl_0_1 cell_2r1w
Xcell_2r1w_115 vdd_uq5 gnd read_bl_0_62 read_bl_1_62 write_bl_0_62 wwl_0_12 rwl_1_12
+ rwl_0_12 cell_2r1w
Xcell_2r1w_104 vdd_uq10 gnd read_bl_0_62 read_bl_1_62 write_bl_0_62 wwl_0_23 rwl_1_23
+ rwl_0_23 cell_2r1w
Xcell_2r1w_2112 vdd_uq30 gnd read_bl_0_30 read_bl_1_30 write_bl_0_30 wwl_0_63 rwl_1_63
+ rwl_0_63 cell_2r1w
Xcell_2r1w_1411 vdd_uq29 gnd read_bl_0_41 read_bl_1_41 write_bl_0_41 wwl_0_60 rwl_1_60
+ rwl_0_60 cell_2r1w
Xcell_2r1w_2123 vdd_uq25 gnd read_bl_0_30 read_bl_1_30 write_bl_0_30 wwl_0_52 rwl_1_52
+ rwl_0_52 cell_2r1w
Xcell_2r1w_2134 vdd_uq19 gnd read_bl_0_30 read_bl_1_30 write_bl_0_30 wwl_0_41 rwl_1_41
+ rwl_0_41 cell_2r1w
Xcell_2r1w_2145 vdd_uq14 gnd read_bl_0_30 read_bl_1_30 write_bl_0_30 wwl_0_30 rwl_1_30
+ rwl_0_30 cell_2r1w
Xcell_2r1w_1400 vdd_uq2 gnd read_bl_0_42 read_bl_1_42 write_bl_0_42 wwl_0_7 rwl_1_7
+ rwl_0_7 cell_2r1w
Xcell_2r1w_2101 vdd_uq4 gnd read_bl_0_31 read_bl_1_31 write_bl_0_31 wwl_0_10 rwl_1_10
+ rwl_0_10 cell_2r1w
Xcell_2r1w_2156 vdd_uq8 gnd read_bl_0_30 read_bl_1_30 write_bl_0_30 wwl_0_19 rwl_1_19
+ rwl_0_19 cell_2r1w
Xcell_2r1w_2178 vdd_uq29 gnd read_bl_0_29 read_bl_1_29 write_bl_0_29 wwl_0_61 rwl_1_61
+ rwl_0_61 cell_2r1w
Xcell_2r1w_1477 vdd_uq28 gnd read_bl_0_40 read_bl_1_40 write_bl_0_40 wwl_0_58 rwl_1_58
+ rwl_0_58 cell_2r1w
Xcell_2r1w_2189 vdd_uq24 gnd read_bl_0_29 read_bl_1_29 write_bl_0_29 wwl_0_50 rwl_1_50
+ rwl_0_50 cell_2r1w
Xcell_2r1w_1422 vdd_uq23 gnd read_bl_0_41 read_bl_1_41 write_bl_0_41 wwl_0_49 rwl_1_49
+ rwl_0_49 cell_2r1w
Xcell_2r1w_1488 vdd_uq22 gnd read_bl_0_40 read_bl_1_40 write_bl_0_40 wwl_0_47 rwl_1_47
+ rwl_0_47 cell_2r1w
Xcell_2r1w_660 vdd_uq20 gnd read_bl_0_53 read_bl_1_53 write_bl_0_53 wwl_0_43 rwl_1_43
+ rwl_0_43 cell_2r1w
Xcell_2r1w_1433 vdd_uq18 gnd read_bl_0_41 read_bl_1_41 write_bl_0_41 wwl_0_38 rwl_1_38
+ rwl_0_38 cell_2r1w
Xcell_2r1w_1499 vdd_uq17 gnd read_bl_0_40 read_bl_1_40 write_bl_0_40 wwl_0_36 rwl_1_36
+ rwl_0_36 cell_2r1w
Xcell_2r1w_671 vdd_uq15 gnd read_bl_0_53 read_bl_1_53 write_bl_0_53 wwl_0_32 rwl_1_32
+ rwl_0_32 cell_2r1w
Xcell_2r1w_1444 vdd_uq12 gnd read_bl_0_41 read_bl_1_41 write_bl_0_41 wwl_0_27 rwl_1_27
+ rwl_0_27 cell_2r1w
Xcell_2r1w_1466 vdd_uq1 gnd read_bl_0_41 read_bl_1_41 write_bl_0_41 wwl_0_5 rwl_1_5
+ rwl_0_5 cell_2r1w
Xcell_2r1w_2167 vdd_uq3 gnd read_bl_0_30 read_bl_1_30 write_bl_0_30 wwl_0_8 rwl_1_8
+ rwl_0_8 cell_2r1w
Xcell_2r1w_693 vdd_uq4 gnd read_bl_0_53 read_bl_1_53 write_bl_0_53 wwl_0_10 rwl_1_10
+ rwl_0_10 cell_2r1w
Xcell_2r1w_1455 vdd_uq7 gnd read_bl_0_41 read_bl_1_41 write_bl_0_41 wwl_0_16 rwl_1_16
+ rwl_0_16 cell_2r1w
Xcell_2r1w_682 vdd_uq9 gnd read_bl_0_53 read_bl_1_53 write_bl_0_53 wwl_0_21 rwl_1_21
+ rwl_0_21 cell_2r1w
Xcell_2r1w_2690 vdd_uq29 gnd read_bl_0_21 read_bl_1_21 write_bl_0_21 wwl_0_61 rwl_1_61
+ rwl_0_61 cell_2r1w
Xcell_2r1w_4070 vdd_uq11 gnd read_bl_0_0 read_bl_1_0 write_bl_0_0 wwl_0_25 rwl_1_25
+ rwl_0_25 cell_2r1w
Xcell_2r1w_4092 vdd gnd read_bl_0_0 read_bl_1_0 write_bl_0_0 wwl_0_3 rwl_1_3 rwl_0_3
+ cell_2r1w
Xcell_2r1w_3391 vdd_uq0 gnd read_bl_0_11 read_bl_1_11 write_bl_0_11 wwl_0_0 rwl_1_0
+ rwl_0_0 cell_2r1w
Xcell_2r1w_3380 vdd_uq4 gnd read_bl_0_11 read_bl_1_11 write_bl_0_11 wwl_0_11 rwl_1_11
+ rwl_0_11 cell_2r1w
Xcell_2r1w_4081 vdd_uq6 gnd read_bl_0_0 read_bl_1_0 write_bl_0_0 wwl_0_14 rwl_1_14
+ rwl_0_14 cell_2r1w
Xcell_2r1w_1230 vdd_uq23 gnd read_bl_0_44 read_bl_1_44 write_bl_0_44 wwl_0_49 rwl_1_49
+ rwl_0_49 cell_2r1w
Xcell_2r1w_1241 vdd_uq18 gnd read_bl_0_44 read_bl_1_44 write_bl_0_44 wwl_0_38 rwl_1_38
+ rwl_0_38 cell_2r1w
Xcell_2r1w_1252 vdd_uq12 gnd read_bl_0_44 read_bl_1_44 write_bl_0_44 wwl_0_27 rwl_1_27
+ rwl_0_27 cell_2r1w
Xcell_2r1w_1285 vdd_uq28 gnd read_bl_0_43 read_bl_1_43 write_bl_0_43 wwl_0_58 rwl_1_58
+ rwl_0_58 cell_2r1w
Xcell_2r1w_1296 vdd_uq22 gnd read_bl_0_43 read_bl_1_43 write_bl_0_43 wwl_0_47 rwl_1_47
+ rwl_0_47 cell_2r1w
Xcell_2r1w_1274 vdd_uq1 gnd read_bl_0_44 read_bl_1_44 write_bl_0_44 wwl_0_5 rwl_1_5
+ rwl_0_5 cell_2r1w
Xcell_2r1w_1263 vdd_uq7 gnd read_bl_0_44 read_bl_1_44 write_bl_0_44 wwl_0_16 rwl_1_16
+ rwl_0_16 cell_2r1w
Xcell_2r1w_490 vdd_uq9 gnd read_bl_0_56 read_bl_1_56 write_bl_0_56 wwl_0_21 rwl_1_21
+ rwl_0_21 cell_2r1w
Xcell_2r1w_1093 vdd_uq28 gnd read_bl_0_46 read_bl_1_46 write_bl_0_46 wwl_0_58 rwl_1_58
+ rwl_0_58 cell_2r1w
Xcell_2r1w_1060 vdd_uq12 gnd read_bl_0_47 read_bl_1_47 write_bl_0_47 wwl_0_27 rwl_1_27
+ rwl_0_27 cell_2r1w
Xcell_2r1w_1082 vdd_uq1 gnd read_bl_0_47 read_bl_1_47 write_bl_0_47 wwl_0_5 rwl_1_5
+ rwl_0_5 cell_2r1w
Xcell_2r1w_1071 vdd_uq7 gnd read_bl_0_47 read_bl_1_47 write_bl_0_47 wwl_0_16 rwl_1_16
+ rwl_0_16 cell_2r1w
Xcell_2r1w_3913 vdd_uq26 gnd read_bl_0_2 read_bl_1_2 write_bl_0_2 wwl_0_54 rwl_1_54
+ rwl_0_54 cell_2r1w
Xcell_2r1w_3924 vdd_uq20 gnd read_bl_0_2 read_bl_1_2 write_bl_0_2 wwl_0_43 rwl_1_43
+ rwl_0_43 cell_2r1w
Xcell_2r1w_3935 vdd_uq15 gnd read_bl_0_2 read_bl_1_2 write_bl_0_2 wwl_0_32 rwl_1_32
+ rwl_0_32 cell_2r1w
Xcell_2r1w_3902 vdd_uq0 gnd read_bl_0_3 read_bl_1_3 write_bl_0_3 wwl_0_1 rwl_1_1 rwl_0_1
+ cell_2r1w
Xcell_2r1w_3946 vdd_uq9 gnd read_bl_0_2 read_bl_1_2 write_bl_0_2 wwl_0_21 rwl_1_21
+ rwl_0_21 cell_2r1w
Xcell_2r1w_3968 vdd_uq30 gnd read_bl_0_1 read_bl_1_1 write_bl_0_1 wwl_0_63 rwl_1_63
+ rwl_0_63 cell_2r1w
Xcell_2r1w_3979 vdd_uq25 gnd read_bl_0_1 read_bl_1_1 write_bl_0_1 wwl_0_52 rwl_1_52
+ rwl_0_52 cell_2r1w
Xcell_2r1w_3957 vdd_uq4 gnd read_bl_0_2 read_bl_1_2 write_bl_0_2 wwl_0_10 rwl_1_10
+ rwl_0_10 cell_2r1w
Xcell_2r1w_3209 vdd_uq26 gnd read_bl_0_13 read_bl_1_13 write_bl_0_13 wwl_0_54 rwl_1_54
+ rwl_0_54 cell_2r1w
Xcell_2r1w_2508 vdd_uq24 gnd read_bl_0_24 read_bl_1_24 write_bl_0_24 wwl_0_51 rwl_1_51
+ rwl_0_51 cell_2r1w
Xcell_2r1w_1807 vdd_uq23 gnd read_bl_0_35 read_bl_1_35 write_bl_0_35 wwl_0_48 rwl_1_48
+ rwl_0_48 cell_2r1w
Xcell_2r1w_2519 vdd_uq19 gnd read_bl_0_24 read_bl_1_24 write_bl_0_24 wwl_0_40 rwl_1_40
+ rwl_0_40 cell_2r1w
Xcell_2r1w_1818 vdd_uq17 gnd read_bl_0_35 read_bl_1_35 write_bl_0_35 wwl_0_37 rwl_1_37
+ rwl_0_37 cell_2r1w
Xcell_2r1w_1829 vdd_uq12 gnd read_bl_0_35 read_bl_1_35 write_bl_0_35 wwl_0_26 rwl_1_26
+ rwl_0_26 cell_2r1w
Xcell_2r1w_3776 vdd_uq30 gnd read_bl_0_4 read_bl_1_4 write_bl_0_4 wwl_0_63 rwl_1_63
+ rwl_0_63 cell_2r1w
Xcell_2r1w_3721 vdd_uq26 gnd read_bl_0_5 read_bl_1_5 write_bl_0_5 wwl_0_54 rwl_1_54
+ rwl_0_54 cell_2r1w
Xcell_2r1w_3787 vdd_uq25 gnd read_bl_0_4 read_bl_1_4 write_bl_0_4 wwl_0_52 rwl_1_52
+ rwl_0_52 cell_2r1w
Xcell_2r1w_3732 vdd_uq20 gnd read_bl_0_5 read_bl_1_5 write_bl_0_5 wwl_0_43 rwl_1_43
+ rwl_0_43 cell_2r1w
Xcell_2r1w_3743 vdd_uq15 gnd read_bl_0_5 read_bl_1_5 write_bl_0_5 wwl_0_32 rwl_1_32
+ rwl_0_32 cell_2r1w
Xcell_2r1w_3710 vdd_uq0 gnd read_bl_0_6 read_bl_1_6 write_bl_0_6 wwl_0_1 rwl_1_1 rwl_0_1
+ cell_2r1w
Xcell_2r1w_3765 vdd_uq4 gnd read_bl_0_5 read_bl_1_5 write_bl_0_5 wwl_0_10 rwl_1_10
+ rwl_0_10 cell_2r1w
Xcell_2r1w_3754 vdd_uq9 gnd read_bl_0_5 read_bl_1_5 write_bl_0_5 wwl_0_21 rwl_1_21
+ rwl_0_21 cell_2r1w
Xcell_2r1w_3798 vdd_uq19 gnd read_bl_0_4 read_bl_1_4 write_bl_0_4 wwl_0_41 rwl_1_41
+ rwl_0_41 cell_2r1w
Xcell_2r1w_319 vdd_uq0 gnd read_bl_0_59 read_bl_1_59 write_bl_0_59 wwl_0_0 rwl_1_0
+ rwl_0_0 cell_2r1w
Xcell_2r1w_308 vdd_uq4 gnd read_bl_0_59 read_bl_1_59 write_bl_0_59 wwl_0_11 rwl_1_11
+ rwl_0_11 cell_2r1w
Xcell_2r1w_2305 vdd_uq30 gnd read_bl_0_27 read_bl_1_27 write_bl_0_27 wwl_0_62 rwl_1_62
+ rwl_0_62 cell_2r1w
Xcell_2r1w_3017 vdd_uq26 gnd read_bl_0_16 read_bl_1_16 write_bl_0_16 wwl_0_54 rwl_1_54
+ rwl_0_54 cell_2r1w
Xcell_2r1w_2316 vdd_uq24 gnd read_bl_0_27 read_bl_1_27 write_bl_0_27 wwl_0_51 rwl_1_51
+ rwl_0_51 cell_2r1w
Xcell_2r1w_3028 vdd_uq20 gnd read_bl_0_16 read_bl_1_16 write_bl_0_16 wwl_0_43 rwl_1_43
+ rwl_0_43 cell_2r1w
Xcell_2r1w_2327 vdd_uq19 gnd read_bl_0_27 read_bl_1_27 write_bl_0_27 wwl_0_40 rwl_1_40
+ rwl_0_40 cell_2r1w
Xcell_2r1w_3039 vdd_uq15 gnd read_bl_0_16 read_bl_1_16 write_bl_0_16 wwl_0_32 rwl_1_32
+ rwl_0_32 cell_2r1w
Xcell_2r1w_2338 vdd_uq13 gnd read_bl_0_27 read_bl_1_27 write_bl_0_27 wwl_0_29 rwl_1_29
+ rwl_0_29 cell_2r1w
Xcell_2r1w_3006 vdd_uq0 gnd read_bl_0_17 read_bl_1_17 write_bl_0_17 wwl_0_1 rwl_1_1
+ rwl_0_1 cell_2r1w
Xcell_2r1w_897 vdd_uq30 gnd read_bl_0_49 read_bl_1_49 write_bl_0_49 wwl_0_62 rwl_1_62
+ rwl_0_62 cell_2r1w
Xcell_2r1w_1604 vdd_uq28 gnd read_bl_0_38 read_bl_1_38 write_bl_0_38 wwl_0_59 rwl_1_59
+ rwl_0_59 cell_2r1w
Xcell_2r1w_842 vdd_uq25 gnd read_bl_0_50 read_bl_1_50 write_bl_0_50 wwl_0_53 rwl_1_53
+ rwl_0_53 cell_2r1w
Xcell_2r1w_1615 vdd_uq23 gnd read_bl_0_38 read_bl_1_38 write_bl_0_38 wwl_0_48 rwl_1_48
+ rwl_0_48 cell_2r1w
Xcell_2r1w_853 vdd_uq20 gnd read_bl_0_50 read_bl_1_50 write_bl_0_50 wwl_0_42 rwl_1_42
+ rwl_0_42 cell_2r1w
Xcell_2r1w_1626 vdd_uq17 gnd read_bl_0_38 read_bl_1_38 write_bl_0_38 wwl_0_37 rwl_1_37
+ rwl_0_37 cell_2r1w
Xcell_2r1w_864 vdd_uq14 gnd read_bl_0_50 read_bl_1_50 write_bl_0_50 wwl_0_31 rwl_1_31
+ rwl_0_31 cell_2r1w
Xcell_2r1w_1637 vdd_uq12 gnd read_bl_0_38 read_bl_1_38 write_bl_0_38 wwl_0_26 rwl_1_26
+ rwl_0_26 cell_2r1w
Xcell_2r1w_1659 vdd_uq1 gnd read_bl_0_38 read_bl_1_38 write_bl_0_38 wwl_0_4 rwl_1_4
+ rwl_0_4 cell_2r1w
Xcell_2r1w_831 vdd_uq0 gnd read_bl_0_51 read_bl_1_51 write_bl_0_51 wwl_0_0 rwl_1_0
+ rwl_0_0 cell_2r1w
Xcell_2r1w_886 vdd_uq3 gnd read_bl_0_50 read_bl_1_50 write_bl_0_50 wwl_0_9 rwl_1_9
+ rwl_0_9 cell_2r1w
Xcell_2r1w_820 vdd_uq4 gnd read_bl_0_51 read_bl_1_51 write_bl_0_51 wwl_0_11 rwl_1_11
+ rwl_0_11 cell_2r1w
Xcell_2r1w_1648 vdd_uq6 gnd read_bl_0_38 read_bl_1_38 write_bl_0_38 wwl_0_15 rwl_1_15
+ rwl_0_15 cell_2r1w
Xcell_2r1w_2349 vdd_uq8 gnd read_bl_0_27 read_bl_1_27 write_bl_0_27 wwl_0_18 rwl_1_18
+ rwl_0_18 cell_2r1w
Xcell_2r1w_875 vdd_uq9 gnd read_bl_0_50 read_bl_1_50 write_bl_0_50 wwl_0_20 rwl_1_20
+ rwl_0_20 cell_2r1w
Xcell_2r1w_3584 vdd_uq30 gnd read_bl_0_7 read_bl_1_7 write_bl_0_7 wwl_0_63 rwl_1_63
+ rwl_0_63 cell_2r1w
Xcell_2r1w_2883 vdd_uq29 gnd read_bl_0_18 read_bl_1_18 write_bl_0_18 wwl_0_60 rwl_1_60
+ rwl_0_60 cell_2r1w
Xcell_2r1w_3595 vdd_uq25 gnd read_bl_0_7 read_bl_1_7 write_bl_0_7 wwl_0_52 rwl_1_52
+ rwl_0_52 cell_2r1w
Xcell_2r1w_2894 vdd_uq23 gnd read_bl_0_18 read_bl_1_18 write_bl_0_18 wwl_0_49 rwl_1_49
+ rwl_0_49 cell_2r1w
Xcell_2r1w_3540 vdd_uq20 gnd read_bl_0_8 read_bl_1_8 write_bl_0_8 wwl_0_43 rwl_1_43
+ rwl_0_43 cell_2r1w
Xcell_2r1w_3551 vdd_uq15 gnd read_bl_0_8 read_bl_1_8 write_bl_0_8 wwl_0_32 rwl_1_32
+ rwl_0_32 cell_2r1w
Xcell_2r1w_2850 vdd_uq13 gnd read_bl_0_19 read_bl_1_19 write_bl_0_19 wwl_0_29 rwl_1_29
+ rwl_0_29 cell_2r1w
Xcell_2r1w_2872 vdd_uq2 gnd read_bl_0_19 read_bl_1_19 write_bl_0_19 wwl_0_7 rwl_1_7
+ rwl_0_7 cell_2r1w
Xcell_2r1w_3573 vdd_uq4 gnd read_bl_0_8 read_bl_1_8 write_bl_0_8 wwl_0_10 rwl_1_10
+ rwl_0_10 cell_2r1w
Xcell_2r1w_2861 vdd_uq8 gnd read_bl_0_19 read_bl_1_19 write_bl_0_19 wwl_0_18 rwl_1_18
+ rwl_0_18 cell_2r1w
Xcell_2r1w_3562 vdd_uq9 gnd read_bl_0_8 read_bl_1_8 write_bl_0_8 wwl_0_21 rwl_1_21
+ rwl_0_21 cell_2r1w
Xcell_2r1w_138 vdd_uq25 gnd read_bl_0_61 read_bl_1_61 write_bl_0_61 wwl_0_53 rwl_1_53
+ rwl_0_53 cell_2r1w
Xcell_2r1w_149 vdd_uq20 gnd read_bl_0_61 read_bl_1_61 write_bl_0_61 wwl_0_42 rwl_1_42
+ rwl_0_42 cell_2r1w
Xcell_2r1w_127 vdd_uq0 gnd read_bl_0_62 read_bl_1_62 write_bl_0_62 wwl_0_0 rwl_1_0
+ rwl_0_0 cell_2r1w
Xcell_2r1w_116 vdd_uq4 gnd read_bl_0_62 read_bl_1_62 write_bl_0_62 wwl_0_11 rwl_1_11
+ rwl_0_11 cell_2r1w
Xcell_2r1w_105 vdd_uq10 gnd read_bl_0_62 read_bl_1_62 write_bl_0_62 wwl_0_22 rwl_1_22
+ rwl_0_22 cell_2r1w
Xcell_2r1w_2113 vdd_uq30 gnd read_bl_0_30 read_bl_1_30 write_bl_0_30 wwl_0_62 rwl_1_62
+ rwl_0_62 cell_2r1w
Xcell_2r1w_2179 vdd_uq29 gnd read_bl_0_29 read_bl_1_29 write_bl_0_29 wwl_0_60 rwl_1_60
+ rwl_0_60 cell_2r1w
Xcell_2r1w_1412 vdd_uq28 gnd read_bl_0_41 read_bl_1_41 write_bl_0_41 wwl_0_59 rwl_1_59
+ rwl_0_59 cell_2r1w
Xcell_2r1w_2124 vdd_uq24 gnd read_bl_0_30 read_bl_1_30 write_bl_0_30 wwl_0_51 rwl_1_51
+ rwl_0_51 cell_2r1w
Xcell_2r1w_1423 vdd_uq23 gnd read_bl_0_41 read_bl_1_41 write_bl_0_41 wwl_0_48 rwl_1_48
+ rwl_0_48 cell_2r1w
Xcell_2r1w_2135 vdd_uq19 gnd read_bl_0_30 read_bl_1_30 write_bl_0_30 wwl_0_40 rwl_1_40
+ rwl_0_40 cell_2r1w
Xcell_2r1w_1434 vdd_uq17 gnd read_bl_0_41 read_bl_1_41 write_bl_0_41 wwl_0_37 rwl_1_37
+ rwl_0_37 cell_2r1w
Xcell_2r1w_2146 vdd_uq13 gnd read_bl_0_30 read_bl_1_30 write_bl_0_30 wwl_0_29 rwl_1_29
+ rwl_0_29 cell_2r1w
Xcell_2r1w_1445 vdd_uq12 gnd read_bl_0_41 read_bl_1_41 write_bl_0_41 wwl_0_26 rwl_1_26
+ rwl_0_26 cell_2r1w
Xcell_2r1w_1401 vdd_uq2 gnd read_bl_0_42 read_bl_1_42 write_bl_0_42 wwl_0_6 rwl_1_6
+ rwl_0_6 cell_2r1w
Xcell_2r1w_2168 vdd_uq2 gnd read_bl_0_30 read_bl_1_30 write_bl_0_30 wwl_0_7 rwl_1_7
+ rwl_0_7 cell_2r1w
Xcell_2r1w_2102 vdd_uq3 gnd read_bl_0_31 read_bl_1_31 write_bl_0_31 wwl_0_9 rwl_1_9
+ rwl_0_9 cell_2r1w
Xcell_2r1w_2157 vdd_uq8 gnd read_bl_0_30 read_bl_1_30 write_bl_0_30 wwl_0_18 rwl_1_18
+ rwl_0_18 cell_2r1w
Xcell_2r1w_1478 vdd_uq27 gnd read_bl_0_40 read_bl_1_40 write_bl_0_40 wwl_0_57 rwl_1_57
+ rwl_0_57 cell_2r1w
Xcell_2r1w_650 vdd_uq25 gnd read_bl_0_53 read_bl_1_53 write_bl_0_53 wwl_0_53 rwl_1_53
+ rwl_0_53 cell_2r1w
Xcell_2r1w_1489 vdd_uq22 gnd read_bl_0_40 read_bl_1_40 write_bl_0_40 wwl_0_46 rwl_1_46
+ rwl_0_46 cell_2r1w
Xcell_2r1w_661 vdd_uq20 gnd read_bl_0_53 read_bl_1_53 write_bl_0_53 wwl_0_42 rwl_1_42
+ rwl_0_42 cell_2r1w
Xcell_2r1w_672 vdd_uq14 gnd read_bl_0_53 read_bl_1_53 write_bl_0_53 wwl_0_31 rwl_1_31
+ rwl_0_31 cell_2r1w
Xcell_2r1w_1467 vdd_uq1 gnd read_bl_0_41 read_bl_1_41 write_bl_0_41 wwl_0_4 rwl_1_4
+ rwl_0_4 cell_2r1w
Xcell_2r1w_694 vdd_uq3 gnd read_bl_0_53 read_bl_1_53 write_bl_0_53 wwl_0_9 rwl_1_9
+ rwl_0_9 cell_2r1w
Xcell_2r1w_1456 vdd_uq6 gnd read_bl_0_41 read_bl_1_41 write_bl_0_41 wwl_0_15 rwl_1_15
+ rwl_0_15 cell_2r1w
Xcell_2r1w_683 vdd_uq9 gnd read_bl_0_53 read_bl_1_53 write_bl_0_53 wwl_0_20 rwl_1_20
+ rwl_0_20 cell_2r1w
Xcell_2r1w_4060 vdd_uq16 gnd read_bl_0_0 read_bl_1_0 write_bl_0_0 wwl_0_35 rwl_1_35
+ rwl_0_35 cell_2r1w
Xcell_2r1w_4071 vdd_uq11 gnd read_bl_0_0 read_bl_1_0 write_bl_0_0 wwl_0_24 rwl_1_24
+ rwl_0_24 cell_2r1w
Xcell_2r1w_4082 vdd_uq5 gnd read_bl_0_0 read_bl_1_0 write_bl_0_0 wwl_0_13 rwl_1_13
+ rwl_0_13 cell_2r1w
Xcell_2r1w_3392 vdd_uq30 gnd read_bl_0_10 read_bl_1_10 write_bl_0_10 wwl_0_63 rwl_1_63
+ rwl_0_63 cell_2r1w
Xcell_2r1w_2691 vdd_uq29 gnd read_bl_0_21 read_bl_1_21 write_bl_0_21 wwl_0_60 rwl_1_60
+ rwl_0_60 cell_2r1w
Xcell_2r1w_1990 vdd_uq27 gnd read_bl_0_32 read_bl_1_32 write_bl_0_32 wwl_0_57 rwl_1_57
+ rwl_0_57 cell_2r1w
Xcell_2r1w_4093 vdd gnd read_bl_0_0 read_bl_1_0 write_bl_0_0 wwl_0_2 rwl_1_2 rwl_0_2
+ cell_2r1w
Xcell_2r1w_2680 vdd_uq2 gnd read_bl_0_22 read_bl_1_22 write_bl_0_22 wwl_0_7 rwl_1_7
+ rwl_0_7 cell_2r1w
Xcell_2r1w_3381 vdd_uq4 gnd read_bl_0_11 read_bl_1_11 write_bl_0_11 wwl_0_10 rwl_1_10
+ rwl_0_10 cell_2r1w
Xcell_2r1w_3370 vdd_uq9 gnd read_bl_0_11 read_bl_1_11 write_bl_0_11 wwl_0_21 rwl_1_21
+ rwl_0_21 cell_2r1w
Xcell_2r1w_1220 vdd_uq28 gnd read_bl_0_44 read_bl_1_44 write_bl_0_44 wwl_0_59 rwl_1_59
+ rwl_0_59 cell_2r1w
Xcell_2r1w_1286 vdd_uq27 gnd read_bl_0_43 read_bl_1_43 write_bl_0_43 wwl_0_57 rwl_1_57
+ rwl_0_57 cell_2r1w
Xcell_2r1w_1231 vdd_uq23 gnd read_bl_0_44 read_bl_1_44 write_bl_0_44 wwl_0_48 rwl_1_48
+ rwl_0_48 cell_2r1w
Xcell_2r1w_1242 vdd_uq17 gnd read_bl_0_44 read_bl_1_44 write_bl_0_44 wwl_0_37 rwl_1_37
+ rwl_0_37 cell_2r1w
Xcell_2r1w_1253 vdd_uq12 gnd read_bl_0_44 read_bl_1_44 write_bl_0_44 wwl_0_26 rwl_1_26
+ rwl_0_26 cell_2r1w
Xcell_2r1w_1275 vdd_uq1 gnd read_bl_0_44 read_bl_1_44 write_bl_0_44 wwl_0_4 rwl_1_4
+ rwl_0_4 cell_2r1w
Xcell_2r1w_1264 vdd_uq6 gnd read_bl_0_44 read_bl_1_44 write_bl_0_44 wwl_0_15 rwl_1_15
+ rwl_0_15 cell_2r1w
Xcell_2r1w_1297 vdd_uq22 gnd read_bl_0_43 read_bl_1_43 write_bl_0_43 wwl_0_46 rwl_1_46
+ rwl_0_46 cell_2r1w
Xcell_2r1w_480 vdd_uq14 gnd read_bl_0_56 read_bl_1_56 write_bl_0_56 wwl_0_31 rwl_1_31
+ rwl_0_31 cell_2r1w
Xcell_2r1w_491 vdd_uq9 gnd read_bl_0_56 read_bl_1_56 write_bl_0_56 wwl_0_20 rwl_1_20
+ rwl_0_20 cell_2r1w
Xcell_2r1w_1094 vdd_uq27 gnd read_bl_0_46 read_bl_1_46 write_bl_0_46 wwl_0_57 rwl_1_57
+ rwl_0_57 cell_2r1w
Xcell_2r1w_1050 vdd_uq17 gnd read_bl_0_47 read_bl_1_47 write_bl_0_47 wwl_0_37 rwl_1_37
+ rwl_0_37 cell_2r1w
Xcell_2r1w_1061 vdd_uq12 gnd read_bl_0_47 read_bl_1_47 write_bl_0_47 wwl_0_26 rwl_1_26
+ rwl_0_26 cell_2r1w
Xcell_2r1w_1083 vdd_uq1 gnd read_bl_0_47 read_bl_1_47 write_bl_0_47 wwl_0_4 rwl_1_4
+ rwl_0_4 cell_2r1w
Xcell_2r1w_1072 vdd_uq6 gnd read_bl_0_47 read_bl_1_47 write_bl_0_47 wwl_0_15 rwl_1_15
+ rwl_0_15 cell_2r1w
Xcell_2r1w_3969 vdd_uq30 gnd read_bl_0_1 read_bl_1_1 write_bl_0_1 wwl_0_62 rwl_1_62
+ rwl_0_62 cell_2r1w
Xcell_2r1w_3914 vdd_uq25 gnd read_bl_0_2 read_bl_1_2 write_bl_0_2 wwl_0_53 rwl_1_53
+ rwl_0_53 cell_2r1w
Xcell_2r1w_3925 vdd_uq20 gnd read_bl_0_2 read_bl_1_2 write_bl_0_2 wwl_0_42 rwl_1_42
+ rwl_0_42 cell_2r1w
Xcell_2r1w_3936 vdd_uq14 gnd read_bl_0_2 read_bl_1_2 write_bl_0_2 wwl_0_31 rwl_1_31
+ rwl_0_31 cell_2r1w
Xcell_2r1w_3903 vdd_uq0 gnd read_bl_0_3 read_bl_1_3 write_bl_0_3 wwl_0_0 rwl_1_0 rwl_0_0
+ cell_2r1w
Xcell_2r1w_3958 vdd_uq3 gnd read_bl_0_2 read_bl_1_2 write_bl_0_2 wwl_0_9 rwl_1_9 rwl_0_9
+ cell_2r1w
Xcell_2r1w_3947 vdd_uq9 gnd read_bl_0_2 read_bl_1_2 write_bl_0_2 wwl_0_20 rwl_1_20
+ rwl_0_20 cell_2r1w
Xcell_2r1w_2509 vdd_uq24 gnd read_bl_0_24 read_bl_1_24 write_bl_0_24 wwl_0_50 rwl_1_50
+ rwl_0_50 cell_2r1w
Xcell_2r1w_1808 vdd_uq22 gnd read_bl_0_35 read_bl_1_35 write_bl_0_35 wwl_0_47 rwl_1_47
+ rwl_0_47 cell_2r1w
Xcell_2r1w_1819 vdd_uq17 gnd read_bl_0_35 read_bl_1_35 write_bl_0_35 wwl_0_36 rwl_1_36
+ rwl_0_36 cell_2r1w
Xcell_2r1w_3777 vdd_uq30 gnd read_bl_0_4 read_bl_1_4 write_bl_0_4 wwl_0_62 rwl_1_62
+ rwl_0_62 cell_2r1w
Xcell_2r1w_3722 vdd_uq25 gnd read_bl_0_5 read_bl_1_5 write_bl_0_5 wwl_0_53 rwl_1_53
+ rwl_0_53 cell_2r1w
Xcell_2r1w_3788 vdd_uq24 gnd read_bl_0_4 read_bl_1_4 write_bl_0_4 wwl_0_51 rwl_1_51
+ rwl_0_51 cell_2r1w
Xcell_2r1w_3733 vdd_uq20 gnd read_bl_0_5 read_bl_1_5 write_bl_0_5 wwl_0_42 rwl_1_42
+ rwl_0_42 cell_2r1w
Xcell_2r1w_3799 vdd_uq19 gnd read_bl_0_4 read_bl_1_4 write_bl_0_4 wwl_0_40 rwl_1_40
+ rwl_0_40 cell_2r1w
Xcell_2r1w_3744 vdd_uq14 gnd read_bl_0_5 read_bl_1_5 write_bl_0_5 wwl_0_31 rwl_1_31
+ rwl_0_31 cell_2r1w
Xcell_2r1w_3711 vdd_uq0 gnd read_bl_0_6 read_bl_1_6 write_bl_0_6 wwl_0_0 rwl_1_0 rwl_0_0
+ cell_2r1w
Xcell_2r1w_3766 vdd_uq3 gnd read_bl_0_5 read_bl_1_5 write_bl_0_5 wwl_0_9 rwl_1_9 rwl_0_9
+ cell_2r1w
Xcell_2r1w_3700 vdd_uq4 gnd read_bl_0_6 read_bl_1_6 write_bl_0_6 wwl_0_11 rwl_1_11
+ rwl_0_11 cell_2r1w
Xcell_2r1w_3755 vdd_uq9 gnd read_bl_0_5 read_bl_1_5 write_bl_0_5 wwl_0_20 rwl_1_20
+ rwl_0_20 cell_2r1w
Xcell_2r1w_309 vdd_uq4 gnd read_bl_0_59 read_bl_1_59 write_bl_0_59 wwl_0_10 rwl_1_10
+ rwl_0_10 cell_2r1w
Xcell_2r1w_2306 vdd_uq29 gnd read_bl_0_27 read_bl_1_27 write_bl_0_27 wwl_0_61 rwl_1_61
+ rwl_0_61 cell_2r1w
Xcell_2r1w_1605 vdd_uq28 gnd read_bl_0_38 read_bl_1_38 write_bl_0_38 wwl_0_58 rwl_1_58
+ rwl_0_58 cell_2r1w
Xcell_2r1w_3018 vdd_uq25 gnd read_bl_0_16 read_bl_1_16 write_bl_0_16 wwl_0_53 rwl_1_53
+ rwl_0_53 cell_2r1w
Xcell_2r1w_2317 vdd_uq24 gnd read_bl_0_27 read_bl_1_27 write_bl_0_27 wwl_0_50 rwl_1_50
+ rwl_0_50 cell_2r1w
Xcell_2r1w_1616 vdd_uq22 gnd read_bl_0_38 read_bl_1_38 write_bl_0_38 wwl_0_47 rwl_1_47
+ rwl_0_47 cell_2r1w
Xcell_2r1w_3029 vdd_uq20 gnd read_bl_0_16 read_bl_1_16 write_bl_0_16 wwl_0_42 rwl_1_42
+ rwl_0_42 cell_2r1w
Xcell_2r1w_2328 vdd_uq18 gnd read_bl_0_27 read_bl_1_27 write_bl_0_27 wwl_0_39 rwl_1_39
+ rwl_0_39 cell_2r1w
Xcell_2r1w_1627 vdd_uq17 gnd read_bl_0_38 read_bl_1_38 write_bl_0_38 wwl_0_36 rwl_1_36
+ rwl_0_36 cell_2r1w
Xcell_2r1w_2339 vdd_uq13 gnd read_bl_0_27 read_bl_1_27 write_bl_0_27 wwl_0_28 rwl_1_28
+ rwl_0_28 cell_2r1w
Xcell_2r1w_3007 vdd_uq0 gnd read_bl_0_17 read_bl_1_17 write_bl_0_17 wwl_0_0 rwl_1_0
+ rwl_0_0 cell_2r1w
Xcell_2r1w_832 vdd_uq30 gnd read_bl_0_50 read_bl_1_50 write_bl_0_50 wwl_0_63 rwl_1_63
+ rwl_0_63 cell_2r1w
Xcell_2r1w_898 vdd_uq29 gnd read_bl_0_49 read_bl_1_49 write_bl_0_49 wwl_0_61 rwl_1_61
+ rwl_0_61 cell_2r1w
Xcell_2r1w_843 vdd_uq25 gnd read_bl_0_50 read_bl_1_50 write_bl_0_50 wwl_0_52 rwl_1_52
+ rwl_0_52 cell_2r1w
Xcell_2r1w_854 vdd_uq19 gnd read_bl_0_50 read_bl_1_50 write_bl_0_50 wwl_0_41 rwl_1_41
+ rwl_0_41 cell_2r1w
Xcell_2r1w_865 vdd_uq14 gnd read_bl_0_50 read_bl_1_50 write_bl_0_50 wwl_0_30 rwl_1_30
+ rwl_0_30 cell_2r1w
Xcell_2r1w_1638 vdd_uq11 gnd read_bl_0_38 read_bl_1_38 write_bl_0_38 wwl_0_25 rwl_1_25
+ rwl_0_25 cell_2r1w
Xcell_2r1w_887 vdd_uq3 gnd read_bl_0_50 read_bl_1_50 write_bl_0_50 wwl_0_8 rwl_1_8
+ rwl_0_8 cell_2r1w
Xcell_2r1w_821 vdd_uq4 gnd read_bl_0_51 read_bl_1_51 write_bl_0_51 wwl_0_10 rwl_1_10
+ rwl_0_10 cell_2r1w
Xcell_2r1w_1649 vdd_uq6 gnd read_bl_0_38 read_bl_1_38 write_bl_0_38 wwl_0_14 rwl_1_14
+ rwl_0_14 cell_2r1w
Xcell_2r1w_876 vdd_uq8 gnd read_bl_0_50 read_bl_1_50 write_bl_0_50 wwl_0_19 rwl_1_19
+ rwl_0_19 cell_2r1w
Xcell_2r1w_810 vdd_uq9 gnd read_bl_0_51 read_bl_1_51 write_bl_0_51 wwl_0_21 rwl_1_21
+ rwl_0_21 cell_2r1w
Xcell_2r1w_3585 vdd_uq30 gnd read_bl_0_7 read_bl_1_7 write_bl_0_7 wwl_0_62 rwl_1_62
+ rwl_0_62 cell_2r1w
Xcell_2r1w_2884 vdd_uq28 gnd read_bl_0_18 read_bl_1_18 write_bl_0_18 wwl_0_59 rwl_1_59
+ rwl_0_59 cell_2r1w
Xcell_2r1w_3530 vdd_uq25 gnd read_bl_0_8 read_bl_1_8 write_bl_0_8 wwl_0_53 rwl_1_53
+ rwl_0_53 cell_2r1w
Xcell_2r1w_3596 vdd_uq24 gnd read_bl_0_7 read_bl_1_7 write_bl_0_7 wwl_0_51 rwl_1_51
+ rwl_0_51 cell_2r1w
Xcell_2r1w_2895 vdd_uq23 gnd read_bl_0_18 read_bl_1_18 write_bl_0_18 wwl_0_48 rwl_1_48
+ rwl_0_48 cell_2r1w
Xcell_2r1w_3541 vdd_uq20 gnd read_bl_0_8 read_bl_1_8 write_bl_0_8 wwl_0_42 rwl_1_42
+ rwl_0_42 cell_2r1w
Xcell_2r1w_2840 vdd_uq18 gnd read_bl_0_19 read_bl_1_19 write_bl_0_19 wwl_0_39 rwl_1_39
+ rwl_0_39 cell_2r1w
Xcell_2r1w_3552 vdd_uq14 gnd read_bl_0_8 read_bl_1_8 write_bl_0_8 wwl_0_31 rwl_1_31
+ rwl_0_31 cell_2r1w
Xcell_2r1w_2851 vdd_uq13 gnd read_bl_0_19 read_bl_1_19 write_bl_0_19 wwl_0_28 rwl_1_28
+ rwl_0_28 cell_2r1w
Xcell_2r1w_2873 vdd_uq2 gnd read_bl_0_19 read_bl_1_19 write_bl_0_19 wwl_0_6 rwl_1_6
+ rwl_0_6 cell_2r1w
Xcell_2r1w_3574 vdd_uq3 gnd read_bl_0_8 read_bl_1_8 write_bl_0_8 wwl_0_9 rwl_1_9 rwl_0_9
+ cell_2r1w
Xcell_2r1w_2862 vdd_uq7 gnd read_bl_0_19 read_bl_1_19 write_bl_0_19 wwl_0_17 rwl_1_17
+ rwl_0_17 cell_2r1w
Xcell_2r1w_3563 vdd_uq9 gnd read_bl_0_8 read_bl_1_8 write_bl_0_8 wwl_0_20 rwl_1_20
+ rwl_0_20 cell_2r1w
Xcell_2r1w_128 vdd_uq30 gnd read_bl_0_61 read_bl_1_61 write_bl_0_61 wwl_0_63 rwl_1_63
+ rwl_0_63 cell_2r1w
Xcell_2r1w_139 vdd_uq25 gnd read_bl_0_61 read_bl_1_61 write_bl_0_61 wwl_0_52 rwl_1_52
+ rwl_0_52 cell_2r1w
Xcell_2r1w_117 vdd_uq4 gnd read_bl_0_62 read_bl_1_62 write_bl_0_62 wwl_0_10 rwl_1_10
+ rwl_0_10 cell_2r1w
Xcell_2r1w_106 vdd_uq9 gnd read_bl_0_62 read_bl_1_62 write_bl_0_62 wwl_0_21 rwl_1_21
+ rwl_0_21 cell_2r1w
Xcell_2r1w_2114 vdd_uq29 gnd read_bl_0_30 read_bl_1_30 write_bl_0_30 wwl_0_61 rwl_1_61
+ rwl_0_61 cell_2r1w
Xcell_2r1w_1413 vdd_uq28 gnd read_bl_0_41 read_bl_1_41 write_bl_0_41 wwl_0_58 rwl_1_58
+ rwl_0_58 cell_2r1w
Xcell_2r1w_2125 vdd_uq24 gnd read_bl_0_30 read_bl_1_30 write_bl_0_30 wwl_0_50 rwl_1_50
+ rwl_0_50 cell_2r1w
Xcell_2r1w_1424 vdd_uq22 gnd read_bl_0_41 read_bl_1_41 write_bl_0_41 wwl_0_47 rwl_1_47
+ rwl_0_47 cell_2r1w
Xcell_2r1w_2136 vdd_uq18 gnd read_bl_0_30 read_bl_1_30 write_bl_0_30 wwl_0_39 rwl_1_39
+ rwl_0_39 cell_2r1w
Xcell_2r1w_1435 vdd_uq17 gnd read_bl_0_41 read_bl_1_41 write_bl_0_41 wwl_0_36 rwl_1_36
+ rwl_0_36 cell_2r1w
Xcell_2r1w_2147 vdd_uq13 gnd read_bl_0_30 read_bl_1_30 write_bl_0_30 wwl_0_28 rwl_1_28
+ rwl_0_28 cell_2r1w
Xcell_2r1w_1446 vdd_uq11 gnd read_bl_0_41 read_bl_1_41 write_bl_0_41 wwl_0_25 rwl_1_25
+ rwl_0_25 cell_2r1w
Xcell_2r1w_1402 vdd_uq1 gnd read_bl_0_42 read_bl_1_42 write_bl_0_42 wwl_0_5 rwl_1_5
+ rwl_0_5 cell_2r1w
Xcell_2r1w_1468 vdd gnd read_bl_0_41 read_bl_1_41 write_bl_0_41 wwl_0_3 rwl_1_3 rwl_0_3
+ cell_2r1w
Xcell_2r1w_2169 vdd_uq2 gnd read_bl_0_30 read_bl_1_30 write_bl_0_30 wwl_0_6 rwl_1_6
+ rwl_0_6 cell_2r1w
Xcell_2r1w_2103 vdd_uq3 gnd read_bl_0_31 read_bl_1_31 write_bl_0_31 wwl_0_8 rwl_1_8
+ rwl_0_8 cell_2r1w
Xcell_2r1w_1457 vdd_uq6 gnd read_bl_0_41 read_bl_1_41 write_bl_0_41 wwl_0_14 rwl_1_14
+ rwl_0_14 cell_2r1w
Xcell_2r1w_2158 vdd_uq7 gnd read_bl_0_30 read_bl_1_30 write_bl_0_30 wwl_0_17 rwl_1_17
+ rwl_0_17 cell_2r1w
Xcell_2r1w_640 vdd_uq30 gnd read_bl_0_53 read_bl_1_53 write_bl_0_53 wwl_0_63 rwl_1_63
+ rwl_0_63 cell_2r1w
Xcell_2r1w_1479 vdd_uq27 gnd read_bl_0_40 read_bl_1_40 write_bl_0_40 wwl_0_56 rwl_1_56
+ rwl_0_56 cell_2r1w
Xcell_2r1w_651 vdd_uq25 gnd read_bl_0_53 read_bl_1_53 write_bl_0_53 wwl_0_52 rwl_1_52
+ rwl_0_52 cell_2r1w
Xcell_2r1w_662 vdd_uq19 gnd read_bl_0_53 read_bl_1_53 write_bl_0_53 wwl_0_41 rwl_1_41
+ rwl_0_41 cell_2r1w
Xcell_2r1w_673 vdd_uq14 gnd read_bl_0_53 read_bl_1_53 write_bl_0_53 wwl_0_30 rwl_1_30
+ rwl_0_30 cell_2r1w
Xcell_2r1w_695 vdd_uq3 gnd read_bl_0_53 read_bl_1_53 write_bl_0_53 wwl_0_8 rwl_1_8
+ rwl_0_8 cell_2r1w
Xcell_2r1w_684 vdd_uq8 gnd read_bl_0_53 read_bl_1_53 write_bl_0_53 wwl_0_19 rwl_1_19
+ rwl_0_19 cell_2r1w
Xcell_2r1w_4050 vdd_uq21 gnd read_bl_0_0 read_bl_1_0 write_bl_0_0 wwl_0_45 rwl_1_45
+ rwl_0_45 cell_2r1w
Xcell_2r1w_4061 vdd_uq16 gnd read_bl_0_0 read_bl_1_0 write_bl_0_0 wwl_0_34 rwl_1_34
+ rwl_0_34 cell_2r1w
Xcell_2r1w_3360 vdd_uq14 gnd read_bl_0_11 read_bl_1_11 write_bl_0_11 wwl_0_31 rwl_1_31
+ rwl_0_31 cell_2r1w
Xcell_2r1w_4094 vdd_uq0 gnd read_bl_0_0 read_bl_1_0 write_bl_0_0 wwl_0_1 rwl_1_1 rwl_0_1
+ cell_2r1w
Xcell_2r1w_4083 vdd_uq5 gnd read_bl_0_0 read_bl_1_0 write_bl_0_0 wwl_0_12 rwl_1_12
+ rwl_0_12 cell_2r1w
Xcell_2r1w_3371 vdd_uq9 gnd read_bl_0_11 read_bl_1_11 write_bl_0_11 wwl_0_20 rwl_1_20
+ rwl_0_20 cell_2r1w
Xcell_2r1w_4072 vdd_uq10 gnd read_bl_0_0 read_bl_1_0 write_bl_0_0 wwl_0_23 rwl_1_23
+ rwl_0_23 cell_2r1w
Xcell_2r1w_3393 vdd_uq30 gnd read_bl_0_10 read_bl_1_10 write_bl_0_10 wwl_0_62 rwl_1_62
+ rwl_0_62 cell_2r1w
Xcell_2r1w_2692 vdd_uq28 gnd read_bl_0_21 read_bl_1_21 write_bl_0_21 wwl_0_59 rwl_1_59
+ rwl_0_59 cell_2r1w
Xcell_2r1w_1991 vdd_uq27 gnd read_bl_0_32 read_bl_1_32 write_bl_0_32 wwl_0_56 rwl_1_56
+ rwl_0_56 cell_2r1w
Xcell_2r1w_1980 vdd gnd read_bl_0_33 read_bl_1_33 write_bl_0_33 wwl_0_3 rwl_1_3 rwl_0_3
+ cell_2r1w
Xcell_2r1w_2681 vdd_uq2 gnd read_bl_0_22 read_bl_1_22 write_bl_0_22 wwl_0_6 rwl_1_6
+ rwl_0_6 cell_2r1w
Xcell_2r1w_3382 vdd_uq3 gnd read_bl_0_11 read_bl_1_11 write_bl_0_11 wwl_0_9 rwl_1_9
+ rwl_0_9 cell_2r1w
Xcell_2r1w_2670 vdd_uq7 gnd read_bl_0_22 read_bl_1_22 write_bl_0_22 wwl_0_17 rwl_1_17
+ rwl_0_17 cell_2r1w
Xcell_2r1w_1221 vdd_uq28 gnd read_bl_0_44 read_bl_1_44 write_bl_0_44 wwl_0_58 rwl_1_58
+ rwl_0_58 cell_2r1w
Xcell_2r1w_1287 vdd_uq27 gnd read_bl_0_43 read_bl_1_43 write_bl_0_43 wwl_0_56 rwl_1_56
+ rwl_0_56 cell_2r1w
Xcell_2r1w_1232 vdd_uq22 gnd read_bl_0_44 read_bl_1_44 write_bl_0_44 wwl_0_47 rwl_1_47
+ rwl_0_47 cell_2r1w
Xcell_2r1w_1298 vdd_uq21 gnd read_bl_0_43 read_bl_1_43 write_bl_0_43 wwl_0_45 rwl_1_45
+ rwl_0_45 cell_2r1w
Xcell_2r1w_470 vdd_uq19 gnd read_bl_0_56 read_bl_1_56 write_bl_0_56 wwl_0_41 rwl_1_41
+ rwl_0_41 cell_2r1w
Xcell_2r1w_1243 vdd_uq17 gnd read_bl_0_44 read_bl_1_44 write_bl_0_44 wwl_0_36 rwl_1_36
+ rwl_0_36 cell_2r1w
Xcell_2r1w_481 vdd_uq14 gnd read_bl_0_56 read_bl_1_56 write_bl_0_56 wwl_0_30 rwl_1_30
+ rwl_0_30 cell_2r1w
Xcell_2r1w_1254 vdd_uq11 gnd read_bl_0_44 read_bl_1_44 write_bl_0_44 wwl_0_25 rwl_1_25
+ rwl_0_25 cell_2r1w
Xcell_2r1w_1210 vdd_uq1 gnd read_bl_0_45 read_bl_1_45 write_bl_0_45 wwl_0_5 rwl_1_5
+ rwl_0_5 cell_2r1w
Xcell_2r1w_1276 vdd gnd read_bl_0_44 read_bl_1_44 write_bl_0_44 wwl_0_3 rwl_1_3 rwl_0_3
+ cell_2r1w
Xcell_2r1w_1265 vdd_uq6 gnd read_bl_0_44 read_bl_1_44 write_bl_0_44 wwl_0_14 rwl_1_14
+ rwl_0_14 cell_2r1w
Xcell_2r1w_492 vdd_uq8 gnd read_bl_0_56 read_bl_1_56 write_bl_0_56 wwl_0_19 rwl_1_19
+ rwl_0_19 cell_2r1w
Xcell_2r1w_3190 vdd_uq3 gnd read_bl_0_14 read_bl_1_14 write_bl_0_14 wwl_0_9 rwl_1_9
+ rwl_0_9 cell_2r1w
Xcell_2r1w_1095 vdd_uq27 gnd read_bl_0_46 read_bl_1_46 write_bl_0_46 wwl_0_56 rwl_1_56
+ rwl_0_56 cell_2r1w
Xcell_2r1w_1040 vdd_uq22 gnd read_bl_0_47 read_bl_1_47 write_bl_0_47 wwl_0_47 rwl_1_47
+ rwl_0_47 cell_2r1w
Xcell_2r1w_1051 vdd_uq17 gnd read_bl_0_47 read_bl_1_47 write_bl_0_47 wwl_0_36 rwl_1_36
+ rwl_0_36 cell_2r1w
Xcell_2r1w_1062 vdd_uq11 gnd read_bl_0_47 read_bl_1_47 write_bl_0_47 wwl_0_25 rwl_1_25
+ rwl_0_25 cell_2r1w
Xcell_2r1w_1084 vdd gnd read_bl_0_47 read_bl_1_47 write_bl_0_47 wwl_0_3 rwl_1_3 rwl_0_3
+ cell_2r1w
Xcell_2r1w_1073 vdd_uq6 gnd read_bl_0_47 read_bl_1_47 write_bl_0_47 wwl_0_14 rwl_1_14
+ rwl_0_14 cell_2r1w
Xcell_2r1w_3904 vdd_uq30 gnd read_bl_0_2 read_bl_1_2 write_bl_0_2 wwl_0_63 rwl_1_63
+ rwl_0_63 cell_2r1w
Xcell_2r1w_3915 vdd_uq25 gnd read_bl_0_2 read_bl_1_2 write_bl_0_2 wwl_0_52 rwl_1_52
+ rwl_0_52 cell_2r1w
Xcell_2r1w_3926 vdd_uq19 gnd read_bl_0_2 read_bl_1_2 write_bl_0_2 wwl_0_41 rwl_1_41
+ rwl_0_41 cell_2r1w
Xcell_2r1w_3937 vdd_uq14 gnd read_bl_0_2 read_bl_1_2 write_bl_0_2 wwl_0_30 rwl_1_30
+ rwl_0_30 cell_2r1w
Xcell_2r1w_3959 vdd_uq3 gnd read_bl_0_2 read_bl_1_2 write_bl_0_2 wwl_0_8 rwl_1_8 rwl_0_8
+ cell_2r1w
Xcell_2r1w_3948 vdd_uq8 gnd read_bl_0_2 read_bl_1_2 write_bl_0_2 wwl_0_19 rwl_1_19
+ rwl_0_19 cell_2r1w
Xcell_2r1w_1809 vdd_uq22 gnd read_bl_0_35 read_bl_1_35 write_bl_0_35 wwl_0_46 rwl_1_46
+ rwl_0_46 cell_2r1w
Xcell_2r1w_3712 vdd_uq30 gnd read_bl_0_5 read_bl_1_5 write_bl_0_5 wwl_0_63 rwl_1_63
+ rwl_0_63 cell_2r1w
Xcell_2r1w_3701 vdd_uq4 gnd read_bl_0_6 read_bl_1_6 write_bl_0_6 wwl_0_10 rwl_1_10
+ rwl_0_10 cell_2r1w
Xcell_2r1w_3778 vdd_uq29 gnd read_bl_0_4 read_bl_1_4 write_bl_0_4 wwl_0_61 rwl_1_61
+ rwl_0_61 cell_2r1w
Xcell_2r1w_3723 vdd_uq25 gnd read_bl_0_5 read_bl_1_5 write_bl_0_5 wwl_0_52 rwl_1_52
+ rwl_0_52 cell_2r1w
Xcell_2r1w_3789 vdd_uq24 gnd read_bl_0_4 read_bl_1_4 write_bl_0_4 wwl_0_50 rwl_1_50
+ rwl_0_50 cell_2r1w
Xcell_2r1w_3734 vdd_uq19 gnd read_bl_0_5 read_bl_1_5 write_bl_0_5 wwl_0_41 rwl_1_41
+ rwl_0_41 cell_2r1w
Xcell_2r1w_3745 vdd_uq14 gnd read_bl_0_5 read_bl_1_5 write_bl_0_5 wwl_0_30 rwl_1_30
+ rwl_0_30 cell_2r1w
Xcell_2r1w_3767 vdd_uq3 gnd read_bl_0_5 read_bl_1_5 write_bl_0_5 wwl_0_8 rwl_1_8 rwl_0_8
+ cell_2r1w
Xcell_2r1w_3756 vdd_uq8 gnd read_bl_0_5 read_bl_1_5 write_bl_0_5 wwl_0_19 rwl_1_19
+ rwl_0_19 cell_2r1w
Xcell_2r1w_3008 vdd_uq30 gnd read_bl_0_16 read_bl_1_16 write_bl_0_16 wwl_0_63 rwl_1_63
+ rwl_0_63 cell_2r1w
Xcell_2r1w_2307 vdd_uq29 gnd read_bl_0_27 read_bl_1_27 write_bl_0_27 wwl_0_60 rwl_1_60
+ rwl_0_60 cell_2r1w
Xcell_2r1w_1606 vdd_uq27 gnd read_bl_0_38 read_bl_1_38 write_bl_0_38 wwl_0_57 rwl_1_57
+ rwl_0_57 cell_2r1w
Xcell_2r1w_3019 vdd_uq25 gnd read_bl_0_16 read_bl_1_16 write_bl_0_16 wwl_0_52 rwl_1_52
+ rwl_0_52 cell_2r1w
Xcell_2r1w_2318 vdd_uq23 gnd read_bl_0_27 read_bl_1_27 write_bl_0_27 wwl_0_49 rwl_1_49
+ rwl_0_49 cell_2r1w
Xcell_2r1w_1617 vdd_uq22 gnd read_bl_0_38 read_bl_1_38 write_bl_0_38 wwl_0_46 rwl_1_46
+ rwl_0_46 cell_2r1w
Xcell_2r1w_2329 vdd_uq18 gnd read_bl_0_27 read_bl_1_27 write_bl_0_27 wwl_0_38 rwl_1_38
+ rwl_0_38 cell_2r1w
Xcell_2r1w_1628 vdd_uq16 gnd read_bl_0_38 read_bl_1_38 write_bl_0_38 wwl_0_35 rwl_1_35
+ rwl_0_35 cell_2r1w
Xcell_2r1w_800 vdd_uq14 gnd read_bl_0_51 read_bl_1_51 write_bl_0_51 wwl_0_31 rwl_1_31
+ rwl_0_31 cell_2r1w
Xcell_2r1w_1639 vdd_uq11 gnd read_bl_0_38 read_bl_1_38 write_bl_0_38 wwl_0_24 rwl_1_24
+ rwl_0_24 cell_2r1w
Xcell_2r1w_822 vdd_uq3 gnd read_bl_0_51 read_bl_1_51 write_bl_0_51 wwl_0_9 rwl_1_9
+ rwl_0_9 cell_2r1w
Xcell_2r1w_811 vdd_uq9 gnd read_bl_0_51 read_bl_1_51 write_bl_0_51 wwl_0_20 rwl_1_20
+ rwl_0_20 cell_2r1w
Xcell_2r1w_833 vdd_uq30 gnd read_bl_0_50 read_bl_1_50 write_bl_0_50 wwl_0_62 rwl_1_62
+ rwl_0_62 cell_2r1w
Xcell_2r1w_899 vdd_uq29 gnd read_bl_0_49 read_bl_1_49 write_bl_0_49 wwl_0_60 rwl_1_60
+ rwl_0_60 cell_2r1w
Xcell_2r1w_844 vdd_uq24 gnd read_bl_0_50 read_bl_1_50 write_bl_0_50 wwl_0_51 rwl_1_51
+ rwl_0_51 cell_2r1w
Xcell_2r1w_855 vdd_uq19 gnd read_bl_0_50 read_bl_1_50 write_bl_0_50 wwl_0_40 rwl_1_40
+ rwl_0_40 cell_2r1w
Xcell_2r1w_866 vdd_uq13 gnd read_bl_0_50 read_bl_1_50 write_bl_0_50 wwl_0_29 rwl_1_29
+ rwl_0_29 cell_2r1w
Xcell_2r1w_888 vdd_uq2 gnd read_bl_0_50 read_bl_1_50 write_bl_0_50 wwl_0_7 rwl_1_7
+ rwl_0_7 cell_2r1w
Xcell_2r1w_877 vdd_uq8 gnd read_bl_0_50 read_bl_1_50 write_bl_0_50 wwl_0_18 rwl_1_18
+ rwl_0_18 cell_2r1w
Xcell_2r1w_3520 vdd_uq30 gnd read_bl_0_8 read_bl_1_8 write_bl_0_8 wwl_0_63 rwl_1_63
+ rwl_0_63 cell_2r1w
Xcell_2r1w_3531 vdd_uq25 gnd read_bl_0_8 read_bl_1_8 write_bl_0_8 wwl_0_52 rwl_1_52
+ rwl_0_52 cell_2r1w
Xcell_2r1w_3542 vdd_uq19 gnd read_bl_0_8 read_bl_1_8 write_bl_0_8 wwl_0_41 rwl_1_41
+ rwl_0_41 cell_2r1w
Xcell_2r1w_3553 vdd_uq14 gnd read_bl_0_8 read_bl_1_8 write_bl_0_8 wwl_0_30 rwl_1_30
+ rwl_0_30 cell_2r1w
Xcell_2r1w_3586 vdd_uq29 gnd read_bl_0_7 read_bl_1_7 write_bl_0_7 wwl_0_61 rwl_1_61
+ rwl_0_61 cell_2r1w
Xcell_2r1w_2885 vdd_uq28 gnd read_bl_0_18 read_bl_1_18 write_bl_0_18 wwl_0_58 rwl_1_58
+ rwl_0_58 cell_2r1w
Xcell_2r1w_3597 vdd_uq24 gnd read_bl_0_7 read_bl_1_7 write_bl_0_7 wwl_0_50 rwl_1_50
+ rwl_0_50 cell_2r1w
Xcell_2r1w_2830 vdd_uq23 gnd read_bl_0_19 read_bl_1_19 write_bl_0_19 wwl_0_49 rwl_1_49
+ rwl_0_49 cell_2r1w
Xcell_2r1w_2896 vdd_uq22 gnd read_bl_0_18 read_bl_1_18 write_bl_0_18 wwl_0_47 rwl_1_47
+ rwl_0_47 cell_2r1w
Xcell_2r1w_2841 vdd_uq18 gnd read_bl_0_19 read_bl_1_19 write_bl_0_19 wwl_0_38 rwl_1_38
+ rwl_0_38 cell_2r1w
Xcell_2r1w_2852 vdd_uq12 gnd read_bl_0_19 read_bl_1_19 write_bl_0_19 wwl_0_27 rwl_1_27
+ rwl_0_27 cell_2r1w
Xcell_2r1w_2874 vdd_uq1 gnd read_bl_0_19 read_bl_1_19 write_bl_0_19 wwl_0_5 rwl_1_5
+ rwl_0_5 cell_2r1w
Xcell_2r1w_3575 vdd_uq3 gnd read_bl_0_8 read_bl_1_8 write_bl_0_8 wwl_0_8 rwl_1_8 rwl_0_8
+ cell_2r1w
Xcell_2r1w_2863 vdd_uq7 gnd read_bl_0_19 read_bl_1_19 write_bl_0_19 wwl_0_16 rwl_1_16
+ rwl_0_16 cell_2r1w
Xcell_2r1w_3564 vdd_uq8 gnd read_bl_0_8 read_bl_1_8 write_bl_0_8 wwl_0_19 rwl_1_19
+ rwl_0_19 cell_2r1w
Xcell_2r1w_107 vdd_uq9 gnd read_bl_0_62 read_bl_1_62 write_bl_0_62 wwl_0_20 rwl_1_20
+ rwl_0_20 cell_2r1w
Xcell_2r1w_129 vdd_uq30 gnd read_bl_0_61 read_bl_1_61 write_bl_0_61 wwl_0_62 rwl_1_62
+ rwl_0_62 cell_2r1w
Xcell_2r1w_118 vdd_uq3 gnd read_bl_0_62 read_bl_1_62 write_bl_0_62 wwl_0_9 rwl_1_9
+ rwl_0_9 cell_2r1w
Xcell_2r1w_2104 vdd_uq2 gnd read_bl_0_31 read_bl_1_31 write_bl_0_31 wwl_0_7 rwl_1_7
+ rwl_0_7 cell_2r1w
Xcell_2r1w_641 vdd_uq30 gnd read_bl_0_53 read_bl_1_53 write_bl_0_53 wwl_0_62 rwl_1_62
+ rwl_0_62 cell_2r1w
Xcell_2r1w_2115 vdd_uq29 gnd read_bl_0_30 read_bl_1_30 write_bl_0_30 wwl_0_60 rwl_1_60
+ rwl_0_60 cell_2r1w
Xcell_2r1w_1414 vdd_uq27 gnd read_bl_0_41 read_bl_1_41 write_bl_0_41 wwl_0_57 rwl_1_57
+ rwl_0_57 cell_2r1w
Xcell_2r1w_652 vdd_uq24 gnd read_bl_0_53 read_bl_1_53 write_bl_0_53 wwl_0_51 rwl_1_51
+ rwl_0_51 cell_2r1w
Xcell_2r1w_2126 vdd_uq23 gnd read_bl_0_30 read_bl_1_30 write_bl_0_30 wwl_0_49 rwl_1_49
+ rwl_0_49 cell_2r1w
Xcell_2r1w_1425 vdd_uq22 gnd read_bl_0_41 read_bl_1_41 write_bl_0_41 wwl_0_46 rwl_1_46
+ rwl_0_46 cell_2r1w
Xcell_2r1w_663 vdd_uq19 gnd read_bl_0_53 read_bl_1_53 write_bl_0_53 wwl_0_40 rwl_1_40
+ rwl_0_40 cell_2r1w
Xcell_2r1w_2137 vdd_uq18 gnd read_bl_0_30 read_bl_1_30 write_bl_0_30 wwl_0_38 rwl_1_38
+ rwl_0_38 cell_2r1w
Xcell_2r1w_1436 vdd_uq16 gnd read_bl_0_41 read_bl_1_41 write_bl_0_41 wwl_0_35 rwl_1_35
+ rwl_0_35 cell_2r1w
Xcell_2r1w_2148 vdd_uq12 gnd read_bl_0_30 read_bl_1_30 write_bl_0_30 wwl_0_27 rwl_1_27
+ rwl_0_27 cell_2r1w
Xcell_2r1w_1447 vdd_uq11 gnd read_bl_0_41 read_bl_1_41 write_bl_0_41 wwl_0_24 rwl_1_24
+ rwl_0_24 cell_2r1w
Xcell_2r1w_1403 vdd_uq1 gnd read_bl_0_42 read_bl_1_42 write_bl_0_42 wwl_0_4 rwl_1_4
+ rwl_0_4 cell_2r1w
Xcell_2r1w_1469 vdd gnd read_bl_0_41 read_bl_1_41 write_bl_0_41 wwl_0_2 rwl_1_2 rwl_0_2
+ cell_2r1w
Xcell_2r1w_630 vdd_uq3 gnd read_bl_0_54 read_bl_1_54 write_bl_0_54 wwl_0_9 rwl_1_9
+ rwl_0_9 cell_2r1w
Xcell_2r1w_1458 vdd_uq5 gnd read_bl_0_41 read_bl_1_41 write_bl_0_41 wwl_0_13 rwl_1_13
+ rwl_0_13 cell_2r1w
Xcell_2r1w_2159 vdd_uq7 gnd read_bl_0_30 read_bl_1_30 write_bl_0_30 wwl_0_16 rwl_1_16
+ rwl_0_16 cell_2r1w
Xcell_2r1w_674 vdd_uq13 gnd read_bl_0_53 read_bl_1_53 write_bl_0_53 wwl_0_29 rwl_1_29
+ rwl_0_29 cell_2r1w
Xcell_2r1w_696 vdd_uq2 gnd read_bl_0_53 read_bl_1_53 write_bl_0_53 wwl_0_7 rwl_1_7
+ rwl_0_7 cell_2r1w
Xcell_2r1w_685 vdd_uq8 gnd read_bl_0_53 read_bl_1_53 write_bl_0_53 wwl_0_18 rwl_1_18
+ rwl_0_18 cell_2r1w
Xcell_2r1w_3394 vdd_uq29 gnd read_bl_0_10 read_bl_1_10 write_bl_0_10 wwl_0_61 rwl_1_61
+ rwl_0_61 cell_2r1w
Xcell_2r1w_4040 vdd_uq26 gnd read_bl_0_0 read_bl_1_0 write_bl_0_0 wwl_0_55 rwl_1_55
+ rwl_0_55 cell_2r1w
Xcell_2r1w_4051 vdd_uq21 gnd read_bl_0_0 read_bl_1_0 write_bl_0_0 wwl_0_44 rwl_1_44
+ rwl_0_44 cell_2r1w
Xcell_2r1w_3350 vdd_uq19 gnd read_bl_0_11 read_bl_1_11 write_bl_0_11 wwl_0_41 rwl_1_41
+ rwl_0_41 cell_2r1w
Xcell_2r1w_4062 vdd_uq15 gnd read_bl_0_0 read_bl_1_0 write_bl_0_0 wwl_0_33 rwl_1_33
+ rwl_0_33 cell_2r1w
Xcell_2r1w_3361 vdd_uq14 gnd read_bl_0_11 read_bl_1_11 write_bl_0_11 wwl_0_30 rwl_1_30
+ rwl_0_30 cell_2r1w
Xcell_2r1w_2660 vdd_uq12 gnd read_bl_0_22 read_bl_1_22 write_bl_0_22 wwl_0_27 rwl_1_27
+ rwl_0_27 cell_2r1w
Xcell_2r1w_4095 vdd_uq0 gnd read_bl_0_0 read_bl_1_0 write_bl_0_0 wwl_0_0 rwl_1_0 rwl_0_0
+ cell_2r1w
Xcell_2r1w_3383 vdd_uq3 gnd read_bl_0_11 read_bl_1_11 write_bl_0_11 wwl_0_8 rwl_1_8
+ rwl_0_8 cell_2r1w
Xcell_2r1w_4084 vdd_uq4 gnd read_bl_0_0 read_bl_1_0 write_bl_0_0 wwl_0_11 rwl_1_11
+ rwl_0_11 cell_2r1w
Xcell_2r1w_3372 vdd_uq8 gnd read_bl_0_11 read_bl_1_11 write_bl_0_11 wwl_0_19 rwl_1_19
+ rwl_0_19 cell_2r1w
Xcell_2r1w_4073 vdd_uq10 gnd read_bl_0_0 read_bl_1_0 write_bl_0_0 wwl_0_22 rwl_1_22
+ rwl_0_22 cell_2r1w
Xcell_2r1w_2693 vdd_uq28 gnd read_bl_0_21 read_bl_1_21 write_bl_0_21 wwl_0_58 rwl_1_58
+ rwl_0_58 cell_2r1w
Xcell_2r1w_1992 vdd_uq26 gnd read_bl_0_32 read_bl_1_32 write_bl_0_32 wwl_0_55 rwl_1_55
+ rwl_0_55 cell_2r1w
Xcell_2r1w_2682 vdd_uq1 gnd read_bl_0_22 read_bl_1_22 write_bl_0_22 wwl_0_5 rwl_1_5
+ rwl_0_5 cell_2r1w
Xcell_2r1w_1981 vdd gnd read_bl_0_33 read_bl_1_33 write_bl_0_33 wwl_0_2 rwl_1_2 rwl_0_2
+ cell_2r1w
Xcell_2r1w_1970 vdd_uq5 gnd read_bl_0_33 read_bl_1_33 write_bl_0_33 wwl_0_13 rwl_1_13
+ rwl_0_13 cell_2r1w
Xcell_2r1w_2671 vdd_uq7 gnd read_bl_0_22 read_bl_1_22 write_bl_0_22 wwl_0_16 rwl_1_16
+ rwl_0_16 cell_2r1w
Xcell_2r1w_1211 vdd_uq1 gnd read_bl_0_45 read_bl_1_45 write_bl_0_45 wwl_0_4 rwl_1_4
+ rwl_0_4 cell_2r1w
Xcell_2r1w_1200 vdd_uq6 gnd read_bl_0_45 read_bl_1_45 write_bl_0_45 wwl_0_15 rwl_1_15
+ rwl_0_15 cell_2r1w
Xcell_2r1w_1222 vdd_uq27 gnd read_bl_0_44 read_bl_1_44 write_bl_0_44 wwl_0_57 rwl_1_57
+ rwl_0_57 cell_2r1w
Xcell_2r1w_1288 vdd_uq26 gnd read_bl_0_43 read_bl_1_43 write_bl_0_43 wwl_0_55 rwl_1_55
+ rwl_0_55 cell_2r1w
Xcell_2r1w_460 vdd_uq24 gnd read_bl_0_56 read_bl_1_56 write_bl_0_56 wwl_0_51 rwl_1_51
+ rwl_0_51 cell_2r1w
Xcell_2r1w_1233 vdd_uq22 gnd read_bl_0_44 read_bl_1_44 write_bl_0_44 wwl_0_46 rwl_1_46
+ rwl_0_46 cell_2r1w
Xcell_2r1w_1299 vdd_uq21 gnd read_bl_0_43 read_bl_1_43 write_bl_0_43 wwl_0_44 rwl_1_44
+ rwl_0_44 cell_2r1w
Xcell_2r1w_471 vdd_uq19 gnd read_bl_0_56 read_bl_1_56 write_bl_0_56 wwl_0_40 rwl_1_40
+ rwl_0_40 cell_2r1w
Xcell_2r1w_1244 vdd_uq16 gnd read_bl_0_44 read_bl_1_44 write_bl_0_44 wwl_0_35 rwl_1_35
+ rwl_0_35 cell_2r1w
Xcell_2r1w_482 vdd_uq13 gnd read_bl_0_56 read_bl_1_56 write_bl_0_56 wwl_0_29 rwl_1_29
+ rwl_0_29 cell_2r1w
Xcell_2r1w_1255 vdd_uq11 gnd read_bl_0_44 read_bl_1_44 write_bl_0_44 wwl_0_24 rwl_1_24
+ rwl_0_24 cell_2r1w
Xcell_2r1w_1277 vdd gnd read_bl_0_44 read_bl_1_44 write_bl_0_44 wwl_0_2 rwl_1_2 rwl_0_2
+ cell_2r1w
Xcell_2r1w_1266 vdd_uq5 gnd read_bl_0_44 read_bl_1_44 write_bl_0_44 wwl_0_13 rwl_1_13
+ rwl_0_13 cell_2r1w
Xcell_2r1w_493 vdd_uq8 gnd read_bl_0_56 read_bl_1_56 write_bl_0_56 wwl_0_18 rwl_1_18
+ rwl_0_18 cell_2r1w
Xcell_2r1w_2490 vdd_uq1 gnd read_bl_0_25 read_bl_1_25 write_bl_0_25 wwl_0_5 rwl_1_5
+ rwl_0_5 cell_2r1w
Xcell_2r1w_3191 vdd_uq3 gnd read_bl_0_14 read_bl_1_14 write_bl_0_14 wwl_0_8 rwl_1_8
+ rwl_0_8 cell_2r1w
Xcell_2r1w_3180 vdd_uq8 gnd read_bl_0_14 read_bl_1_14 write_bl_0_14 wwl_0_19 rwl_1_19
+ rwl_0_19 cell_2r1w
Xcell_2r1w_1030 vdd_uq27 gnd read_bl_0_47 read_bl_1_47 write_bl_0_47 wwl_0_57 rwl_1_57
+ rwl_0_57 cell_2r1w
Xcell_2r1w_1041 vdd_uq22 gnd read_bl_0_47 read_bl_1_47 write_bl_0_47 wwl_0_46 rwl_1_46
+ rwl_0_46 cell_2r1w
Xcell_2r1w_1052 vdd_uq16 gnd read_bl_0_47 read_bl_1_47 write_bl_0_47 wwl_0_35 rwl_1_35
+ rwl_0_35 cell_2r1w
Xcell_2r1w_1096 vdd_uq26 gnd read_bl_0_46 read_bl_1_46 write_bl_0_46 wwl_0_55 rwl_1_55
+ rwl_0_55 cell_2r1w
Xcell_2r1w_290 vdd_uq13 gnd read_bl_0_59 read_bl_1_59 write_bl_0_59 wwl_0_29 rwl_1_29
+ rwl_0_29 cell_2r1w
Xcell_2r1w_1063 vdd_uq11 gnd read_bl_0_47 read_bl_1_47 write_bl_0_47 wwl_0_24 rwl_1_24
+ rwl_0_24 cell_2r1w
Xcell_2r1w_1085 vdd gnd read_bl_0_47 read_bl_1_47 write_bl_0_47 wwl_0_2 rwl_1_2 rwl_0_2
+ cell_2r1w
Xcell_2r1w_1074 vdd_uq5 gnd read_bl_0_47 read_bl_1_47 write_bl_0_47 wwl_0_13 rwl_1_13
+ rwl_0_13 cell_2r1w
Xcell_2r1w_3905 vdd_uq30 gnd read_bl_0_2 read_bl_1_2 write_bl_0_2 wwl_0_62 rwl_1_62
+ rwl_0_62 cell_2r1w
Xcell_2r1w_3916 vdd_uq24 gnd read_bl_0_2 read_bl_1_2 write_bl_0_2 wwl_0_51 rwl_1_51
+ rwl_0_51 cell_2r1w
Xcell_2r1w_3927 vdd_uq19 gnd read_bl_0_2 read_bl_1_2 write_bl_0_2 wwl_0_40 rwl_1_40
+ rwl_0_40 cell_2r1w
Xcell_2r1w_3938 vdd_uq13 gnd read_bl_0_2 read_bl_1_2 write_bl_0_2 wwl_0_29 rwl_1_29
+ rwl_0_29 cell_2r1w
Xcell_2r1w_3949 vdd_uq8 gnd read_bl_0_2 read_bl_1_2 write_bl_0_2 wwl_0_18 rwl_1_18
+ rwl_0_18 cell_2r1w
Xcell_2r1w_3713 vdd_uq30 gnd read_bl_0_5 read_bl_1_5 write_bl_0_5 wwl_0_62 rwl_1_62
+ rwl_0_62 cell_2r1w
Xcell_2r1w_3724 vdd_uq24 gnd read_bl_0_5 read_bl_1_5 write_bl_0_5 wwl_0_51 rwl_1_51
+ rwl_0_51 cell_2r1w
Xcell_2r1w_3735 vdd_uq19 gnd read_bl_0_5 read_bl_1_5 write_bl_0_5 wwl_0_40 rwl_1_40
+ rwl_0_40 cell_2r1w
Xcell_2r1w_3702 vdd_uq3 gnd read_bl_0_6 read_bl_1_6 write_bl_0_6 wwl_0_9 rwl_1_9 rwl_0_9
+ cell_2r1w
Xcell_2r1w_3779 vdd_uq29 gnd read_bl_0_4 read_bl_1_4 write_bl_0_4 wwl_0_60 rwl_1_60
+ rwl_0_60 cell_2r1w
Xcell_2r1w_3746 vdd_uq13 gnd read_bl_0_5 read_bl_1_5 write_bl_0_5 wwl_0_29 rwl_1_29
+ rwl_0_29 cell_2r1w
Xcell_2r1w_3768 vdd_uq2 gnd read_bl_0_5 read_bl_1_5 write_bl_0_5 wwl_0_7 rwl_1_7 rwl_0_7
+ cell_2r1w
Xcell_2r1w_3757 vdd_uq8 gnd read_bl_0_5 read_bl_1_5 write_bl_0_5 wwl_0_18 rwl_1_18
+ rwl_0_18 cell_2r1w
Xcell_2r1w_3009 vdd_uq30 gnd read_bl_0_16 read_bl_1_16 write_bl_0_16 wwl_0_62 rwl_1_62
+ rwl_0_62 cell_2r1w
Xcell_2r1w_834 vdd_uq29 gnd read_bl_0_50 read_bl_1_50 write_bl_0_50 wwl_0_61 rwl_1_61
+ rwl_0_61 cell_2r1w
Xcell_2r1w_2308 vdd_uq28 gnd read_bl_0_27 read_bl_1_27 write_bl_0_27 wwl_0_59 rwl_1_59
+ rwl_0_59 cell_2r1w
Xcell_2r1w_1607 vdd_uq27 gnd read_bl_0_38 read_bl_1_38 write_bl_0_38 wwl_0_56 rwl_1_56
+ rwl_0_56 cell_2r1w
Xcell_2r1w_845 vdd_uq24 gnd read_bl_0_50 read_bl_1_50 write_bl_0_50 wwl_0_50 rwl_1_50
+ rwl_0_50 cell_2r1w
Xcell_2r1w_2319 vdd_uq23 gnd read_bl_0_27 read_bl_1_27 write_bl_0_27 wwl_0_48 rwl_1_48
+ rwl_0_48 cell_2r1w
Xcell_2r1w_1618 vdd_uq21 gnd read_bl_0_38 read_bl_1_38 write_bl_0_38 wwl_0_45 rwl_1_45
+ rwl_0_45 cell_2r1w
Xcell_2r1w_1629 vdd_uq16 gnd read_bl_0_38 read_bl_1_38 write_bl_0_38 wwl_0_34 rwl_1_34
+ rwl_0_34 cell_2r1w
Xcell_2r1w_801 vdd_uq14 gnd read_bl_0_51 read_bl_1_51 write_bl_0_51 wwl_0_30 rwl_1_30
+ rwl_0_30 cell_2r1w
Xcell_2r1w_823 vdd_uq3 gnd read_bl_0_51 read_bl_1_51 write_bl_0_51 wwl_0_8 rwl_1_8
+ rwl_0_8 cell_2r1w
Xcell_2r1w_812 vdd_uq8 gnd read_bl_0_51 read_bl_1_51 write_bl_0_51 wwl_0_19 rwl_1_19
+ rwl_0_19 cell_2r1w
Xcell_2r1w_856 vdd_uq18 gnd read_bl_0_50 read_bl_1_50 write_bl_0_50 wwl_0_39 rwl_1_39
+ rwl_0_39 cell_2r1w
Xcell_2r1w_867 vdd_uq13 gnd read_bl_0_50 read_bl_1_50 write_bl_0_50 wwl_0_28 rwl_1_28
+ rwl_0_28 cell_2r1w
Xcell_2r1w_889 vdd_uq2 gnd read_bl_0_50 read_bl_1_50 write_bl_0_50 wwl_0_6 rwl_1_6
+ rwl_0_6 cell_2r1w
Xcell_2r1w_878 vdd_uq7 gnd read_bl_0_50 read_bl_1_50 write_bl_0_50 wwl_0_17 rwl_1_17
+ rwl_0_17 cell_2r1w
Xcell_2r1w_3521 vdd_uq30 gnd read_bl_0_8 read_bl_1_8 write_bl_0_8 wwl_0_62 rwl_1_62
+ rwl_0_62 cell_2r1w
Xcell_2r1w_3587 vdd_uq29 gnd read_bl_0_7 read_bl_1_7 write_bl_0_7 wwl_0_60 rwl_1_60
+ rwl_0_60 cell_2r1w
Xcell_2r1w_2820 vdd_uq28 gnd read_bl_0_19 read_bl_1_19 write_bl_0_19 wwl_0_59 rwl_1_59
+ rwl_0_59 cell_2r1w
Xcell_2r1w_3532 vdd_uq24 gnd read_bl_0_8 read_bl_1_8 write_bl_0_8 wwl_0_51 rwl_1_51
+ rwl_0_51 cell_2r1w
Xcell_2r1w_2831 vdd_uq23 gnd read_bl_0_19 read_bl_1_19 write_bl_0_19 wwl_0_48 rwl_1_48
+ rwl_0_48 cell_2r1w
Xcell_2r1w_3543 vdd_uq19 gnd read_bl_0_8 read_bl_1_8 write_bl_0_8 wwl_0_40 rwl_1_40
+ rwl_0_40 cell_2r1w
Xcell_2r1w_2842 vdd_uq17 gnd read_bl_0_19 read_bl_1_19 write_bl_0_19 wwl_0_37 rwl_1_37
+ rwl_0_37 cell_2r1w
Xcell_2r1w_3554 vdd_uq13 gnd read_bl_0_8 read_bl_1_8 write_bl_0_8 wwl_0_29 rwl_1_29
+ rwl_0_29 cell_2r1w
Xcell_2r1w_3576 vdd_uq2 gnd read_bl_0_8 read_bl_1_8 write_bl_0_8 wwl_0_7 rwl_1_7 rwl_0_7
+ cell_2r1w
Xcell_2r1w_3510 vdd_uq3 gnd read_bl_0_9 read_bl_1_9 write_bl_0_9 wwl_0_9 rwl_1_9 rwl_0_9
+ cell_2r1w
Xcell_2r1w_3565 vdd_uq8 gnd read_bl_0_8 read_bl_1_8 write_bl_0_8 wwl_0_18 rwl_1_18
+ rwl_0_18 cell_2r1w
Xcell_2r1w_2886 vdd_uq27 gnd read_bl_0_18 read_bl_1_18 write_bl_0_18 wwl_0_57 rwl_1_57
+ rwl_0_57 cell_2r1w
Xcell_2r1w_3598 vdd_uq23 gnd read_bl_0_7 read_bl_1_7 write_bl_0_7 wwl_0_49 rwl_1_49
+ rwl_0_49 cell_2r1w
Xcell_2r1w_2897 vdd_uq22 gnd read_bl_0_18 read_bl_1_18 write_bl_0_18 wwl_0_46 rwl_1_46
+ rwl_0_46 cell_2r1w
Xcell_2r1w_2853 vdd_uq12 gnd read_bl_0_19 read_bl_1_19 write_bl_0_19 wwl_0_26 rwl_1_26
+ rwl_0_26 cell_2r1w
Xcell_2r1w_2875 vdd_uq1 gnd read_bl_0_19 read_bl_1_19 write_bl_0_19 wwl_0_4 rwl_1_4
+ rwl_0_4 cell_2r1w
Xcell_2r1w_2864 vdd_uq6 gnd read_bl_0_19 read_bl_1_19 write_bl_0_19 wwl_0_15 rwl_1_15
+ rwl_0_15 cell_2r1w
Xcell_2r1w_119 vdd_uq3 gnd read_bl_0_62 read_bl_1_62 write_bl_0_62 wwl_0_8 rwl_1_8
+ rwl_0_8 cell_2r1w
Xcell_2r1w_108 vdd_uq8 gnd read_bl_0_62 read_bl_1_62 write_bl_0_62 wwl_0_19 rwl_1_19
+ rwl_0_19 cell_2r1w
Xcell_2r1w_2116 vdd_uq28 gnd read_bl_0_30 read_bl_1_30 write_bl_0_30 wwl_0_59 rwl_1_59
+ rwl_0_59 cell_2r1w
Xcell_2r1w_2127 vdd_uq23 gnd read_bl_0_30 read_bl_1_30 write_bl_0_30 wwl_0_48 rwl_1_48
+ rwl_0_48 cell_2r1w
Xcell_2r1w_2138 vdd_uq17 gnd read_bl_0_30 read_bl_1_30 write_bl_0_30 wwl_0_37 rwl_1_37
+ rwl_0_37 cell_2r1w
Xcell_2r1w_2105 vdd_uq2 gnd read_bl_0_31 read_bl_1_31 write_bl_0_31 wwl_0_6 rwl_1_6
+ rwl_0_6 cell_2r1w
Xcell_2r1w_642 vdd_uq29 gnd read_bl_0_53 read_bl_1_53 write_bl_0_53 wwl_0_61 rwl_1_61
+ rwl_0_61 cell_2r1w
Xcell_2r1w_1415 vdd_uq27 gnd read_bl_0_41 read_bl_1_41 write_bl_0_41 wwl_0_56 rwl_1_56
+ rwl_0_56 cell_2r1w
Xcell_2r1w_653 vdd_uq24 gnd read_bl_0_53 read_bl_1_53 write_bl_0_53 wwl_0_50 rwl_1_50
+ rwl_0_50 cell_2r1w
Xcell_2r1w_1426 vdd_uq21 gnd read_bl_0_41 read_bl_1_41 write_bl_0_41 wwl_0_45 rwl_1_45
+ rwl_0_45 cell_2r1w
Xcell_2r1w_664 vdd_uq18 gnd read_bl_0_53 read_bl_1_53 write_bl_0_53 wwl_0_39 rwl_1_39
+ rwl_0_39 cell_2r1w
Xcell_2r1w_1437 vdd_uq16 gnd read_bl_0_41 read_bl_1_41 write_bl_0_41 wwl_0_34 rwl_1_34
+ rwl_0_34 cell_2r1w
Xcell_2r1w_675 vdd_uq13 gnd read_bl_0_53 read_bl_1_53 write_bl_0_53 wwl_0_28 rwl_1_28
+ rwl_0_28 cell_2r1w
Xcell_2r1w_2149 vdd_uq12 gnd read_bl_0_30 read_bl_1_30 write_bl_0_30 wwl_0_26 rwl_1_26
+ rwl_0_26 cell_2r1w
Xcell_2r1w_1404 vdd gnd read_bl_0_42 read_bl_1_42 write_bl_0_42 wwl_0_3 rwl_1_3 rwl_0_3
+ cell_2r1w
Xcell_2r1w_697 vdd_uq2 gnd read_bl_0_53 read_bl_1_53 write_bl_0_53 wwl_0_6 rwl_1_6
+ rwl_0_6 cell_2r1w
Xcell_2r1w_631 vdd_uq3 gnd read_bl_0_54 read_bl_1_54 write_bl_0_54 wwl_0_8 rwl_1_8
+ rwl_0_8 cell_2r1w
Xcell_2r1w_1459 vdd_uq5 gnd read_bl_0_41 read_bl_1_41 write_bl_0_41 wwl_0_12 rwl_1_12
+ rwl_0_12 cell_2r1w
Xcell_2r1w_686 vdd_uq7 gnd read_bl_0_53 read_bl_1_53 write_bl_0_53 wwl_0_17 rwl_1_17
+ rwl_0_17 cell_2r1w
Xcell_2r1w_620 vdd_uq8 gnd read_bl_0_54 read_bl_1_54 write_bl_0_54 wwl_0_19 rwl_1_19
+ rwl_0_19 cell_2r1w
Xcell_2r1w_1448 vdd_uq10 gnd read_bl_0_41 read_bl_1_41 write_bl_0_41 wwl_0_23 rwl_1_23
+ rwl_0_23 cell_2r1w
Xcell_2r1w_4030 vdd_uq0 gnd read_bl_0_1 read_bl_1_1 write_bl_0_1 wwl_0_1 rwl_1_1 rwl_0_1
+ cell_2r1w
Xcell_2r1w_3395 vdd_uq29 gnd read_bl_0_10 read_bl_1_10 write_bl_0_10 wwl_0_60 rwl_1_60
+ rwl_0_60 cell_2r1w
Xcell_2r1w_2694 vdd_uq27 gnd read_bl_0_21 read_bl_1_21 write_bl_0_21 wwl_0_57 rwl_1_57
+ rwl_0_57 cell_2r1w
Xcell_2r1w_4041 vdd_uq26 gnd read_bl_0_0 read_bl_1_0 write_bl_0_0 wwl_0_54 rwl_1_54
+ rwl_0_54 cell_2r1w
Xcell_2r1w_3340 vdd_uq24 gnd read_bl_0_11 read_bl_1_11 write_bl_0_11 wwl_0_51 rwl_1_51
+ rwl_0_51 cell_2r1w
Xcell_2r1w_4052 vdd_uq20 gnd read_bl_0_0 read_bl_1_0 write_bl_0_0 wwl_0_43 rwl_1_43
+ rwl_0_43 cell_2r1w
Xcell_2r1w_3351 vdd_uq19 gnd read_bl_0_11 read_bl_1_11 write_bl_0_11 wwl_0_40 rwl_1_40
+ rwl_0_40 cell_2r1w
Xcell_2r1w_2650 vdd_uq17 gnd read_bl_0_22 read_bl_1_22 write_bl_0_22 wwl_0_37 rwl_1_37
+ rwl_0_37 cell_2r1w
Xcell_2r1w_4063 vdd_uq15 gnd read_bl_0_0 read_bl_1_0 write_bl_0_0 wwl_0_32 rwl_1_32
+ rwl_0_32 cell_2r1w
Xcell_2r1w_3362 vdd_uq13 gnd read_bl_0_11 read_bl_1_11 write_bl_0_11 wwl_0_29 rwl_1_29
+ rwl_0_29 cell_2r1w
Xcell_2r1w_2661 vdd_uq12 gnd read_bl_0_22 read_bl_1_22 write_bl_0_22 wwl_0_26 rwl_1_26
+ rwl_0_26 cell_2r1w
Xcell_2r1w_2683 vdd_uq1 gnd read_bl_0_22 read_bl_1_22 write_bl_0_22 wwl_0_4 rwl_1_4
+ rwl_0_4 cell_2r1w
Xcell_2r1w_3384 vdd_uq2 gnd read_bl_0_11 read_bl_1_11 write_bl_0_11 wwl_0_7 rwl_1_7
+ rwl_0_7 cell_2r1w
Xcell_2r1w_4085 vdd_uq4 gnd read_bl_0_0 read_bl_1_0 write_bl_0_0 wwl_0_10 rwl_1_10
+ rwl_0_10 cell_2r1w
Xcell_2r1w_2672 vdd_uq6 gnd read_bl_0_22 read_bl_1_22 write_bl_0_22 wwl_0_15 rwl_1_15
+ rwl_0_15 cell_2r1w
Xcell_2r1w_3373 vdd_uq8 gnd read_bl_0_11 read_bl_1_11 write_bl_0_11 wwl_0_18 rwl_1_18
+ rwl_0_18 cell_2r1w
Xcell_2r1w_4074 vdd_uq9 gnd read_bl_0_0 read_bl_1_0 write_bl_0_0 wwl_0_21 rwl_1_21
+ rwl_0_21 cell_2r1w
Xcell_2r1w_1993 vdd_uq26 gnd read_bl_0_32 read_bl_1_32 write_bl_0_32 wwl_0_54 rwl_1_54
+ rwl_0_54 cell_2r1w
Xcell_2r1w_1982 vdd_uq0 gnd read_bl_0_33 read_bl_1_33 write_bl_0_33 wwl_0_1 rwl_1_1
+ rwl_0_1 cell_2r1w
Xcell_2r1w_1971 vdd_uq5 gnd read_bl_0_33 read_bl_1_33 write_bl_0_33 wwl_0_12 rwl_1_12
+ rwl_0_12 cell_2r1w
Xcell_2r1w_1960 vdd_uq10 gnd read_bl_0_33 read_bl_1_33 write_bl_0_33 wwl_0_23 rwl_1_23
+ rwl_0_23 cell_2r1w
Xcell_2r1w_1223 vdd_uq27 gnd read_bl_0_44 read_bl_1_44 write_bl_0_44 wwl_0_56 rwl_1_56
+ rwl_0_56 cell_2r1w
Xcell_2r1w_1234 vdd_uq21 gnd read_bl_0_44 read_bl_1_44 write_bl_0_44 wwl_0_45 rwl_1_45
+ rwl_0_45 cell_2r1w
Xcell_2r1w_1212 vdd gnd read_bl_0_45 read_bl_1_45 write_bl_0_45 wwl_0_3 rwl_1_3 rwl_0_3
+ cell_2r1w
Xcell_2r1w_1201 vdd_uq6 gnd read_bl_0_45 read_bl_1_45 write_bl_0_45 wwl_0_14 rwl_1_14
+ rwl_0_14 cell_2r1w
Xcell_2r1w_450 vdd_uq29 gnd read_bl_0_56 read_bl_1_56 write_bl_0_56 wwl_0_61 rwl_1_61
+ rwl_0_61 cell_2r1w
Xcell_2r1w_1289 vdd_uq26 gnd read_bl_0_43 read_bl_1_43 write_bl_0_43 wwl_0_54 rwl_1_54
+ rwl_0_54 cell_2r1w
Xcell_2r1w_461 vdd_uq24 gnd read_bl_0_56 read_bl_1_56 write_bl_0_56 wwl_0_50 rwl_1_50
+ rwl_0_50 cell_2r1w
Xcell_2r1w_472 vdd_uq18 gnd read_bl_0_56 read_bl_1_56 write_bl_0_56 wwl_0_39 rwl_1_39
+ rwl_0_39 cell_2r1w
Xcell_2r1w_1245 vdd_uq16 gnd read_bl_0_44 read_bl_1_44 write_bl_0_44 wwl_0_34 rwl_1_34
+ rwl_0_34 cell_2r1w
Xcell_2r1w_483 vdd_uq13 gnd read_bl_0_56 read_bl_1_56 write_bl_0_56 wwl_0_28 rwl_1_28
+ rwl_0_28 cell_2r1w
Xcell_2r1w_1278 vdd_uq0 gnd read_bl_0_44 read_bl_1_44 write_bl_0_44 wwl_0_1 rwl_1_1
+ rwl_0_1 cell_2r1w
Xcell_2r1w_1267 vdd_uq5 gnd read_bl_0_44 read_bl_1_44 write_bl_0_44 wwl_0_12 rwl_1_12
+ rwl_0_12 cell_2r1w
Xcell_2r1w_494 vdd_uq7 gnd read_bl_0_56 read_bl_1_56 write_bl_0_56 wwl_0_17 rwl_1_17
+ rwl_0_17 cell_2r1w
Xcell_2r1w_1256 vdd_uq10 gnd read_bl_0_44 read_bl_1_44 write_bl_0_44 wwl_0_23 rwl_1_23
+ rwl_0_23 cell_2r1w
Xcell_2r1w_3170 vdd_uq13 gnd read_bl_0_14 read_bl_1_14 write_bl_0_14 wwl_0_29 rwl_1_29
+ rwl_0_29 cell_2r1w
Xcell_2r1w_2491 vdd_uq1 gnd read_bl_0_25 read_bl_1_25 write_bl_0_25 wwl_0_4 rwl_1_4
+ rwl_0_4 cell_2r1w
Xcell_2r1w_1790 vdd_uq0 gnd read_bl_0_36 read_bl_1_36 write_bl_0_36 wwl_0_1 rwl_1_1
+ rwl_0_1 cell_2r1w
Xcell_2r1w_3192 vdd_uq2 gnd read_bl_0_14 read_bl_1_14 write_bl_0_14 wwl_0_7 rwl_1_7
+ rwl_0_7 cell_2r1w
Xcell_2r1w_2480 vdd_uq6 gnd read_bl_0_25 read_bl_1_25 write_bl_0_25 wwl_0_15 rwl_1_15
+ rwl_0_15 cell_2r1w
Xcell_2r1w_3181 vdd_uq8 gnd read_bl_0_14 read_bl_1_14 write_bl_0_14 wwl_0_18 rwl_1_18
+ rwl_0_18 cell_2r1w
Xcell_2r1w_1031 vdd_uq27 gnd read_bl_0_47 read_bl_1_47 write_bl_0_47 wwl_0_56 rwl_1_56
+ rwl_0_56 cell_2r1w
Xcell_2r1w_1042 vdd_uq21 gnd read_bl_0_47 read_bl_1_47 write_bl_0_47 wwl_0_45 rwl_1_45
+ rwl_0_45 cell_2r1w
Xcell_2r1w_1053 vdd_uq16 gnd read_bl_0_47 read_bl_1_47 write_bl_0_47 wwl_0_34 rwl_1_34
+ rwl_0_34 cell_2r1w
Xcell_2r1w_1020 vdd gnd read_bl_0_48 read_bl_1_48 write_bl_0_48 wwl_0_3 rwl_1_3 rwl_0_3
+ cell_2r1w
Xcell_2r1w_1086 vdd_uq0 gnd read_bl_0_47 read_bl_1_47 write_bl_0_47 wwl_0_1 rwl_1_1
+ rwl_0_1 cell_2r1w
Xcell_2r1w_1075 vdd_uq5 gnd read_bl_0_47 read_bl_1_47 write_bl_0_47 wwl_0_12 rwl_1_12
+ rwl_0_12 cell_2r1w
Xcell_2r1w_1064 vdd_uq10 gnd read_bl_0_47 read_bl_1_47 write_bl_0_47 wwl_0_23 rwl_1_23
+ rwl_0_23 cell_2r1w
Xcell_2r1w_1097 vdd_uq26 gnd read_bl_0_46 read_bl_1_46 write_bl_0_46 wwl_0_54 rwl_1_54
+ rwl_0_54 cell_2r1w
Xcell_2r1w_280 vdd_uq18 gnd read_bl_0_59 read_bl_1_59 write_bl_0_59 wwl_0_39 rwl_1_39
+ rwl_0_39 cell_2r1w
Xcell_2r1w_291 vdd_uq13 gnd read_bl_0_59 read_bl_1_59 write_bl_0_59 wwl_0_28 rwl_1_28
+ rwl_0_28 cell_2r1w
Xcell_2r1w_3906 vdd_uq29 gnd read_bl_0_2 read_bl_1_2 write_bl_0_2 wwl_0_61 rwl_1_61
+ rwl_0_61 cell_2r1w
Xcell_2r1w_3917 vdd_uq24 gnd read_bl_0_2 read_bl_1_2 write_bl_0_2 wwl_0_50 rwl_1_50
+ rwl_0_50 cell_2r1w
Xcell_2r1w_3928 vdd_uq18 gnd read_bl_0_2 read_bl_1_2 write_bl_0_2 wwl_0_39 rwl_1_39
+ rwl_0_39 cell_2r1w
Xcell_2r1w_3939 vdd_uq13 gnd read_bl_0_2 read_bl_1_2 write_bl_0_2 wwl_0_28 rwl_1_28
+ rwl_0_28 cell_2r1w
Xcell_2r1w_3714 vdd_uq29 gnd read_bl_0_5 read_bl_1_5 write_bl_0_5 wwl_0_61 rwl_1_61
+ rwl_0_61 cell_2r1w
Xcell_2r1w_3725 vdd_uq24 gnd read_bl_0_5 read_bl_1_5 write_bl_0_5 wwl_0_50 rwl_1_50
+ rwl_0_50 cell_2r1w
Xcell_2r1w_3736 vdd_uq18 gnd read_bl_0_5 read_bl_1_5 write_bl_0_5 wwl_0_39 rwl_1_39
+ rwl_0_39 cell_2r1w
Xcell_2r1w_3747 vdd_uq13 gnd read_bl_0_5 read_bl_1_5 write_bl_0_5 wwl_0_28 rwl_1_28
+ rwl_0_28 cell_2r1w
Xcell_2r1w_3769 vdd_uq2 gnd read_bl_0_5 read_bl_1_5 write_bl_0_5 wwl_0_6 rwl_1_6 rwl_0_6
+ cell_2r1w
Xcell_2r1w_3703 vdd_uq3 gnd read_bl_0_6 read_bl_1_6 write_bl_0_6 wwl_0_8 rwl_1_8 rwl_0_8
+ cell_2r1w
Xcell_2r1w_3758 vdd_uq7 gnd read_bl_0_5 read_bl_1_5 write_bl_0_5 wwl_0_17 rwl_1_17
+ rwl_0_17 cell_2r1w
Xcell_2r1w_2309 vdd_uq28 gnd read_bl_0_27 read_bl_1_27 write_bl_0_27 wwl_0_58 rwl_1_58
+ rwl_0_58 cell_2r1w
Xcell_2r1w_835 vdd_uq29 gnd read_bl_0_50 read_bl_1_50 write_bl_0_50 wwl_0_60 rwl_1_60
+ rwl_0_60 cell_2r1w
Xcell_2r1w_1608 vdd_uq26 gnd read_bl_0_38 read_bl_1_38 write_bl_0_38 wwl_0_55 rwl_1_55
+ rwl_0_55 cell_2r1w
Xcell_2r1w_846 vdd_uq23 gnd read_bl_0_50 read_bl_1_50 write_bl_0_50 wwl_0_49 rwl_1_49
+ rwl_0_49 cell_2r1w
Xcell_2r1w_1619 vdd_uq21 gnd read_bl_0_38 read_bl_1_38 write_bl_0_38 wwl_0_44 rwl_1_44
+ rwl_0_44 cell_2r1w
Xcell_2r1w_857 vdd_uq18 gnd read_bl_0_50 read_bl_1_50 write_bl_0_50 wwl_0_38 rwl_1_38
+ rwl_0_38 cell_2r1w
Xcell_2r1w_802 vdd_uq13 gnd read_bl_0_51 read_bl_1_51 write_bl_0_51 wwl_0_29 rwl_1_29
+ rwl_0_29 cell_2r1w
Xcell_2r1w_868 vdd_uq12 gnd read_bl_0_50 read_bl_1_50 write_bl_0_50 wwl_0_27 rwl_1_27
+ rwl_0_27 cell_2r1w
Xcell_2r1w_824 vdd_uq2 gnd read_bl_0_51 read_bl_1_51 write_bl_0_51 wwl_0_7 rwl_1_7
+ rwl_0_7 cell_2r1w
Xcell_2r1w_879 vdd_uq7 gnd read_bl_0_50 read_bl_1_50 write_bl_0_50 wwl_0_16 rwl_1_16
+ rwl_0_16 cell_2r1w
Xcell_2r1w_813 vdd_uq8 gnd read_bl_0_51 read_bl_1_51 write_bl_0_51 wwl_0_18 rwl_1_18
+ rwl_0_18 cell_2r1w
Xcell_2r1w_3522 vdd_uq29 gnd read_bl_0_8 read_bl_1_8 write_bl_0_8 wwl_0_61 rwl_1_61
+ rwl_0_61 cell_2r1w
Xcell_2r1w_3588 vdd_uq28 gnd read_bl_0_7 read_bl_1_7 write_bl_0_7 wwl_0_59 rwl_1_59
+ rwl_0_59 cell_2r1w
Xcell_2r1w_2821 vdd_uq28 gnd read_bl_0_19 read_bl_1_19 write_bl_0_19 wwl_0_58 rwl_1_58
+ rwl_0_58 cell_2r1w
Xcell_2r1w_3533 vdd_uq24 gnd read_bl_0_8 read_bl_1_8 write_bl_0_8 wwl_0_50 rwl_1_50
+ rwl_0_50 cell_2r1w
Xcell_2r1w_3599 vdd_uq23 gnd read_bl_0_7 read_bl_1_7 write_bl_0_7 wwl_0_48 rwl_1_48
+ rwl_0_48 cell_2r1w
Xcell_2r1w_2832 vdd_uq22 gnd read_bl_0_19 read_bl_1_19 write_bl_0_19 wwl_0_47 rwl_1_47
+ rwl_0_47 cell_2r1w
Xcell_2r1w_3544 vdd_uq18 gnd read_bl_0_8 read_bl_1_8 write_bl_0_8 wwl_0_39 rwl_1_39
+ rwl_0_39 cell_2r1w
Xcell_2r1w_2843 vdd_uq17 gnd read_bl_0_19 read_bl_1_19 write_bl_0_19 wwl_0_36 rwl_1_36
+ rwl_0_36 cell_2r1w
Xcell_2r1w_3555 vdd_uq13 gnd read_bl_0_8 read_bl_1_8 write_bl_0_8 wwl_0_28 rwl_1_28
+ rwl_0_28 cell_2r1w
Xcell_2r1w_2854 vdd_uq11 gnd read_bl_0_19 read_bl_1_19 write_bl_0_19 wwl_0_25 rwl_1_25
+ rwl_0_25 cell_2r1w
Xcell_2r1w_2810 vdd_uq1 gnd read_bl_0_20 read_bl_1_20 write_bl_0_20 wwl_0_5 rwl_1_5
+ rwl_0_5 cell_2r1w
Xcell_2r1w_2876 vdd gnd read_bl_0_19 read_bl_1_19 write_bl_0_19 wwl_0_3 rwl_1_3 rwl_0_3
+ cell_2r1w
Xcell_2r1w_3577 vdd_uq2 gnd read_bl_0_8 read_bl_1_8 write_bl_0_8 wwl_0_6 rwl_1_6 rwl_0_6
+ cell_2r1w
Xcell_2r1w_3511 vdd_uq3 gnd read_bl_0_9 read_bl_1_9 write_bl_0_9 wwl_0_8 rwl_1_8 rwl_0_8
+ cell_2r1w
Xcell_2r1w_2865 vdd_uq6 gnd read_bl_0_19 read_bl_1_19 write_bl_0_19 wwl_0_14 rwl_1_14
+ rwl_0_14 cell_2r1w
Xcell_2r1w_3566 vdd_uq7 gnd read_bl_0_8 read_bl_1_8 write_bl_0_8 wwl_0_17 rwl_1_17
+ rwl_0_17 cell_2r1w
Xcell_2r1w_3500 vdd_uq8 gnd read_bl_0_9 read_bl_1_9 write_bl_0_9 wwl_0_19 rwl_1_19
+ rwl_0_19 cell_2r1w
Xcell_2r1w_2887 vdd_uq27 gnd read_bl_0_18 read_bl_1_18 write_bl_0_18 wwl_0_56 rwl_1_56
+ rwl_0_56 cell_2r1w
Xcell_2r1w_2898 vdd_uq21 gnd read_bl_0_18 read_bl_1_18 write_bl_0_18 wwl_0_45 rwl_1_45
+ rwl_0_45 cell_2r1w
Xcell_2r1w_109 vdd_uq8 gnd read_bl_0_62 read_bl_1_62 write_bl_0_62 wwl_0_18 rwl_1_18
+ rwl_0_18 cell_2r1w
Xcell_2r1w_2117 vdd_uq28 gnd read_bl_0_30 read_bl_1_30 write_bl_0_30 wwl_0_58 rwl_1_58
+ rwl_0_58 cell_2r1w
Xcell_2r1w_1416 vdd_uq26 gnd read_bl_0_41 read_bl_1_41 write_bl_0_41 wwl_0_55 rwl_1_55
+ rwl_0_55 cell_2r1w
Xcell_2r1w_2128 vdd_uq22 gnd read_bl_0_30 read_bl_1_30 write_bl_0_30 wwl_0_47 rwl_1_47
+ rwl_0_47 cell_2r1w
Xcell_2r1w_1427 vdd_uq21 gnd read_bl_0_41 read_bl_1_41 write_bl_0_41 wwl_0_44 rwl_1_44
+ rwl_0_44 cell_2r1w
Xcell_2r1w_2139 vdd_uq17 gnd read_bl_0_30 read_bl_1_30 write_bl_0_30 wwl_0_36 rwl_1_36
+ rwl_0_36 cell_2r1w
Xcell_2r1w_2106 vdd_uq1 gnd read_bl_0_31 read_bl_1_31 write_bl_0_31 wwl_0_5 rwl_1_5
+ rwl_0_5 cell_2r1w
Xcell_2r1w_1405 vdd gnd read_bl_0_42 read_bl_1_42 write_bl_0_42 wwl_0_2 rwl_1_2 rwl_0_2
+ cell_2r1w
Xcell_2r1w_643 vdd_uq29 gnd read_bl_0_53 read_bl_1_53 write_bl_0_53 wwl_0_60 rwl_1_60
+ rwl_0_60 cell_2r1w
Xcell_2r1w_654 vdd_uq23 gnd read_bl_0_53 read_bl_1_53 write_bl_0_53 wwl_0_49 rwl_1_49
+ rwl_0_49 cell_2r1w
Xcell_2r1w_665 vdd_uq18 gnd read_bl_0_53 read_bl_1_53 write_bl_0_53 wwl_0_38 rwl_1_38
+ rwl_0_38 cell_2r1w
Xcell_2r1w_1438 vdd_uq15 gnd read_bl_0_41 read_bl_1_41 write_bl_0_41 wwl_0_33 rwl_1_33
+ rwl_0_33 cell_2r1w
Xcell_2r1w_610 vdd_uq13 gnd read_bl_0_54 read_bl_1_54 write_bl_0_54 wwl_0_29 rwl_1_29
+ rwl_0_29 cell_2r1w
Xcell_2r1w_676 vdd_uq12 gnd read_bl_0_53 read_bl_1_53 write_bl_0_53 wwl_0_27 rwl_1_27
+ rwl_0_27 cell_2r1w
Xcell_2r1w_698 vdd_uq1 gnd read_bl_0_53 read_bl_1_53 write_bl_0_53 wwl_0_5 rwl_1_5
+ rwl_0_5 cell_2r1w
Xcell_2r1w_632 vdd_uq2 gnd read_bl_0_54 read_bl_1_54 write_bl_0_54 wwl_0_7 rwl_1_7
+ rwl_0_7 cell_2r1w
Xcell_2r1w_687 vdd_uq7 gnd read_bl_0_53 read_bl_1_53 write_bl_0_53 wwl_0_16 rwl_1_16
+ rwl_0_16 cell_2r1w
Xcell_2r1w_621 vdd_uq8 gnd read_bl_0_54 read_bl_1_54 write_bl_0_54 wwl_0_18 rwl_1_18
+ rwl_0_18 cell_2r1w
Xcell_2r1w_1449 vdd_uq10 gnd read_bl_0_41 read_bl_1_41 write_bl_0_41 wwl_0_22 rwl_1_22
+ rwl_0_22 cell_2r1w
Xcell_2r1w_4042 vdd_uq25 gnd read_bl_0_0 read_bl_1_0 write_bl_0_0 wwl_0_53 rwl_1_53
+ rwl_0_53 cell_2r1w
Xcell_2r1w_4053 vdd_uq20 gnd read_bl_0_0 read_bl_1_0 write_bl_0_0 wwl_0_42 rwl_1_42
+ rwl_0_42 cell_2r1w
Xcell_2r1w_4064 vdd_uq14 gnd read_bl_0_0 read_bl_1_0 write_bl_0_0 wwl_0_31 rwl_1_31
+ rwl_0_31 cell_2r1w
Xcell_2r1w_4031 vdd_uq0 gnd read_bl_0_1 read_bl_1_1 write_bl_0_1 wwl_0_0 rwl_1_0 rwl_0_0
+ cell_2r1w
Xcell_2r1w_4020 vdd_uq4 gnd read_bl_0_1 read_bl_1_1 write_bl_0_1 wwl_0_11 rwl_1_11
+ rwl_0_11 cell_2r1w
Xcell_2r1w_3330 vdd_uq29 gnd read_bl_0_11 read_bl_1_11 write_bl_0_11 wwl_0_61 rwl_1_61
+ rwl_0_61 cell_2r1w
Xcell_2r1w_3396 vdd_uq28 gnd read_bl_0_10 read_bl_1_10 write_bl_0_10 wwl_0_59 rwl_1_59
+ rwl_0_59 cell_2r1w
Xcell_2r1w_2695 vdd_uq27 gnd read_bl_0_21 read_bl_1_21 write_bl_0_21 wwl_0_56 rwl_1_56
+ rwl_0_56 cell_2r1w
Xcell_2r1w_3341 vdd_uq24 gnd read_bl_0_11 read_bl_1_11 write_bl_0_11 wwl_0_50 rwl_1_50
+ rwl_0_50 cell_2r1w
Xcell_2r1w_2640 vdd_uq22 gnd read_bl_0_22 read_bl_1_22 write_bl_0_22 wwl_0_47 rwl_1_47
+ rwl_0_47 cell_2r1w
Xcell_2r1w_3352 vdd_uq18 gnd read_bl_0_11 read_bl_1_11 write_bl_0_11 wwl_0_39 rwl_1_39
+ rwl_0_39 cell_2r1w
Xcell_2r1w_2651 vdd_uq17 gnd read_bl_0_22 read_bl_1_22 write_bl_0_22 wwl_0_36 rwl_1_36
+ rwl_0_36 cell_2r1w
Xcell_2r1w_1950 vdd_uq15 gnd read_bl_0_33 read_bl_1_33 write_bl_0_33 wwl_0_33 rwl_1_33
+ rwl_0_33 cell_2r1w
Xcell_2r1w_3363 vdd_uq13 gnd read_bl_0_11 read_bl_1_11 write_bl_0_11 wwl_0_28 rwl_1_28
+ rwl_0_28 cell_2r1w
Xcell_2r1w_2662 vdd_uq11 gnd read_bl_0_22 read_bl_1_22 write_bl_0_22 wwl_0_25 rwl_1_25
+ rwl_0_25 cell_2r1w
Xcell_2r1w_2684 vdd gnd read_bl_0_22 read_bl_1_22 write_bl_0_22 wwl_0_3 rwl_1_3 rwl_0_3
+ cell_2r1w
Xcell_2r1w_3385 vdd_uq2 gnd read_bl_0_11 read_bl_1_11 write_bl_0_11 wwl_0_6 rwl_1_6
+ rwl_0_6 cell_2r1w
Xcell_2r1w_4086 vdd_uq3 gnd read_bl_0_0 read_bl_1_0 write_bl_0_0 wwl_0_9 rwl_1_9 rwl_0_9
+ cell_2r1w
Xcell_2r1w_1972 vdd_uq4 gnd read_bl_0_33 read_bl_1_33 write_bl_0_33 wwl_0_11 rwl_1_11
+ rwl_0_11 cell_2r1w
Xcell_2r1w_2673 vdd_uq6 gnd read_bl_0_22 read_bl_1_22 write_bl_0_22 wwl_0_14 rwl_1_14
+ rwl_0_14 cell_2r1w
Xcell_2r1w_3374 vdd_uq7 gnd read_bl_0_11 read_bl_1_11 write_bl_0_11 wwl_0_17 rwl_1_17
+ rwl_0_17 cell_2r1w
Xcell_2r1w_4075 vdd_uq9 gnd read_bl_0_0 read_bl_1_0 write_bl_0_0 wwl_0_20 rwl_1_20
+ rwl_0_20 cell_2r1w
Xcell_2r1w_1961 vdd_uq10 gnd read_bl_0_33 read_bl_1_33 write_bl_0_33 wwl_0_22 rwl_1_22
+ rwl_0_22 cell_2r1w
Xcell_2r1w_1994 vdd_uq25 gnd read_bl_0_32 read_bl_1_32 write_bl_0_32 wwl_0_53 rwl_1_53
+ rwl_0_53 cell_2r1w
Xcell_2r1w_1983 vdd_uq0 gnd read_bl_0_33 read_bl_1_33 write_bl_0_33 wwl_0_0 rwl_1_0
+ rwl_0_0 cell_2r1w
Xcell_2r1w_1224 vdd_uq26 gnd read_bl_0_44 read_bl_1_44 write_bl_0_44 wwl_0_55 rwl_1_55
+ rwl_0_55 cell_2r1w
Xcell_2r1w_1235 vdd_uq21 gnd read_bl_0_44 read_bl_1_44 write_bl_0_44 wwl_0_44 rwl_1_44
+ rwl_0_44 cell_2r1w
Xcell_2r1w_1246 vdd_uq15 gnd read_bl_0_44 read_bl_1_44 write_bl_0_44 wwl_0_33 rwl_1_33
+ rwl_0_33 cell_2r1w
Xcell_2r1w_1213 vdd gnd read_bl_0_45 read_bl_1_45 write_bl_0_45 wwl_0_2 rwl_1_2 rwl_0_2
+ cell_2r1w
Xcell_2r1w_1268 vdd_uq4 gnd read_bl_0_44 read_bl_1_44 write_bl_0_44 wwl_0_11 rwl_1_11
+ rwl_0_11 cell_2r1w
Xcell_2r1w_1202 vdd_uq5 gnd read_bl_0_45 read_bl_1_45 write_bl_0_45 wwl_0_13 rwl_1_13
+ rwl_0_13 cell_2r1w
Xcell_2r1w_1257 vdd_uq10 gnd read_bl_0_44 read_bl_1_44 write_bl_0_44 wwl_0_22 rwl_1_22
+ rwl_0_22 cell_2r1w
Xcell_2r1w_451 vdd_uq29 gnd read_bl_0_56 read_bl_1_56 write_bl_0_56 wwl_0_60 rwl_1_60
+ rwl_0_60 cell_2r1w
Xcell_2r1w_462 vdd_uq23 gnd read_bl_0_56 read_bl_1_56 write_bl_0_56 wwl_0_49 rwl_1_49
+ rwl_0_49 cell_2r1w
Xcell_2r1w_473 vdd_uq18 gnd read_bl_0_56 read_bl_1_56 write_bl_0_56 wwl_0_38 rwl_1_38
+ rwl_0_38 cell_2r1w
Xcell_2r1w_484 vdd_uq12 gnd read_bl_0_56 read_bl_1_56 write_bl_0_56 wwl_0_27 rwl_1_27
+ rwl_0_27 cell_2r1w
Xcell_2r1w_1279 vdd_uq0 gnd read_bl_0_44 read_bl_1_44 write_bl_0_44 wwl_0_0 rwl_1_0
+ rwl_0_0 cell_2r1w
Xcell_2r1w_440 vdd_uq2 gnd read_bl_0_57 read_bl_1_57 write_bl_0_57 wwl_0_7 rwl_1_7
+ rwl_0_7 cell_2r1w
Xcell_2r1w_495 vdd_uq7 gnd read_bl_0_56 read_bl_1_56 write_bl_0_56 wwl_0_16 rwl_1_16
+ rwl_0_16 cell_2r1w
Xcell_2r1w_3160 vdd_uq18 gnd read_bl_0_14 read_bl_1_14 write_bl_0_14 wwl_0_39 rwl_1_39
+ rwl_0_39 cell_2r1w
Xcell_2r1w_3171 vdd_uq13 gnd read_bl_0_14 read_bl_1_14 write_bl_0_14 wwl_0_28 rwl_1_28
+ rwl_0_28 cell_2r1w
Xcell_2r1w_2470 vdd_uq11 gnd read_bl_0_25 read_bl_1_25 write_bl_0_25 wwl_0_25 rwl_1_25
+ rwl_0_25 cell_2r1w
Xcell_2r1w_2492 vdd gnd read_bl_0_25 read_bl_1_25 write_bl_0_25 wwl_0_3 rwl_1_3 rwl_0_3
+ cell_2r1w
Xcell_2r1w_1791 vdd_uq0 gnd read_bl_0_36 read_bl_1_36 write_bl_0_36 wwl_0_0 rwl_1_0
+ rwl_0_0 cell_2r1w
Xcell_2r1w_3193 vdd_uq2 gnd read_bl_0_14 read_bl_1_14 write_bl_0_14 wwl_0_6 rwl_1_6
+ rwl_0_6 cell_2r1w
Xcell_2r1w_1780 vdd_uq4 gnd read_bl_0_36 read_bl_1_36 write_bl_0_36 wwl_0_11 rwl_1_11
+ rwl_0_11 cell_2r1w
Xcell_2r1w_2481 vdd_uq6 gnd read_bl_0_25 read_bl_1_25 write_bl_0_25 wwl_0_14 rwl_1_14
+ rwl_0_14 cell_2r1w
Xcell_2r1w_3182 vdd_uq7 gnd read_bl_0_14 read_bl_1_14 write_bl_0_14 wwl_0_17 rwl_1_17
+ rwl_0_17 cell_2r1w
Xcell_2r1w_1032 vdd_uq26 gnd read_bl_0_47 read_bl_1_47 write_bl_0_47 wwl_0_55 rwl_1_55
+ rwl_0_55 cell_2r1w
Xcell_2r1w_1098 vdd_uq25 gnd read_bl_0_46 read_bl_1_46 write_bl_0_46 wwl_0_53 rwl_1_53
+ rwl_0_53 cell_2r1w
Xcell_2r1w_270 vdd_uq23 gnd read_bl_0_59 read_bl_1_59 write_bl_0_59 wwl_0_49 rwl_1_49
+ rwl_0_49 cell_2r1w
Xcell_2r1w_1043 vdd_uq21 gnd read_bl_0_47 read_bl_1_47 write_bl_0_47 wwl_0_44 rwl_1_44
+ rwl_0_44 cell_2r1w
Xcell_2r1w_281 vdd_uq18 gnd read_bl_0_59 read_bl_1_59 write_bl_0_59 wwl_0_38 rwl_1_38
+ rwl_0_38 cell_2r1w
Xcell_2r1w_1054 vdd_uq15 gnd read_bl_0_47 read_bl_1_47 write_bl_0_47 wwl_0_33 rwl_1_33
+ rwl_0_33 cell_2r1w
Xcell_2r1w_1021 vdd gnd read_bl_0_48 read_bl_1_48 write_bl_0_48 wwl_0_2 rwl_1_2 rwl_0_2
+ cell_2r1w
Xcell_2r1w_1087 vdd_uq0 gnd read_bl_0_47 read_bl_1_47 write_bl_0_47 wwl_0_0 rwl_1_0
+ rwl_0_0 cell_2r1w
Xcell_2r1w_1076 vdd_uq4 gnd read_bl_0_47 read_bl_1_47 write_bl_0_47 wwl_0_11 rwl_1_11
+ rwl_0_11 cell_2r1w
Xcell_2r1w_1010 vdd_uq5 gnd read_bl_0_48 read_bl_1_48 write_bl_0_48 wwl_0_13 rwl_1_13
+ rwl_0_13 cell_2r1w
Xcell_2r1w_1065 vdd_uq10 gnd read_bl_0_47 read_bl_1_47 write_bl_0_47 wwl_0_22 rwl_1_22
+ rwl_0_22 cell_2r1w
Xcell_2r1w_292 vdd_uq12 gnd read_bl_0_59 read_bl_1_59 write_bl_0_59 wwl_0_27 rwl_1_27
+ rwl_0_27 cell_2r1w
Xcell_2r1w_3907 vdd_uq29 gnd read_bl_0_2 read_bl_1_2 write_bl_0_2 wwl_0_60 rwl_1_60
+ rwl_0_60 cell_2r1w
Xcell_2r1w_3918 vdd_uq23 gnd read_bl_0_2 read_bl_1_2 write_bl_0_2 wwl_0_49 rwl_1_49
+ rwl_0_49 cell_2r1w
Xcell_2r1w_3929 vdd_uq18 gnd read_bl_0_2 read_bl_1_2 write_bl_0_2 wwl_0_38 rwl_1_38
+ rwl_0_38 cell_2r1w
Xcell_2r1w_3715 vdd_uq29 gnd read_bl_0_5 read_bl_1_5 write_bl_0_5 wwl_0_60 rwl_1_60
+ rwl_0_60 cell_2r1w
Xcell_2r1w_3726 vdd_uq23 gnd read_bl_0_5 read_bl_1_5 write_bl_0_5 wwl_0_49 rwl_1_49
+ rwl_0_49 cell_2r1w
Xcell_2r1w_3737 vdd_uq18 gnd read_bl_0_5 read_bl_1_5 write_bl_0_5 wwl_0_38 rwl_1_38
+ rwl_0_38 cell_2r1w
Xcell_2r1w_3748 vdd_uq12 gnd read_bl_0_5 read_bl_1_5 write_bl_0_5 wwl_0_27 rwl_1_27
+ rwl_0_27 cell_2r1w
Xcell_2r1w_3704 vdd_uq2 gnd read_bl_0_6 read_bl_1_6 write_bl_0_6 wwl_0_7 rwl_1_7 rwl_0_7
+ cell_2r1w
Xcell_2r1w_3759 vdd_uq7 gnd read_bl_0_5 read_bl_1_5 write_bl_0_5 wwl_0_16 rwl_1_16
+ rwl_0_16 cell_2r1w
Xcell_2r1w_1609 vdd_uq26 gnd read_bl_0_38 read_bl_1_38 write_bl_0_38 wwl_0_54 rwl_1_54
+ rwl_0_54 cell_2r1w
Xcell_2r1w_836 vdd_uq28 gnd read_bl_0_50 read_bl_1_50 write_bl_0_50 wwl_0_59 rwl_1_59
+ rwl_0_59 cell_2r1w
Xcell_2r1w_847 vdd_uq23 gnd read_bl_0_50 read_bl_1_50 write_bl_0_50 wwl_0_48 rwl_1_48
+ rwl_0_48 cell_2r1w
Xcell_2r1w_858 vdd_uq17 gnd read_bl_0_50 read_bl_1_50 write_bl_0_50 wwl_0_37 rwl_1_37
+ rwl_0_37 cell_2r1w
Xcell_2r1w_803 vdd_uq13 gnd read_bl_0_51 read_bl_1_51 write_bl_0_51 wwl_0_28 rwl_1_28
+ rwl_0_28 cell_2r1w
Xcell_2r1w_869 vdd_uq12 gnd read_bl_0_50 read_bl_1_50 write_bl_0_50 wwl_0_26 rwl_1_26
+ rwl_0_26 cell_2r1w
Xcell_2r1w_825 vdd_uq2 gnd read_bl_0_51 read_bl_1_51 write_bl_0_51 wwl_0_6 rwl_1_6
+ rwl_0_6 cell_2r1w
Xcell_2r1w_814 vdd_uq7 gnd read_bl_0_51 read_bl_1_51 write_bl_0_51 wwl_0_17 rwl_1_17
+ rwl_0_17 cell_2r1w
Xcell_2r1w_3501 vdd_uq8 gnd read_bl_0_9 read_bl_1_9 write_bl_0_9 wwl_0_18 rwl_1_18
+ rwl_0_18 cell_2r1w
Xcell_2r1w_3523 vdd_uq29 gnd read_bl_0_8 read_bl_1_8 write_bl_0_8 wwl_0_60 rwl_1_60
+ rwl_0_60 cell_2r1w
Xcell_2r1w_3589 vdd_uq28 gnd read_bl_0_7 read_bl_1_7 write_bl_0_7 wwl_0_58 rwl_1_58
+ rwl_0_58 cell_2r1w
Xcell_2r1w_2822 vdd_uq27 gnd read_bl_0_19 read_bl_1_19 write_bl_0_19 wwl_0_57 rwl_1_57
+ rwl_0_57 cell_2r1w
Xcell_2r1w_2888 vdd_uq26 gnd read_bl_0_18 read_bl_1_18 write_bl_0_18 wwl_0_55 rwl_1_55
+ rwl_0_55 cell_2r1w
Xcell_2r1w_3534 vdd_uq23 gnd read_bl_0_8 read_bl_1_8 write_bl_0_8 wwl_0_49 rwl_1_49
+ rwl_0_49 cell_2r1w
Xcell_2r1w_2833 vdd_uq22 gnd read_bl_0_19 read_bl_1_19 write_bl_0_19 wwl_0_46 rwl_1_46
+ rwl_0_46 cell_2r1w
Xcell_2r1w_2899 vdd_uq21 gnd read_bl_0_18 read_bl_1_18 write_bl_0_18 wwl_0_44 rwl_1_44
+ rwl_0_44 cell_2r1w
Xcell_2r1w_3545 vdd_uq18 gnd read_bl_0_8 read_bl_1_8 write_bl_0_8 wwl_0_38 rwl_1_38
+ rwl_0_38 cell_2r1w
Xcell_2r1w_2844 vdd_uq16 gnd read_bl_0_19 read_bl_1_19 write_bl_0_19 wwl_0_35 rwl_1_35
+ rwl_0_35 cell_2r1w
Xcell_2r1w_3556 vdd_uq12 gnd read_bl_0_8 read_bl_1_8 write_bl_0_8 wwl_0_27 rwl_1_27
+ rwl_0_27 cell_2r1w
Xcell_2r1w_2855 vdd_uq11 gnd read_bl_0_19 read_bl_1_19 write_bl_0_19 wwl_0_24 rwl_1_24
+ rwl_0_24 cell_2r1w
Xcell_2r1w_3578 vdd_uq1 gnd read_bl_0_8 read_bl_1_8 write_bl_0_8 wwl_0_5 rwl_1_5 rwl_0_5
+ cell_2r1w
Xcell_2r1w_2811 vdd_uq1 gnd read_bl_0_20 read_bl_1_20 write_bl_0_20 wwl_0_4 rwl_1_4
+ rwl_0_4 cell_2r1w
Xcell_2r1w_2877 vdd gnd read_bl_0_19 read_bl_1_19 write_bl_0_19 wwl_0_2 rwl_1_2 rwl_0_2
+ cell_2r1w
Xcell_2r1w_3512 vdd_uq2 gnd read_bl_0_9 read_bl_1_9 write_bl_0_9 wwl_0_7 rwl_1_7 rwl_0_7
+ cell_2r1w
Xcell_2r1w_2866 vdd_uq5 gnd read_bl_0_19 read_bl_1_19 write_bl_0_19 wwl_0_13 rwl_1_13
+ rwl_0_13 cell_2r1w
Xcell_2r1w_2800 vdd_uq6 gnd read_bl_0_20 read_bl_1_20 write_bl_0_20 wwl_0_15 rwl_1_15
+ rwl_0_15 cell_2r1w
Xcell_2r1w_3567 vdd_uq7 gnd read_bl_0_8 read_bl_1_8 write_bl_0_8 wwl_0_16 rwl_1_16
+ rwl_0_16 cell_2r1w
Xcell_2r1w_2118 vdd_uq27 gnd read_bl_0_30 read_bl_1_30 write_bl_0_30 wwl_0_57 rwl_1_57
+ rwl_0_57 cell_2r1w
Xcell_2r1w_1417 vdd_uq26 gnd read_bl_0_41 read_bl_1_41 write_bl_0_41 wwl_0_54 rwl_1_54
+ rwl_0_54 cell_2r1w
Xcell_2r1w_2129 vdd_uq22 gnd read_bl_0_30 read_bl_1_30 write_bl_0_30 wwl_0_46 rwl_1_46
+ rwl_0_46 cell_2r1w
Xcell_2r1w_1428 vdd_uq20 gnd read_bl_0_41 read_bl_1_41 write_bl_0_41 wwl_0_43 rwl_1_43
+ rwl_0_43 cell_2r1w
Xcell_2r1w_600 vdd_uq18 gnd read_bl_0_54 read_bl_1_54 write_bl_0_54 wwl_0_39 rwl_1_39
+ rwl_0_39 cell_2r1w
Xcell_2r1w_1439 vdd_uq15 gnd read_bl_0_41 read_bl_1_41 write_bl_0_41 wwl_0_32 rwl_1_32
+ rwl_0_32 cell_2r1w
Xcell_2r1w_611 vdd_uq13 gnd read_bl_0_54 read_bl_1_54 write_bl_0_54 wwl_0_28 rwl_1_28
+ rwl_0_28 cell_2r1w
Xcell_2r1w_2107 vdd_uq1 gnd read_bl_0_31 read_bl_1_31 write_bl_0_31 wwl_0_4 rwl_1_4
+ rwl_0_4 cell_2r1w
Xcell_2r1w_1406 vdd_uq0 gnd read_bl_0_42 read_bl_1_42 write_bl_0_42 wwl_0_1 rwl_1_1
+ rwl_0_1 cell_2r1w
Xcell_2r1w_644 vdd_uq28 gnd read_bl_0_53 read_bl_1_53 write_bl_0_53 wwl_0_59 rwl_1_59
+ rwl_0_59 cell_2r1w
Xcell_2r1w_655 vdd_uq23 gnd read_bl_0_53 read_bl_1_53 write_bl_0_53 wwl_0_48 rwl_1_48
+ rwl_0_48 cell_2r1w
Xcell_2r1w_666 vdd_uq17 gnd read_bl_0_53 read_bl_1_53 write_bl_0_53 wwl_0_37 rwl_1_37
+ rwl_0_37 cell_2r1w
Xcell_2r1w_677 vdd_uq12 gnd read_bl_0_53 read_bl_1_53 write_bl_0_53 wwl_0_26 rwl_1_26
+ rwl_0_26 cell_2r1w
Xcell_2r1w_699 vdd_uq1 gnd read_bl_0_53 read_bl_1_53 write_bl_0_53 wwl_0_4 rwl_1_4
+ rwl_0_4 cell_2r1w
Xcell_2r1w_633 vdd_uq2 gnd read_bl_0_54 read_bl_1_54 write_bl_0_54 wwl_0_6 rwl_1_6
+ rwl_0_6 cell_2r1w
Xcell_2r1w_688 vdd_uq6 gnd read_bl_0_53 read_bl_1_53 write_bl_0_53 wwl_0_15 rwl_1_15
+ rwl_0_15 cell_2r1w
Xcell_2r1w_622 vdd_uq7 gnd read_bl_0_54 read_bl_1_54 write_bl_0_54 wwl_0_17 rwl_1_17
+ rwl_0_17 cell_2r1w
Xcell_2r1w_4032 vdd_uq30 gnd read_bl_0_0 read_bl_1_0 write_bl_0_0 wwl_0_63 rwl_1_63
+ rwl_0_63 cell_2r1w
Xcell_2r1w_3331 vdd_uq29 gnd read_bl_0_11 read_bl_1_11 write_bl_0_11 wwl_0_60 rwl_1_60
+ rwl_0_60 cell_2r1w
Xcell_2r1w_4043 vdd_uq25 gnd read_bl_0_0 read_bl_1_0 write_bl_0_0 wwl_0_52 rwl_1_52
+ rwl_0_52 cell_2r1w
Xcell_2r1w_3342 vdd_uq23 gnd read_bl_0_11 read_bl_1_11 write_bl_0_11 wwl_0_49 rwl_1_49
+ rwl_0_49 cell_2r1w
Xcell_2r1w_4054 vdd_uq19 gnd read_bl_0_0 read_bl_1_0 write_bl_0_0 wwl_0_41 rwl_1_41
+ rwl_0_41 cell_2r1w
Xcell_2r1w_3353 vdd_uq18 gnd read_bl_0_11 read_bl_1_11 write_bl_0_11 wwl_0_38 rwl_1_38
+ rwl_0_38 cell_2r1w
Xcell_2r1w_4065 vdd_uq14 gnd read_bl_0_0 read_bl_1_0 write_bl_0_0 wwl_0_30 rwl_1_30
+ rwl_0_30 cell_2r1w
Xcell_2r1w_3320 vdd_uq2 gnd read_bl_0_12 read_bl_1_12 write_bl_0_12 wwl_0_7 rwl_1_7
+ rwl_0_7 cell_2r1w
Xcell_2r1w_4087 vdd_uq3 gnd read_bl_0_0 read_bl_1_0 write_bl_0_0 wwl_0_8 rwl_1_8 rwl_0_8
+ cell_2r1w
Xcell_2r1w_4021 vdd_uq4 gnd read_bl_0_1 read_bl_1_1 write_bl_0_1 wwl_0_10 rwl_1_10
+ rwl_0_10 cell_2r1w
Xcell_2r1w_4076 vdd_uq8 gnd read_bl_0_0 read_bl_1_0 write_bl_0_0 wwl_0_19 rwl_1_19
+ rwl_0_19 cell_2r1w
Xcell_2r1w_4010 vdd_uq9 gnd read_bl_0_1 read_bl_1_1 write_bl_0_1 wwl_0_21 rwl_1_21
+ rwl_0_21 cell_2r1w
Xcell_2r1w_1984 vdd_uq30 gnd read_bl_0_32 read_bl_1_32 write_bl_0_32 wwl_0_63 rwl_1_63
+ rwl_0_63 cell_2r1w
Xcell_2r1w_3397 vdd_uq28 gnd read_bl_0_10 read_bl_1_10 write_bl_0_10 wwl_0_58 rwl_1_58
+ rwl_0_58 cell_2r1w
Xcell_2r1w_2630 vdd_uq27 gnd read_bl_0_22 read_bl_1_22 write_bl_0_22 wwl_0_57 rwl_1_57
+ rwl_0_57 cell_2r1w
Xcell_2r1w_2696 vdd_uq26 gnd read_bl_0_21 read_bl_1_21 write_bl_0_21 wwl_0_55 rwl_1_55
+ rwl_0_55 cell_2r1w
Xcell_2r1w_1995 vdd_uq25 gnd read_bl_0_32 read_bl_1_32 write_bl_0_32 wwl_0_52 rwl_1_52
+ rwl_0_52 cell_2r1w
Xcell_2r1w_2641 vdd_uq22 gnd read_bl_0_22 read_bl_1_22 write_bl_0_22 wwl_0_46 rwl_1_46
+ rwl_0_46 cell_2r1w
Xcell_2r1w_1940 vdd_uq20 gnd read_bl_0_33 read_bl_1_33 write_bl_0_33 wwl_0_43 rwl_1_43
+ rwl_0_43 cell_2r1w
Xcell_2r1w_2652 vdd_uq16 gnd read_bl_0_22 read_bl_1_22 write_bl_0_22 wwl_0_35 rwl_1_35
+ rwl_0_35 cell_2r1w
Xcell_2r1w_1951 vdd_uq15 gnd read_bl_0_33 read_bl_1_33 write_bl_0_33 wwl_0_32 rwl_1_32
+ rwl_0_32 cell_2r1w
Xcell_2r1w_3364 vdd_uq12 gnd read_bl_0_11 read_bl_1_11 write_bl_0_11 wwl_0_27 rwl_1_27
+ rwl_0_27 cell_2r1w
Xcell_2r1w_2663 vdd_uq11 gnd read_bl_0_22 read_bl_1_22 write_bl_0_22 wwl_0_24 rwl_1_24
+ rwl_0_24 cell_2r1w
Xcell_2r1w_3386 vdd_uq1 gnd read_bl_0_11 read_bl_1_11 write_bl_0_11 wwl_0_5 rwl_1_5
+ rwl_0_5 cell_2r1w
Xcell_2r1w_2685 vdd gnd read_bl_0_22 read_bl_1_22 write_bl_0_22 wwl_0_2 rwl_1_2 rwl_0_2
+ cell_2r1w
Xcell_2r1w_1973 vdd_uq4 gnd read_bl_0_33 read_bl_1_33 write_bl_0_33 wwl_0_10 rwl_1_10
+ rwl_0_10 cell_2r1w
Xcell_2r1w_2674 vdd_uq5 gnd read_bl_0_22 read_bl_1_22 write_bl_0_22 wwl_0_13 rwl_1_13
+ rwl_0_13 cell_2r1w
Xcell_2r1w_3375 vdd_uq7 gnd read_bl_0_11 read_bl_1_11 write_bl_0_11 wwl_0_16 rwl_1_16
+ rwl_0_16 cell_2r1w
Xcell_2r1w_1962 vdd_uq9 gnd read_bl_0_33 read_bl_1_33 write_bl_0_33 wwl_0_21 rwl_1_21
+ rwl_0_21 cell_2r1w
Xcell_2r1w_452 vdd_uq28 gnd read_bl_0_56 read_bl_1_56 write_bl_0_56 wwl_0_59 rwl_1_59
+ rwl_0_59 cell_2r1w
Xcell_2r1w_1225 vdd_uq26 gnd read_bl_0_44 read_bl_1_44 write_bl_0_44 wwl_0_54 rwl_1_54
+ rwl_0_54 cell_2r1w
Xcell_2r1w_463 vdd_uq23 gnd read_bl_0_56 read_bl_1_56 write_bl_0_56 wwl_0_48 rwl_1_48
+ rwl_0_48 cell_2r1w
Xcell_2r1w_1236 vdd_uq20 gnd read_bl_0_44 read_bl_1_44 write_bl_0_44 wwl_0_43 rwl_1_43
+ rwl_0_43 cell_2r1w
Xcell_2r1w_1247 vdd_uq15 gnd read_bl_0_44 read_bl_1_44 write_bl_0_44 wwl_0_32 rwl_1_32
+ rwl_0_32 cell_2r1w
Xcell_2r1w_1214 vdd_uq0 gnd read_bl_0_45 read_bl_1_45 write_bl_0_45 wwl_0_1 rwl_1_1
+ rwl_0_1 cell_2r1w
Xcell_2r1w_441 vdd_uq2 gnd read_bl_0_57 read_bl_1_57 write_bl_0_57 wwl_0_6 rwl_1_6
+ rwl_0_6 cell_2r1w
Xcell_2r1w_1269 vdd_uq4 gnd read_bl_0_44 read_bl_1_44 write_bl_0_44 wwl_0_10 rwl_1_10
+ rwl_0_10 cell_2r1w
Xcell_2r1w_1203 vdd_uq5 gnd read_bl_0_45 read_bl_1_45 write_bl_0_45 wwl_0_12 rwl_1_12
+ rwl_0_12 cell_2r1w
Xcell_2r1w_430 vdd_uq7 gnd read_bl_0_57 read_bl_1_57 write_bl_0_57 wwl_0_17 rwl_1_17
+ rwl_0_17 cell_2r1w
Xcell_2r1w_1258 vdd_uq9 gnd read_bl_0_44 read_bl_1_44 write_bl_0_44 wwl_0_21 rwl_1_21
+ rwl_0_21 cell_2r1w
Xcell_2r1w_474 vdd_uq17 gnd read_bl_0_56 read_bl_1_56 write_bl_0_56 wwl_0_37 rwl_1_37
+ rwl_0_37 cell_2r1w
Xcell_2r1w_485 vdd_uq12 gnd read_bl_0_56 read_bl_1_56 write_bl_0_56 wwl_0_26 rwl_1_26
+ rwl_0_26 cell_2r1w
Xcell_2r1w_496 vdd_uq6 gnd read_bl_0_56 read_bl_1_56 write_bl_0_56 wwl_0_15 rwl_1_15
+ rwl_0_15 cell_2r1w
Xcell_2r1w_3150 vdd_uq23 gnd read_bl_0_14 read_bl_1_14 write_bl_0_14 wwl_0_49 rwl_1_49
+ rwl_0_49 cell_2r1w
Xcell_2r1w_3161 vdd_uq18 gnd read_bl_0_14 read_bl_1_14 write_bl_0_14 wwl_0_38 rwl_1_38
+ rwl_0_38 cell_2r1w
Xcell_2r1w_3172 vdd_uq12 gnd read_bl_0_14 read_bl_1_14 write_bl_0_14 wwl_0_27 rwl_1_27
+ rwl_0_27 cell_2r1w
Xcell_2r1w_3194 vdd_uq1 gnd read_bl_0_14 read_bl_1_14 write_bl_0_14 wwl_0_5 rwl_1_5
+ rwl_0_5 cell_2r1w
Xcell_2r1w_3183 vdd_uq7 gnd read_bl_0_14 read_bl_1_14 write_bl_0_14 wwl_0_16 rwl_1_16
+ rwl_0_16 cell_2r1w
Xcell_2r1w_1792 vdd_uq30 gnd read_bl_0_35 read_bl_1_35 write_bl_0_35 wwl_0_63 rwl_1_63
+ rwl_0_63 cell_2r1w
Xcell_2r1w_2460 vdd_uq16 gnd read_bl_0_25 read_bl_1_25 write_bl_0_25 wwl_0_35 rwl_1_35
+ rwl_0_35 cell_2r1w
Xcell_2r1w_2471 vdd_uq11 gnd read_bl_0_25 read_bl_1_25 write_bl_0_25 wwl_0_24 rwl_1_24
+ rwl_0_24 cell_2r1w
Xcell_2r1w_2493 vdd gnd read_bl_0_25 read_bl_1_25 write_bl_0_25 wwl_0_2 rwl_1_2 rwl_0_2
+ cell_2r1w
Xcell_2r1w_1781 vdd_uq4 gnd read_bl_0_36 read_bl_1_36 write_bl_0_36 wwl_0_10 rwl_1_10
+ rwl_0_10 cell_2r1w
Xcell_2r1w_2482 vdd_uq5 gnd read_bl_0_25 read_bl_1_25 write_bl_0_25 wwl_0_13 rwl_1_13
+ rwl_0_13 cell_2r1w
Xcell_2r1w_1770 vdd_uq9 gnd read_bl_0_36 read_bl_1_36 write_bl_0_36 wwl_0_21 rwl_1_21
+ rwl_0_21 cell_2r1w
Xcell_2r1w_1000 vdd_uq10 gnd read_bl_0_48 read_bl_1_48 write_bl_0_48 wwl_0_23 rwl_1_23
+ rwl_0_23 cell_2r1w
Xcell_2r1w_1088 vdd_uq30 gnd read_bl_0_46 read_bl_1_46 write_bl_0_46 wwl_0_63 rwl_1_63
+ rwl_0_63 cell_2r1w
Xcell_2r1w_260 vdd_uq28 gnd read_bl_0_59 read_bl_1_59 write_bl_0_59 wwl_0_59 rwl_1_59
+ rwl_0_59 cell_2r1w
Xcell_2r1w_1033 vdd_uq26 gnd read_bl_0_47 read_bl_1_47 write_bl_0_47 wwl_0_54 rwl_1_54
+ rwl_0_54 cell_2r1w
Xcell_2r1w_1099 vdd_uq25 gnd read_bl_0_46 read_bl_1_46 write_bl_0_46 wwl_0_52 rwl_1_52
+ rwl_0_52 cell_2r1w
Xcell_2r1w_271 vdd_uq23 gnd read_bl_0_59 read_bl_1_59 write_bl_0_59 wwl_0_48 rwl_1_48
+ rwl_0_48 cell_2r1w
Xcell_2r1w_1044 vdd_uq20 gnd read_bl_0_47 read_bl_1_47 write_bl_0_47 wwl_0_43 rwl_1_43
+ rwl_0_43 cell_2r1w
Xcell_2r1w_282 vdd_uq17 gnd read_bl_0_59 read_bl_1_59 write_bl_0_59 wwl_0_37 rwl_1_37
+ rwl_0_37 cell_2r1w
Xcell_2r1w_1055 vdd_uq15 gnd read_bl_0_47 read_bl_1_47 write_bl_0_47 wwl_0_32 rwl_1_32
+ rwl_0_32 cell_2r1w
Xcell_2r1w_293 vdd_uq12 gnd read_bl_0_59 read_bl_1_59 write_bl_0_59 wwl_0_26 rwl_1_26
+ rwl_0_26 cell_2r1w
Xcell_2r1w_1022 vdd_uq0 gnd read_bl_0_48 read_bl_1_48 write_bl_0_48 wwl_0_1 rwl_1_1
+ rwl_0_1 cell_2r1w
Xcell_2r1w_1077 vdd_uq4 gnd read_bl_0_47 read_bl_1_47 write_bl_0_47 wwl_0_10 rwl_1_10
+ rwl_0_10 cell_2r1w
Xcell_2r1w_1011 vdd_uq5 gnd read_bl_0_48 read_bl_1_48 write_bl_0_48 wwl_0_12 rwl_1_12
+ rwl_0_12 cell_2r1w
Xcell_2r1w_1066 vdd_uq9 gnd read_bl_0_47 read_bl_1_47 write_bl_0_47 wwl_0_21 rwl_1_21
+ rwl_0_21 cell_2r1w
Xcell_2r1w_2290 vdd_uq5 gnd read_bl_0_28 read_bl_1_28 write_bl_0_28 wwl_0_13 rwl_1_13
+ rwl_0_13 cell_2r1w
Xcell_2r1w_3908 vdd_uq28 gnd read_bl_0_2 read_bl_1_2 write_bl_0_2 wwl_0_59 rwl_1_59
+ rwl_0_59 cell_2r1w
Xcell_2r1w_3919 vdd_uq23 gnd read_bl_0_2 read_bl_1_2 write_bl_0_2 wwl_0_48 rwl_1_48
+ rwl_0_48 cell_2r1w
Xcell_2r1w_3716 vdd_uq28 gnd read_bl_0_5 read_bl_1_5 write_bl_0_5 wwl_0_59 rwl_1_59
+ rwl_0_59 cell_2r1w
Xcell_2r1w_3727 vdd_uq23 gnd read_bl_0_5 read_bl_1_5 write_bl_0_5 wwl_0_48 rwl_1_48
+ rwl_0_48 cell_2r1w
Xcell_2r1w_3738 vdd_uq17 gnd read_bl_0_5 read_bl_1_5 write_bl_0_5 wwl_0_37 rwl_1_37
+ rwl_0_37 cell_2r1w
Xcell_2r1w_3749 vdd_uq12 gnd read_bl_0_5 read_bl_1_5 write_bl_0_5 wwl_0_26 rwl_1_26
+ rwl_0_26 cell_2r1w
Xcell_2r1w_3705 vdd_uq2 gnd read_bl_0_6 read_bl_1_6 write_bl_0_6 wwl_0_6 rwl_1_6 rwl_0_6
+ cell_2r1w
Xcell_2r1w_804 vdd_uq12 gnd read_bl_0_51 read_bl_1_51 write_bl_0_51 wwl_0_27 rwl_1_27
+ rwl_0_27 cell_2r1w
Xcell_2r1w_837 vdd_uq28 gnd read_bl_0_50 read_bl_1_50 write_bl_0_50 wwl_0_58 rwl_1_58
+ rwl_0_58 cell_2r1w
Xcell_2r1w_848 vdd_uq22 gnd read_bl_0_50 read_bl_1_50 write_bl_0_50 wwl_0_47 rwl_1_47
+ rwl_0_47 cell_2r1w
Xcell_2r1w_859 vdd_uq17 gnd read_bl_0_50 read_bl_1_50 write_bl_0_50 wwl_0_36 rwl_1_36
+ rwl_0_36 cell_2r1w
Xcell_2r1w_826 vdd_uq1 gnd read_bl_0_51 read_bl_1_51 write_bl_0_51 wwl_0_5 rwl_1_5
+ rwl_0_5 cell_2r1w
Xcell_2r1w_815 vdd_uq7 gnd read_bl_0_51 read_bl_1_51 write_bl_0_51 wwl_0_16 rwl_1_16
+ rwl_0_16 cell_2r1w
Xcell_2r1w_3524 vdd_uq28 gnd read_bl_0_8 read_bl_1_8 write_bl_0_8 wwl_0_59 rwl_1_59
+ rwl_0_59 cell_2r1w
Xcell_2r1w_3535 vdd_uq23 gnd read_bl_0_8 read_bl_1_8 write_bl_0_8 wwl_0_48 rwl_1_48
+ rwl_0_48 cell_2r1w
Xcell_2r1w_3513 vdd_uq2 gnd read_bl_0_9 read_bl_1_9 write_bl_0_9 wwl_0_6 rwl_1_6 rwl_0_6
+ cell_2r1w
Xcell_2r1w_3502 vdd_uq7 gnd read_bl_0_9 read_bl_1_9 write_bl_0_9 wwl_0_17 rwl_1_17
+ rwl_0_17 cell_2r1w
Xcell_2r1w_2823 vdd_uq27 gnd read_bl_0_19 read_bl_1_19 write_bl_0_19 wwl_0_56 rwl_1_56
+ rwl_0_56 cell_2r1w
Xcell_2r1w_2889 vdd_uq26 gnd read_bl_0_18 read_bl_1_18 write_bl_0_18 wwl_0_54 rwl_1_54
+ rwl_0_54 cell_2r1w
Xcell_2r1w_2834 vdd_uq21 gnd read_bl_0_19 read_bl_1_19 write_bl_0_19 wwl_0_45 rwl_1_45
+ rwl_0_45 cell_2r1w
Xcell_2r1w_3546 vdd_uq17 gnd read_bl_0_8 read_bl_1_8 write_bl_0_8 wwl_0_37 rwl_1_37
+ rwl_0_37 cell_2r1w
Xcell_2r1w_2845 vdd_uq16 gnd read_bl_0_19 read_bl_1_19 write_bl_0_19 wwl_0_34 rwl_1_34
+ rwl_0_34 cell_2r1w
Xcell_2r1w_3557 vdd_uq12 gnd read_bl_0_8 read_bl_1_8 write_bl_0_8 wwl_0_26 rwl_1_26
+ rwl_0_26 cell_2r1w
Xcell_2r1w_3579 vdd_uq1 gnd read_bl_0_8 read_bl_1_8 write_bl_0_8 wwl_0_4 rwl_1_4 rwl_0_4
+ cell_2r1w
Xcell_2r1w_2812 vdd gnd read_bl_0_20 read_bl_1_20 write_bl_0_20 wwl_0_3 rwl_1_3 rwl_0_3
+ cell_2r1w
Xcell_2r1w_2878 vdd_uq0 gnd read_bl_0_19 read_bl_1_19 write_bl_0_19 wwl_0_1 rwl_1_1
+ rwl_0_1 cell_2r1w
Xcell_2r1w_2867 vdd_uq5 gnd read_bl_0_19 read_bl_1_19 write_bl_0_19 wwl_0_12 rwl_1_12
+ rwl_0_12 cell_2r1w
Xcell_2r1w_2801 vdd_uq6 gnd read_bl_0_20 read_bl_1_20 write_bl_0_20 wwl_0_14 rwl_1_14
+ rwl_0_14 cell_2r1w
Xcell_2r1w_3568 vdd_uq6 gnd read_bl_0_8 read_bl_1_8 write_bl_0_8 wwl_0_15 rwl_1_15
+ rwl_0_15 cell_2r1w
Xcell_2r1w_2856 vdd_uq10 gnd read_bl_0_19 read_bl_1_19 write_bl_0_19 wwl_0_23 rwl_1_23
+ rwl_0_23 cell_2r1w
Xcell_2r1w_645 vdd_uq28 gnd read_bl_0_53 read_bl_1_53 write_bl_0_53 wwl_0_58 rwl_1_58
+ rwl_0_58 cell_2r1w
Xcell_2r1w_2119 vdd_uq27 gnd read_bl_0_30 read_bl_1_30 write_bl_0_30 wwl_0_56 rwl_1_56
+ rwl_0_56 cell_2r1w
Xcell_2r1w_1418 vdd_uq25 gnd read_bl_0_41 read_bl_1_41 write_bl_0_41 wwl_0_53 rwl_1_53
+ rwl_0_53 cell_2r1w
Xcell_2r1w_1429 vdd_uq20 gnd read_bl_0_41 read_bl_1_41 write_bl_0_41 wwl_0_42 rwl_1_42
+ rwl_0_42 cell_2r1w
Xcell_2r1w_601 vdd_uq18 gnd read_bl_0_54 read_bl_1_54 write_bl_0_54 wwl_0_38 rwl_1_38
+ rwl_0_38 cell_2r1w
Xcell_2r1w_612 vdd_uq12 gnd read_bl_0_54 read_bl_1_54 write_bl_0_54 wwl_0_27 rwl_1_27
+ rwl_0_27 cell_2r1w
Xcell_2r1w_634 vdd_uq1 gnd read_bl_0_54 read_bl_1_54 write_bl_0_54 wwl_0_5 rwl_1_5
+ rwl_0_5 cell_2r1w
Xcell_2r1w_2108 vdd gnd read_bl_0_31 read_bl_1_31 write_bl_0_31 wwl_0_3 rwl_1_3 rwl_0_3
+ cell_2r1w
Xcell_2r1w_1407 vdd_uq0 gnd read_bl_0_42 read_bl_1_42 write_bl_0_42 wwl_0_0 rwl_1_0
+ rwl_0_0 cell_2r1w
Xcell_2r1w_623 vdd_uq7 gnd read_bl_0_54 read_bl_1_54 write_bl_0_54 wwl_0_16 rwl_1_16
+ rwl_0_16 cell_2r1w
Xcell_2r1w_656 vdd_uq22 gnd read_bl_0_53 read_bl_1_53 write_bl_0_53 wwl_0_47 rwl_1_47
+ rwl_0_47 cell_2r1w
Xcell_2r1w_667 vdd_uq17 gnd read_bl_0_53 read_bl_1_53 write_bl_0_53 wwl_0_36 rwl_1_36
+ rwl_0_36 cell_2r1w
Xcell_2r1w_678 vdd_uq11 gnd read_bl_0_53 read_bl_1_53 write_bl_0_53 wwl_0_25 rwl_1_25
+ rwl_0_25 cell_2r1w
Xcell_2r1w_689 vdd_uq6 gnd read_bl_0_53 read_bl_1_53 write_bl_0_53 wwl_0_14 rwl_1_14
+ rwl_0_14 cell_2r1w
Xcell_2r1w_4033 vdd_uq30 gnd read_bl_0_0 read_bl_1_0 write_bl_0_0 wwl_0_62 rwl_1_62
+ rwl_0_62 cell_2r1w
Xcell_2r1w_3332 vdd_uq28 gnd read_bl_0_11 read_bl_1_11 write_bl_0_11 wwl_0_59 rwl_1_59
+ rwl_0_59 cell_2r1w
Xcell_2r1w_2631 vdd_uq27 gnd read_bl_0_22 read_bl_1_22 write_bl_0_22 wwl_0_56 rwl_1_56
+ rwl_0_56 cell_2r1w
Xcell_2r1w_4044 vdd_uq24 gnd read_bl_0_0 read_bl_1_0 write_bl_0_0 wwl_0_51 rwl_1_51
+ rwl_0_51 cell_2r1w
Xcell_2r1w_3343 vdd_uq23 gnd read_bl_0_11 read_bl_1_11 write_bl_0_11 wwl_0_48 rwl_1_48
+ rwl_0_48 cell_2r1w
Xcell_2r1w_2642 vdd_uq21 gnd read_bl_0_22 read_bl_1_22 write_bl_0_22 wwl_0_45 rwl_1_45
+ rwl_0_45 cell_2r1w
Xcell_2r1w_4055 vdd_uq19 gnd read_bl_0_0 read_bl_1_0 write_bl_0_0 wwl_0_40 rwl_1_40
+ rwl_0_40 cell_2r1w
Xcell_2r1w_3354 vdd_uq17 gnd read_bl_0_11 read_bl_1_11 write_bl_0_11 wwl_0_37 rwl_1_37
+ rwl_0_37 cell_2r1w
Xcell_2r1w_4000 vdd_uq14 gnd read_bl_0_1 read_bl_1_1 write_bl_0_1 wwl_0_31 rwl_1_31
+ rwl_0_31 cell_2r1w
Xcell_2r1w_4066 vdd_uq13 gnd read_bl_0_0 read_bl_1_0 write_bl_0_0 wwl_0_29 rwl_1_29
+ rwl_0_29 cell_2r1w
Xcell_2r1w_3365 vdd_uq12 gnd read_bl_0_11 read_bl_1_11 write_bl_0_11 wwl_0_26 rwl_1_26
+ rwl_0_26 cell_2r1w
Xcell_2r1w_3387 vdd_uq1 gnd read_bl_0_11 read_bl_1_11 write_bl_0_11 wwl_0_4 rwl_1_4
+ rwl_0_4 cell_2r1w
Xcell_2r1w_2620 vdd gnd read_bl_0_23 read_bl_1_23 write_bl_0_23 wwl_0_3 rwl_1_3 rwl_0_3
+ cell_2r1w
Xcell_2r1w_3321 vdd_uq2 gnd read_bl_0_12 read_bl_1_12 write_bl_0_12 wwl_0_6 rwl_1_6
+ rwl_0_6 cell_2r1w
Xcell_2r1w_4088 vdd_uq2 gnd read_bl_0_0 read_bl_1_0 write_bl_0_0 wwl_0_7 rwl_1_7 rwl_0_7
+ cell_2r1w
Xcell_2r1w_4022 vdd_uq3 gnd read_bl_0_1 read_bl_1_1 write_bl_0_1 wwl_0_9 rwl_1_9 rwl_0_9
+ cell_2r1w
Xcell_2r1w_3376 vdd_uq6 gnd read_bl_0_11 read_bl_1_11 write_bl_0_11 wwl_0_15 rwl_1_15
+ rwl_0_15 cell_2r1w
Xcell_2r1w_3310 vdd_uq7 gnd read_bl_0_12 read_bl_1_12 write_bl_0_12 wwl_0_17 rwl_1_17
+ rwl_0_17 cell_2r1w
Xcell_2r1w_4077 vdd_uq8 gnd read_bl_0_0 read_bl_1_0 write_bl_0_0 wwl_0_18 rwl_1_18
+ rwl_0_18 cell_2r1w
Xcell_2r1w_4011 vdd_uq9 gnd read_bl_0_1 read_bl_1_1 write_bl_0_1 wwl_0_20 rwl_1_20
+ rwl_0_20 cell_2r1w
Xcell_2r1w_1985 vdd_uq30 gnd read_bl_0_32 read_bl_1_32 write_bl_0_32 wwl_0_62 rwl_1_62
+ rwl_0_62 cell_2r1w
Xcell_2r1w_3398 vdd_uq27 gnd read_bl_0_10 read_bl_1_10 write_bl_0_10 wwl_0_57 rwl_1_57
+ rwl_0_57 cell_2r1w
Xcell_2r1w_2697 vdd_uq26 gnd read_bl_0_21 read_bl_1_21 write_bl_0_21 wwl_0_54 rwl_1_54
+ rwl_0_54 cell_2r1w
Xcell_2r1w_1930 vdd_uq25 gnd read_bl_0_33 read_bl_1_33 write_bl_0_33 wwl_0_53 rwl_1_53
+ rwl_0_53 cell_2r1w
Xcell_2r1w_1996 vdd_uq24 gnd read_bl_0_32 read_bl_1_32 write_bl_0_32 wwl_0_51 rwl_1_51
+ rwl_0_51 cell_2r1w
Xcell_2r1w_1941 vdd_uq20 gnd read_bl_0_33 read_bl_1_33 write_bl_0_33 wwl_0_42 rwl_1_42
+ rwl_0_42 cell_2r1w
Xcell_2r1w_2653 vdd_uq16 gnd read_bl_0_22 read_bl_1_22 write_bl_0_22 wwl_0_34 rwl_1_34
+ rwl_0_34 cell_2r1w
Xcell_2r1w_1952 vdd_uq14 gnd read_bl_0_33 read_bl_1_33 write_bl_0_33 wwl_0_31 rwl_1_31
+ rwl_0_31 cell_2r1w
Xcell_2r1w_2686 vdd_uq0 gnd read_bl_0_22 read_bl_1_22 write_bl_0_22 wwl_0_1 rwl_1_1
+ rwl_0_1 cell_2r1w
Xcell_2r1w_1974 vdd_uq3 gnd read_bl_0_33 read_bl_1_33 write_bl_0_33 wwl_0_9 rwl_1_9
+ rwl_0_9 cell_2r1w
Xcell_2r1w_2675 vdd_uq5 gnd read_bl_0_22 read_bl_1_22 write_bl_0_22 wwl_0_12 rwl_1_12
+ rwl_0_12 cell_2r1w
Xcell_2r1w_1963 vdd_uq9 gnd read_bl_0_33 read_bl_1_33 write_bl_0_33 wwl_0_20 rwl_1_20
+ rwl_0_20 cell_2r1w
Xcell_2r1w_2664 vdd_uq10 gnd read_bl_0_22 read_bl_1_22 write_bl_0_22 wwl_0_23 rwl_1_23
+ rwl_0_23 cell_2r1w
Xcell_2r1w_453 vdd_uq28 gnd read_bl_0_56 read_bl_1_56 write_bl_0_56 wwl_0_58 rwl_1_58
+ rwl_0_58 cell_2r1w
Xcell_2r1w_1226 vdd_uq25 gnd read_bl_0_44 read_bl_1_44 write_bl_0_44 wwl_0_53 rwl_1_53
+ rwl_0_53 cell_2r1w
Xcell_2r1w_464 vdd_uq22 gnd read_bl_0_56 read_bl_1_56 write_bl_0_56 wwl_0_47 rwl_1_47
+ rwl_0_47 cell_2r1w
Xcell_2r1w_1237 vdd_uq20 gnd read_bl_0_44 read_bl_1_44 write_bl_0_44 wwl_0_42 rwl_1_42
+ rwl_0_42 cell_2r1w
Xcell_2r1w_475 vdd_uq17 gnd read_bl_0_56 read_bl_1_56 write_bl_0_56 wwl_0_36 rwl_1_36
+ rwl_0_36 cell_2r1w
Xcell_2r1w_1248 vdd_uq14 gnd read_bl_0_44 read_bl_1_44 write_bl_0_44 wwl_0_31 rwl_1_31
+ rwl_0_31 cell_2r1w
Xcell_2r1w_420 vdd_uq12 gnd read_bl_0_57 read_bl_1_57 write_bl_0_57 wwl_0_27 rwl_1_27
+ rwl_0_27 cell_2r1w
Xcell_2r1w_486 vdd_uq11 gnd read_bl_0_56 read_bl_1_56 write_bl_0_56 wwl_0_25 rwl_1_25
+ rwl_0_25 cell_2r1w
Xcell_2r1w_442 vdd_uq1 gnd read_bl_0_57 read_bl_1_57 write_bl_0_57 wwl_0_5 rwl_1_5
+ rwl_0_5 cell_2r1w
Xcell_2r1w_1215 vdd_uq0 gnd read_bl_0_45 read_bl_1_45 write_bl_0_45 wwl_0_0 rwl_1_0
+ rwl_0_0 cell_2r1w
Xcell_2r1w_1204 vdd_uq4 gnd read_bl_0_45 read_bl_1_45 write_bl_0_45 wwl_0_11 rwl_1_11
+ rwl_0_11 cell_2r1w
Xcell_2r1w_497 vdd_uq6 gnd read_bl_0_56 read_bl_1_56 write_bl_0_56 wwl_0_14 rwl_1_14
+ rwl_0_14 cell_2r1w
Xcell_2r1w_431 vdd_uq7 gnd read_bl_0_57 read_bl_1_57 write_bl_0_57 wwl_0_16 rwl_1_16
+ rwl_0_16 cell_2r1w
Xcell_2r1w_1259 vdd_uq9 gnd read_bl_0_44 read_bl_1_44 write_bl_0_44 wwl_0_20 rwl_1_20
+ rwl_0_20 cell_2r1w
Xcell_2r1w_3140 vdd_uq28 gnd read_bl_0_14 read_bl_1_14 write_bl_0_14 wwl_0_59 rwl_1_59
+ rwl_0_59 cell_2r1w
Xcell_2r1w_3151 vdd_uq23 gnd read_bl_0_14 read_bl_1_14 write_bl_0_14 wwl_0_48 rwl_1_48
+ rwl_0_48 cell_2r1w
Xcell_2r1w_2450 vdd_uq21 gnd read_bl_0_25 read_bl_1_25 write_bl_0_25 wwl_0_45 rwl_1_45
+ rwl_0_45 cell_2r1w
Xcell_2r1w_3162 vdd_uq17 gnd read_bl_0_14 read_bl_1_14 write_bl_0_14 wwl_0_37 rwl_1_37
+ rwl_0_37 cell_2r1w
Xcell_2r1w_2461 vdd_uq16 gnd read_bl_0_25 read_bl_1_25 write_bl_0_25 wwl_0_34 rwl_1_34
+ rwl_0_34 cell_2r1w
Xcell_2r1w_3173 vdd_uq12 gnd read_bl_0_14 read_bl_1_14 write_bl_0_14 wwl_0_26 rwl_1_26
+ rwl_0_26 cell_2r1w
Xcell_2r1w_3195 vdd_uq1 gnd read_bl_0_14 read_bl_1_14 write_bl_0_14 wwl_0_4 rwl_1_4
+ rwl_0_4 cell_2r1w
Xcell_2r1w_2483 vdd_uq5 gnd read_bl_0_25 read_bl_1_25 write_bl_0_25 wwl_0_12 rwl_1_12
+ rwl_0_12 cell_2r1w
Xcell_2r1w_3184 vdd_uq6 gnd read_bl_0_14 read_bl_1_14 write_bl_0_14 wwl_0_15 rwl_1_15
+ rwl_0_15 cell_2r1w
Xcell_2r1w_2472 vdd_uq10 gnd read_bl_0_25 read_bl_1_25 write_bl_0_25 wwl_0_23 rwl_1_23
+ rwl_0_23 cell_2r1w
Xcell_2r1w_1793 vdd_uq30 gnd read_bl_0_35 read_bl_1_35 write_bl_0_35 wwl_0_62 rwl_1_62
+ rwl_0_62 cell_2r1w
Xcell_2r1w_1760 vdd_uq14 gnd read_bl_0_36 read_bl_1_36 write_bl_0_36 wwl_0_31 rwl_1_31
+ rwl_0_31 cell_2r1w
Xcell_2r1w_2494 vdd_uq0 gnd read_bl_0_25 read_bl_1_25 write_bl_0_25 wwl_0_1 rwl_1_1
+ rwl_0_1 cell_2r1w
Xcell_2r1w_1782 vdd_uq3 gnd read_bl_0_36 read_bl_1_36 write_bl_0_36 wwl_0_9 rwl_1_9
+ rwl_0_9 cell_2r1w
Xcell_2r1w_1771 vdd_uq9 gnd read_bl_0_36 read_bl_1_36 write_bl_0_36 wwl_0_20 rwl_1_20
+ rwl_0_20 cell_2r1w
Xcell_2r1w_1034 vdd_uq25 gnd read_bl_0_47 read_bl_1_47 write_bl_0_47 wwl_0_53 rwl_1_53
+ rwl_0_53 cell_2r1w
Xcell_2r1w_1023 vdd_uq0 gnd read_bl_0_48 read_bl_1_48 write_bl_0_48 wwl_0_0 rwl_1_0
+ rwl_0_0 cell_2r1w
Xcell_2r1w_1012 vdd_uq4 gnd read_bl_0_48 read_bl_1_48 write_bl_0_48 wwl_0_11 rwl_1_11
+ rwl_0_11 cell_2r1w
Xcell_2r1w_1001 vdd_uq10 gnd read_bl_0_48 read_bl_1_48 write_bl_0_48 wwl_0_22 rwl_1_22
+ rwl_0_22 cell_2r1w
Xcell_2r1w_1089 vdd_uq30 gnd read_bl_0_46 read_bl_1_46 write_bl_0_46 wwl_0_62 rwl_1_62
+ rwl_0_62 cell_2r1w
Xcell_2r1w_261 vdd_uq28 gnd read_bl_0_59 read_bl_1_59 write_bl_0_59 wwl_0_58 rwl_1_58
+ rwl_0_58 cell_2r1w
Xcell_2r1w_272 vdd_uq22 gnd read_bl_0_59 read_bl_1_59 write_bl_0_59 wwl_0_47 rwl_1_47
+ rwl_0_47 cell_2r1w
Xcell_2r1w_1045 vdd_uq20 gnd read_bl_0_47 read_bl_1_47 write_bl_0_47 wwl_0_42 rwl_1_42
+ rwl_0_42 cell_2r1w
Xcell_2r1w_283 vdd_uq17 gnd read_bl_0_59 read_bl_1_59 write_bl_0_59 wwl_0_36 rwl_1_36
+ rwl_0_36 cell_2r1w
Xcell_2r1w_1056 vdd_uq14 gnd read_bl_0_47 read_bl_1_47 write_bl_0_47 wwl_0_31 rwl_1_31
+ rwl_0_31 cell_2r1w
Xcell_2r1w_294 vdd_uq11 gnd read_bl_0_59 read_bl_1_59 write_bl_0_59 wwl_0_25 rwl_1_25
+ rwl_0_25 cell_2r1w
Xcell_2r1w_250 vdd_uq1 gnd read_bl_0_60 read_bl_1_60 write_bl_0_60 wwl_0_5 rwl_1_5
+ rwl_0_5 cell_2r1w
Xcell_2r1w_1078 vdd_uq3 gnd read_bl_0_47 read_bl_1_47 write_bl_0_47 wwl_0_9 rwl_1_9
+ rwl_0_9 cell_2r1w
Xcell_2r1w_1067 vdd_uq9 gnd read_bl_0_47 read_bl_1_47 write_bl_0_47 wwl_0_20 rwl_1_20
+ rwl_0_20 cell_2r1w
Xcell_2r1w_1590 vdd_uq3 gnd read_bl_0_39 read_bl_1_39 write_bl_0_39 wwl_0_9 rwl_1_9
+ rwl_0_9 cell_2r1w
Xcell_2r1w_2291 vdd_uq5 gnd read_bl_0_28 read_bl_1_28 write_bl_0_28 wwl_0_12 rwl_1_12
+ rwl_0_12 cell_2r1w
Xcell_2r1w_2280 vdd_uq10 gnd read_bl_0_28 read_bl_1_28 write_bl_0_28 wwl_0_23 rwl_1_23
+ rwl_0_23 cell_2r1w
Xcell_2r1w_3909 vdd_uq28 gnd read_bl_0_2 read_bl_1_2 write_bl_0_2 wwl_0_58 rwl_1_58
+ rwl_0_58 cell_2r1w
Xcell_2r1w_3717 vdd_uq28 gnd read_bl_0_5 read_bl_1_5 write_bl_0_5 wwl_0_58 rwl_1_58
+ rwl_0_58 cell_2r1w
Xcell_2r1w_3706 vdd_uq1 gnd read_bl_0_6 read_bl_1_6 write_bl_0_6 wwl_0_5 rwl_1_5 rwl_0_5
+ cell_2r1w
Xcell_2r1w_3728 vdd_uq22 gnd read_bl_0_5 read_bl_1_5 write_bl_0_5 wwl_0_47 rwl_1_47
+ rwl_0_47 cell_2r1w
Xcell_2r1w_3739 vdd_uq17 gnd read_bl_0_5 read_bl_1_5 write_bl_0_5 wwl_0_36 rwl_1_36
+ rwl_0_36 cell_2r1w
Xcell_2r1w_805 vdd_uq12 gnd read_bl_0_51 read_bl_1_51 write_bl_0_51 wwl_0_26 rwl_1_26
+ rwl_0_26 cell_2r1w
Xcell_2r1w_827 vdd_uq1 gnd read_bl_0_51 read_bl_1_51 write_bl_0_51 wwl_0_4 rwl_1_4
+ rwl_0_4 cell_2r1w
Xcell_2r1w_816 vdd_uq6 gnd read_bl_0_51 read_bl_1_51 write_bl_0_51 wwl_0_15 rwl_1_15
+ rwl_0_15 cell_2r1w
Xcell_2r1w_838 vdd_uq27 gnd read_bl_0_50 read_bl_1_50 write_bl_0_50 wwl_0_57 rwl_1_57
+ rwl_0_57 cell_2r1w
Xcell_2r1w_849 vdd_uq22 gnd read_bl_0_50 read_bl_1_50 write_bl_0_50 wwl_0_46 rwl_1_46
+ rwl_0_46 cell_2r1w
Xcell_2r1w_3525 vdd_uq28 gnd read_bl_0_8 read_bl_1_8 write_bl_0_8 wwl_0_58 rwl_1_58
+ rwl_0_58 cell_2r1w
Xcell_2r1w_2824 vdd_uq26 gnd read_bl_0_19 read_bl_1_19 write_bl_0_19 wwl_0_55 rwl_1_55
+ rwl_0_55 cell_2r1w
Xcell_2r1w_3536 vdd_uq22 gnd read_bl_0_8 read_bl_1_8 write_bl_0_8 wwl_0_47 rwl_1_47
+ rwl_0_47 cell_2r1w
Xcell_2r1w_3547 vdd_uq17 gnd read_bl_0_8 read_bl_1_8 write_bl_0_8 wwl_0_36 rwl_1_36
+ rwl_0_36 cell_2r1w
Xcell_2r1w_3558 vdd_uq11 gnd read_bl_0_8 read_bl_1_8 write_bl_0_8 wwl_0_25 rwl_1_25
+ rwl_0_25 cell_2r1w
Xcell_2r1w_3514 vdd_uq1 gnd read_bl_0_9 read_bl_1_9 write_bl_0_9 wwl_0_5 rwl_1_5 rwl_0_5
+ cell_2r1w
Xcell_2r1w_2813 vdd gnd read_bl_0_20 read_bl_1_20 write_bl_0_20 wwl_0_2 rwl_1_2 rwl_0_2
+ cell_2r1w
Xcell_2r1w_3569 vdd_uq6 gnd read_bl_0_8 read_bl_1_8 write_bl_0_8 wwl_0_14 rwl_1_14
+ rwl_0_14 cell_2r1w
Xcell_2r1w_2802 vdd_uq5 gnd read_bl_0_20 read_bl_1_20 write_bl_0_20 wwl_0_13 rwl_1_13
+ rwl_0_13 cell_2r1w
Xcell_2r1w_3503 vdd_uq7 gnd read_bl_0_9 read_bl_1_9 write_bl_0_9 wwl_0_16 rwl_1_16
+ rwl_0_16 cell_2r1w
Xcell_2r1w_2835 vdd_uq21 gnd read_bl_0_19 read_bl_1_19 write_bl_0_19 wwl_0_44 rwl_1_44
+ rwl_0_44 cell_2r1w
Xcell_2r1w_2846 vdd_uq15 gnd read_bl_0_19 read_bl_1_19 write_bl_0_19 wwl_0_33 rwl_1_33
+ rwl_0_33 cell_2r1w
Xcell_2r1w_2879 vdd_uq0 gnd read_bl_0_19 read_bl_1_19 write_bl_0_19 wwl_0_0 rwl_1_0
+ rwl_0_0 cell_2r1w
Xcell_2r1w_2868 vdd_uq4 gnd read_bl_0_19 read_bl_1_19 write_bl_0_19 wwl_0_11 rwl_1_11
+ rwl_0_11 cell_2r1w
Xcell_2r1w_2857 vdd_uq10 gnd read_bl_0_19 read_bl_1_19 write_bl_0_19 wwl_0_22 rwl_1_22
+ rwl_0_22 cell_2r1w
Xcell_2r1w_2109 vdd gnd read_bl_0_31 read_bl_1_31 write_bl_0_31 wwl_0_2 rwl_1_2 rwl_0_2
+ cell_2r1w
Xcell_2r1w_1408 vdd_uq30 gnd read_bl_0_41 read_bl_1_41 write_bl_0_41 wwl_0_63 rwl_1_63
+ rwl_0_63 cell_2r1w
Xcell_2r1w_646 vdd_uq27 gnd read_bl_0_53 read_bl_1_53 write_bl_0_53 wwl_0_57 rwl_1_57
+ rwl_0_57 cell_2r1w
Xcell_2r1w_1419 vdd_uq25 gnd read_bl_0_41 read_bl_1_41 write_bl_0_41 wwl_0_52 rwl_1_52
+ rwl_0_52 cell_2r1w
Xcell_2r1w_657 vdd_uq22 gnd read_bl_0_53 read_bl_1_53 write_bl_0_53 wwl_0_46 rwl_1_46
+ rwl_0_46 cell_2r1w
Xcell_2r1w_602 vdd_uq17 gnd read_bl_0_54 read_bl_1_54 write_bl_0_54 wwl_0_37 rwl_1_37
+ rwl_0_37 cell_2r1w
Xcell_2r1w_668 vdd_uq16 gnd read_bl_0_53 read_bl_1_53 write_bl_0_53 wwl_0_35 rwl_1_35
+ rwl_0_35 cell_2r1w
Xcell_2r1w_613 vdd_uq12 gnd read_bl_0_54 read_bl_1_54 write_bl_0_54 wwl_0_26 rwl_1_26
+ rwl_0_26 cell_2r1w
Xcell_2r1w_679 vdd_uq11 gnd read_bl_0_53 read_bl_1_53 write_bl_0_53 wwl_0_24 rwl_1_24
+ rwl_0_24 cell_2r1w
Xcell_2r1w_635 vdd_uq1 gnd read_bl_0_54 read_bl_1_54 write_bl_0_54 wwl_0_4 rwl_1_4
+ rwl_0_4 cell_2r1w
Xcell_2r1w_624 vdd_uq6 gnd read_bl_0_54 read_bl_1_54 write_bl_0_54 wwl_0_15 rwl_1_15
+ rwl_0_15 cell_2r1w
Xcell_2r1w_4001 vdd_uq14 gnd read_bl_0_1 read_bl_1_1 write_bl_0_1 wwl_0_30 rwl_1_30
+ rwl_0_30 cell_2r1w
Xcell_2r1w_4012 vdd_uq8 gnd read_bl_0_1 read_bl_1_1 write_bl_0_1 wwl_0_19 rwl_1_19
+ rwl_0_19 cell_2r1w
Xcell_2r1w_1920 vdd_uq30 gnd read_bl_0_33 read_bl_1_33 write_bl_0_33 wwl_0_63 rwl_1_63
+ rwl_0_63 cell_2r1w
Xcell_2r1w_4034 vdd_uq29 gnd read_bl_0_0 read_bl_1_0 write_bl_0_0 wwl_0_61 rwl_1_61
+ rwl_0_61 cell_2r1w
Xcell_2r1w_3333 vdd_uq28 gnd read_bl_0_11 read_bl_1_11 write_bl_0_11 wwl_0_58 rwl_1_58
+ rwl_0_58 cell_2r1w
Xcell_2r1w_2632 vdd_uq26 gnd read_bl_0_22 read_bl_1_22 write_bl_0_22 wwl_0_55 rwl_1_55
+ rwl_0_55 cell_2r1w
Xcell_2r1w_3399 vdd_uq27 gnd read_bl_0_10 read_bl_1_10 write_bl_0_10 wwl_0_56 rwl_1_56
+ rwl_0_56 cell_2r1w
Xcell_2r1w_1931 vdd_uq25 gnd read_bl_0_33 read_bl_1_33 write_bl_0_33 wwl_0_52 rwl_1_52
+ rwl_0_52 cell_2r1w
Xcell_2r1w_4045 vdd_uq24 gnd read_bl_0_0 read_bl_1_0 write_bl_0_0 wwl_0_50 rwl_1_50
+ rwl_0_50 cell_2r1w
Xcell_2r1w_3344 vdd_uq22 gnd read_bl_0_11 read_bl_1_11 write_bl_0_11 wwl_0_47 rwl_1_47
+ rwl_0_47 cell_2r1w
Xcell_2r1w_2643 vdd_uq21 gnd read_bl_0_22 read_bl_1_22 write_bl_0_22 wwl_0_44 rwl_1_44
+ rwl_0_44 cell_2r1w
Xcell_2r1w_4056 vdd_uq18 gnd read_bl_0_0 read_bl_1_0 write_bl_0_0 wwl_0_39 rwl_1_39
+ rwl_0_39 cell_2r1w
Xcell_2r1w_3355 vdd_uq17 gnd read_bl_0_11 read_bl_1_11 write_bl_0_11 wwl_0_36 rwl_1_36
+ rwl_0_36 cell_2r1w
Xcell_2r1w_2654 vdd_uq15 gnd read_bl_0_22 read_bl_1_22 write_bl_0_22 wwl_0_33 rwl_1_33
+ rwl_0_33 cell_2r1w
Xcell_2r1w_3300 vdd_uq12 gnd read_bl_0_12 read_bl_1_12 write_bl_0_12 wwl_0_27 rwl_1_27
+ rwl_0_27 cell_2r1w
Xcell_2r1w_4067 vdd_uq13 gnd read_bl_0_0 read_bl_1_0 write_bl_0_0 wwl_0_28 rwl_1_28
+ rwl_0_28 cell_2r1w
Xcell_2r1w_3366 vdd_uq11 gnd read_bl_0_11 read_bl_1_11 write_bl_0_11 wwl_0_25 rwl_1_25
+ rwl_0_25 cell_2r1w
Xcell_2r1w_3322 vdd_uq1 gnd read_bl_0_12 read_bl_1_12 write_bl_0_12 wwl_0_5 rwl_1_5
+ rwl_0_5 cell_2r1w
Xcell_2r1w_3388 vdd gnd read_bl_0_11 read_bl_1_11 write_bl_0_11 wwl_0_3 rwl_1_3 rwl_0_3
+ cell_2r1w
Xcell_2r1w_2621 vdd gnd read_bl_0_23 read_bl_1_23 write_bl_0_23 wwl_0_2 rwl_1_2 rwl_0_2
+ cell_2r1w
Xcell_2r1w_4089 vdd_uq2 gnd read_bl_0_0 read_bl_1_0 write_bl_0_0 wwl_0_6 rwl_1_6 rwl_0_6
+ cell_2r1w
Xcell_2r1w_4023 vdd_uq3 gnd read_bl_0_1 read_bl_1_1 write_bl_0_1 wwl_0_8 rwl_1_8 rwl_0_8
+ cell_2r1w
Xcell_2r1w_3377 vdd_uq6 gnd read_bl_0_11 read_bl_1_11 write_bl_0_11 wwl_0_14 rwl_1_14
+ rwl_0_14 cell_2r1w
Xcell_2r1w_2610 vdd_uq5 gnd read_bl_0_23 read_bl_1_23 write_bl_0_23 wwl_0_13 rwl_1_13
+ rwl_0_13 cell_2r1w
Xcell_2r1w_3311 vdd_uq7 gnd read_bl_0_12 read_bl_1_12 write_bl_0_12 wwl_0_16 rwl_1_16
+ rwl_0_16 cell_2r1w
Xcell_2r1w_4078 vdd_uq7 gnd read_bl_0_0 read_bl_1_0 write_bl_0_0 wwl_0_17 rwl_1_17
+ rwl_0_17 cell_2r1w
Xcell_2r1w_2665 vdd_uq10 gnd read_bl_0_22 read_bl_1_22 write_bl_0_22 wwl_0_22 rwl_1_22
+ rwl_0_22 cell_2r1w
Xcell_2r1w_1986 vdd_uq29 gnd read_bl_0_32 read_bl_1_32 write_bl_0_32 wwl_0_61 rwl_1_61
+ rwl_0_61 cell_2r1w
Xcell_2r1w_2698 vdd_uq25 gnd read_bl_0_21 read_bl_1_21 write_bl_0_21 wwl_0_53 rwl_1_53
+ rwl_0_53 cell_2r1w
Xcell_2r1w_1997 vdd_uq24 gnd read_bl_0_32 read_bl_1_32 write_bl_0_32 wwl_0_50 rwl_1_50
+ rwl_0_50 cell_2r1w
Xcell_2r1w_1942 vdd_uq19 gnd read_bl_0_33 read_bl_1_33 write_bl_0_33 wwl_0_41 rwl_1_41
+ rwl_0_41 cell_2r1w
Xcell_2r1w_1953 vdd_uq14 gnd read_bl_0_33 read_bl_1_33 write_bl_0_33 wwl_0_30 rwl_1_30
+ rwl_0_30 cell_2r1w
Xcell_2r1w_2687 vdd_uq0 gnd read_bl_0_22 read_bl_1_22 write_bl_0_22 wwl_0_0 rwl_1_0
+ rwl_0_0 cell_2r1w
Xcell_2r1w_1975 vdd_uq3 gnd read_bl_0_33 read_bl_1_33 write_bl_0_33 wwl_0_8 rwl_1_8
+ rwl_0_8 cell_2r1w
Xcell_2r1w_2676 vdd_uq4 gnd read_bl_0_22 read_bl_1_22 write_bl_0_22 wwl_0_11 rwl_1_11
+ rwl_0_11 cell_2r1w
Xcell_2r1w_1964 vdd_uq8 gnd read_bl_0_33 read_bl_1_33 write_bl_0_33 wwl_0_19 rwl_1_19
+ rwl_0_19 cell_2r1w
Xcell_2r1w_1216 vdd_uq30 gnd read_bl_0_44 read_bl_1_44 write_bl_0_44 wwl_0_63 rwl_1_63
+ rwl_0_63 cell_2r1w
Xcell_2r1w_1205 vdd_uq4 gnd read_bl_0_45 read_bl_1_45 write_bl_0_45 wwl_0_10 rwl_1_10
+ rwl_0_10 cell_2r1w
Xcell_2r1w_454 vdd_uq27 gnd read_bl_0_56 read_bl_1_56 write_bl_0_56 wwl_0_57 rwl_1_57
+ rwl_0_57 cell_2r1w
Xcell_2r1w_1227 vdd_uq25 gnd read_bl_0_44 read_bl_1_44 write_bl_0_44 wwl_0_52 rwl_1_52
+ rwl_0_52 cell_2r1w
Xcell_2r1w_465 vdd_uq22 gnd read_bl_0_56 read_bl_1_56 write_bl_0_56 wwl_0_46 rwl_1_46
+ rwl_0_46 cell_2r1w
Xcell_2r1w_1238 vdd_uq19 gnd read_bl_0_44 read_bl_1_44 write_bl_0_44 wwl_0_41 rwl_1_41
+ rwl_0_41 cell_2r1w
Xcell_2r1w_410 vdd_uq17 gnd read_bl_0_57 read_bl_1_57 write_bl_0_57 wwl_0_37 rwl_1_37
+ rwl_0_37 cell_2r1w
Xcell_2r1w_476 vdd_uq16 gnd read_bl_0_56 read_bl_1_56 write_bl_0_56 wwl_0_35 rwl_1_35
+ rwl_0_35 cell_2r1w
Xcell_2r1w_1249 vdd_uq14 gnd read_bl_0_44 read_bl_1_44 write_bl_0_44 wwl_0_30 rwl_1_30
+ rwl_0_30 cell_2r1w
Xcell_2r1w_421 vdd_uq12 gnd read_bl_0_57 read_bl_1_57 write_bl_0_57 wwl_0_26 rwl_1_26
+ rwl_0_26 cell_2r1w
Xcell_2r1w_487 vdd_uq11 gnd read_bl_0_56 read_bl_1_56 write_bl_0_56 wwl_0_24 rwl_1_24
+ rwl_0_24 cell_2r1w
Xcell_2r1w_443 vdd_uq1 gnd read_bl_0_57 read_bl_1_57 write_bl_0_57 wwl_0_4 rwl_1_4
+ rwl_0_4 cell_2r1w
Xcell_2r1w_498 vdd_uq5 gnd read_bl_0_56 read_bl_1_56 write_bl_0_56 wwl_0_13 rwl_1_13
+ rwl_0_13 cell_2r1w
Xcell_2r1w_432 vdd_uq6 gnd read_bl_0_57 read_bl_1_57 write_bl_0_57 wwl_0_15 rwl_1_15
+ rwl_0_15 cell_2r1w
Xcell_2r1w_3141 vdd_uq28 gnd read_bl_0_14 read_bl_1_14 write_bl_0_14 wwl_0_58 rwl_1_58
+ rwl_0_58 cell_2r1w
Xcell_2r1w_2440 vdd_uq26 gnd read_bl_0_25 read_bl_1_25 write_bl_0_25 wwl_0_55 rwl_1_55
+ rwl_0_55 cell_2r1w
Xcell_2r1w_3152 vdd_uq22 gnd read_bl_0_14 read_bl_1_14 write_bl_0_14 wwl_0_47 rwl_1_47
+ rwl_0_47 cell_2r1w
Xcell_2r1w_2451 vdd_uq21 gnd read_bl_0_25 read_bl_1_25 write_bl_0_25 wwl_0_44 rwl_1_44
+ rwl_0_44 cell_2r1w
Xcell_2r1w_1750 vdd_uq19 gnd read_bl_0_36 read_bl_1_36 write_bl_0_36 wwl_0_41 rwl_1_41
+ rwl_0_41 cell_2r1w
Xcell_2r1w_3163 vdd_uq17 gnd read_bl_0_14 read_bl_1_14 write_bl_0_14 wwl_0_36 rwl_1_36
+ rwl_0_36 cell_2r1w
Xcell_2r1w_2462 vdd_uq15 gnd read_bl_0_25 read_bl_1_25 write_bl_0_25 wwl_0_33 rwl_1_33
+ rwl_0_33 cell_2r1w
Xcell_2r1w_1761 vdd_uq14 gnd read_bl_0_36 read_bl_1_36 write_bl_0_36 wwl_0_30 rwl_1_30
+ rwl_0_30 cell_2r1w
Xcell_2r1w_3174 vdd_uq11 gnd read_bl_0_14 read_bl_1_14 write_bl_0_14 wwl_0_25 rwl_1_25
+ rwl_0_25 cell_2r1w
Xcell_2r1w_3130 vdd_uq1 gnd read_bl_0_15 read_bl_1_15 write_bl_0_15 wwl_0_5 rwl_1_5
+ rwl_0_5 cell_2r1w
Xcell_2r1w_3196 vdd gnd read_bl_0_14 read_bl_1_14 write_bl_0_14 wwl_0_3 rwl_1_3 rwl_0_3
+ cell_2r1w
Xcell_2r1w_2495 vdd_uq0 gnd read_bl_0_25 read_bl_1_25 write_bl_0_25 wwl_0_0 rwl_1_0
+ rwl_0_0 cell_2r1w
Xcell_2r1w_2484 vdd_uq4 gnd read_bl_0_25 read_bl_1_25 write_bl_0_25 wwl_0_11 rwl_1_11
+ rwl_0_11 cell_2r1w
Xcell_2r1w_3185 vdd_uq6 gnd read_bl_0_14 read_bl_1_14 write_bl_0_14 wwl_0_14 rwl_1_14
+ rwl_0_14 cell_2r1w
Xcell_2r1w_1772 vdd_uq8 gnd read_bl_0_36 read_bl_1_36 write_bl_0_36 wwl_0_19 rwl_1_19
+ rwl_0_19 cell_2r1w
Xcell_2r1w_2473 vdd_uq10 gnd read_bl_0_25 read_bl_1_25 write_bl_0_25 wwl_0_22 rwl_1_22
+ rwl_0_22 cell_2r1w
Xcell_2r1w_1794 vdd_uq29 gnd read_bl_0_35 read_bl_1_35 write_bl_0_35 wwl_0_61 rwl_1_61
+ rwl_0_61 cell_2r1w
Xcell_2r1w_1783 vdd_uq3 gnd read_bl_0_36 read_bl_1_36 write_bl_0_36 wwl_0_8 rwl_1_8
+ rwl_0_8 cell_2r1w
Xcell_2r1w_1024 vdd_uq30 gnd read_bl_0_47 read_bl_1_47 write_bl_0_47 wwl_0_63 rwl_1_63
+ rwl_0_63 cell_2r1w
Xcell_2r1w_1035 vdd_uq25 gnd read_bl_0_47 read_bl_1_47 write_bl_0_47 wwl_0_52 rwl_1_52
+ rwl_0_52 cell_2r1w
Xcell_2r1w_1046 vdd_uq19 gnd read_bl_0_47 read_bl_1_47 write_bl_0_47 wwl_0_41 rwl_1_41
+ rwl_0_41 cell_2r1w
Xcell_2r1w_1057 vdd_uq14 gnd read_bl_0_47 read_bl_1_47 write_bl_0_47 wwl_0_30 rwl_1_30
+ rwl_0_30 cell_2r1w
Xcell_2r1w_1013 vdd_uq4 gnd read_bl_0_48 read_bl_1_48 write_bl_0_48 wwl_0_10 rwl_1_10
+ rwl_0_10 cell_2r1w
Xcell_2r1w_1068 vdd_uq8 gnd read_bl_0_47 read_bl_1_47 write_bl_0_47 wwl_0_19 rwl_1_19
+ rwl_0_19 cell_2r1w
Xcell_2r1w_1002 vdd_uq9 gnd read_bl_0_48 read_bl_1_48 write_bl_0_48 wwl_0_21 rwl_1_21
+ rwl_0_21 cell_2r1w
Xcell_2r1w_262 vdd_uq27 gnd read_bl_0_59 read_bl_1_59 write_bl_0_59 wwl_0_57 rwl_1_57
+ rwl_0_57 cell_2r1w
Xcell_2r1w_273 vdd_uq22 gnd read_bl_0_59 read_bl_1_59 write_bl_0_59 wwl_0_46 rwl_1_46
+ rwl_0_46 cell_2r1w
Xcell_2r1w_284 vdd_uq16 gnd read_bl_0_59 read_bl_1_59 write_bl_0_59 wwl_0_35 rwl_1_35
+ rwl_0_35 cell_2r1w
Xcell_2r1w_295 vdd_uq11 gnd read_bl_0_59 read_bl_1_59 write_bl_0_59 wwl_0_24 rwl_1_24
+ rwl_0_24 cell_2r1w
Xcell_2r1w_251 vdd_uq1 gnd read_bl_0_60 read_bl_1_60 write_bl_0_60 wwl_0_4 rwl_1_4
+ rwl_0_4 cell_2r1w
Xcell_2r1w_1079 vdd_uq3 gnd read_bl_0_47 read_bl_1_47 write_bl_0_47 wwl_0_8 rwl_1_8
+ rwl_0_8 cell_2r1w
Xcell_2r1w_240 vdd_uq6 gnd read_bl_0_60 read_bl_1_60 write_bl_0_60 wwl_0_15 rwl_1_15
+ rwl_0_15 cell_2r1w
Xcell_2r1w_2270 vdd_uq15 gnd read_bl_0_28 read_bl_1_28 write_bl_0_28 wwl_0_33 rwl_1_33
+ rwl_0_33 cell_2r1w
Xcell_2r1w_1591 vdd_uq3 gnd read_bl_0_39 read_bl_1_39 write_bl_0_39 wwl_0_8 rwl_1_8
+ rwl_0_8 cell_2r1w
Xcell_2r1w_2292 vdd_uq4 gnd read_bl_0_28 read_bl_1_28 write_bl_0_28 wwl_0_11 rwl_1_11
+ rwl_0_11 cell_2r1w
Xcell_2r1w_1580 vdd_uq8 gnd read_bl_0_39 read_bl_1_39 write_bl_0_39 wwl_0_19 rwl_1_19
+ rwl_0_19 cell_2r1w
Xcell_2r1w_2281 vdd_uq10 gnd read_bl_0_28 read_bl_1_28 write_bl_0_28 wwl_0_22 rwl_1_22
+ rwl_0_22 cell_2r1w
Xcell_2r1w_3718 vdd_uq27 gnd read_bl_0_5 read_bl_1_5 write_bl_0_5 wwl_0_57 rwl_1_57
+ rwl_0_57 cell_2r1w
Xcell_2r1w_3729 vdd_uq22 gnd read_bl_0_5 read_bl_1_5 write_bl_0_5 wwl_0_46 rwl_1_46
+ rwl_0_46 cell_2r1w
Xcell_2r1w_3707 vdd_uq1 gnd read_bl_0_6 read_bl_1_6 write_bl_0_6 wwl_0_4 rwl_1_4 rwl_0_4
+ cell_2r1w
Xcell_2r1w_839 vdd_uq27 gnd read_bl_0_50 read_bl_1_50 write_bl_0_50 wwl_0_56 rwl_1_56
+ rwl_0_56 cell_2r1w
Xcell_2r1w_806 vdd_uq11 gnd read_bl_0_51 read_bl_1_51 write_bl_0_51 wwl_0_25 rwl_1_25
+ rwl_0_25 cell_2r1w
Xcell_2r1w_828 vdd gnd read_bl_0_51 read_bl_1_51 write_bl_0_51 wwl_0_3 rwl_1_3 rwl_0_3
+ cell_2r1w
Xcell_2r1w_817 vdd_uq6 gnd read_bl_0_51 read_bl_1_51 write_bl_0_51 wwl_0_14 rwl_1_14
+ rwl_0_14 cell_2r1w
Xcell_2r1w_3526 vdd_uq27 gnd read_bl_0_8 read_bl_1_8 write_bl_0_8 wwl_0_57 rwl_1_57
+ rwl_0_57 cell_2r1w
Xcell_2r1w_2825 vdd_uq26 gnd read_bl_0_19 read_bl_1_19 write_bl_0_19 wwl_0_54 rwl_1_54
+ rwl_0_54 cell_2r1w
Xcell_2r1w_3537 vdd_uq22 gnd read_bl_0_8 read_bl_1_8 write_bl_0_8 wwl_0_46 rwl_1_46
+ rwl_0_46 cell_2r1w
Xcell_2r1w_2836 vdd_uq20 gnd read_bl_0_19 read_bl_1_19 write_bl_0_19 wwl_0_43 rwl_1_43
+ rwl_0_43 cell_2r1w
Xcell_2r1w_3548 vdd_uq16 gnd read_bl_0_8 read_bl_1_8 write_bl_0_8 wwl_0_35 rwl_1_35
+ rwl_0_35 cell_2r1w
Xcell_2r1w_2847 vdd_uq15 gnd read_bl_0_19 read_bl_1_19 write_bl_0_19 wwl_0_32 rwl_1_32
+ rwl_0_32 cell_2r1w
Xcell_2r1w_3559 vdd_uq11 gnd read_bl_0_8 read_bl_1_8 write_bl_0_8 wwl_0_24 rwl_1_24
+ rwl_0_24 cell_2r1w
Xcell_2r1w_3515 vdd_uq1 gnd read_bl_0_9 read_bl_1_9 write_bl_0_9 wwl_0_4 rwl_1_4 rwl_0_4
+ cell_2r1w
Xcell_2r1w_2814 vdd_uq0 gnd read_bl_0_20 read_bl_1_20 write_bl_0_20 wwl_0_1 rwl_1_1
+ rwl_0_1 cell_2r1w
Xcell_2r1w_2803 vdd_uq5 gnd read_bl_0_20 read_bl_1_20 write_bl_0_20 wwl_0_12 rwl_1_12
+ rwl_0_12 cell_2r1w
Xcell_2r1w_3504 vdd_uq6 gnd read_bl_0_9 read_bl_1_9 write_bl_0_9 wwl_0_15 rwl_1_15
+ rwl_0_15 cell_2r1w
Xcell_2r1w_2858 vdd_uq9 gnd read_bl_0_19 read_bl_1_19 write_bl_0_19 wwl_0_21 rwl_1_21
+ rwl_0_21 cell_2r1w
Xcell_2r1w_2869 vdd_uq4 gnd read_bl_0_19 read_bl_1_19 write_bl_0_19 wwl_0_10 rwl_1_10
+ rwl_0_10 cell_2r1w
Xcell_2r1w_1409 vdd_uq30 gnd read_bl_0_41 read_bl_1_41 write_bl_0_41 wwl_0_62 rwl_1_62
+ rwl_0_62 cell_2r1w
Xcell_2r1w_647 vdd_uq27 gnd read_bl_0_53 read_bl_1_53 write_bl_0_53 wwl_0_56 rwl_1_56
+ rwl_0_56 cell_2r1w
Xcell_2r1w_658 vdd_uq21 gnd read_bl_0_53 read_bl_1_53 write_bl_0_53 wwl_0_45 rwl_1_45
+ rwl_0_45 cell_2r1w
Xcell_2r1w_603 vdd_uq17 gnd read_bl_0_54 read_bl_1_54 write_bl_0_54 wwl_0_36 rwl_1_36
+ rwl_0_36 cell_2r1w
Xcell_2r1w_669 vdd_uq16 gnd read_bl_0_53 read_bl_1_53 write_bl_0_53 wwl_0_34 rwl_1_34
+ rwl_0_34 cell_2r1w
Xcell_2r1w_614 vdd_uq11 gnd read_bl_0_54 read_bl_1_54 write_bl_0_54 wwl_0_25 rwl_1_25
+ rwl_0_25 cell_2r1w
Xcell_2r1w_636 vdd gnd read_bl_0_54 read_bl_1_54 write_bl_0_54 wwl_0_3 rwl_1_3 rwl_0_3
+ cell_2r1w
Xcell_2r1w_625 vdd_uq6 gnd read_bl_0_54 read_bl_1_54 write_bl_0_54 wwl_0_14 rwl_1_14
+ rwl_0_14 cell_2r1w
Xcell_2r1w_4035 vdd_uq29 gnd read_bl_0_0 read_bl_1_0 write_bl_0_0 wwl_0_60 rwl_1_60
+ rwl_0_60 cell_2r1w
Xcell_2r1w_4046 vdd_uq23 gnd read_bl_0_0 read_bl_1_0 write_bl_0_0 wwl_0_49 rwl_1_49
+ rwl_0_49 cell_2r1w
Xcell_2r1w_4002 vdd_uq13 gnd read_bl_0_1 read_bl_1_1 write_bl_0_1 wwl_0_29 rwl_1_29
+ rwl_0_29 cell_2r1w
Xcell_2r1w_3301 vdd_uq12 gnd read_bl_0_12 read_bl_1_12 write_bl_0_12 wwl_0_26 rwl_1_26
+ rwl_0_26 cell_2r1w
Xcell_2r1w_4024 vdd_uq2 gnd read_bl_0_1 read_bl_1_1 write_bl_0_1 wwl_0_7 rwl_1_7 rwl_0_7
+ cell_2r1w
Xcell_2r1w_4013 vdd_uq8 gnd read_bl_0_1 read_bl_1_1 write_bl_0_1 wwl_0_18 rwl_1_18
+ rwl_0_18 cell_2r1w
Xcell_2r1w_2688 vdd_uq30 gnd read_bl_0_21 read_bl_1_21 write_bl_0_21 wwl_0_63 rwl_1_63
+ rwl_0_63 cell_2r1w
Xcell_2r1w_1921 vdd_uq30 gnd read_bl_0_33 read_bl_1_33 write_bl_0_33 wwl_0_62 rwl_1_62
+ rwl_0_62 cell_2r1w
Xcell_2r1w_3334 vdd_uq27 gnd read_bl_0_11 read_bl_1_11 write_bl_0_11 wwl_0_57 rwl_1_57
+ rwl_0_57 cell_2r1w
Xcell_2r1w_2633 vdd_uq26 gnd read_bl_0_22 read_bl_1_22 write_bl_0_22 wwl_0_54 rwl_1_54
+ rwl_0_54 cell_2r1w
Xcell_2r1w_2699 vdd_uq25 gnd read_bl_0_21 read_bl_1_21 write_bl_0_21 wwl_0_52 rwl_1_52
+ rwl_0_52 cell_2r1w
Xcell_2r1w_1932 vdd_uq24 gnd read_bl_0_33 read_bl_1_33 write_bl_0_33 wwl_0_51 rwl_1_51
+ rwl_0_51 cell_2r1w
Xcell_2r1w_3345 vdd_uq22 gnd read_bl_0_11 read_bl_1_11 write_bl_0_11 wwl_0_46 rwl_1_46
+ rwl_0_46 cell_2r1w
Xcell_2r1w_2644 vdd_uq20 gnd read_bl_0_22 read_bl_1_22 write_bl_0_22 wwl_0_43 rwl_1_43
+ rwl_0_43 cell_2r1w
Xcell_2r1w_1943 vdd_uq19 gnd read_bl_0_33 read_bl_1_33 write_bl_0_33 wwl_0_40 rwl_1_40
+ rwl_0_40 cell_2r1w
Xcell_2r1w_4057 vdd_uq18 gnd read_bl_0_0 read_bl_1_0 write_bl_0_0 wwl_0_38 rwl_1_38
+ rwl_0_38 cell_2r1w
Xcell_2r1w_3356 vdd_uq16 gnd read_bl_0_11 read_bl_1_11 write_bl_0_11 wwl_0_35 rwl_1_35
+ rwl_0_35 cell_2r1w
Xcell_2r1w_2655 vdd_uq15 gnd read_bl_0_22 read_bl_1_22 write_bl_0_22 wwl_0_32 rwl_1_32
+ rwl_0_32 cell_2r1w
Xcell_2r1w_1954 vdd_uq13 gnd read_bl_0_33 read_bl_1_33 write_bl_0_33 wwl_0_29 rwl_1_29
+ rwl_0_29 cell_2r1w
Xcell_2r1w_4068 vdd_uq12 gnd read_bl_0_0 read_bl_1_0 write_bl_0_0 wwl_0_27 rwl_1_27
+ rwl_0_27 cell_2r1w
Xcell_2r1w_3367 vdd_uq11 gnd read_bl_0_11 read_bl_1_11 write_bl_0_11 wwl_0_24 rwl_1_24
+ rwl_0_24 cell_2r1w
Xcell_2r1w_3323 vdd_uq1 gnd read_bl_0_12 read_bl_1_12 write_bl_0_12 wwl_0_4 rwl_1_4
+ rwl_0_4 cell_2r1w
Xcell_2r1w_3389 vdd gnd read_bl_0_11 read_bl_1_11 write_bl_0_11 wwl_0_2 rwl_1_2 rwl_0_2
+ cell_2r1w
Xcell_2r1w_2622 vdd_uq0 gnd read_bl_0_23 read_bl_1_23 write_bl_0_23 wwl_0_1 rwl_1_1
+ rwl_0_1 cell_2r1w
Xcell_2r1w_1910 vdd_uq3 gnd read_bl_0_34 read_bl_1_34 write_bl_0_34 wwl_0_9 rwl_1_9
+ rwl_0_9 cell_2r1w
Xcell_2r1w_2677 vdd_uq4 gnd read_bl_0_22 read_bl_1_22 write_bl_0_22 wwl_0_10 rwl_1_10
+ rwl_0_10 cell_2r1w
Xcell_2r1w_2611 vdd_uq5 gnd read_bl_0_23 read_bl_1_23 write_bl_0_23 wwl_0_12 rwl_1_12
+ rwl_0_12 cell_2r1w
Xcell_2r1w_3378 vdd_uq5 gnd read_bl_0_11 read_bl_1_11 write_bl_0_11 wwl_0_13 rwl_1_13
+ rwl_0_13 cell_2r1w
Xcell_2r1w_3312 vdd_uq6 gnd read_bl_0_12 read_bl_1_12 write_bl_0_12 wwl_0_15 rwl_1_15
+ rwl_0_15 cell_2r1w
Xcell_2r1w_4079 vdd_uq7 gnd read_bl_0_0 read_bl_1_0 write_bl_0_0 wwl_0_16 rwl_1_16
+ rwl_0_16 cell_2r1w
Xcell_2r1w_2666 vdd_uq9 gnd read_bl_0_22 read_bl_1_22 write_bl_0_22 wwl_0_21 rwl_1_21
+ rwl_0_21 cell_2r1w
Xcell_2r1w_2600 vdd_uq10 gnd read_bl_0_23 read_bl_1_23 write_bl_0_23 wwl_0_23 rwl_1_23
+ rwl_0_23 cell_2r1w
Xcell_2r1w_1987 vdd_uq29 gnd read_bl_0_32 read_bl_1_32 write_bl_0_32 wwl_0_60 rwl_1_60
+ rwl_0_60 cell_2r1w
Xcell_2r1w_1998 vdd_uq23 gnd read_bl_0_32 read_bl_1_32 write_bl_0_32 wwl_0_49 rwl_1_49
+ rwl_0_49 cell_2r1w
Xcell_2r1w_1976 vdd_uq2 gnd read_bl_0_33 read_bl_1_33 write_bl_0_33 wwl_0_7 rwl_1_7
+ rwl_0_7 cell_2r1w
Xcell_2r1w_1965 vdd_uq8 gnd read_bl_0_33 read_bl_1_33 write_bl_0_33 wwl_0_18 rwl_1_18
+ rwl_0_18 cell_2r1w
Xcell_2r1w_3890 vdd_uq5 gnd read_bl_0_3 read_bl_1_3 write_bl_0_3 wwl_0_13 rwl_1_13
+ rwl_0_13 cell_2r1w
Xcell_2r1w_1217 vdd_uq30 gnd read_bl_0_44 read_bl_1_44 write_bl_0_44 wwl_0_62 rwl_1_62
+ rwl_0_62 cell_2r1w
Xcell_2r1w_1228 vdd_uq24 gnd read_bl_0_44 read_bl_1_44 write_bl_0_44 wwl_0_51 rwl_1_51
+ rwl_0_51 cell_2r1w
Xcell_2r1w_400 vdd_uq22 gnd read_bl_0_57 read_bl_1_57 write_bl_0_57 wwl_0_47 rwl_1_47
+ rwl_0_47 cell_2r1w
Xcell_2r1w_1239 vdd_uq19 gnd read_bl_0_44 read_bl_1_44 write_bl_0_44 wwl_0_40 rwl_1_40
+ rwl_0_40 cell_2r1w
Xcell_2r1w_411 vdd_uq17 gnd read_bl_0_57 read_bl_1_57 write_bl_0_57 wwl_0_36 rwl_1_36
+ rwl_0_36 cell_2r1w
Xcell_2r1w_1206 vdd_uq3 gnd read_bl_0_45 read_bl_1_45 write_bl_0_45 wwl_0_9 rwl_1_9
+ rwl_0_9 cell_2r1w
Xcell_2r1w_455 vdd_uq27 gnd read_bl_0_56 read_bl_1_56 write_bl_0_56 wwl_0_56 rwl_1_56
+ rwl_0_56 cell_2r1w
Xcell_2r1w_466 vdd_uq21 gnd read_bl_0_56 read_bl_1_56 write_bl_0_56 wwl_0_45 rwl_1_45
+ rwl_0_45 cell_2r1w
Xcell_2r1w_477 vdd_uq16 gnd read_bl_0_56 read_bl_1_56 write_bl_0_56 wwl_0_34 rwl_1_34
+ rwl_0_34 cell_2r1w
Xcell_2r1w_422 vdd_uq11 gnd read_bl_0_57 read_bl_1_57 write_bl_0_57 wwl_0_25 rwl_1_25
+ rwl_0_25 cell_2r1w
Xcell_2r1w_444 vdd gnd read_bl_0_57 read_bl_1_57 write_bl_0_57 wwl_0_3 rwl_1_3 rwl_0_3
+ cell_2r1w
Xcell_2r1w_499 vdd_uq5 gnd read_bl_0_56 read_bl_1_56 write_bl_0_56 wwl_0_12 rwl_1_12
+ rwl_0_12 cell_2r1w
Xcell_2r1w_433 vdd_uq6 gnd read_bl_0_57 read_bl_1_57 write_bl_0_57 wwl_0_14 rwl_1_14
+ rwl_0_14 cell_2r1w
Xcell_2r1w_488 vdd_uq10 gnd read_bl_0_56 read_bl_1_56 write_bl_0_56 wwl_0_23 rwl_1_23
+ rwl_0_23 cell_2r1w
Xcell_2r1w_3142 vdd_uq27 gnd read_bl_0_14 read_bl_1_14 write_bl_0_14 wwl_0_57 rwl_1_57
+ rwl_0_57 cell_2r1w
Xcell_2r1w_3131 vdd_uq1 gnd read_bl_0_15 read_bl_1_15 write_bl_0_15 wwl_0_4 rwl_1_4
+ rwl_0_4 cell_2r1w
Xcell_2r1w_3120 vdd_uq6 gnd read_bl_0_15 read_bl_1_15 write_bl_0_15 wwl_0_15 rwl_1_15
+ rwl_0_15 cell_2r1w
Xcell_2r1w_2496 vdd_uq30 gnd read_bl_0_24 read_bl_1_24 write_bl_0_24 wwl_0_63 rwl_1_63
+ rwl_0_63 cell_2r1w
Xcell_2r1w_1795 vdd_uq29 gnd read_bl_0_35 read_bl_1_35 write_bl_0_35 wwl_0_60 rwl_1_60
+ rwl_0_60 cell_2r1w
Xcell_2r1w_2441 vdd_uq26 gnd read_bl_0_25 read_bl_1_25 write_bl_0_25 wwl_0_54 rwl_1_54
+ rwl_0_54 cell_2r1w
Xcell_2r1w_1740 vdd_uq24 gnd read_bl_0_36 read_bl_1_36 write_bl_0_36 wwl_0_51 rwl_1_51
+ rwl_0_51 cell_2r1w
Xcell_2r1w_3153 vdd_uq22 gnd read_bl_0_14 read_bl_1_14 write_bl_0_14 wwl_0_46 rwl_1_46
+ rwl_0_46 cell_2r1w
Xcell_2r1w_2452 vdd_uq20 gnd read_bl_0_25 read_bl_1_25 write_bl_0_25 wwl_0_43 rwl_1_43
+ rwl_0_43 cell_2r1w
Xcell_2r1w_1751 vdd_uq19 gnd read_bl_0_36 read_bl_1_36 write_bl_0_36 wwl_0_40 rwl_1_40
+ rwl_0_40 cell_2r1w
Xcell_2r1w_3164 vdd_uq16 gnd read_bl_0_14 read_bl_1_14 write_bl_0_14 wwl_0_35 rwl_1_35
+ rwl_0_35 cell_2r1w
Xcell_2r1w_2463 vdd_uq15 gnd read_bl_0_25 read_bl_1_25 write_bl_0_25 wwl_0_32 rwl_1_32
+ rwl_0_32 cell_2r1w
Xcell_2r1w_1762 vdd_uq13 gnd read_bl_0_36 read_bl_1_36 write_bl_0_36 wwl_0_29 rwl_1_29
+ rwl_0_29 cell_2r1w
Xcell_2r1w_3175 vdd_uq11 gnd read_bl_0_14 read_bl_1_14 write_bl_0_14 wwl_0_24 rwl_1_24
+ rwl_0_24 cell_2r1w
Xcell_2r1w_3197 vdd gnd read_bl_0_14 read_bl_1_14 write_bl_0_14 wwl_0_2 rwl_1_2 rwl_0_2
+ cell_2r1w
Xcell_2r1w_2430 vdd_uq0 gnd read_bl_0_26 read_bl_1_26 write_bl_0_26 wwl_0_1 rwl_1_1
+ rwl_0_1 cell_2r1w
Xcell_2r1w_1784 vdd_uq2 gnd read_bl_0_36 read_bl_1_36 write_bl_0_36 wwl_0_7 rwl_1_7
+ rwl_0_7 cell_2r1w
Xcell_2r1w_2485 vdd_uq4 gnd read_bl_0_25 read_bl_1_25 write_bl_0_25 wwl_0_10 rwl_1_10
+ rwl_0_10 cell_2r1w
Xcell_2r1w_3186 vdd_uq5 gnd read_bl_0_14 read_bl_1_14 write_bl_0_14 wwl_0_13 rwl_1_13
+ rwl_0_13 cell_2r1w
Xcell_2r1w_1773 vdd_uq8 gnd read_bl_0_36 read_bl_1_36 write_bl_0_36 wwl_0_18 rwl_1_18
+ rwl_0_18 cell_2r1w
Xcell_2r1w_2474 vdd_uq9 gnd read_bl_0_25 read_bl_1_25 write_bl_0_25 wwl_0_21 rwl_1_21
+ rwl_0_21 cell_2r1w
Xcell_2r1w_90 vdd_uq17 gnd read_bl_0_62 read_bl_1_62 write_bl_0_62 wwl_0_37 rwl_1_37
+ rwl_0_37 cell_2r1w
Xcell_2r1w_1025 vdd_uq30 gnd read_bl_0_47 read_bl_1_47 write_bl_0_47 wwl_0_62 rwl_1_62
+ rwl_0_62 cell_2r1w
Xcell_2r1w_263 vdd_uq27 gnd read_bl_0_59 read_bl_1_59 write_bl_0_59 wwl_0_56 rwl_1_56
+ rwl_0_56 cell_2r1w
Xcell_2r1w_1036 vdd_uq24 gnd read_bl_0_47 read_bl_1_47 write_bl_0_47 wwl_0_51 rwl_1_51
+ rwl_0_51 cell_2r1w
Xcell_2r1w_1047 vdd_uq19 gnd read_bl_0_47 read_bl_1_47 write_bl_0_47 wwl_0_40 rwl_1_40
+ rwl_0_40 cell_2r1w
Xcell_2r1w_1058 vdd_uq13 gnd read_bl_0_47 read_bl_1_47 write_bl_0_47 wwl_0_29 rwl_1_29
+ rwl_0_29 cell_2r1w
Xcell_2r1w_230 vdd_uq11 gnd read_bl_0_60 read_bl_1_60 write_bl_0_60 wwl_0_25 rwl_1_25
+ rwl_0_25 cell_2r1w
Xcell_2r1w_252 vdd gnd read_bl_0_60 read_bl_1_60 write_bl_0_60 wwl_0_3 rwl_1_3 rwl_0_3
+ cell_2r1w
Xcell_2r1w_1014 vdd_uq3 gnd read_bl_0_48 read_bl_1_48 write_bl_0_48 wwl_0_9 rwl_1_9
+ rwl_0_9 cell_2r1w
Xcell_2r1w_241 vdd_uq6 gnd read_bl_0_60 read_bl_1_60 write_bl_0_60 wwl_0_14 rwl_1_14
+ rwl_0_14 cell_2r1w
Xcell_2r1w_1069 vdd_uq8 gnd read_bl_0_47 read_bl_1_47 write_bl_0_47 wwl_0_18 rwl_1_18
+ rwl_0_18 cell_2r1w
Xcell_2r1w_1003 vdd_uq9 gnd read_bl_0_48 read_bl_1_48 write_bl_0_48 wwl_0_20 rwl_1_20
+ rwl_0_20 cell_2r1w
Xcell_2r1w_274 vdd_uq21 gnd read_bl_0_59 read_bl_1_59 write_bl_0_59 wwl_0_45 rwl_1_45
+ rwl_0_45 cell_2r1w
Xcell_2r1w_285 vdd_uq16 gnd read_bl_0_59 read_bl_1_59 write_bl_0_59 wwl_0_34 rwl_1_34
+ rwl_0_34 cell_2r1w
Xcell_2r1w_296 vdd_uq10 gnd read_bl_0_59 read_bl_1_59 write_bl_0_59 wwl_0_23 rwl_1_23
+ rwl_0_23 cell_2r1w
Xcell_2r1w_2260 vdd_uq20 gnd read_bl_0_28 read_bl_1_28 write_bl_0_28 wwl_0_43 rwl_1_43
+ rwl_0_43 cell_2r1w
Xcell_2r1w_2271 vdd_uq15 gnd read_bl_0_28 read_bl_1_28 write_bl_0_28 wwl_0_32 rwl_1_32
+ rwl_0_32 cell_2r1w
Xcell_2r1w_1570 vdd_uq13 gnd read_bl_0_39 read_bl_1_39 write_bl_0_39 wwl_0_29 rwl_1_29
+ rwl_0_29 cell_2r1w
Xcell_2r1w_1592 vdd_uq2 gnd read_bl_0_39 read_bl_1_39 write_bl_0_39 wwl_0_7 rwl_1_7
+ rwl_0_7 cell_2r1w
Xcell_2r1w_2293 vdd_uq4 gnd read_bl_0_28 read_bl_1_28 write_bl_0_28 wwl_0_10 rwl_1_10
+ rwl_0_10 cell_2r1w
Xcell_2r1w_1581 vdd_uq8 gnd read_bl_0_39 read_bl_1_39 write_bl_0_39 wwl_0_18 rwl_1_18
+ rwl_0_18 cell_2r1w
Xcell_2r1w_2282 vdd_uq9 gnd read_bl_0_28 read_bl_1_28 write_bl_0_28 wwl_0_21 rwl_1_21
+ rwl_0_21 cell_2r1w
Xcell_2r1w_2090 vdd_uq9 gnd read_bl_0_31 read_bl_1_31 write_bl_0_31 wwl_0_21 rwl_1_21
+ rwl_0_21 cell_2r1w
Xcell_2r1w_3719 vdd_uq27 gnd read_bl_0_5 read_bl_1_5 write_bl_0_5 wwl_0_56 rwl_1_56
+ rwl_0_56 cell_2r1w
Xcell_2r1w_3708 vdd gnd read_bl_0_6 read_bl_1_6 write_bl_0_6 wwl_0_3 rwl_1_3 rwl_0_3
+ cell_2r1w
Xcell_2r1w_807 vdd_uq11 gnd read_bl_0_51 read_bl_1_51 write_bl_0_51 wwl_0_24 rwl_1_24
+ rwl_0_24 cell_2r1w
Xcell_2r1w_829 vdd gnd read_bl_0_51 read_bl_1_51 write_bl_0_51 wwl_0_2 rwl_1_2 rwl_0_2
+ cell_2r1w
Xcell_2r1w_818 vdd_uq5 gnd read_bl_0_51 read_bl_1_51 write_bl_0_51 wwl_0_13 rwl_1_13
+ rwl_0_13 cell_2r1w
Xcell_2r1w_3527 vdd_uq27 gnd read_bl_0_8 read_bl_1_8 write_bl_0_8 wwl_0_56 rwl_1_56
+ rwl_0_56 cell_2r1w
Xcell_2r1w_2826 vdd_uq25 gnd read_bl_0_19 read_bl_1_19 write_bl_0_19 wwl_0_53 rwl_1_53
+ rwl_0_53 cell_2r1w
Xcell_2r1w_3538 vdd_uq21 gnd read_bl_0_8 read_bl_1_8 write_bl_0_8 wwl_0_45 rwl_1_45
+ rwl_0_45 cell_2r1w
Xcell_2r1w_2837 vdd_uq20 gnd read_bl_0_19 read_bl_1_19 write_bl_0_19 wwl_0_42 rwl_1_42
+ rwl_0_42 cell_2r1w
Xcell_2r1w_3549 vdd_uq16 gnd read_bl_0_8 read_bl_1_8 write_bl_0_8 wwl_0_34 rwl_1_34
+ rwl_0_34 cell_2r1w
Xcell_2r1w_2848 vdd_uq14 gnd read_bl_0_19 read_bl_1_19 write_bl_0_19 wwl_0_31 rwl_1_31
+ rwl_0_31 cell_2r1w
Xcell_2r1w_3516 vdd gnd read_bl_0_9 read_bl_1_9 write_bl_0_9 wwl_0_3 rwl_1_3 rwl_0_3
+ cell_2r1w
Xcell_2r1w_2815 vdd_uq0 gnd read_bl_0_20 read_bl_1_20 write_bl_0_20 wwl_0_0 rwl_1_0
+ rwl_0_0 cell_2r1w
Xcell_2r1w_2804 vdd_uq4 gnd read_bl_0_20 read_bl_1_20 write_bl_0_20 wwl_0_11 rwl_1_11
+ rwl_0_11 cell_2r1w
Xcell_2r1w_3505 vdd_uq6 gnd read_bl_0_9 read_bl_1_9 write_bl_0_9 wwl_0_14 rwl_1_14
+ rwl_0_14 cell_2r1w
Xcell_2r1w_2859 vdd_uq9 gnd read_bl_0_19 read_bl_1_19 write_bl_0_19 wwl_0_20 rwl_1_20
+ rwl_0_20 cell_2r1w
Xcell_2r1w_648 vdd_uq26 gnd read_bl_0_53 read_bl_1_53 write_bl_0_53 wwl_0_55 rwl_1_55
+ rwl_0_55 cell_2r1w
Xcell_2r1w_659 vdd_uq21 gnd read_bl_0_53 read_bl_1_53 write_bl_0_53 wwl_0_44 rwl_1_44
+ rwl_0_44 cell_2r1w
Xcell_2r1w_604 vdd_uq16 gnd read_bl_0_54 read_bl_1_54 write_bl_0_54 wwl_0_35 rwl_1_35
+ rwl_0_35 cell_2r1w
Xcell_2r1w_615 vdd_uq11 gnd read_bl_0_54 read_bl_1_54 write_bl_0_54 wwl_0_24 rwl_1_24
+ rwl_0_24 cell_2r1w
Xcell_2r1w_637 vdd gnd read_bl_0_54 read_bl_1_54 write_bl_0_54 wwl_0_2 rwl_1_2 rwl_0_2
+ cell_2r1w
Xcell_2r1w_626 vdd_uq5 gnd read_bl_0_54 read_bl_1_54 write_bl_0_54 wwl_0_13 rwl_1_13
+ rwl_0_13 cell_2r1w
Xcell_2r1w_4036 vdd_uq28 gnd read_bl_0_0 read_bl_1_0 write_bl_0_0 wwl_0_59 rwl_1_59
+ rwl_0_59 cell_2r1w
Xcell_2r1w_3335 vdd_uq27 gnd read_bl_0_11 read_bl_1_11 write_bl_0_11 wwl_0_56 rwl_1_56
+ rwl_0_56 cell_2r1w
Xcell_2r1w_4047 vdd_uq23 gnd read_bl_0_0 read_bl_1_0 write_bl_0_0 wwl_0_48 rwl_1_48
+ rwl_0_48 cell_2r1w
Xcell_2r1w_4058 vdd_uq17 gnd read_bl_0_0 read_bl_1_0 write_bl_0_0 wwl_0_37 rwl_1_37
+ rwl_0_37 cell_2r1w
Xcell_2r1w_4003 vdd_uq13 gnd read_bl_0_1 read_bl_1_1 write_bl_0_1 wwl_0_28 rwl_1_28
+ rwl_0_28 cell_2r1w
Xcell_2r1w_4069 vdd_uq12 gnd read_bl_0_0 read_bl_1_0 write_bl_0_0 wwl_0_26 rwl_1_26
+ rwl_0_26 cell_2r1w
Xcell_2r1w_3302 vdd_uq11 gnd read_bl_0_12 read_bl_1_12 write_bl_0_12 wwl_0_25 rwl_1_25
+ rwl_0_25 cell_2r1w
Xcell_2r1w_3324 vdd gnd read_bl_0_12 read_bl_1_12 write_bl_0_12 wwl_0_3 rwl_1_3 rwl_0_3
+ cell_2r1w
Xcell_2r1w_4025 vdd_uq2 gnd read_bl_0_1 read_bl_1_1 write_bl_0_1 wwl_0_6 rwl_1_6 rwl_0_6
+ cell_2r1w
Xcell_2r1w_3313 vdd_uq6 gnd read_bl_0_12 read_bl_1_12 write_bl_0_12 wwl_0_14 rwl_1_14
+ rwl_0_14 cell_2r1w
Xcell_2r1w_4014 vdd_uq7 gnd read_bl_0_1 read_bl_1_1 write_bl_0_1 wwl_0_17 rwl_1_17
+ rwl_0_17 cell_2r1w
Xcell_2r1w_2689 vdd_uq30 gnd read_bl_0_21 read_bl_1_21 write_bl_0_21 wwl_0_62 rwl_1_62
+ rwl_0_62 cell_2r1w
Xcell_2r1w_1922 vdd_uq29 gnd read_bl_0_33 read_bl_1_33 write_bl_0_33 wwl_0_61 rwl_1_61
+ rwl_0_61 cell_2r1w
Xcell_2r1w_1988 vdd_uq28 gnd read_bl_0_32 read_bl_1_32 write_bl_0_32 wwl_0_59 rwl_1_59
+ rwl_0_59 cell_2r1w
Xcell_2r1w_2634 vdd_uq25 gnd read_bl_0_22 read_bl_1_22 write_bl_0_22 wwl_0_53 rwl_1_53
+ rwl_0_53 cell_2r1w
Xcell_2r1w_1933 vdd_uq24 gnd read_bl_0_33 read_bl_1_33 write_bl_0_33 wwl_0_50 rwl_1_50
+ rwl_0_50 cell_2r1w
Xcell_2r1w_3346 vdd_uq21 gnd read_bl_0_11 read_bl_1_11 write_bl_0_11 wwl_0_45 rwl_1_45
+ rwl_0_45 cell_2r1w
Xcell_2r1w_2645 vdd_uq20 gnd read_bl_0_22 read_bl_1_22 write_bl_0_22 wwl_0_42 rwl_1_42
+ rwl_0_42 cell_2r1w
Xcell_2r1w_1944 vdd_uq18 gnd read_bl_0_33 read_bl_1_33 write_bl_0_33 wwl_0_39 rwl_1_39
+ rwl_0_39 cell_2r1w
Xcell_2r1w_3357 vdd_uq16 gnd read_bl_0_11 read_bl_1_11 write_bl_0_11 wwl_0_34 rwl_1_34
+ rwl_0_34 cell_2r1w
Xcell_2r1w_2656 vdd_uq14 gnd read_bl_0_22 read_bl_1_22 write_bl_0_22 wwl_0_31 rwl_1_31
+ rwl_0_31 cell_2r1w
Xcell_2r1w_1955 vdd_uq13 gnd read_bl_0_33 read_bl_1_33 write_bl_0_33 wwl_0_28 rwl_1_28
+ rwl_0_28 cell_2r1w
Xcell_2r1w_2623 vdd_uq0 gnd read_bl_0_23 read_bl_1_23 write_bl_0_23 wwl_0_0 rwl_1_0
+ rwl_0_0 cell_2r1w
Xcell_2r1w_1977 vdd_uq2 gnd read_bl_0_33 read_bl_1_33 write_bl_0_33 wwl_0_6 rwl_1_6
+ rwl_0_6 cell_2r1w
Xcell_2r1w_1911 vdd_uq3 gnd read_bl_0_34 read_bl_1_34 write_bl_0_34 wwl_0_8 rwl_1_8
+ rwl_0_8 cell_2r1w
Xcell_2r1w_2678 vdd_uq3 gnd read_bl_0_22 read_bl_1_22 write_bl_0_22 wwl_0_9 rwl_1_9
+ rwl_0_9 cell_2r1w
Xcell_2r1w_2612 vdd_uq4 gnd read_bl_0_23 read_bl_1_23 write_bl_0_23 wwl_0_11 rwl_1_11
+ rwl_0_11 cell_2r1w
Xcell_2r1w_3379 vdd_uq5 gnd read_bl_0_11 read_bl_1_11 write_bl_0_11 wwl_0_12 rwl_1_12
+ rwl_0_12 cell_2r1w
Xcell_2r1w_1966 vdd_uq7 gnd read_bl_0_33 read_bl_1_33 write_bl_0_33 wwl_0_17 rwl_1_17
+ rwl_0_17 cell_2r1w
Xcell_2r1w_1900 vdd_uq8 gnd read_bl_0_34 read_bl_1_34 write_bl_0_34 wwl_0_19 rwl_1_19
+ rwl_0_19 cell_2r1w
Xcell_2r1w_2667 vdd_uq9 gnd read_bl_0_22 read_bl_1_22 write_bl_0_22 wwl_0_20 rwl_1_20
+ rwl_0_20 cell_2r1w
Xcell_2r1w_2601 vdd_uq10 gnd read_bl_0_23 read_bl_1_23 write_bl_0_23 wwl_0_22 rwl_1_22
+ rwl_0_22 cell_2r1w
Xcell_2r1w_3368 vdd_uq10 gnd read_bl_0_11 read_bl_1_11 write_bl_0_11 wwl_0_23 rwl_1_23
+ rwl_0_23 cell_2r1w
Xcell_2r1w_1999 vdd_uq23 gnd read_bl_0_32 read_bl_1_32 write_bl_0_32 wwl_0_48 rwl_1_48
+ rwl_0_48 cell_2r1w
Xcell_2r1w_3891 vdd_uq5 gnd read_bl_0_3 read_bl_1_3 write_bl_0_3 wwl_0_12 rwl_1_12
+ rwl_0_12 cell_2r1w
Xcell_2r1w_3880 vdd_uq10 gnd read_bl_0_3 read_bl_1_3 write_bl_0_3 wwl_0_23 rwl_1_23
+ rwl_0_23 cell_2r1w
Xcell_2r1w_1218 vdd_uq29 gnd read_bl_0_44 read_bl_1_44 write_bl_0_44 wwl_0_61 rwl_1_61
+ rwl_0_61 cell_2r1w
Xcell_2r1w_1229 vdd_uq24 gnd read_bl_0_44 read_bl_1_44 write_bl_0_44 wwl_0_50 rwl_1_50
+ rwl_0_50 cell_2r1w
Xcell_2r1w_401 vdd_uq22 gnd read_bl_0_57 read_bl_1_57 write_bl_0_57 wwl_0_46 rwl_1_46
+ rwl_0_46 cell_2r1w
Xcell_2r1w_412 vdd_uq16 gnd read_bl_0_57 read_bl_1_57 write_bl_0_57 wwl_0_35 rwl_1_35
+ rwl_0_35 cell_2r1w
Xcell_2r1w_423 vdd_uq11 gnd read_bl_0_57 read_bl_1_57 write_bl_0_57 wwl_0_24 rwl_1_24
+ rwl_0_24 cell_2r1w
Xcell_2r1w_445 vdd gnd read_bl_0_57 read_bl_1_57 write_bl_0_57 wwl_0_2 rwl_1_2 rwl_0_2
+ cell_2r1w
Xcell_2r1w_1207 vdd_uq3 gnd read_bl_0_45 read_bl_1_45 write_bl_0_45 wwl_0_8 rwl_1_8
+ rwl_0_8 cell_2r1w
Xcell_2r1w_434 vdd_uq5 gnd read_bl_0_57 read_bl_1_57 write_bl_0_57 wwl_0_13 rwl_1_13
+ rwl_0_13 cell_2r1w
Xcell_2r1w_456 vdd_uq26 gnd read_bl_0_56 read_bl_1_56 write_bl_0_56 wwl_0_55 rwl_1_55
+ rwl_0_55 cell_2r1w
Xcell_2r1w_467 vdd_uq21 gnd read_bl_0_56 read_bl_1_56 write_bl_0_56 wwl_0_44 rwl_1_44
+ rwl_0_44 cell_2r1w
Xcell_2r1w_478 vdd_uq15 gnd read_bl_0_56 read_bl_1_56 write_bl_0_56 wwl_0_33 rwl_1_33
+ rwl_0_33 cell_2r1w
Xcell_2r1w_489 vdd_uq10 gnd read_bl_0_56 read_bl_1_56 write_bl_0_56 wwl_0_22 rwl_1_22
+ rwl_0_22 cell_2r1w
Xcell_2r1w_3143 vdd_uq27 gnd read_bl_0_14 read_bl_1_14 write_bl_0_14 wwl_0_56 rwl_1_56
+ rwl_0_56 cell_2r1w
Xcell_2r1w_3154 vdd_uq21 gnd read_bl_0_14 read_bl_1_14 write_bl_0_14 wwl_0_45 rwl_1_45
+ rwl_0_45 cell_2r1w
Xcell_2r1w_3165 vdd_uq16 gnd read_bl_0_14 read_bl_1_14 write_bl_0_14 wwl_0_34 rwl_1_34
+ rwl_0_34 cell_2r1w
Xcell_2r1w_3110 vdd_uq11 gnd read_bl_0_15 read_bl_1_15 write_bl_0_15 wwl_0_25 rwl_1_25
+ rwl_0_25 cell_2r1w
Xcell_2r1w_3132 vdd gnd read_bl_0_15 read_bl_1_15 write_bl_0_15 wwl_0_3 rwl_1_3 rwl_0_3
+ cell_2r1w
Xcell_2r1w_2431 vdd_uq0 gnd read_bl_0_26 read_bl_1_26 write_bl_0_26 wwl_0_0 rwl_1_0
+ rwl_0_0 cell_2r1w
Xcell_2r1w_2420 vdd_uq4 gnd read_bl_0_26 read_bl_1_26 write_bl_0_26 wwl_0_11 rwl_1_11
+ rwl_0_11 cell_2r1w
Xcell_2r1w_3121 vdd_uq6 gnd read_bl_0_15 read_bl_1_15 write_bl_0_15 wwl_0_14 rwl_1_14
+ rwl_0_14 cell_2r1w
Xcell_2r1w_3176 vdd_uq10 gnd read_bl_0_14 read_bl_1_14 write_bl_0_14 wwl_0_23 rwl_1_23
+ rwl_0_23 cell_2r1w
Xcell_2r1w_2497 vdd_uq30 gnd read_bl_0_24 read_bl_1_24 write_bl_0_24 wwl_0_62 rwl_1_62
+ rwl_0_62 cell_2r1w
Xcell_2r1w_1730 vdd_uq29 gnd read_bl_0_36 read_bl_1_36 write_bl_0_36 wwl_0_61 rwl_1_61
+ rwl_0_61 cell_2r1w
Xcell_2r1w_1796 vdd_uq28 gnd read_bl_0_35 read_bl_1_35 write_bl_0_35 wwl_0_59 rwl_1_59
+ rwl_0_59 cell_2r1w
Xcell_2r1w_2442 vdd_uq25 gnd read_bl_0_25 read_bl_1_25 write_bl_0_25 wwl_0_53 rwl_1_53
+ rwl_0_53 cell_2r1w
Xcell_2r1w_1741 vdd_uq24 gnd read_bl_0_36 read_bl_1_36 write_bl_0_36 wwl_0_50 rwl_1_50
+ rwl_0_50 cell_2r1w
Xcell_2r1w_2453 vdd_uq20 gnd read_bl_0_25 read_bl_1_25 write_bl_0_25 wwl_0_42 rwl_1_42
+ rwl_0_42 cell_2r1w
Xcell_2r1w_1752 vdd_uq18 gnd read_bl_0_36 read_bl_1_36 write_bl_0_36 wwl_0_39 rwl_1_39
+ rwl_0_39 cell_2r1w
Xcell_2r1w_990 vdd_uq15 gnd read_bl_0_48 read_bl_1_48 write_bl_0_48 wwl_0_33 rwl_1_33
+ rwl_0_33 cell_2r1w
Xcell_2r1w_2464 vdd_uq14 gnd read_bl_0_25 read_bl_1_25 write_bl_0_25 wwl_0_31 rwl_1_31
+ rwl_0_31 cell_2r1w
Xcell_2r1w_1763 vdd_uq13 gnd read_bl_0_36 read_bl_1_36 write_bl_0_36 wwl_0_28 rwl_1_28
+ rwl_0_28 cell_2r1w
Xcell_2r1w_3198 vdd_uq0 gnd read_bl_0_14 read_bl_1_14 write_bl_0_14 wwl_0_1 rwl_1_1
+ rwl_0_1 cell_2r1w
Xcell_2r1w_1785 vdd_uq2 gnd read_bl_0_36 read_bl_1_36 write_bl_0_36 wwl_0_6 rwl_1_6
+ rwl_0_6 cell_2r1w
Xcell_2r1w_2486 vdd_uq3 gnd read_bl_0_25 read_bl_1_25 write_bl_0_25 wwl_0_9 rwl_1_9
+ rwl_0_9 cell_2r1w
Xcell_2r1w_3187 vdd_uq5 gnd read_bl_0_14 read_bl_1_14 write_bl_0_14 wwl_0_12 rwl_1_12
+ rwl_0_12 cell_2r1w
Xcell_2r1w_1774 vdd_uq7 gnd read_bl_0_36 read_bl_1_36 write_bl_0_36 wwl_0_17 rwl_1_17
+ rwl_0_17 cell_2r1w
Xcell_2r1w_2475 vdd_uq9 gnd read_bl_0_25 read_bl_1_25 write_bl_0_25 wwl_0_20 rwl_1_20
+ rwl_0_20 cell_2r1w
Xcell_2r1w_80 vdd_uq22 gnd read_bl_0_62 read_bl_1_62 write_bl_0_62 wwl_0_47 rwl_1_47
+ rwl_0_47 cell_2r1w
Xcell_2r1w_91 vdd_uq17 gnd read_bl_0_62 read_bl_1_62 write_bl_0_62 wwl_0_36 rwl_1_36
+ rwl_0_36 cell_2r1w
Xcell_2r1w_1026 vdd_uq29 gnd read_bl_0_47 read_bl_1_47 write_bl_0_47 wwl_0_61 rwl_1_61
+ rwl_0_61 cell_2r1w
Xcell_2r1w_264 vdd_uq26 gnd read_bl_0_59 read_bl_1_59 write_bl_0_59 wwl_0_55 rwl_1_55
+ rwl_0_55 cell_2r1w
Xcell_2r1w_1037 vdd_uq24 gnd read_bl_0_47 read_bl_1_47 write_bl_0_47 wwl_0_50 rwl_1_50
+ rwl_0_50 cell_2r1w
Xcell_2r1w_275 vdd_uq21 gnd read_bl_0_59 read_bl_1_59 write_bl_0_59 wwl_0_44 rwl_1_44
+ rwl_0_44 cell_2r1w
Xcell_2r1w_1048 vdd_uq18 gnd read_bl_0_47 read_bl_1_47 write_bl_0_47 wwl_0_39 rwl_1_39
+ rwl_0_39 cell_2r1w
Xcell_2r1w_220 vdd_uq16 gnd read_bl_0_60 read_bl_1_60 write_bl_0_60 wwl_0_35 rwl_1_35
+ rwl_0_35 cell_2r1w
Xcell_2r1w_286 vdd_uq15 gnd read_bl_0_59 read_bl_1_59 write_bl_0_59 wwl_0_33 rwl_1_33
+ rwl_0_33 cell_2r1w
Xcell_2r1w_1059 vdd_uq13 gnd read_bl_0_47 read_bl_1_47 write_bl_0_47 wwl_0_28 rwl_1_28
+ rwl_0_28 cell_2r1w
Xcell_2r1w_231 vdd_uq11 gnd read_bl_0_60 read_bl_1_60 write_bl_0_60 wwl_0_24 rwl_1_24
+ rwl_0_24 cell_2r1w
Xcell_2r1w_253 vdd gnd read_bl_0_60 read_bl_1_60 write_bl_0_60 wwl_0_2 rwl_1_2 rwl_0_2
+ cell_2r1w
Xcell_2r1w_1015 vdd_uq3 gnd read_bl_0_48 read_bl_1_48 write_bl_0_48 wwl_0_8 rwl_1_8
+ rwl_0_8 cell_2r1w
Xcell_2r1w_242 vdd_uq5 gnd read_bl_0_60 read_bl_1_60 write_bl_0_60 wwl_0_13 rwl_1_13
+ rwl_0_13 cell_2r1w
Xcell_2r1w_1004 vdd_uq8 gnd read_bl_0_48 read_bl_1_48 write_bl_0_48 wwl_0_19 rwl_1_19
+ rwl_0_19 cell_2r1w
Xcell_2r1w_297 vdd_uq10 gnd read_bl_0_59 read_bl_1_59 write_bl_0_59 wwl_0_22 rwl_1_22
+ rwl_0_22 cell_2r1w
Xcell_2r1w_2250 vdd_uq25 gnd read_bl_0_28 read_bl_1_28 write_bl_0_28 wwl_0_53 rwl_1_53
+ rwl_0_53 cell_2r1w
Xcell_2r1w_2261 vdd_uq20 gnd read_bl_0_28 read_bl_1_28 write_bl_0_28 wwl_0_42 rwl_1_42
+ rwl_0_42 cell_2r1w
Xcell_2r1w_2272 vdd_uq14 gnd read_bl_0_28 read_bl_1_28 write_bl_0_28 wwl_0_31 rwl_1_31
+ rwl_0_31 cell_2r1w
Xcell_2r1w_2283 vdd_uq9 gnd read_bl_0_28 read_bl_1_28 write_bl_0_28 wwl_0_20 rwl_1_20
+ rwl_0_20 cell_2r1w
Xcell_2r1w_1560 vdd_uq18 gnd read_bl_0_39 read_bl_1_39 write_bl_0_39 wwl_0_39 rwl_1_39
+ rwl_0_39 cell_2r1w
Xcell_2r1w_1571 vdd_uq13 gnd read_bl_0_39 read_bl_1_39 write_bl_0_39 wwl_0_28 rwl_1_28
+ rwl_0_28 cell_2r1w
Xcell_2r1w_1593 vdd_uq2 gnd read_bl_0_39 read_bl_1_39 write_bl_0_39 wwl_0_6 rwl_1_6
+ rwl_0_6 cell_2r1w
Xcell_2r1w_2294 vdd_uq3 gnd read_bl_0_28 read_bl_1_28 write_bl_0_28 wwl_0_9 rwl_1_9
+ rwl_0_9 cell_2r1w
Xcell_2r1w_1582 vdd_uq7 gnd read_bl_0_39 read_bl_1_39 write_bl_0_39 wwl_0_17 rwl_1_17
+ rwl_0_17 cell_2r1w
Xcell_2r1w_2080 vdd_uq14 gnd read_bl_0_31 read_bl_1_31 write_bl_0_31 wwl_0_31 rwl_1_31
+ rwl_0_31 cell_2r1w
Xcell_2r1w_1390 vdd_uq7 gnd read_bl_0_42 read_bl_1_42 write_bl_0_42 wwl_0_17 rwl_1_17
+ rwl_0_17 cell_2r1w
Xcell_2r1w_2091 vdd_uq9 gnd read_bl_0_31 read_bl_1_31 write_bl_0_31 wwl_0_20 rwl_1_20
+ rwl_0_20 cell_2r1w
Xcell_2r1w_3709 vdd gnd read_bl_0_6 read_bl_1_6 write_bl_0_6 wwl_0_2 rwl_1_2 rwl_0_2
+ cell_2r1w
Xcell_2r1w_819 vdd_uq5 gnd read_bl_0_51 read_bl_1_51 write_bl_0_51 wwl_0_12 rwl_1_12
+ rwl_0_12 cell_2r1w
Xcell_2r1w_808 vdd_uq10 gnd read_bl_0_51 read_bl_1_51 write_bl_0_51 wwl_0_23 rwl_1_23
+ rwl_0_23 cell_2r1w
Xcell_2r1w_3517 vdd gnd read_bl_0_9 read_bl_1_9 write_bl_0_9 wwl_0_2 rwl_1_2 rwl_0_2
+ cell_2r1w
Xcell_2r1w_3506 vdd_uq5 gnd read_bl_0_9 read_bl_1_9 write_bl_0_9 wwl_0_13 rwl_1_13
+ rwl_0_13 cell_2r1w
Xcell_2r1w_2816 vdd_uq30 gnd read_bl_0_19 read_bl_1_19 write_bl_0_19 wwl_0_63 rwl_1_63
+ rwl_0_63 cell_2r1w
Xcell_2r1w_3528 vdd_uq26 gnd read_bl_0_8 read_bl_1_8 write_bl_0_8 wwl_0_55 rwl_1_55
+ rwl_0_55 cell_2r1w
Xcell_2r1w_2827 vdd_uq25 gnd read_bl_0_19 read_bl_1_19 write_bl_0_19 wwl_0_52 rwl_1_52
+ rwl_0_52 cell_2r1w
Xcell_2r1w_3539 vdd_uq21 gnd read_bl_0_8 read_bl_1_8 write_bl_0_8 wwl_0_44 rwl_1_44
+ rwl_0_44 cell_2r1w
Xcell_2r1w_2838 vdd_uq19 gnd read_bl_0_19 read_bl_1_19 write_bl_0_19 wwl_0_41 rwl_1_41
+ rwl_0_41 cell_2r1w
Xcell_2r1w_2849 vdd_uq14 gnd read_bl_0_19 read_bl_1_19 write_bl_0_19 wwl_0_30 rwl_1_30
+ rwl_0_30 cell_2r1w
Xcell_2r1w_2805 vdd_uq4 gnd read_bl_0_20 read_bl_1_20 write_bl_0_20 wwl_0_10 rwl_1_10
+ rwl_0_10 cell_2r1w
Xcell_2r1w_605 vdd_uq16 gnd read_bl_0_54 read_bl_1_54 write_bl_0_54 wwl_0_34 rwl_1_34
+ rwl_0_34 cell_2r1w
Xcell_2r1w_627 vdd_uq5 gnd read_bl_0_54 read_bl_1_54 write_bl_0_54 wwl_0_12 rwl_1_12
+ rwl_0_12 cell_2r1w
Xcell_2r1w_616 vdd_uq10 gnd read_bl_0_54 read_bl_1_54 write_bl_0_54 wwl_0_23 rwl_1_23
+ rwl_0_23 cell_2r1w
Xcell_2r1w_649 vdd_uq26 gnd read_bl_0_53 read_bl_1_53 write_bl_0_53 wwl_0_54 rwl_1_54
+ rwl_0_54 cell_2r1w
Xcell_2r1w_638 vdd_uq0 gnd read_bl_0_54 read_bl_1_54 write_bl_0_54 wwl_0_1 rwl_1_1
+ rwl_0_1 cell_2r1w
Xcell_2r1w_2624 vdd_uq30 gnd read_bl_0_22 read_bl_1_22 write_bl_0_22 wwl_0_63 rwl_1_63
+ rwl_0_63 cell_2r1w
Xcell_2r1w_4037 vdd_uq28 gnd read_bl_0_0 read_bl_1_0 write_bl_0_0 wwl_0_58 rwl_1_58
+ rwl_0_58 cell_2r1w
Xcell_2r1w_3336 vdd_uq26 gnd read_bl_0_11 read_bl_1_11 write_bl_0_11 wwl_0_55 rwl_1_55
+ rwl_0_55 cell_2r1w
Xcell_2r1w_4048 vdd_uq22 gnd read_bl_0_0 read_bl_1_0 write_bl_0_0 wwl_0_47 rwl_1_47
+ rwl_0_47 cell_2r1w
Xcell_2r1w_3347 vdd_uq21 gnd read_bl_0_11 read_bl_1_11 write_bl_0_11 wwl_0_44 rwl_1_44
+ rwl_0_44 cell_2r1w
Xcell_2r1w_4059 vdd_uq17 gnd read_bl_0_0 read_bl_1_0 write_bl_0_0 wwl_0_36 rwl_1_36
+ rwl_0_36 cell_2r1w
Xcell_2r1w_3358 vdd_uq15 gnd read_bl_0_11 read_bl_1_11 write_bl_0_11 wwl_0_33 rwl_1_33
+ rwl_0_33 cell_2r1w
Xcell_2r1w_4004 vdd_uq12 gnd read_bl_0_1 read_bl_1_1 write_bl_0_1 wwl_0_27 rwl_1_27
+ rwl_0_27 cell_2r1w
Xcell_2r1w_3303 vdd_uq11 gnd read_bl_0_12 read_bl_1_12 write_bl_0_12 wwl_0_24 rwl_1_24
+ rwl_0_24 cell_2r1w
Xcell_2r1w_4026 vdd_uq1 gnd read_bl_0_1 read_bl_1_1 write_bl_0_1 wwl_0_5 rwl_1_5 rwl_0_5
+ cell_2r1w
Xcell_2r1w_3325 vdd gnd read_bl_0_12 read_bl_1_12 write_bl_0_12 wwl_0_2 rwl_1_2 rwl_0_2
+ cell_2r1w
Xcell_2r1w_2613 vdd_uq4 gnd read_bl_0_23 read_bl_1_23 write_bl_0_23 wwl_0_10 rwl_1_10
+ rwl_0_10 cell_2r1w
Xcell_2r1w_3314 vdd_uq5 gnd read_bl_0_12 read_bl_1_12 write_bl_0_12 wwl_0_13 rwl_1_13
+ rwl_0_13 cell_2r1w
Xcell_2r1w_4015 vdd_uq7 gnd read_bl_0_1 read_bl_1_1 write_bl_0_1 wwl_0_16 rwl_1_16
+ rwl_0_16 cell_2r1w
Xcell_2r1w_2602 vdd_uq9 gnd read_bl_0_23 read_bl_1_23 write_bl_0_23 wwl_0_21 rwl_1_21
+ rwl_0_21 cell_2r1w
Xcell_2r1w_3369 vdd_uq10 gnd read_bl_0_11 read_bl_1_11 write_bl_0_11 wwl_0_22 rwl_1_22
+ rwl_0_22 cell_2r1w
Xcell_2r1w_1923 vdd_uq29 gnd read_bl_0_33 read_bl_1_33 write_bl_0_33 wwl_0_60 rwl_1_60
+ rwl_0_60 cell_2r1w
Xcell_2r1w_1989 vdd_uq28 gnd read_bl_0_32 read_bl_1_32 write_bl_0_32 wwl_0_58 rwl_1_58
+ rwl_0_58 cell_2r1w
Xcell_2r1w_2635 vdd_uq25 gnd read_bl_0_22 read_bl_1_22 write_bl_0_22 wwl_0_52 rwl_1_52
+ rwl_0_52 cell_2r1w
Xcell_2r1w_1934 vdd_uq23 gnd read_bl_0_33 read_bl_1_33 write_bl_0_33 wwl_0_49 rwl_1_49
+ rwl_0_49 cell_2r1w
Xcell_2r1w_2646 vdd_uq19 gnd read_bl_0_22 read_bl_1_22 write_bl_0_22 wwl_0_41 rwl_1_41
+ rwl_0_41 cell_2r1w
Xcell_2r1w_1945 vdd_uq18 gnd read_bl_0_33 read_bl_1_33 write_bl_0_33 wwl_0_38 rwl_1_38
+ rwl_0_38 cell_2r1w
Xcell_2r1w_2657 vdd_uq14 gnd read_bl_0_22 read_bl_1_22 write_bl_0_22 wwl_0_30 rwl_1_30
+ rwl_0_30 cell_2r1w
Xcell_2r1w_1956 vdd_uq12 gnd read_bl_0_33 read_bl_1_33 write_bl_0_33 wwl_0_27 rwl_1_27
+ rwl_0_27 cell_2r1w
Xcell_2r1w_1978 vdd_uq1 gnd read_bl_0_33 read_bl_1_33 write_bl_0_33 wwl_0_5 rwl_1_5
+ rwl_0_5 cell_2r1w
Xcell_2r1w_1912 vdd_uq2 gnd read_bl_0_34 read_bl_1_34 write_bl_0_34 wwl_0_7 rwl_1_7
+ rwl_0_7 cell_2r1w
Xcell_2r1w_2679 vdd_uq3 gnd read_bl_0_22 read_bl_1_22 write_bl_0_22 wwl_0_8 rwl_1_8
+ rwl_0_8 cell_2r1w
Xcell_2r1w_1967 vdd_uq7 gnd read_bl_0_33 read_bl_1_33 write_bl_0_33 wwl_0_16 rwl_1_16
+ rwl_0_16 cell_2r1w
Xcell_2r1w_1901 vdd_uq8 gnd read_bl_0_34 read_bl_1_34 write_bl_0_34 wwl_0_18 rwl_1_18
+ rwl_0_18 cell_2r1w
Xcell_2r1w_2668 vdd_uq8 gnd read_bl_0_22 read_bl_1_22 write_bl_0_22 wwl_0_19 rwl_1_19
+ rwl_0_19 cell_2r1w
Xcell_2r1w_3870 vdd_uq15 gnd read_bl_0_3 read_bl_1_3 write_bl_0_3 wwl_0_33 rwl_1_33
+ rwl_0_33 cell_2r1w
Xcell_2r1w_3892 vdd_uq4 gnd read_bl_0_3 read_bl_1_3 write_bl_0_3 wwl_0_11 rwl_1_11
+ rwl_0_11 cell_2r1w
Xcell_2r1w_3881 vdd_uq10 gnd read_bl_0_3 read_bl_1_3 write_bl_0_3 wwl_0_22 rwl_1_22
+ rwl_0_22 cell_2r1w
Xcell_2r1w_1219 vdd_uq29 gnd read_bl_0_44 read_bl_1_44 write_bl_0_44 wwl_0_60 rwl_1_60
+ rwl_0_60 cell_2r1w
Xcell_2r1w_457 vdd_uq26 gnd read_bl_0_56 read_bl_1_56 write_bl_0_56 wwl_0_54 rwl_1_54
+ rwl_0_54 cell_2r1w
Xcell_2r1w_402 vdd_uq21 gnd read_bl_0_57 read_bl_1_57 write_bl_0_57 wwl_0_45 rwl_1_45
+ rwl_0_45 cell_2r1w
Xcell_2r1w_468 vdd_uq20 gnd read_bl_0_56 read_bl_1_56 write_bl_0_56 wwl_0_43 rwl_1_43
+ rwl_0_43 cell_2r1w
Xcell_2r1w_413 vdd_uq16 gnd read_bl_0_57 read_bl_1_57 write_bl_0_57 wwl_0_34 rwl_1_34
+ rwl_0_34 cell_2r1w
Xcell_2r1w_479 vdd_uq15 gnd read_bl_0_56 read_bl_1_56 write_bl_0_56 wwl_0_32 rwl_1_32
+ rwl_0_32 cell_2r1w
Xcell_2r1w_446 vdd_uq0 gnd read_bl_0_57 read_bl_1_57 write_bl_0_57 wwl_0_1 rwl_1_1
+ rwl_0_1 cell_2r1w
Xcell_2r1w_1208 vdd_uq2 gnd read_bl_0_45 read_bl_1_45 write_bl_0_45 wwl_0_7 rwl_1_7
+ rwl_0_7 cell_2r1w
Xcell_2r1w_435 vdd_uq5 gnd read_bl_0_57 read_bl_1_57 write_bl_0_57 wwl_0_12 rwl_1_12
+ rwl_0_12 cell_2r1w
Xcell_2r1w_424 vdd_uq10 gnd read_bl_0_57 read_bl_1_57 write_bl_0_57 wwl_0_23 rwl_1_23
+ rwl_0_23 cell_2r1w
Xcell_2r1w_2432 vdd_uq30 gnd read_bl_0_25 read_bl_1_25 write_bl_0_25 wwl_0_63 rwl_1_63
+ rwl_0_63 cell_2r1w
Xcell_2r1w_3144 vdd_uq26 gnd read_bl_0_14 read_bl_1_14 write_bl_0_14 wwl_0_55 rwl_1_55
+ rwl_0_55 cell_2r1w
Xcell_2r1w_2443 vdd_uq25 gnd read_bl_0_25 read_bl_1_25 write_bl_0_25 wwl_0_52 rwl_1_52
+ rwl_0_52 cell_2r1w
Xcell_2r1w_3155 vdd_uq21 gnd read_bl_0_14 read_bl_1_14 write_bl_0_14 wwl_0_44 rwl_1_44
+ rwl_0_44 cell_2r1w
Xcell_2r1w_2454 vdd_uq19 gnd read_bl_0_25 read_bl_1_25 write_bl_0_25 wwl_0_41 rwl_1_41
+ rwl_0_41 cell_2r1w
Xcell_2r1w_3100 vdd_uq16 gnd read_bl_0_15 read_bl_1_15 write_bl_0_15 wwl_0_35 rwl_1_35
+ rwl_0_35 cell_2r1w
Xcell_2r1w_3166 vdd_uq15 gnd read_bl_0_14 read_bl_1_14 write_bl_0_14 wwl_0_33 rwl_1_33
+ rwl_0_33 cell_2r1w
Xcell_2r1w_2465 vdd_uq14 gnd read_bl_0_25 read_bl_1_25 write_bl_0_25 wwl_0_30 rwl_1_30
+ rwl_0_30 cell_2r1w
Xcell_2r1w_3111 vdd_uq11 gnd read_bl_0_15 read_bl_1_15 write_bl_0_15 wwl_0_24 rwl_1_24
+ rwl_0_24 cell_2r1w
Xcell_2r1w_3133 vdd gnd read_bl_0_15 read_bl_1_15 write_bl_0_15 wwl_0_2 rwl_1_2 rwl_0_2
+ cell_2r1w
Xcell_2r1w_3199 vdd_uq0 gnd read_bl_0_14 read_bl_1_14 write_bl_0_14 wwl_0_0 rwl_1_0
+ rwl_0_0 cell_2r1w
Xcell_2r1w_1720 vdd_uq2 gnd read_bl_0_37 read_bl_1_37 write_bl_0_37 wwl_0_7 rwl_1_7
+ rwl_0_7 cell_2r1w
Xcell_2r1w_2421 vdd_uq4 gnd read_bl_0_26 read_bl_1_26 write_bl_0_26 wwl_0_10 rwl_1_10
+ rwl_0_10 cell_2r1w
Xcell_2r1w_3188 vdd_uq4 gnd read_bl_0_14 read_bl_1_14 write_bl_0_14 wwl_0_11 rwl_1_11
+ rwl_0_11 cell_2r1w
Xcell_2r1w_3122 vdd_uq5 gnd read_bl_0_15 read_bl_1_15 write_bl_0_15 wwl_0_13 rwl_1_13
+ rwl_0_13 cell_2r1w
Xcell_2r1w_2410 vdd_uq9 gnd read_bl_0_26 read_bl_1_26 write_bl_0_26 wwl_0_21 rwl_1_21
+ rwl_0_21 cell_2r1w
Xcell_2r1w_3177 vdd_uq10 gnd read_bl_0_14 read_bl_1_14 write_bl_0_14 wwl_0_22 rwl_1_22
+ rwl_0_22 cell_2r1w
Xcell_2r1w_2498 vdd_uq29 gnd read_bl_0_24 read_bl_1_24 write_bl_0_24 wwl_0_61 rwl_1_61
+ rwl_0_61 cell_2r1w
Xcell_2r1w_1731 vdd_uq29 gnd read_bl_0_36 read_bl_1_36 write_bl_0_36 wwl_0_60 rwl_1_60
+ rwl_0_60 cell_2r1w
Xcell_2r1w_1797 vdd_uq28 gnd read_bl_0_35 read_bl_1_35 write_bl_0_35 wwl_0_58 rwl_1_58
+ rwl_0_58 cell_2r1w
Xcell_2r1w_1742 vdd_uq23 gnd read_bl_0_36 read_bl_1_36 write_bl_0_36 wwl_0_49 rwl_1_49
+ rwl_0_49 cell_2r1w
Xcell_2r1w_980 vdd_uq20 gnd read_bl_0_48 read_bl_1_48 write_bl_0_48 wwl_0_43 rwl_1_43
+ rwl_0_43 cell_2r1w
Xcell_2r1w_1753 vdd_uq18 gnd read_bl_0_36 read_bl_1_36 write_bl_0_36 wwl_0_38 rwl_1_38
+ rwl_0_38 cell_2r1w
Xcell_2r1w_991 vdd_uq15 gnd read_bl_0_48 read_bl_1_48 write_bl_0_48 wwl_0_32 rwl_1_32
+ rwl_0_32 cell_2r1w
Xcell_2r1w_1764 vdd_uq12 gnd read_bl_0_36 read_bl_1_36 write_bl_0_36 wwl_0_27 rwl_1_27
+ rwl_0_27 cell_2r1w
Xcell_2r1w_1786 vdd_uq1 gnd read_bl_0_36 read_bl_1_36 write_bl_0_36 wwl_0_5 rwl_1_5
+ rwl_0_5 cell_2r1w
Xcell_2r1w_2487 vdd_uq3 gnd read_bl_0_25 read_bl_1_25 write_bl_0_25 wwl_0_8 rwl_1_8
+ rwl_0_8 cell_2r1w
Xcell_2r1w_1775 vdd_uq7 gnd read_bl_0_36 read_bl_1_36 write_bl_0_36 wwl_0_16 rwl_1_16
+ rwl_0_16 cell_2r1w
Xcell_2r1w_2476 vdd_uq8 gnd read_bl_0_25 read_bl_1_25 write_bl_0_25 wwl_0_19 rwl_1_19
+ rwl_0_19 cell_2r1w
Xcell_2r1w_70 vdd_uq27 gnd read_bl_0_62 read_bl_1_62 write_bl_0_62 wwl_0_57 rwl_1_57
+ rwl_0_57 cell_2r1w
Xcell_2r1w_81 vdd_uq22 gnd read_bl_0_62 read_bl_1_62 write_bl_0_62 wwl_0_46 rwl_1_46
+ rwl_0_46 cell_2r1w
Xcell_2r1w_92 vdd_uq16 gnd read_bl_0_62 read_bl_1_62 write_bl_0_62 wwl_0_35 rwl_1_35
+ rwl_0_35 cell_2r1w
Xcell_2r1w_1016 vdd_uq2 gnd read_bl_0_48 read_bl_1_48 write_bl_0_48 wwl_0_7 rwl_1_7
+ rwl_0_7 cell_2r1w
Xcell_2r1w_1005 vdd_uq8 gnd read_bl_0_48 read_bl_1_48 write_bl_0_48 wwl_0_18 rwl_1_18
+ rwl_0_18 cell_2r1w
Xcell_2r1w_1027 vdd_uq29 gnd read_bl_0_47 read_bl_1_47 write_bl_0_47 wwl_0_60 rwl_1_60
+ rwl_0_60 cell_2r1w
Xcell_2r1w_265 vdd_uq26 gnd read_bl_0_59 read_bl_1_59 write_bl_0_59 wwl_0_54 rwl_1_54
+ rwl_0_54 cell_2r1w
Xcell_2r1w_1038 vdd_uq23 gnd read_bl_0_47 read_bl_1_47 write_bl_0_47 wwl_0_49 rwl_1_49
+ rwl_0_49 cell_2r1w
Xcell_2r1w_210 vdd_uq21 gnd read_bl_0_60 read_bl_1_60 write_bl_0_60 wwl_0_45 rwl_1_45
+ rwl_0_45 cell_2r1w
Xcell_2r1w_276 vdd_uq20 gnd read_bl_0_59 read_bl_1_59 write_bl_0_59 wwl_0_43 rwl_1_43
+ rwl_0_43 cell_2r1w
Xcell_2r1w_1049 vdd_uq18 gnd read_bl_0_47 read_bl_1_47 write_bl_0_47 wwl_0_38 rwl_1_38
+ rwl_0_38 cell_2r1w
Xcell_2r1w_221 vdd_uq16 gnd read_bl_0_60 read_bl_1_60 write_bl_0_60 wwl_0_34 rwl_1_34
+ rwl_0_34 cell_2r1w
Xcell_2r1w_287 vdd_uq15 gnd read_bl_0_59 read_bl_1_59 write_bl_0_59 wwl_0_32 rwl_1_32
+ rwl_0_32 cell_2r1w
Xcell_2r1w_254 vdd_uq0 gnd read_bl_0_60 read_bl_1_60 write_bl_0_60 wwl_0_1 rwl_1_1
+ rwl_0_1 cell_2r1w
Xcell_2r1w_243 vdd_uq5 gnd read_bl_0_60 read_bl_1_60 write_bl_0_60 wwl_0_12 rwl_1_12
+ rwl_0_12 cell_2r1w
Xcell_2r1w_298 vdd_uq9 gnd read_bl_0_59 read_bl_1_59 write_bl_0_59 wwl_0_21 rwl_1_21
+ rwl_0_21 cell_2r1w
Xcell_2r1w_232 vdd_uq10 gnd read_bl_0_60 read_bl_1_60 write_bl_0_60 wwl_0_23 rwl_1_23
+ rwl_0_23 cell_2r1w
Xcell_2r1w_2240 vdd_uq30 gnd read_bl_0_28 read_bl_1_28 write_bl_0_28 wwl_0_63 rwl_1_63
+ rwl_0_63 cell_2r1w
Xcell_2r1w_2251 vdd_uq25 gnd read_bl_0_28 read_bl_1_28 write_bl_0_28 wwl_0_52 rwl_1_52
+ rwl_0_52 cell_2r1w
Xcell_2r1w_1550 vdd_uq23 gnd read_bl_0_39 read_bl_1_39 write_bl_0_39 wwl_0_49 rwl_1_49
+ rwl_0_49 cell_2r1w
Xcell_2r1w_2262 vdd_uq19 gnd read_bl_0_28 read_bl_1_28 write_bl_0_28 wwl_0_41 rwl_1_41
+ rwl_0_41 cell_2r1w
Xcell_2r1w_1561 vdd_uq18 gnd read_bl_0_39 read_bl_1_39 write_bl_0_39 wwl_0_38 rwl_1_38
+ rwl_0_38 cell_2r1w
Xcell_2r1w_2273 vdd_uq14 gnd read_bl_0_28 read_bl_1_28 write_bl_0_28 wwl_0_30 rwl_1_30
+ rwl_0_30 cell_2r1w
Xcell_2r1w_1572 vdd_uq12 gnd read_bl_0_39 read_bl_1_39 write_bl_0_39 wwl_0_27 rwl_1_27
+ rwl_0_27 cell_2r1w
Xcell_2r1w_2295 vdd_uq3 gnd read_bl_0_28 read_bl_1_28 write_bl_0_28 wwl_0_8 rwl_1_8
+ rwl_0_8 cell_2r1w
Xcell_2r1w_2284 vdd_uq8 gnd read_bl_0_28 read_bl_1_28 write_bl_0_28 wwl_0_19 rwl_1_19
+ rwl_0_19 cell_2r1w
Xcell_2r1w_1594 vdd_uq1 gnd read_bl_0_39 read_bl_1_39 write_bl_0_39 wwl_0_5 rwl_1_5
+ rwl_0_5 cell_2r1w
Xcell_2r1w_1583 vdd_uq7 gnd read_bl_0_39 read_bl_1_39 write_bl_0_39 wwl_0_16 rwl_1_16
+ rwl_0_16 cell_2r1w
Xcell_2r1w_2070 vdd_uq19 gnd read_bl_0_31 read_bl_1_31 write_bl_0_31 wwl_0_41 rwl_1_41
+ rwl_0_41 cell_2r1w
Xcell_2r1w_2081 vdd_uq14 gnd read_bl_0_31 read_bl_1_31 write_bl_0_31 wwl_0_30 rwl_1_30
+ rwl_0_30 cell_2r1w
Xcell_2r1w_1380 vdd_uq12 gnd read_bl_0_42 read_bl_1_42 write_bl_0_42 wwl_0_27 rwl_1_27
+ rwl_0_27 cell_2r1w
Xcell_2r1w_1391 vdd_uq7 gnd read_bl_0_42 read_bl_1_42 write_bl_0_42 wwl_0_16 rwl_1_16
+ rwl_0_16 cell_2r1w
Xcell_2r1w_2092 vdd_uq8 gnd read_bl_0_31 read_bl_1_31 write_bl_0_31 wwl_0_19 rwl_1_19
+ rwl_0_19 cell_2r1w
Xcell_2r1w_809 vdd_uq10 gnd read_bl_0_51 read_bl_1_51 write_bl_0_51 wwl_0_22 rwl_1_22
+ rwl_0_22 cell_2r1w
Xcell_2r1w_3529 vdd_uq26 gnd read_bl_0_8 read_bl_1_8 write_bl_0_8 wwl_0_54 rwl_1_54
+ rwl_0_54 cell_2r1w
Xcell_2r1w_3518 vdd_uq0 gnd read_bl_0_9 read_bl_1_9 write_bl_0_9 wwl_0_1 rwl_1_1 rwl_0_1
+ cell_2r1w
Xcell_2r1w_2806 vdd_uq3 gnd read_bl_0_20 read_bl_1_20 write_bl_0_20 wwl_0_9 rwl_1_9
+ rwl_0_9 cell_2r1w
Xcell_2r1w_3507 vdd_uq5 gnd read_bl_0_9 read_bl_1_9 write_bl_0_9 wwl_0_12 rwl_1_12
+ rwl_0_12 cell_2r1w
Xcell_2r1w_2817 vdd_uq30 gnd read_bl_0_19 read_bl_1_19 write_bl_0_19 wwl_0_62 rwl_1_62
+ rwl_0_62 cell_2r1w
Xcell_2r1w_2828 vdd_uq24 gnd read_bl_0_19 read_bl_1_19 write_bl_0_19 wwl_0_51 rwl_1_51
+ rwl_0_51 cell_2r1w
Xcell_2r1w_2839 vdd_uq19 gnd read_bl_0_19 read_bl_1_19 write_bl_0_19 wwl_0_40 rwl_1_40
+ rwl_0_40 cell_2r1w
Xcell_2r1w_606 vdd_uq15 gnd read_bl_0_54 read_bl_1_54 write_bl_0_54 wwl_0_33 rwl_1_33
+ rwl_0_33 cell_2r1w
Xcell_2r1w_639 vdd_uq0 gnd read_bl_0_54 read_bl_1_54 write_bl_0_54 wwl_0_0 rwl_1_0
+ rwl_0_0 cell_2r1w
Xcell_2r1w_628 vdd_uq4 gnd read_bl_0_54 read_bl_1_54 write_bl_0_54 wwl_0_11 rwl_1_11
+ rwl_0_11 cell_2r1w
Xcell_2r1w_617 vdd_uq10 gnd read_bl_0_54 read_bl_1_54 write_bl_0_54 wwl_0_22 rwl_1_22
+ rwl_0_22 cell_2r1w
Xcell_2r1w_2625 vdd_uq30 gnd read_bl_0_22 read_bl_1_22 write_bl_0_22 wwl_0_62 rwl_1_62
+ rwl_0_62 cell_2r1w
Xcell_2r1w_4038 vdd_uq27 gnd read_bl_0_0 read_bl_1_0 write_bl_0_0 wwl_0_57 rwl_1_57
+ rwl_0_57 cell_2r1w
Xcell_2r1w_3337 vdd_uq26 gnd read_bl_0_11 read_bl_1_11 write_bl_0_11 wwl_0_54 rwl_1_54
+ rwl_0_54 cell_2r1w
Xcell_2r1w_2636 vdd_uq24 gnd read_bl_0_22 read_bl_1_22 write_bl_0_22 wwl_0_51 rwl_1_51
+ rwl_0_51 cell_2r1w
Xcell_2r1w_4049 vdd_uq22 gnd read_bl_0_0 read_bl_1_0 write_bl_0_0 wwl_0_46 rwl_1_46
+ rwl_0_46 cell_2r1w
Xcell_2r1w_3348 vdd_uq20 gnd read_bl_0_11 read_bl_1_11 write_bl_0_11 wwl_0_43 rwl_1_43
+ rwl_0_43 cell_2r1w
Xcell_2r1w_2647 vdd_uq19 gnd read_bl_0_22 read_bl_1_22 write_bl_0_22 wwl_0_40 rwl_1_40
+ rwl_0_40 cell_2r1w
Xcell_2r1w_3359 vdd_uq15 gnd read_bl_0_11 read_bl_1_11 write_bl_0_11 wwl_0_32 rwl_1_32
+ rwl_0_32 cell_2r1w
Xcell_2r1w_4005 vdd_uq12 gnd read_bl_0_1 read_bl_1_1 write_bl_0_1 wwl_0_26 rwl_1_26
+ rwl_0_26 cell_2r1w
Xcell_2r1w_4027 vdd_uq1 gnd read_bl_0_1 read_bl_1_1 write_bl_0_1 wwl_0_4 rwl_1_4 rwl_0_4
+ cell_2r1w
Xcell_2r1w_3326 vdd_uq0 gnd read_bl_0_12 read_bl_1_12 write_bl_0_12 wwl_0_1 rwl_1_1
+ rwl_0_1 cell_2r1w
Xcell_2r1w_1913 vdd_uq2 gnd read_bl_0_34 read_bl_1_34 write_bl_0_34 wwl_0_6 rwl_1_6
+ rwl_0_6 cell_2r1w
Xcell_2r1w_2614 vdd_uq3 gnd read_bl_0_23 read_bl_1_23 write_bl_0_23 wwl_0_9 rwl_1_9
+ rwl_0_9 cell_2r1w
Xcell_2r1w_3315 vdd_uq5 gnd read_bl_0_12 read_bl_1_12 write_bl_0_12 wwl_0_12 rwl_1_12
+ rwl_0_12 cell_2r1w
Xcell_2r1w_4016 vdd_uq6 gnd read_bl_0_1 read_bl_1_1 write_bl_0_1 wwl_0_15 rwl_1_15
+ rwl_0_15 cell_2r1w
Xcell_2r1w_1902 vdd_uq7 gnd read_bl_0_34 read_bl_1_34 write_bl_0_34 wwl_0_17 rwl_1_17
+ rwl_0_17 cell_2r1w
Xcell_2r1w_2603 vdd_uq9 gnd read_bl_0_23 read_bl_1_23 write_bl_0_23 wwl_0_20 rwl_1_20
+ rwl_0_20 cell_2r1w
Xcell_2r1w_3304 vdd_uq10 gnd read_bl_0_12 read_bl_1_12 write_bl_0_12 wwl_0_23 rwl_1_23
+ rwl_0_23 cell_2r1w
.ends

.subckt replica_bitcell_array rwl_1_28 rwl_0_61 rwl_0_38 wwl_0_40 wwl_0_51 wwl_0_62
+ rwl_0_5 rwl_1_61 rwl_1_38 wwl_0_30 wwl_0_41 wwl_0_52 wwl_0_63 rwl_0_48 rwl_1_5 rwl_0_15
+ wwl_0_20 wwl_0_31 wwl_0_42 wwl_0_53 rwl_1_48 rwl_0_58 rwl_1_15 wwl_0_10 wwl_0_21
+ wwl_0_32 wwl_0_43 wwl_0_54 rwl_0_25 rwl_0_2 rwl_1_58 wwl_0_11 wwl_0_22 wwl_0_33
+ wwl_0_44 wwl_0_55 rwl_1_25 rwl_1_2 rwl_0_35 rwl_0_12 wwl_0_12 wwl_0_23 wwl_0_34
+ wwl_0_45 wwl_0_56 rwl_1_35 rwl_1_12 rwl_0_45 rwl_0_22 wwl_0_13 wwl_0_24 wwl_0_35
+ wwl_0_46 wwl_0_57 wwl_0_0 rwl_1_45 rwl_1_22 wwl_0_14 wwl_0_25 wwl_0_36 wwl_0_47
+ wwl_0_58 rwl_0_55 rwl_0_32 rwl_0_9 wwl_0_15 wwl_0_26 wwl_0_37 rwl_1_55 wwl_0_48
+ wwl_0_59 rwl_1_32 rwl_1_9 rwl_0_42 rwl_0_19 wwl_0_16 wwl_0_27 wwl_0_38 wwl_0_49
+ rwl_1_42 rwl_1_19 rwl_0_52 rwl_0_29 rwl_0_6 wwl_0_17 wwl_0_28 wwl_0_39 rwl_1_52
+ rwl_1_29 rwl_1_6 rwl_0_62 wwl_0_18 wwl_0_29 rwl_0_39 rwl_0_16 rwl_1_62 wwl_0_19
+ rwl_1_39 rwl_1_16 rwl_0_49 rwl_0_26 rwl_1_49 rwl_1_26 rwl_0_59 rwl_0_36 rwl_0_3
+ rwl_1_59 rwl_1_36 rwl_0_46 rwl_1_3 rwl_0_13 rwl_1_46 rwl_0_56 rwl_1_13 rwl_0_23
+ rwl_0_0 wwl_0_1 rwl_1_56 rwl_1_23 rwl_1_0 rwl_0_33 rwl_0_10 rwl_1_33 rwl_1_10 rwl_0_43
+ rwl_0_20 rwl_1_43 rwl_1_20 rwl_0_53 rwl_0_30 rwl_0_7 rwl_1_53 rwl_1_30 rwl_1_7 rwl_0_63
+ rwl_0_40 rwl_0_17 rwl_1_63 rwl_1_40 rwl_1_17 rwl_0_50 rwl_0_27 gnd rwl_1_50 rwl_1_27
+ rwl_0_60 rwl_0_37 rwl_0_4 rwl_1_60 rwl_1_37 rwl_0_47 rwl_1_4 rwl_0_14 rwl_1_47 rwl_0_57
+ rwl_1_14 rwl_0_24 rwl_0_1 wwl_0_2 rwl_1_57 rwl_1_24 rwl_1_1 rwl_0_34 wwl_0_3 rwl_0_11
+ rwl_1_34 wwl_0_4 rwl_1_11 rwl_0_44 rwl_0_21 wwl_0_5 rwl_1_44 rwl_1_21 rwl_0_54 rwl_0_31
+ rwl_0_8 wwl_0_6 rwl_1_54 rwl_1_31 rwl_1_8 rwl_0_41 wwl_0_7 rwl_0_18 wwl_0_60 rwl_1_41
+ wwl_0_8 rwl_1_18 rwl_0_51 rwl_0_28 wwl_0_50 wwl_0_61 wwl_0_9 rwl_1_51
Xbitcell_array_0 write_bl_0_56 wwl_0_1 read_bl_1_29 read_bl_0_0 rwl_0_0 write_bl_0_44
+ read_bl_0_24 wwl_0_57 rwl_0_47 write_bl_0_53 wwl_0_43 read_bl_0_51 read_bl_1_26
+ read_bl_0_22 write_bl_0_5 wwl_0_35 read_bl_0_39 read_bl_0_2 read_bl_0_48 wwl_0_56
+ wwl_0_37 write_bl_0_3 read_bl_0_37 write_bl_0_20 rwl_1_12 read_bl_0_60 rwl_0_11
+ wwl_0_20 write_bl_0_15 read_bl_0_31 write_bl_0_32 read_bl_0_58 write_bl_0_61 read_bl_0_63
+ read_bl_0_47 rwl_0_24 write_bl_0_12 read_bl_1_21 write_bl_0_30 read_bl_0_29 read_bl_0_10
+ write_bl_0_37 rwl_0_2 read_bl_1_19 read_bl_1_36 read_bl_0_7 write_bl_0_34 read_bl_1_34
+ read_bl_1_57 rwl_1_43 rwl_1_5 wwl_0_42 rwl_0_46 read_bl_1_28 rwl_1_35 write_bl_0_0
+ read_bl_1_55 rwl_1_21 read_bl_0_41 rwl_1_47 read_bl_1_44 read_bl_1_7 wwl_0_55 read_bl_0_50
+ rwl_1_13 write_bl_0_22 write_bl_0_42 read_bl_0_20 rwl_1_15 rwl_1_60 write_bl_0_49
+ wwl_0_33 read_bl_1_4 rwl_0_3 rwl_0_40 read_bl_0_17 rwl_1_57 read_bl_0_12 write_bl_0_58
+ write_bl_0_63 read_bl_1_14 rwl_0_1 read_bl_0_46 read_bl_0_27 read_bl_0_9 read_bl_0_34
+ read_bl_0_25 read_bl_1_30 rwl_0_45 rwl_1_20 read_bl_1_46 rwl_1_46 rwl_0_23 read_bl_1_9
+ rwl_1_24 rwl_1_59 write_bl_0_51 wwl_0_6 wwl_0_32 read_bl_1_6 write_bl_0_39 write_bl_0_2
+ read_bl_0_19 rwl_1_37 write_bl_0_48 rwl_1_56 wwl_0_10 read_bl_1_16 wwl_0_50 rwl_1_34
+ wwl_0_28 read_bl_1_49 wwl_0_54 rwl_1_39 write_bl_0_47 read_bl_1_38 write_bl_0_10
+ wwl_0_3 rwl_0_58 write_bl_0_7 read_bl_1_48 rwl_0_22 wwl_0_5 read_bl_1_56 wwl_0_47
+ read_bl_1_45 rwl_1_58 read_bl_1_8 read_bl_1_54 write_bl_0_41 rwl_1_10 read_bl_0_21
+ rwl_1_36 rwl_0_9 write_bl_0_50 read_bl_0_36 rwl_1_33 wwl_0_40 wwl_0_62 wwl_0_51
+ wwl_0_41 write_bl_0_60 wwl_0_27 read_bl_1_40 rwl_1_32 wwl_0_19 read_bl_0_55 rwl_1_16
+ write_bl_0_46 rwl_0_57 rwl_0_31 read_bl_1_18 read_bl_0_26 write_bl_0_9 read_bl_0_44
+ read_bl_0_53 rwl_0_6 read_bl_0_4 rwl_1_9 read_bl_1_47 wwl_0_24 read_bl_1_25 rwl_0_50
+ write_bl_0_52 read_bl_0_14 rwl_0_34 read_bl_0_42 read_bl_1_52 read_bl_1_23 rwl_0_28
+ write_bl_0_19 read_bl_1_50 rwl_1_19 read_bl_1_62 wwl_0_18 write_bl_0_17 wwl_0_4
+ rwl_0_30 rwl_0_56 write_bl_0_29 read_bl_0_28 write_bl_0_11 read_bl_1_59 write_bl_0_57
+ rwl_0_8 wwl_0_17 write_bl_0_62 write_bl_0_27 read_bl_0_6 wwl_0_59 rwl_1_50 read_bl_0_16
+ rwl_0_44 rwl_0_27 read_bl_0_49 write_bl_0_21 read_bl_0_38 read_bl_1_3 read_bl_1_61
+ rwl_0_21 read_bl_0_57 rwl_0_7 read_bl_0_45 wwl_0_16 read_bl_0_8 write_bl_0_55 read_bl_1_11
+ wwl_0_58 read_bl_0_54 write_bl_0_26 rwl_0_20 rwl_0_62 read_bl_1_33 write_bl_0_4
+ rwl_0_43 wwl_0_26 rwl_1_27 write_bl_0_16 read_bl_1_42 rwl_0_4 write_bl_0_14 write_bl_0_38
+ read_bl_1_51 wwl_0_46 read_bl_0_35 write_bl_0_36 write_bl_0_31 read_bl_1_13 write_bl_0_28
+ rwl_0_19 rwl_1_62 read_bl_0_52 wwl_0_9 read_bl_1_35 rwl_0_61 write_bl_0_43 write_bl_0_6
+ read_bl_0_23 wwl_0_48 read_bl_0_62 read_bl_1_1 wwl_0_45 rwl_1_42 read_bl_0_59 read_bl_1_5
+ rwl_0_49 read_bl_0_18 rwl_1_55 read_bl_1_20 read_bl_1_32 read_bl_1_15 rwl_0_60 read_bl_1_12
+ write_bl_0_45 write_bl_0_8 wwl_0_21 rwl_0_38 rwl_0_12 write_bl_0_24 read_bl_0_3
+ read_bl_0_1 read_bl_0_61 wwl_0_22 read_bl_0_13 rwl_0_48 rwl_1_54 read_bl_0_11 write_bl_0_35
+ read_bl_0_33 rwl_0_37 wwl_0_49 read_bl_1_10 rwl_1_25 write_bl_0_23 read_bl_0_40
+ read_bl_1_0 rwl_0_33 rwl_1_0 read_bl_1_24 rwl_0_25 rwl_1_31 read_bl_1_22 read_bl_1_39
+ write_bl_0_18 read_bl_1_37 read_bl_1_60 write_bl_0_33 rwl_1_49 read_bl_1_31 wwl_0_61
+ rwl_1_41 rwl_1_53 read_bl_1_63 read_bl_1_58 rwl_0_52 write_bl_0_54 write_bl_0_25
+ read_bl_0_5 rwl_1_2 rwl_1_4 write_bl_0_1 read_bl_0_15 wwl_0_7 rwl_0_10 read_bl_1_41
+ read_bl_0_30 write_bl_0_59 read_bl_1_17 rwl_1_40 rwl_1_26 wwl_0_38 rwl_1_18 read_bl_1_27
+ rwl_1_1 rwl_1_45 rwl_1_23 wwl_0_31 write_bl_0_13 rwl_0_35 read_bl_1_2 rwl_0_13 rwl_1_3
+ wwl_0_53 rwl_1_22 read_bl_0_32 wwl_0_8 read_bl_0_56 wwl_0_30 wwl_0_63 wwl_0_52 read_bl_1_53
+ read_bl_0_43 rwl_0_55 rwl_1_30 rwl_1_8 write_bl_0_40 rwl_1_44 wwl_0_13 rwl_0_32
+ rwl_1_7 wwl_0_29 wwl_0_15 rwl_0_41 rwl_0_16 wwl_0_34 wwl_0_14 rwl_0_18 rwl_0_54
+ wwl_0_11 rwl_1_6 rwl_0_17 rwl_0_53 rwl_0_14 rwl_1_52 rwl_0_59 rwl_0_5 rwl_1_51 rwl_1_63
+ rwl_1_29 rwl_1_28 rwl_1_14 rwl_1_11 wwl_0_23 rwl_0_42 rwl_1_17 read_bl_1_43 wwl_0_39
+ wwl_0_25 rwl_0_51 rwl_0_29 wwl_0_0 rwl_0_26 wwl_0_2 wwl_0_44 rwl_0_63 rwl_1_61 rwl_1_38
+ wwl_0_36 rwl_0_39 rwl_0_36 wwl_0_12 rwl_0_15 rwl_1_48 wwl_0_60 gnd bitcell_array
.ends

.subckt bank addr2 vdd_uq243 vdd_uq232 vdd_uq221 vdd_uq210 gnd dout1_19 wl_en vdd_uq233
+ vdd_uq211 vdd_uq175 addr3 vdd_uq121 vdd_uq244 vdd_uq222 vdd_uq200 dout1_30 vdd_uq235
+ vdd_uq213 vdd_uq179 addr4 vdd_uq234 vdd_uq223 vdd_uq212 vdd_uq201 dout1_20 dout1_31
+ vdd_uq237 vdd_uq215 vdd_uq183 p_en_bar addr5 vdd_uq224 vdd_uq203 vdd_uq89 vdd vdd_uq71
+ dout1_10 dout1_21 vdd_uq239 vdd_uq217 vdd_uq187 addr6 vdd_uq236 vdd_uq225 vdd_uq214
+ dout1_11 dout1_22 vdd_uq241 vdd_uq219 vdd_uq189 addr7 vdd_uq226 vdd_uq204 dout1_12
+ dout1_23 vdd_uq193 addr8 vdd_uq238 vdd_uq227 vdd_uq216 vdd_uq205 dout1_13 dout1_24
+ vdd_uq197 vdd_uq228 vdd_uq206 dout1_14 dout1_25 vdd_uq161 vdd_uq229 vdd_uq218 vdd_uq207
+ dout1_15 dout1_26 dout1_0 vdd_uq208 dout1_16 dout1_27 dout1_1 vdd_uq209 dout1_17
+ dout1_28 dout1_2 dout1_18 dout1_29 vdd_uq191 dout1_3 vdd_uq181 dout1_4 vdd_uq192
+ vdd_uq170 dout1_5 vdd_uq160 vdd_uq171 vdd_uq182 dout1_6 vdd_uq195 vdd_uq150 vdd_uq173
+ dout1_7 vdd_uq240 w_en vdd_uq91 vdd_uq140 vdd_uq151 vdd_uq163 vdd_uq185 dout1_8
+ vdd_uq196 vdd_uq81 vdd_uq130 vdd_uq141 vdd_uq152 vdd_uq174 dout1_9 vdd_uq93 vdd_uq131
+ vdd_uq142 vdd_uq153 vdd_uq164 vdd_uq186 vdd_uq83 vdd_uq111 vdd_uq132 vdd_uq143 vdd_uq154
+ vdd_uq199 vdd_uq165 vdd_uq177 vdd_uq188 vdd_uq73 vdd_uq95 vdd_uq101 vdd_uq123 vdd_uq133
+ vdd_uq144 vdd_uq155 vdd_uq167 vdd_uq85 vdd_uq113 vdd_uq134 vdd_uq145 vdd_uq156 vdd_uq178
+ vdd_uq75 vdd_uq97 vdd_uq103 vdd_uq125 vdd_uq135 vdd_uq146 vdd_uq157 vdd_uq168 addr1
+ vdd_uq65 vdd_uq87 vdd_uq115 vdd_uq136 vdd_uq147 vdd_uq158 vdd_uq169 vdd_uq77 vdd_uq99
+ vdd_uq105 vdd_uq127 vdd_uq137 vdd_uq148 vdd_uq159 vdd_uq67 vdd_uq117 vdd_uq138 vdd_uq149
+ vdd_uq79 vdd_uq107 vdd_uq128 vdd_uq139 vdd_uq69 vdd_uq119 vdd_uq129 vdd_uq109 vdd_uq230
+ vdd_uq242 vdd_uq231 vdd_uq220
Xport_data_0 din0_15 din0_26 dout1_19 din0_6 din0_16 din0_27 p_en_bar din0_7 dout1_30
+ din0_17 din0_28 gnd pinvbuf_0/Z din0_8 dout1_20 dout1_31 din0_18 din0_29 din0_9
+ vdd dout1_10 dout1_21 din0_19 dout1_11 dout1_22 dout1_12 dout1_23 dout1_13 dout1_24
+ w_en dout1_14 dout1_25 dout1_15 dout1_26 dout1_0 dout1_16 dout1_27 dout1_1 dout1_17
+ dout1_28 dout1_2 dout1_18 dout1_29 dout1_3 dout1_4 dout1_5 dout1_6 vdd_uq150 dout1_7
+ vdd_uq91 vdd_uq140 vdd_uq151 dout1_8 vdd_uq81 vdd_uq130 vdd_uq141 vdd_uq152 dout1_9
+ vdd_uq71 vdd_uq93 vdd_uq121 vdd_uq131 vdd_uq142 vdd_uq153 vdd_uq83 vdd_uq111 vdd_uq132
+ vdd_uq143 vdd_uq154 vdd_uq73 vdd_uq95 vdd_uq101 vdd_uq123 vdd_uq133 vdd_uq144 vdd_uq155
+ vdd_uq85 vdd_uq113 vdd_uq134 vdd_uq145 vdd_uq156 vdd_uq125 vdd_uq75 vdd_uq97 vdd_uq103
+ vdd_uq135 vdd_uq146 vdd_uq157 p_en_bar vdd_uq65 vdd_uq87 vdd_uq115 vdd_uq136 vdd_uq147
+ vdd_uq158 vdd_uq77 vdd_uq99 vdd_uq105 vdd_uq127 vdd_uq137 vdd_uq148 vdd_uq159 din0_21
+ vdd_uq67 vdd_uq89 vdd_uq117 vdd_uq138 vdd_uq149 vdd_uq107 vdd_uq79 vdd_uq128 vdd_uq139
+ pinvbuf_0/Z vdd_uq69 vdd_uq119 vdd_uq129 vdd_uq109 din0_30 din0_20 din0_31 din0_0
+ din0_10 din0_1 din0_11 din0_22 din0_2 din0_12 din0_23 din0_3 din0_13 din0_24 din0_4
+ din0_14 din0_25 din0_5 port_data
Xpinvbuf_0 pinvbuf_0/Z pinvbuf_0/Z pinvbuf_0/Z gnd vdd_uq244 addr0 pinvbuf
Xport_address_0 addr3 wl_en port_address_0/wwl0_0 port_address_0/rwl1_0 port_address_0/rwl1_55
+ port_address_0/rwl1_44 port_address_0/rwl1_11 port_address_0/rwl1_22 port_address_0/rwl1_33
+ addr4 gnd port_address_0/rwl1_1 port_address_0/wwl0_1 vdd_uq160 port_address_0/rwl1_56
+ port_address_0/rwl1_45 port_address_0/rwl1_34 port_address_0/rwl1_12 port_address_0/rwl1_23
+ addr5 vdd_uq243 port_address_0/rwl1_2 port_address_0/wwl0_2 vdd_uq163 port_address_0/rwl1_13
+ port_address_0/rwl1_24 port_address_0/rwl1_57 port_address_0/rwl1_46 port_address_0/rwl1_35
+ addr6 vdd_uq223 port_address_0/rwl1_3 port_address_0/wwl0_3 port_address_0/rwl1_58
+ port_address_0/rwl1_47 port_address_0/rwl1_36 port_address_0/rwl1_14 port_address_0/rwl1_25
+ addr7 vdd_uq225 vdd_uq201 port_address_0/wwl0_4 port_address_0/rwl1_4 vdd_uq164
+ port_address_0/rwl1_59 port_address_0/rwl1_48 port_address_0/rwl1_37 port_address_0/rwl1_15
+ port_address_0/rwl1_26 addr8 vdd_uq227 vdd_uq205 vdd_uq165 port_address_0/rwl1_5
+ port_address_0/wwl0_5 port_address_0/rwl1_49 port_address_0/rwl1_38 port_address_0/rwl1_16
+ port_address_0/rwl1_27 vdd_uq229 vdd_uq207 vdd_uq169 port_address_0/rwl1_6 port_address_0/wwl0_6
+ vdd_uq167 port_address_0/rwl1_39 port_address_0/rwl1_17 port_address_0/rwl1_28 vdd_uq231
+ vdd_uq209 vdd_uq171 port_address_0/rwl1_7 port_address_0/wwl0_7 port_address_0/rwl1_18
+ port_address_0/rwl1_29 vdd_uq233 vdd_uq211 vdd_uq175 port_address_0/rwl1_8 port_address_0/wwl0_8
+ vdd_uq168 port_address_0/rwl1_19 vdd_uq235 vdd_uq213 vdd_uq179 port_address_0/rwl1_9
+ port_address_0/wwl0_9 vdd_uq237 vdd_uq215 vdd_uq183 vdd_uq170 vdd_uq239 vdd_uq217
+ vdd_uq187 port_address_0/wwl0_60 vdd_uq241 vdd_uq219 vdd_uq189 port_address_0/wwl0_61
+ port_address_0/wwl0_50 vdd_uq221 vdd_uq193 port_address_0/wwl0_62 port_address_0/wwl0_51
+ port_address_0/wwl0_40 vdd_uq197 port_address_0/wwl0_63 port_address_0/wwl0_52 port_address_0/wwl0_41
+ port_address_0/wwl0_30 vdd_uq161 port_address_0/wwl0_53 port_address_0/wwl0_42 port_address_0/wwl0_20
+ port_address_0/wwl0_31 addr1 port_address_0/wwl0_54 port_address_0/wwl0_43 port_address_0/wwl0_10
+ port_address_0/wwl0_21 port_address_0/wwl0_32 addr2 port_address_0/wwl0_55 port_address_0/wwl0_44
+ port_address_0/wwl0_33 port_address_0/wwl0_11 port_address_0/wwl0_22 port_address_0/wwl0_60
+ vdd_uq242 port_address_0/wwl0_56 port_address_0/wwl0_45 port_address_0/wwl0_34 port_address_0/wwl0_12
+ port_address_0/wwl0_23 port_address_0/wwl0_61 port_address_0/rwl0_50 vdd_uq232 port_address_0/rwl0_0
+ port_address_0/wwl0_57 port_address_0/wwl0_46 port_address_0/wwl0_35 port_address_0/wwl0_13
+ port_address_0/wwl0_24 vdd_uq240 port_address_0/rwl0_40 port_address_0/wwl0_62 port_address_0/wwl0_51
+ vdd_uq222 port_address_0/rwl0_1 port_address_0/wwl0_58 port_address_0/wwl0_47 port_address_0/wwl0_36
+ port_address_0/wwl0_14 port_address_0/wwl0_25 port_address_0/wwl0_63 port_address_0/rwl0_52
+ port_address_0/rwl0_41 port_address_0/rwl0_30 vdd_uq212 vdd_uq234 port_address_0/rwl0_2
+ port_address_0/wwl0_59 port_address_0/wwl0_48 port_address_0/wwl0_37 port_address_0/wwl0_15
+ port_address_0/wwl0_26 port_address_0/wwl0_53 port_address_0/rwl0_42 port_address_0/rwl0_20
+ port_address_0/rwl0_31 vdd_uq203 vdd_uq191 vdd_uq224 port_address_0/rwl0_3 port_address_0/wwl0_49
+ port_address_0/wwl0_38 port_address_0/wwl0_16 port_address_0/wwl0_27 port_address_0/wwl0_54
+ port_address_0/rwl0_43 port_address_0/rwl0_10 port_address_0/rwl0_21 port_address_0/rwl0_32
+ vdd_uq192 vdd_uq181 vdd_uq214 vdd_uq236 port_address_0/rwl0_4 port_address_0/wwl0_39
+ port_address_0/wwl0_17 port_address_0/wwl0_28 port_address_0/wwl0_55 port_address_0/rwl0_44
+ port_address_0/rwl0_33 port_address_0/rwl0_11 port_address_0/rwl0_22 vdd_uq182 vdd_uq204
+ vdd_uq226 port_address_0/rwl0_5 port_address_0/wwl0_18 port_address_0/wwl0_29 port_address_0/wwl0_56
+ port_address_0/wwl0_45 port_address_0/rwl0_34 port_address_0/rwl0_12 port_address_0/rwl0_23
+ vdd_uq173 vdd_uq195 vdd_uq216 vdd_uq238 port_address_0/rwl0_6 port_address_0/wwl0_19
+ port_address_0/wwl0_57 port_address_0/rwl0_46 port_address_0/rwl0_35 port_address_0/rwl0_13
+ port_address_0/rwl0_24 vdd_uq185 vdd_uq206 vdd_uq228 port_address_0/rwl0_7 port_address_0/wwl0_58
+ port_address_0/wwl0_47 port_address_0/rwl0_36 port_address_0/rwl0_14 port_address_0/rwl0_25
+ vdd_uq196 vdd_uq174 vdd_uq218 port_address_0/rwl0_8 port_address_0/wwl0_59 port_address_0/rwl0_48
+ port_address_0/rwl0_37 port_address_0/rwl0_15 port_address_0/rwl0_26 vdd_uq186 vdd_uq208
+ vdd_uq230 port_address_0/rwl0_9 port_address_0/wwl0_49 port_address_0/rwl0_38 port_address_0/rwl0_16
+ port_address_0/rwl0_27 vdd_uq199 vdd_uq177 vdd_uq220 port_address_0/rwl0_39 port_address_0/rwl0_17
+ port_address_0/rwl0_28 port_address_0/rwl1_60 vdd_uq188 vdd_uq210 port_address_0/rwl0_18
+ port_address_0/rwl0_29 port_address_0/rwl1_61 port_address_0/rwl1_50 vdd_uq200 vdd_uq178
+ port_address_0/rwl0_19 port_address_0/rwl1_62 port_address_0/rwl1_51 port_address_0/rwl1_40
+ port_address_0/rwl1_63 port_address_0/rwl1_52 port_address_0/rwl1_41 port_address_0/rwl1_30
+ port_address_0/rwl1_53 port_address_0/rwl1_42 port_address_0/rwl1_20 port_address_0/rwl1_31
+ port_address_0/rwl1_54 port_address_0/rwl1_43 port_address_0/rwl1_10 port_address_0/rwl1_21
+ port_address_0/rwl1_32 port_address
Xreplica_bitcell_array_0 port_address_0/rwl1_28 port_address_0/wwl0_61 port_address_0/rwl0_38
+ port_address_0/wwl0_40 port_address_0/wwl0_51 port_address_0/wwl0_62 port_address_0/rwl0_5
+ port_address_0/rwl1_61 port_address_0/rwl1_38 port_address_0/wwl0_30 port_address_0/wwl0_41
+ port_address_0/wwl0_52 port_address_0/wwl0_63 port_address_0/rwl0_48 port_address_0/rwl1_5
+ port_address_0/rwl0_15 port_address_0/wwl0_20 port_address_0/wwl0_31 port_address_0/wwl0_42
+ port_address_0/wwl0_53 port_address_0/rwl1_48 port_address_0/wwl0_58 port_address_0/rwl1_15
+ port_address_0/wwl0_10 port_address_0/wwl0_21 port_address_0/wwl0_32 port_address_0/wwl0_43
+ port_address_0/wwl0_54 port_address_0/rwl0_25 port_address_0/rwl0_2 port_address_0/rwl1_58
+ port_address_0/wwl0_11 port_address_0/wwl0_22 port_address_0/wwl0_33 port_address_0/wwl0_44
+ port_address_0/wwl0_55 port_address_0/rwl1_25 port_address_0/rwl1_2 port_address_0/rwl0_35
+ port_address_0/rwl0_12 port_address_0/wwl0_12 port_address_0/wwl0_23 port_address_0/wwl0_34
+ port_address_0/wwl0_45 port_address_0/wwl0_56 port_address_0/rwl1_35 port_address_0/rwl1_12
+ port_address_0/wwl0_45 port_address_0/rwl0_22 port_address_0/wwl0_13 port_address_0/wwl0_24
+ port_address_0/wwl0_35 port_address_0/wwl0_46 port_address_0/wwl0_57 port_address_0/wwl0_0
+ port_address_0/rwl1_45 port_address_0/rwl1_22 port_address_0/wwl0_14 port_address_0/wwl0_25
+ port_address_0/wwl0_36 port_address_0/wwl0_47 port_address_0/wwl0_58 port_address_0/wwl0_55
+ port_address_0/rwl0_32 port_address_0/rwl0_9 port_address_0/wwl0_15 port_address_0/wwl0_26
+ port_address_0/wwl0_37 port_address_0/rwl1_55 port_address_0/wwl0_48 port_address_0/wwl0_59
+ port_address_0/rwl1_32 port_address_0/rwl1_9 port_address_0/rwl0_42 port_address_0/rwl0_19
+ port_address_0/wwl0_16 port_address_0/wwl0_27 port_address_0/wwl0_38 port_address_0/wwl0_49
+ port_address_0/rwl1_42 port_address_0/rwl1_19 port_address_0/rwl0_52 port_address_0/rwl0_29
+ port_address_0/rwl0_6 port_address_0/wwl0_17 port_address_0/wwl0_28 port_address_0/wwl0_39
+ port_address_0/rwl1_52 port_address_0/rwl1_29 port_address_0/rwl1_6 port_address_0/wwl0_62
+ port_address_0/wwl0_18 port_address_0/wwl0_29 port_address_0/rwl0_39 port_address_0/rwl0_16
+ port_address_0/rwl1_62 port_address_0/wwl0_19 port_address_0/rwl1_39 port_address_0/rwl1_16
+ port_address_0/wwl0_49 port_address_0/rwl0_26 port_address_0/rwl1_49 port_address_0/rwl1_26
+ port_address_0/wwl0_59 port_address_0/rwl0_36 port_address_0/rwl0_3 port_address_0/rwl1_59
+ port_address_0/rwl1_36 port_address_0/rwl0_46 port_address_0/rwl1_3 port_address_0/rwl0_13
+ port_address_0/rwl1_46 port_address_0/wwl0_56 port_address_0/rwl1_13 port_address_0/rwl0_23
+ port_address_0/rwl0_0 port_address_0/wwl0_1 port_address_0/rwl1_56 port_address_0/rwl1_23
+ port_address_0/rwl1_0 port_address_0/rwl0_33 port_address_0/rwl0_10 port_address_0/rwl1_33
+ port_address_0/rwl1_10 port_address_0/rwl0_43 port_address_0/rwl0_20 port_address_0/rwl1_43
+ port_address_0/rwl1_20 port_address_0/wwl0_53 port_address_0/rwl0_30 port_address_0/rwl0_7
+ port_address_0/rwl1_53 port_address_0/rwl1_30 port_address_0/rwl1_7 port_address_0/wwl0_63
+ port_address_0/rwl0_40 port_address_0/rwl0_17 port_address_0/rwl1_63 port_address_0/rwl1_40
+ port_address_0/rwl1_17 port_address_0/rwl0_50 port_address_0/rwl0_27 gnd port_address_0/rwl1_50
+ port_address_0/rwl1_27 port_address_0/wwl0_60 port_address_0/rwl0_37 port_address_0/rwl0_4
+ port_address_0/rwl1_60 port_address_0/rwl1_37 port_address_0/wwl0_47 port_address_0/rwl1_4
+ port_address_0/rwl0_14 port_address_0/rwl1_47 port_address_0/wwl0_57 port_address_0/rwl1_14
+ port_address_0/rwl0_24 port_address_0/rwl0_1 port_address_0/wwl0_2 port_address_0/rwl1_57
+ port_address_0/rwl1_24 port_address_0/rwl1_1 port_address_0/rwl0_34 port_address_0/wwl0_3
+ port_address_0/rwl0_11 port_address_0/rwl1_34 port_address_0/wwl0_4 port_address_0/rwl1_11
+ port_address_0/rwl0_44 port_address_0/rwl0_21 port_address_0/wwl0_5 port_address_0/rwl1_44
+ port_address_0/rwl1_21 port_address_0/wwl0_54 port_address_0/rwl0_31 port_address_0/rwl0_8
+ port_address_0/wwl0_6 port_address_0/rwl1_54 port_address_0/rwl1_31 port_address_0/rwl1_8
+ port_address_0/rwl0_41 port_address_0/wwl0_7 port_address_0/rwl0_18 port_address_0/wwl0_60
+ port_address_0/rwl1_41 port_address_0/wwl0_8 port_address_0/rwl1_18 port_address_0/wwl0_51
+ port_address_0/rwl0_28 port_address_0/wwl0_50 port_address_0/wwl0_61 port_address_0/wwl0_9
+ port_address_0/rwl1_51 replica_bitcell_array
.ends

.subckt sram_0rw2r1w_32_128_sky130A
Xcontrol_logic_multiport_0 vdd clk web vdd csb vdd vdd control_logic_multiport
Xdata_dff_0 vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd
+ vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd data_dff
Xcol_addr_dff_0 vdd vdd vdd vdd col_addr_dff
Xrow_addr_dff_0 addr1[8] vdd vdd vdd vdd vdd bank_0/addr1 bank_0/addr2 bank_0/addr4
+ bank_0/addr3 vdd bank_0/addr5 bank_0/addr6 bank_0/addr7 bank_0/addr8 vdd vdd addr1[2]
+ addr1[3] addr1[4] addr1[5] addr1[6] addr1[7] row_addr_dff
Xbank_0 bank_0/addr2 vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd bank_0/addr3 vdd vdd
+ vdd vdd vdd vdd vdd vdd bank_0/addr4 vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd bank_0/addr5
+ vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd bank_0/addr6 vdd vdd vdd vdd vdd vdd vdd
+ vdd bank_0/addr7 vdd vdd vdd vdd vdd bank_0/addr8 vdd vdd vdd vdd vdd vdd vdd vdd
+ vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd
+ vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd
+ vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd
+ vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd
+ vdd vdd vdd vdd vdd vdd vdd bank_0/addr1 vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd
+ vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd
+ bank
.ends

