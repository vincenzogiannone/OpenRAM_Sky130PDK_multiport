magic
tech sky130A
timestamp 1644951705
<< checkpaint >>
rect -630 -630 631 631
<< properties >>
string GDS_FILE sram_0rw2r1w_16_128_sky130A.gds
string GDS_END 1452188
string GDS_START 1451736
<< end >>
