magic
tech sky130A
magscale 1 2
timestamp 1643593061
<< checkpaint >>
rect -1260 -1260 14784 29884
<< metal1 >>
rect 6547 27848 6688 27876
rect 6547 27836 6575 27848
rect 6398 27808 6575 27836
rect 6547 27722 6688 27750
rect 6547 27710 6575 27722
rect 6398 27682 6575 27710
rect 6547 27496 6688 27524
rect 6547 27484 6575 27496
rect 6398 27456 6575 27484
rect 6547 26444 6688 26464
rect 6398 26436 6688 26444
rect 6398 26416 6575 26436
rect 6547 26218 6688 26238
rect 6398 26210 6688 26218
rect 6398 26190 6575 26210
rect 6547 26092 6688 26112
rect 6398 26084 6688 26092
rect 6398 26064 6575 26084
rect 6547 24768 6688 24796
rect 6547 24760 6575 24768
rect 6398 24732 6575 24760
rect 6547 24642 6688 24670
rect 6547 24634 6575 24642
rect 6398 24606 6575 24634
rect 6547 24416 6688 24444
rect 6547 24408 6575 24416
rect 6398 24380 6575 24408
rect 6547 23368 6688 23384
rect 6398 23356 6688 23368
rect 6398 23340 6575 23356
rect 6547 23142 6688 23158
rect 6398 23130 6688 23142
rect 6398 23114 6575 23130
rect 6547 23016 6688 23032
rect 6398 23004 6688 23016
rect 6398 22988 6575 23004
rect 6547 21688 6688 21716
rect 6547 21684 6575 21688
rect 6398 21656 6575 21684
rect 6547 21562 6688 21590
rect 6547 21558 6575 21562
rect 6398 21530 6575 21558
rect 6547 21336 6688 21364
rect 6547 21332 6575 21336
rect 6398 21304 6575 21332
rect 6547 20292 6688 20304
rect 6398 20276 6688 20292
rect 6398 20264 6575 20276
rect 6547 20066 6688 20078
rect 6398 20050 6688 20066
rect 6398 20038 6575 20050
rect 6547 19940 6688 19952
rect 6398 19924 6688 19940
rect 6398 19912 6575 19924
rect 6547 18608 6688 18636
rect 6398 18580 6575 18608
rect 6547 18482 6688 18510
rect 6398 18454 6575 18482
rect 6547 18256 6688 18284
rect 6398 18228 6575 18256
rect 6547 17216 6688 17224
rect 6398 17196 6688 17216
rect 6398 17188 6575 17196
rect 6547 16990 6688 16998
rect 6398 16970 6688 16990
rect 6398 16962 6575 16970
rect 6547 16864 6688 16872
rect 6398 16844 6688 16864
rect 6398 16836 6575 16844
rect 6547 15532 6688 15556
rect 6398 15528 6688 15532
rect 6398 15504 6575 15528
rect 6547 15406 6688 15430
rect 6398 15402 6688 15406
rect 6398 15378 6575 15402
rect 6547 15180 6688 15204
rect 6398 15176 6688 15180
rect 6398 15152 6575 15176
rect 6547 14140 6688 14144
rect 6398 14116 6688 14140
rect 6398 14112 6575 14116
rect 6547 13914 6688 13918
rect 6398 13890 6688 13914
rect 6398 13886 6575 13890
rect 6547 13788 6688 13792
rect 6398 13764 6688 13788
rect 6398 13760 6575 13764
rect 6547 12456 6688 12476
rect 6398 12448 6688 12456
rect 6398 12428 6575 12448
rect 6547 12330 6688 12350
rect 6398 12322 6688 12330
rect 6398 12302 6575 12322
rect 6547 12104 6688 12124
rect 6398 12096 6688 12104
rect 6398 12076 6575 12096
rect 6398 11036 6688 11064
rect 6398 10810 6688 10838
rect 6398 10684 6688 10712
rect 6547 9380 6688 9396
rect 6398 9368 6688 9380
rect 6398 9352 6575 9368
rect 6547 9254 6688 9270
rect 6398 9242 6688 9254
rect 6398 9226 6575 9242
rect 6547 9028 6688 9044
rect 6398 9016 6688 9028
rect 6398 9000 6575 9016
rect 6398 7984 6575 7988
rect 6398 7960 6688 7984
rect 6547 7956 6688 7960
rect 6398 7758 6575 7762
rect 6398 7734 6688 7758
rect 6547 7730 6688 7734
rect 6398 7632 6575 7636
rect 6398 7608 6688 7632
rect 6547 7604 6688 7608
rect 6547 6304 6688 6316
rect 6398 6288 6688 6304
rect 6398 6276 6575 6288
rect 6547 6178 6688 6190
rect 6398 6162 6688 6178
rect 6398 6150 6575 6162
rect 6547 5952 6688 5964
rect 6398 5936 6688 5952
rect 6398 5924 6575 5936
rect 6398 4904 6575 4912
rect 6398 4884 6688 4904
rect 6547 4876 6688 4884
rect 6398 4678 6575 4686
rect 6398 4658 6688 4678
rect 6547 4650 6688 4658
rect 6398 4552 6575 4560
rect 6398 4532 6688 4552
rect 6547 4524 6688 4532
rect 6310 3400 6316 3452
rect 6368 3440 6374 3452
rect 6368 3412 7426 3440
rect 6368 3400 6374 3412
rect 8526 1279 8532 1291
rect 7855 1251 8532 1279
rect 8526 1239 8532 1251
rect 8584 1239 8590 1291
<< via1 >>
rect 6316 3400 6368 3452
rect 8532 1239 8584 1291
<< metal2 >>
rect 18 3880 46 28512
rect 102 3880 130 28512
rect 186 3880 214 28512
rect 270 3880 298 28512
rect 354 3880 382 28512
rect 438 3880 466 28512
rect 5194 28474 5222 28502
rect 6328 3452 6356 3796
rect 6884 3496 6938 3524
rect 7662 3496 7716 3524
rect 6328 0 6356 3400
rect 8544 1291 8572 28624
rect 11438 2352 11466 2592
rect 11898 2352 11926 2592
rect 8544 0 8572 1239
<< metal3 >>
rect 828 28482 888 28542
rect 1700 28482 1760 28542
rect 6368 28458 6428 28518
rect 5164 28074 5224 28134
rect 828 26942 888 27002
rect 1700 26942 1760 27002
rect 6368 26920 6428 26980
rect 5164 26560 5224 26620
rect 828 25402 888 25462
rect 1700 25402 1760 25462
rect 6368 25382 6428 25442
rect 5164 25046 5224 25106
rect 828 23862 888 23922
rect 1700 23862 1760 23922
rect 6368 23844 6428 23904
rect 5164 23532 5224 23592
rect 828 22322 888 22382
rect 1700 22322 1760 22382
rect 6368 22306 6428 22366
rect 5164 22018 5224 22078
rect 6368 20768 6428 20828
rect 5164 20504 5224 20564
rect 828 19246 888 19306
rect 1700 19246 1760 19306
rect 6368 19230 6428 19290
rect 5164 18990 5224 19050
rect 828 17706 888 17766
rect 1700 17706 1760 17766
rect 6368 17692 6428 17752
rect 5164 17476 5224 17536
rect 828 16166 888 16226
rect 1700 16166 1760 16226
rect 6368 16154 6428 16214
rect 5164 15962 5224 16022
rect 828 14626 888 14686
rect 1700 14626 1760 14686
rect 6368 14616 6428 14676
rect 5164 14448 5224 14508
rect 828 13086 888 13146
rect 1700 13086 1760 13146
rect 6368 13078 6428 13138
rect 5164 12934 5224 12994
rect 6368 11540 6428 11600
rect 5164 11420 5224 11480
rect 828 10010 888 10070
rect 1700 10010 1760 10070
rect 6368 10002 6428 10062
rect 5164 9906 5224 9966
rect 828 8470 888 8530
rect 1700 8470 1760 8530
rect 6368 8464 6428 8524
rect 5164 8392 5224 8452
rect 828 6930 888 6990
rect 1700 6930 1760 6990
rect 5164 6878 5224 6938
rect 6368 6926 6428 6986
rect 828 5390 888 5450
rect 1700 5390 1760 5450
rect 5164 5364 5224 5424
rect 6368 5388 6428 5448
rect 828 3850 888 3910
rect 1700 3850 1760 3910
rect 5164 3850 5224 3910
rect 6368 3850 6428 3910
rect 7007 3724 7067 3784
rect 7785 3724 7845 3784
rect 7007 2892 7067 2952
rect 7785 2892 7845 2952
rect 11342 2528 11402 2588
rect 11802 2528 11862 2588
rect 12898 2528 12958 2588
rect 13358 2528 13418 2588
rect 11342 1582 11402 1642
rect 11802 1582 11862 1642
rect 12898 1582 12958 1642
rect 13358 1582 13418 1642
rect 6851 332 6911 392
rect 7629 332 7689 392
rect 8407 332 8467 392
use contact_17  contact_17_0
timestamp 1643593061
transform 1 0 8526 0 1 1239
box 0 0 1 1
use contact_17  contact_17_1
timestamp 1643593061
transform 1 0 6310 0 1 3400
box 0 0 1 1
use port_address  port_address_0
timestamp 1643593061
transform 1 0 0 0 1 3880
box 0 -42 6430 24662
use port_data  port_data_0
timestamp 1643593061
transform 1 0 6688 0 1 0
box 0 238 6836 3796
use replica_bitcell_array  replica_bitcell_array_0
timestamp 1643593061
transform 1 0 6688 0 1 3880
box 0 -42 1556 24682
<< labels >>
rlabel metal2 s 6328 0 6356 3796 4 w_en
rlabel metal2 s 5194 28474 5222 28502 4 wl_en
rlabel metal2 s 8544 0 8572 28624 4 p_en_bar
rlabel metal2 s 6884 3496 6938 3524 4 din0_0
rlabel metal2 s 7662 3496 7716 3524 4 din0_1
rlabel metal2 s 11438 2352 11466 2592 4 dout0_0
rlabel metal2 s 11452 2472 11452 2472 4 dout1_0
rlabel metal2 s 11898 2352 11926 2592 4 dout0_1
rlabel metal2 s 11912 2472 11912 2472 4 dout1_1
rlabel metal2 s 18 3880 46 28512 4 addr0
rlabel metal2 s 102 3880 130 28512 4 addr1
rlabel metal2 s 186 3880 214 28512 4 addr2
rlabel metal2 s 270 3880 298 28512 4 addr3
rlabel metal2 s 354 3880 382 28512 4 addr4
rlabel metal2 s 438 3880 466 28512 4 addr5
rlabel metal3 s 6368 11540 6428 11600 4 vdd
rlabel metal3 s 13358 1582 13418 1642 4 vdd
rlabel metal3 s 11342 1582 11402 1642 4 vdd
rlabel metal3 s 828 26942 888 27002 4 vdd
rlabel metal3 s 6368 20768 6428 20828 4 vdd
rlabel metal3 s 11802 1582 11862 1642 4 vdd
rlabel metal3 s 1700 8470 1760 8530 4 vdd
rlabel metal3 s 6368 17692 6428 17752 4 vdd
rlabel metal3 s 828 23862 888 23922 4 vdd
rlabel metal3 s 7006 2892 7066 2952 4 vdd
rlabel metal3 s 828 5390 888 5450 4 vdd
rlabel metal3 s 6368 26920 6428 26980 4 vdd
rlabel metal3 s 12898 1582 12958 1642 4 vdd
rlabel metal3 s 5164 23532 5224 23592 4 vdd
rlabel metal3 s 5164 5364 5224 5424 4 vdd
rlabel metal3 s 6368 8464 6428 8524 4 vdd
rlabel metal3 s 5164 8392 5224 8452 4 vdd
rlabel metal3 s 8406 332 8466 392 4 vdd
rlabel metal3 s 1700 23862 1760 23922 4 vdd
rlabel metal3 s 5164 26560 5224 26620 4 vdd
rlabel metal3 s 5164 14448 5224 14508 4 vdd
rlabel metal3 s 1700 5390 1760 5450 4 vdd
rlabel metal3 s 5164 17476 5224 17536 4 vdd
rlabel metal3 s 1700 14626 1760 14686 4 vdd
rlabel metal3 s 1700 17706 1760 17766 4 vdd
rlabel metal3 s 5164 20504 5224 20564 4 vdd
rlabel metal3 s 5164 11420 5224 11480 4 vdd
rlabel metal3 s 828 14626 888 14686 4 vdd
rlabel metal3 s 6368 14616 6428 14676 4 vdd
rlabel metal3 s 6368 23844 6428 23904 4 vdd
rlabel metal3 s 828 17706 888 17766 4 vdd
rlabel metal3 s 1700 26942 1760 27002 4 vdd
rlabel metal3 s 6850 332 6910 392 4 vdd
rlabel metal3 s 7628 332 7688 392 4 vdd
rlabel metal3 s 7784 2892 7844 2952 4 vdd
rlabel metal3 s 6368 5388 6428 5448 4 vdd
rlabel metal3 s 828 8470 888 8530 4 vdd
rlabel metal3 s 11802 2528 11862 2588 4 gnd
rlabel metal3 s 6368 22306 6428 22366 4 gnd
rlabel metal3 s 1700 22322 1760 22382 4 gnd
rlabel metal3 s 6368 13078 6428 13138 4 gnd
rlabel metal3 s 1700 6930 1760 6990 4 gnd
rlabel metal3 s 5164 3850 5224 3910 4 gnd
rlabel metal3 s 1700 28482 1760 28542 4 gnd
rlabel metal3 s 6368 10002 6428 10062 4 gnd
rlabel metal3 s 5164 9906 5224 9966 4 gnd
rlabel metal3 s 6368 16154 6428 16214 4 gnd
rlabel metal3 s 828 25402 888 25462 4 gnd
rlabel metal3 s 828 3850 888 3910 4 gnd
rlabel metal3 s 6368 19230 6428 19290 4 gnd
rlabel metal3 s 1700 19246 1760 19306 4 gnd
rlabel metal3 s 6368 28458 6428 28518 4 gnd
rlabel metal3 s 5164 25046 5224 25106 4 gnd
rlabel metal3 s 5164 15962 5224 16022 4 gnd
rlabel metal3 s 6368 25382 6428 25442 4 gnd
rlabel metal3 s 828 22322 888 22382 4 gnd
rlabel metal3 s 828 28482 888 28542 4 gnd
rlabel metal3 s 828 10010 888 10070 4 gnd
rlabel metal3 s 828 13086 888 13146 4 gnd
rlabel metal3 s 7006 3724 7066 3784 4 gnd
rlabel metal3 s 5164 12934 5224 12994 4 gnd
rlabel metal3 s 5164 6878 5224 6938 4 gnd
rlabel metal3 s 6368 3850 6428 3910 4 gnd
rlabel metal3 s 828 19246 888 19306 4 gnd
rlabel metal3 s 11342 2528 11402 2588 4 gnd
rlabel metal3 s 828 16166 888 16226 4 gnd
rlabel metal3 s 1700 13086 1760 13146 4 gnd
rlabel metal3 s 5164 22018 5224 22078 4 gnd
rlabel metal3 s 5164 28074 5224 28134 4 gnd
rlabel metal3 s 6368 6926 6428 6986 4 gnd
rlabel metal3 s 13358 2528 13418 2588 4 gnd
rlabel metal3 s 7784 3724 7844 3784 4 gnd
rlabel metal3 s 1700 3850 1760 3910 4 gnd
rlabel metal3 s 1700 25402 1760 25462 4 gnd
rlabel metal3 s 5164 18990 5224 19050 4 gnd
rlabel metal3 s 12898 2528 12958 2588 4 gnd
rlabel metal3 s 1700 16166 1760 16226 4 gnd
rlabel metal3 s 1700 10010 1760 10070 4 gnd
rlabel metal3 s 828 6930 888 6990 4 gnd
<< properties >>
string FIXED_BBOX 0 0 13608 28624
string GDS_FILE sram_0rw2r1w_2_16_sky130A.gds
string GDS_END 181528
string GDS_START 148748
<< end >>
