magic
tech sky130A
magscale 1 2
timestamp 1643678851
<< checkpaint >>
rect -1296 -1277 9558 2155
<< nwell >>
rect -36 402 8298 895
<< locali >>
rect 0 821 8262 855
rect 48 344 114 410
rect 196 360 432 394
rect 547 360 783 394
rect 902 360 1242 394
rect 1558 354 2025 388
rect 2775 352 3780 386
rect 5934 352 5968 386
rect 0 -17 8262 17
use pinv_10  pinv_10_0
timestamp 1643678851
transform 1 0 3699 0 1 0
box -36 -17 4599 895
use pinv_9  pinv_9_0
timestamp 1643678851
transform 1 0 1944 0 1 0
box -36 -17 1791 895
use pinv_8  pinv_8_0
timestamp 1643678851
transform 1 0 1161 0 1 0
box -36 -17 819 895
use pinv_7  pinv_7_0
timestamp 1643678851
transform 1 0 702 0 1 0
box -36 -17 495 895
use pinv_0  pinv_0_0
timestamp 1643678851
transform 1 0 351 0 1 0
box -36 -17 387 895
use pinv_0  pinv_0_1
timestamp 1643678851
transform 1 0 0 0 1 0
box -36 -17 387 895
<< labels >>
rlabel locali s 5951 369 5951 369 4 Z
rlabel locali s 81 377 81 377 4 A
rlabel locali s 4131 0 4131 0 4 gnd
rlabel locali s 4131 838 4131 838 4 vdd
<< properties >>
string FIXED_BBOX 0 0 8262 838
string GDS_FILE sram_0rw2r1w_16_128_sky130A.gds
string GDS_END 2047248
string GDS_START 2045646
<< end >>
