magic
tech sky130A
timestamp 1643671299
<< checkpaint >>
rect -630 -651 13078 12971
<< metal1 >>
rect 0 11984 12448 11998
rect 0 11921 12448 11935
rect 0 11808 12448 11822
rect 0 11278 12448 11292
rect 0 11165 12448 11179
rect 0 11102 12448 11116
rect 0 10444 12448 10458
rect 0 10381 12448 10395
rect 0 10268 12448 10282
rect 0 9738 12448 9752
rect 0 9625 12448 9639
rect 0 9562 12448 9576
rect 0 8904 12448 8918
rect 0 8841 12448 8855
rect 0 8728 12448 8742
rect 0 8198 12448 8212
rect 0 8085 12448 8099
rect 0 8022 12448 8036
rect 0 7364 12448 7378
rect 0 7301 12448 7315
rect 0 7188 12448 7202
rect 0 6658 12448 6672
rect 0 6545 12448 6559
rect 0 6482 12448 6496
rect 0 5824 12448 5838
rect 0 5761 12448 5775
rect 0 5648 12448 5662
rect 0 5118 12448 5132
rect 0 5005 12448 5019
rect 0 4942 12448 4956
rect 0 4284 12448 4298
rect 0 4221 12448 4235
rect 0 4108 12448 4122
rect 0 3578 12448 3592
rect 0 3465 12448 3479
rect 0 3402 12448 3416
rect 0 2744 12448 2758
rect 0 2681 12448 2695
rect 0 2568 12448 2582
rect 0 2038 12448 2052
rect 0 1925 12448 1939
rect 0 1862 12448 1876
rect 0 1204 12448 1218
rect 0 1141 12448 1155
rect 0 1028 12448 1042
rect 0 498 12448 512
rect 0 385 12448 399
rect 0 322 12448 336
<< metal2 >>
rect 96 0 110 12320
rect 222 0 236 12320
rect 313 0 327 12320
rect 485 0 499 12320
rect 611 0 625 12320
rect 702 0 716 12320
rect 874 0 888 12320
rect 1000 0 1014 12320
rect 1091 0 1105 12320
rect 1263 0 1277 12320
rect 1389 0 1403 12320
rect 1480 0 1494 12320
rect 1652 0 1666 12320
rect 1778 0 1792 12320
rect 1869 0 1883 12320
rect 2041 0 2055 12320
rect 2167 0 2181 12320
rect 2258 0 2272 12320
rect 2430 0 2444 12320
rect 2556 0 2570 12320
rect 2647 0 2661 12320
rect 2819 0 2833 12320
rect 2945 0 2959 12320
rect 3036 0 3050 12320
rect 3208 0 3222 12320
rect 3334 0 3348 12320
rect 3425 0 3439 12320
rect 3597 0 3611 12320
rect 3723 0 3737 12320
rect 3814 0 3828 12320
rect 3986 0 4000 12320
rect 4112 0 4126 12320
rect 4203 0 4217 12320
rect 4375 0 4389 12320
rect 4501 0 4515 12320
rect 4592 0 4606 12320
rect 4764 0 4778 12320
rect 4890 0 4904 12320
rect 4981 0 4995 12320
rect 5153 0 5167 12320
rect 5279 0 5293 12320
rect 5370 0 5384 12320
rect 5542 0 5556 12320
rect 5668 0 5682 12320
rect 5759 0 5773 12320
rect 5931 0 5945 12320
rect 6057 0 6071 12320
rect 6148 0 6162 12320
rect 6320 0 6334 12320
rect 6446 0 6460 12320
rect 6537 0 6551 12320
rect 6709 0 6723 12320
rect 6835 0 6849 12320
rect 6926 0 6940 12320
rect 7098 0 7112 12320
rect 7224 0 7238 12320
rect 7315 0 7329 12320
rect 7487 0 7501 12320
rect 7613 0 7627 12320
rect 7704 0 7718 12320
rect 7876 0 7890 12320
rect 8002 0 8016 12320
rect 8093 0 8107 12320
rect 8265 0 8279 12320
rect 8391 0 8405 12320
rect 8482 0 8496 12320
rect 8654 0 8668 12320
rect 8780 0 8794 12320
rect 8871 0 8885 12320
rect 9043 0 9057 12320
rect 9169 0 9183 12320
rect 9260 0 9274 12320
rect 9432 0 9446 12320
rect 9558 0 9572 12320
rect 9649 0 9663 12320
rect 9821 0 9835 12320
rect 9947 0 9961 12320
rect 10038 0 10052 12320
rect 10210 0 10224 12320
rect 10336 0 10350 12320
rect 10427 0 10441 12320
rect 10599 0 10613 12320
rect 10725 0 10739 12320
rect 10816 0 10830 12320
rect 10988 0 11002 12320
rect 11114 0 11128 12320
rect 11205 0 11219 12320
rect 11377 0 11391 12320
rect 11503 0 11517 12320
rect 11594 0 11608 12320
rect 11766 0 11780 12320
rect 11892 0 11906 12320
rect 11983 0 11997 12320
rect 12155 0 12169 12320
rect 12281 0 12295 12320
rect 12372 0 12386 12320
use bitcell_array  bitcell_array_0
timestamp 1643671299
transform 1 0 0 0 1 0
box 0 -21 12448 12341
<< labels >>
rlabel metal1 s 0 385 12448 399 4 rwl_0_0
rlabel metal1 s 0 498 12448 512 4 rwl_1_0
rlabel metal1 s 0 322 12448 336 4 wwl_0_0
rlabel metal1 s 0 1141 12448 1155 4 rwl_0_1
rlabel metal1 s 0 1028 12448 1042 4 rwl_1_1
rlabel metal1 s 0 1204 12448 1218 4 wwl_0_1
rlabel metal1 s 0 1925 12448 1939 4 rwl_0_2
rlabel metal1 s 0 2038 12448 2052 4 rwl_1_2
rlabel metal1 s 0 1862 12448 1876 4 wwl_0_2
rlabel metal1 s 0 2681 12448 2695 4 rwl_0_3
rlabel metal1 s 0 2568 12448 2582 4 rwl_1_3
rlabel metal1 s 0 2744 12448 2758 4 wwl_0_3
rlabel metal1 s 0 3465 12448 3479 4 rwl_0_4
rlabel metal1 s 0 3578 12448 3592 4 rwl_1_4
rlabel metal1 s 0 3402 12448 3416 4 wwl_0_4
rlabel metal1 s 0 4221 12448 4235 4 rwl_0_5
rlabel metal1 s 0 4108 12448 4122 4 rwl_1_5
rlabel metal1 s 0 4284 12448 4298 4 wwl_0_5
rlabel metal1 s 0 5005 12448 5019 4 rwl_0_6
rlabel metal1 s 0 5118 12448 5132 4 rwl_1_6
rlabel metal1 s 0 4942 12448 4956 4 wwl_0_6
rlabel metal1 s 0 5761 12448 5775 4 rwl_0_7
rlabel metal1 s 0 5648 12448 5662 4 rwl_1_7
rlabel metal1 s 0 5824 12448 5838 4 wwl_0_7
rlabel metal1 s 0 6545 12448 6559 4 rwl_0_8
rlabel metal1 s 0 6658 12448 6672 4 rwl_1_8
rlabel metal1 s 0 6482 12448 6496 4 wwl_0_8
rlabel metal1 s 0 7301 12448 7315 4 rwl_0_9
rlabel metal1 s 0 7188 12448 7202 4 rwl_1_9
rlabel metal1 s 0 7364 12448 7378 4 wwl_0_9
rlabel metal1 s 0 8085 12448 8099 4 rwl_0_10
rlabel metal1 s 0 8198 12448 8212 4 rwl_1_10
rlabel metal1 s 0 8022 12448 8036 4 wwl_0_10
rlabel metal1 s 0 8841 12448 8855 4 rwl_0_11
rlabel metal1 s 0 8728 12448 8742 4 rwl_1_11
rlabel metal1 s 0 8904 12448 8918 4 wwl_0_11
rlabel metal1 s 0 9625 12448 9639 4 rwl_0_12
rlabel metal1 s 0 9738 12448 9752 4 rwl_1_12
rlabel metal1 s 0 9562 12448 9576 4 wwl_0_12
rlabel metal1 s 0 10381 12448 10395 4 rwl_0_13
rlabel metal1 s 0 10268 12448 10282 4 rwl_1_13
rlabel metal1 s 0 10444 12448 10458 4 wwl_0_13
rlabel metal1 s 0 11165 12448 11179 4 rwl_0_14
rlabel metal1 s 0 11278 12448 11292 4 rwl_1_14
rlabel metal1 s 0 11102 12448 11116 4 wwl_0_14
rlabel metal1 s 0 11921 12448 11935 4 rwl_0_15
rlabel metal1 s 0 11808 12448 11822 4 rwl_1_15
rlabel metal1 s 0 11984 12448 11998 4 wwl_0_15
rlabel metal2 s 96 0 110 12320 4 read_bl_0_0
rlabel metal2 s 485 0 499 12320 4 read_bl_0_1
rlabel metal2 s 874 0 888 12320 4 read_bl_0_2
rlabel metal2 s 1263 0 1277 12320 4 read_bl_0_3
rlabel metal2 s 1652 0 1666 12320 4 read_bl_0_4
rlabel metal2 s 2041 0 2055 12320 4 read_bl_0_5
rlabel metal2 s 2430 0 2444 12320 4 read_bl_0_6
rlabel metal2 s 2819 0 2833 12320 4 read_bl_0_7
rlabel metal2 s 3208 0 3222 12320 4 read_bl_0_8
rlabel metal2 s 3597 0 3611 12320 4 read_bl_0_9
rlabel metal2 s 3986 0 4000 12320 4 read_bl_0_10
rlabel metal2 s 4375 0 4389 12320 4 read_bl_0_11
rlabel metal2 s 4764 0 4778 12320 4 read_bl_0_12
rlabel metal2 s 5153 0 5167 12320 4 read_bl_0_13
rlabel metal2 s 5542 0 5556 12320 4 read_bl_0_14
rlabel metal2 s 5931 0 5945 12320 4 read_bl_0_15
rlabel metal2 s 6320 0 6334 12320 4 read_bl_0_16
rlabel metal2 s 6709 0 6723 12320 4 read_bl_0_17
rlabel metal2 s 7098 0 7112 12320 4 read_bl_0_18
rlabel metal2 s 7487 0 7501 12320 4 read_bl_0_19
rlabel metal2 s 7876 0 7890 12320 4 read_bl_0_20
rlabel metal2 s 8265 0 8279 12320 4 read_bl_0_21
rlabel metal2 s 8654 0 8668 12320 4 read_bl_0_22
rlabel metal2 s 9043 0 9057 12320 4 read_bl_0_23
rlabel metal2 s 9432 0 9446 12320 4 read_bl_0_24
rlabel metal2 s 9821 0 9835 12320 4 read_bl_0_25
rlabel metal2 s 10210 0 10224 12320 4 read_bl_0_26
rlabel metal2 s 10599 0 10613 12320 4 read_bl_0_27
rlabel metal2 s 10988 0 11002 12320 4 read_bl_0_28
rlabel metal2 s 11377 0 11391 12320 4 read_bl_0_29
rlabel metal2 s 11766 0 11780 12320 4 read_bl_0_30
rlabel metal2 s 12155 0 12169 12320 4 read_bl_0_31
rlabel metal2 s 222 0 236 12320 4 read_bl_1_0
rlabel metal2 s 611 0 625 12320 4 read_bl_1_1
rlabel metal2 s 1000 0 1014 12320 4 read_bl_1_2
rlabel metal2 s 1389 0 1403 12320 4 read_bl_1_3
rlabel metal2 s 1778 0 1792 12320 4 read_bl_1_4
rlabel metal2 s 2167 0 2181 12320 4 read_bl_1_5
rlabel metal2 s 2556 0 2570 12320 4 read_bl_1_6
rlabel metal2 s 2945 0 2959 12320 4 read_bl_1_7
rlabel metal2 s 3334 0 3348 12320 4 read_bl_1_8
rlabel metal2 s 3723 0 3737 12320 4 read_bl_1_9
rlabel metal2 s 4112 0 4126 12320 4 read_bl_1_10
rlabel metal2 s 4501 0 4515 12320 4 read_bl_1_11
rlabel metal2 s 4890 0 4904 12320 4 read_bl_1_12
rlabel metal2 s 5279 0 5293 12320 4 read_bl_1_13
rlabel metal2 s 5668 0 5682 12320 4 read_bl_1_14
rlabel metal2 s 6057 0 6071 12320 4 read_bl_1_15
rlabel metal2 s 6446 0 6460 12320 4 read_bl_1_16
rlabel metal2 s 6835 0 6849 12320 4 read_bl_1_17
rlabel metal2 s 7224 0 7238 12320 4 read_bl_1_18
rlabel metal2 s 7613 0 7627 12320 4 read_bl_1_19
rlabel metal2 s 8002 0 8016 12320 4 read_bl_1_20
rlabel metal2 s 8391 0 8405 12320 4 read_bl_1_21
rlabel metal2 s 8780 0 8794 12320 4 read_bl_1_22
rlabel metal2 s 9169 0 9183 12320 4 read_bl_1_23
rlabel metal2 s 9558 0 9572 12320 4 read_bl_1_24
rlabel metal2 s 9947 0 9961 12320 4 read_bl_1_25
rlabel metal2 s 10336 0 10350 12320 4 read_bl_1_26
rlabel metal2 s 10725 0 10739 12320 4 read_bl_1_27
rlabel metal2 s 11114 0 11128 12320 4 read_bl_1_28
rlabel metal2 s 11503 0 11517 12320 4 read_bl_1_29
rlabel metal2 s 11892 0 11906 12320 4 read_bl_1_30
rlabel metal2 s 12281 0 12295 12320 4 read_bl_1_31
rlabel metal2 s 313 0 327 12320 4 write_bl_0_0
rlabel metal2 s 702 0 716 12320 4 write_bl_0_1
rlabel metal2 s 1091 0 1105 12320 4 write_bl_0_2
rlabel metal2 s 1480 0 1494 12320 4 write_bl_0_3
rlabel metal2 s 1869 0 1883 12320 4 write_bl_0_4
rlabel metal2 s 2258 0 2272 12320 4 write_bl_0_5
rlabel metal2 s 2647 0 2661 12320 4 write_bl_0_6
rlabel metal2 s 3036 0 3050 12320 4 write_bl_0_7
rlabel metal2 s 3425 0 3439 12320 4 write_bl_0_8
rlabel metal2 s 3814 0 3828 12320 4 write_bl_0_9
rlabel metal2 s 4203 0 4217 12320 4 write_bl_0_10
rlabel metal2 s 4592 0 4606 12320 4 write_bl_0_11
rlabel metal2 s 4981 0 4995 12320 4 write_bl_0_12
rlabel metal2 s 5370 0 5384 12320 4 write_bl_0_13
rlabel metal2 s 5759 0 5773 12320 4 write_bl_0_14
rlabel metal2 s 6148 0 6162 12320 4 write_bl_0_15
rlabel metal2 s 6537 0 6551 12320 4 write_bl_0_16
rlabel metal2 s 6926 0 6940 12320 4 write_bl_0_17
rlabel metal2 s 7315 0 7329 12320 4 write_bl_0_18
rlabel metal2 s 7704 0 7718 12320 4 write_bl_0_19
rlabel metal2 s 8093 0 8107 12320 4 write_bl_0_20
rlabel metal2 s 8482 0 8496 12320 4 write_bl_0_21
rlabel metal2 s 8871 0 8885 12320 4 write_bl_0_22
rlabel metal2 s 9260 0 9274 12320 4 write_bl_0_23
rlabel metal2 s 9649 0 9663 12320 4 write_bl_0_24
rlabel metal2 s 10038 0 10052 12320 4 write_bl_0_25
rlabel metal2 s 10427 0 10441 12320 4 write_bl_0_26
rlabel metal2 s 10816 0 10830 12320 4 write_bl_0_27
rlabel metal2 s 11205 0 11219 12320 4 write_bl_0_28
rlabel metal2 s 11594 0 11608 12320 4 write_bl_0_29
rlabel metal2 s 11983 0 11997 12320 4 write_bl_0_30
rlabel metal2 s 12372 0 12386 12320 4 write_bl_0_31
<< properties >>
string FIXED_BBOX 0 0 24896 24640
string GDS_FILE sram_0rw2r1w_16_32_sky130A.gds
string GDS_END 417044
string GDS_START 389080
<< end >>
