magic
tech sky130A
magscale 1 2
timestamp 1644951705
<< checkpaint >>
rect -1260 -1284 49027 2212
<< metal1 >>
rect 712 900 764 906
rect 712 842 764 848
rect 3824 900 3876 906
rect 3824 842 3876 848
rect 6936 900 6988 906
rect 6936 842 6988 848
rect 10048 900 10100 906
rect 10048 842 10100 848
rect 13160 900 13212 906
rect 13160 842 13212 848
rect 16272 900 16324 906
rect 16272 842 16324 848
rect 19384 900 19436 906
rect 19384 842 19436 848
rect 22496 900 22548 906
rect 22496 842 22548 848
rect 25608 900 25660 906
rect 25608 842 25660 848
rect 28720 900 28772 906
rect 28720 842 28772 848
rect 31832 900 31884 906
rect 31832 842 31884 848
rect 34944 900 34996 906
rect 34944 842 34996 848
rect 38056 900 38108 906
rect 38056 842 38108 848
rect 41168 900 41220 906
rect 41168 842 41220 848
rect 44280 900 44332 906
rect 44280 842 44332 848
rect 47392 900 47444 906
rect 47392 842 47444 848
rect 0 356 47767 384
rect 712 68 764 74
rect 712 10 764 16
rect 3824 68 3876 74
rect 3824 10 3876 16
rect 6936 68 6988 74
rect 6936 10 6988 16
rect 10048 68 10100 74
rect 10048 10 10100 16
rect 13160 68 13212 74
rect 13160 10 13212 16
rect 16272 68 16324 74
rect 16272 10 16324 16
rect 19384 68 19436 74
rect 19384 10 19436 16
rect 22496 68 22548 74
rect 22496 10 22548 16
rect 25608 68 25660 74
rect 25608 10 25660 16
rect 28720 68 28772 74
rect 28720 10 28772 16
rect 31832 68 31884 74
rect 31832 10 31884 16
rect 34944 68 34996 74
rect 34944 10 34996 16
rect 38056 68 38108 74
rect 38056 10 38108 16
rect 41168 68 41220 74
rect 41168 10 41220 16
rect 44280 68 44332 74
rect 44280 10 44332 16
rect 47392 68 47444 74
rect 47392 10 47444 16
<< via1 >>
rect 712 848 764 900
rect 3824 848 3876 900
rect 6936 848 6988 900
rect 10048 848 10100 900
rect 13160 848 13212 900
rect 16272 848 16324 900
rect 19384 848 19436 900
rect 22496 848 22548 900
rect 25608 848 25660 900
rect 28720 848 28772 900
rect 31832 848 31884 900
rect 34944 848 34996 900
rect 38056 848 38108 900
rect 41168 848 41220 900
rect 44280 848 44332 900
rect 47392 848 47444 900
rect 712 16 764 68
rect 3824 16 3876 68
rect 6936 16 6988 68
rect 10048 16 10100 68
rect 13160 16 13212 68
rect 16272 16 16324 68
rect 19384 16 19436 68
rect 22496 16 22548 68
rect 25608 16 25660 68
rect 28720 16 28772 68
rect 31832 16 31884 68
rect 34944 16 34996 68
rect 38056 16 38108 68
rect 41168 16 41220 68
rect 44280 16 44332 68
rect 47392 16 47444 68
<< metal2 >>
rect 710 902 766 911
rect 710 837 766 846
rect 1019 322 1047 952
rect 3822 902 3878 911
rect 3822 837 3878 846
rect 4131 322 4159 952
rect 6934 902 6990 911
rect 6934 837 6990 846
rect 7243 322 7271 952
rect 10046 902 10102 911
rect 10046 837 10102 846
rect 10355 322 10383 952
rect 13158 902 13214 911
rect 13158 837 13214 846
rect 13467 322 13495 952
rect 16270 902 16326 911
rect 16270 837 16326 846
rect 16579 322 16607 952
rect 19382 902 19438 911
rect 19382 837 19438 846
rect 19691 322 19719 952
rect 22494 902 22550 911
rect 22494 837 22550 846
rect 22803 322 22831 952
rect 25606 902 25662 911
rect 25606 837 25662 846
rect 25915 322 25943 952
rect 28718 902 28774 911
rect 28718 837 28774 846
rect 29027 322 29055 952
rect 31830 902 31886 911
rect 31830 837 31886 846
rect 32139 322 32167 952
rect 34942 902 34998 911
rect 34942 837 34998 846
rect 35251 322 35279 952
rect 38054 902 38110 911
rect 38054 837 38110 846
rect 38363 322 38391 952
rect 41166 902 41222 911
rect 41166 837 41222 846
rect 41475 322 41503 952
rect 44278 902 44334 911
rect 44278 837 44334 846
rect 44587 322 44615 952
rect 47390 902 47446 911
rect 47390 837 47446 846
rect 47699 322 47727 952
rect 585 272 639 300
rect 3697 272 3751 300
rect 6809 272 6863 300
rect 9921 272 9975 300
rect 13033 272 13087 300
rect 16145 272 16199 300
rect 19257 272 19311 300
rect 22369 272 22423 300
rect 25481 272 25535 300
rect 28593 272 28647 300
rect 31705 272 31759 300
rect 34817 272 34871 300
rect 37929 272 37983 300
rect 41041 272 41095 300
rect 44153 272 44207 300
rect 47265 272 47319 300
rect 710 70 766 79
rect 710 5 766 14
rect 3822 70 3878 79
rect 3822 5 3878 14
rect 6934 70 6990 79
rect 6934 5 6990 14
rect 10046 70 10102 79
rect 10046 5 10102 14
rect 13158 70 13214 79
rect 13158 5 13214 14
rect 16270 70 16326 79
rect 16270 5 16326 14
rect 19382 70 19438 79
rect 19382 5 19438 14
rect 22494 70 22550 79
rect 22494 5 22550 14
rect 25606 70 25662 79
rect 25606 5 25662 14
rect 28718 70 28774 79
rect 28718 5 28774 14
rect 31830 70 31886 79
rect 31830 5 31886 14
rect 34942 70 34998 79
rect 34942 5 34998 14
rect 38054 70 38110 79
rect 38054 5 38110 14
rect 41166 70 41222 79
rect 41166 5 41222 14
rect 44278 70 44334 79
rect 44278 5 44334 14
rect 47390 70 47446 79
rect 47390 5 47446 14
<< via2 >>
rect 710 900 766 902
rect 710 848 712 900
rect 712 848 764 900
rect 764 848 766 900
rect 710 846 766 848
rect 3822 900 3878 902
rect 3822 848 3824 900
rect 3824 848 3876 900
rect 3876 848 3878 900
rect 3822 846 3878 848
rect 6934 900 6990 902
rect 6934 848 6936 900
rect 6936 848 6988 900
rect 6988 848 6990 900
rect 6934 846 6990 848
rect 10046 900 10102 902
rect 10046 848 10048 900
rect 10048 848 10100 900
rect 10100 848 10102 900
rect 10046 846 10102 848
rect 13158 900 13214 902
rect 13158 848 13160 900
rect 13160 848 13212 900
rect 13212 848 13214 900
rect 13158 846 13214 848
rect 16270 900 16326 902
rect 16270 848 16272 900
rect 16272 848 16324 900
rect 16324 848 16326 900
rect 16270 846 16326 848
rect 19382 900 19438 902
rect 19382 848 19384 900
rect 19384 848 19436 900
rect 19436 848 19438 900
rect 19382 846 19438 848
rect 22494 900 22550 902
rect 22494 848 22496 900
rect 22496 848 22548 900
rect 22548 848 22550 900
rect 22494 846 22550 848
rect 25606 900 25662 902
rect 25606 848 25608 900
rect 25608 848 25660 900
rect 25660 848 25662 900
rect 25606 846 25662 848
rect 28718 900 28774 902
rect 28718 848 28720 900
rect 28720 848 28772 900
rect 28772 848 28774 900
rect 28718 846 28774 848
rect 31830 900 31886 902
rect 31830 848 31832 900
rect 31832 848 31884 900
rect 31884 848 31886 900
rect 31830 846 31886 848
rect 34942 900 34998 902
rect 34942 848 34944 900
rect 34944 848 34996 900
rect 34996 848 34998 900
rect 34942 846 34998 848
rect 38054 900 38110 902
rect 38054 848 38056 900
rect 38056 848 38108 900
rect 38108 848 38110 900
rect 38054 846 38110 848
rect 41166 900 41222 902
rect 41166 848 41168 900
rect 41168 848 41220 900
rect 41220 848 41222 900
rect 41166 846 41222 848
rect 44278 900 44334 902
rect 44278 848 44280 900
rect 44280 848 44332 900
rect 44332 848 44334 900
rect 44278 846 44334 848
rect 47390 900 47446 902
rect 47390 848 47392 900
rect 47392 848 47444 900
rect 47444 848 47446 900
rect 47390 846 47446 848
rect 710 68 766 70
rect 710 16 712 68
rect 712 16 764 68
rect 764 16 766 68
rect 710 14 766 16
rect 3822 68 3878 70
rect 3822 16 3824 68
rect 3824 16 3876 68
rect 3876 16 3878 68
rect 3822 14 3878 16
rect 6934 68 6990 70
rect 6934 16 6936 68
rect 6936 16 6988 68
rect 6988 16 6990 68
rect 6934 14 6990 16
rect 10046 68 10102 70
rect 10046 16 10048 68
rect 10048 16 10100 68
rect 10100 16 10102 68
rect 10046 14 10102 16
rect 13158 68 13214 70
rect 13158 16 13160 68
rect 13160 16 13212 68
rect 13212 16 13214 68
rect 13158 14 13214 16
rect 16270 68 16326 70
rect 16270 16 16272 68
rect 16272 16 16324 68
rect 16324 16 16326 68
rect 16270 14 16326 16
rect 19382 68 19438 70
rect 19382 16 19384 68
rect 19384 16 19436 68
rect 19436 16 19438 68
rect 19382 14 19438 16
rect 22494 68 22550 70
rect 22494 16 22496 68
rect 22496 16 22548 68
rect 22548 16 22550 68
rect 22494 14 22550 16
rect 25606 68 25662 70
rect 25606 16 25608 68
rect 25608 16 25660 68
rect 25660 16 25662 68
rect 25606 14 25662 16
rect 28718 68 28774 70
rect 28718 16 28720 68
rect 28720 16 28772 68
rect 28772 16 28774 68
rect 28718 14 28774 16
rect 31830 68 31886 70
rect 31830 16 31832 68
rect 31832 16 31884 68
rect 31884 16 31886 68
rect 31830 14 31886 16
rect 34942 68 34998 70
rect 34942 16 34944 68
rect 34944 16 34996 68
rect 34996 16 34998 68
rect 34942 14 34998 16
rect 38054 68 38110 70
rect 38054 16 38056 68
rect 38056 16 38108 68
rect 38108 16 38110 68
rect 38054 14 38110 16
rect 41166 68 41222 70
rect 41166 16 41168 68
rect 41168 16 41220 68
rect 41220 16 41222 68
rect 41166 14 41222 16
rect 44278 68 44334 70
rect 44278 16 44280 68
rect 44280 16 44332 68
rect 44332 16 44334 68
rect 44278 14 44334 16
rect 47390 68 47446 70
rect 47390 16 47392 68
rect 47392 16 47444 68
rect 47444 16 47446 68
rect 47390 14 47446 16
<< metal3 >>
rect 705 902 771 940
rect 705 846 710 902
rect 766 846 771 902
rect 705 808 771 846
rect 3817 902 3883 940
rect 3817 846 3822 902
rect 3878 846 3883 902
rect 3817 808 3883 846
rect 6929 902 6995 940
rect 6929 846 6934 902
rect 6990 846 6995 902
rect 6929 808 6995 846
rect 10041 902 10107 940
rect 10041 846 10046 902
rect 10102 846 10107 902
rect 10041 808 10107 846
rect 13153 902 13219 940
rect 13153 846 13158 902
rect 13214 846 13219 902
rect 13153 808 13219 846
rect 16265 902 16331 940
rect 16265 846 16270 902
rect 16326 846 16331 902
rect 16265 808 16331 846
rect 19377 902 19443 940
rect 19377 846 19382 902
rect 19438 846 19443 902
rect 19377 808 19443 846
rect 22489 902 22555 940
rect 22489 846 22494 902
rect 22550 846 22555 902
rect 22489 808 22555 846
rect 25601 902 25667 940
rect 25601 846 25606 902
rect 25662 846 25667 902
rect 25601 808 25667 846
rect 28713 902 28779 940
rect 28713 846 28718 902
rect 28774 846 28779 902
rect 28713 808 28779 846
rect 31825 902 31891 940
rect 31825 846 31830 902
rect 31886 846 31891 902
rect 31825 808 31891 846
rect 34937 902 35003 940
rect 34937 846 34942 902
rect 34998 846 35003 902
rect 34937 808 35003 846
rect 38049 902 38115 940
rect 38049 846 38054 902
rect 38110 846 38115 902
rect 38049 808 38115 846
rect 41161 902 41227 940
rect 41161 846 41166 902
rect 41222 846 41227 902
rect 41161 808 41227 846
rect 44273 902 44339 940
rect 44273 846 44278 902
rect 44334 846 44339 902
rect 44273 808 44339 846
rect 47385 902 47451 940
rect 47385 846 47390 902
rect 47446 846 47451 902
rect 47385 808 47451 846
rect 705 70 771 108
rect 705 14 710 70
rect 766 14 771 70
rect 705 -24 771 14
rect 3817 70 3883 108
rect 3817 14 3822 70
rect 3878 14 3883 70
rect 3817 -24 3883 14
rect 6929 70 6995 108
rect 6929 14 6934 70
rect 6990 14 6995 70
rect 6929 -24 6995 14
rect 10041 70 10107 108
rect 10041 14 10046 70
rect 10102 14 10107 70
rect 10041 -24 10107 14
rect 13153 70 13219 108
rect 13153 14 13158 70
rect 13214 14 13219 70
rect 13153 -24 13219 14
rect 16265 70 16331 108
rect 16265 14 16270 70
rect 16326 14 16331 70
rect 16265 -24 16331 14
rect 19377 70 19443 108
rect 19377 14 19382 70
rect 19438 14 19443 70
rect 19377 -24 19443 14
rect 22489 70 22555 108
rect 22489 14 22494 70
rect 22550 14 22555 70
rect 22489 -24 22555 14
rect 25601 70 25667 108
rect 25601 14 25606 70
rect 25662 14 25667 70
rect 25601 -24 25667 14
rect 28713 70 28779 108
rect 28713 14 28718 70
rect 28774 14 28779 70
rect 28713 -24 28779 14
rect 31825 70 31891 108
rect 31825 14 31830 70
rect 31886 14 31891 70
rect 31825 -24 31891 14
rect 34937 70 35003 108
rect 34937 14 34942 70
rect 34998 14 35003 70
rect 34937 -24 35003 14
rect 38049 70 38115 108
rect 38049 14 38054 70
rect 38110 14 38115 70
rect 38049 -24 38115 14
rect 41161 70 41227 108
rect 41161 14 41166 70
rect 41222 14 41227 70
rect 41161 -24 41227 14
rect 44273 70 44339 108
rect 44273 14 44278 70
rect 44334 14 44339 70
rect 44273 -24 44339 14
rect 47385 70 47451 108
rect 47385 14 47390 70
rect 47446 14 47451 70
rect 47385 -24 47451 14
use contact_23  contact_23_0
timestamp 1644951705
transform 1 0 47385 0 1 -24
box 0 0 1 1
use contact_22  contact_22_0
timestamp 1644951705
transform 1 0 47392 0 1 10
box 0 0 1 1
use contact_23  contact_23_1
timestamp 1644951705
transform 1 0 47385 0 1 808
box 0 0 1 1
use contact_22  contact_22_1
timestamp 1644951705
transform 1 0 47392 0 1 842
box 0 0 1 1
use contact_23  contact_23_2
timestamp 1644951705
transform 1 0 44273 0 1 -24
box 0 0 1 1
use contact_22  contact_22_2
timestamp 1644951705
transform 1 0 44280 0 1 10
box 0 0 1 1
use contact_23  contact_23_3
timestamp 1644951705
transform 1 0 44273 0 1 808
box 0 0 1 1
use contact_22  contact_22_3
timestamp 1644951705
transform 1 0 44280 0 1 842
box 0 0 1 1
use contact_23  contact_23_4
timestamp 1644951705
transform 1 0 41161 0 1 -24
box 0 0 1 1
use contact_22  contact_22_4
timestamp 1644951705
transform 1 0 41168 0 1 10
box 0 0 1 1
use contact_23  contact_23_5
timestamp 1644951705
transform 1 0 41161 0 1 808
box 0 0 1 1
use contact_22  contact_22_5
timestamp 1644951705
transform 1 0 41168 0 1 842
box 0 0 1 1
use contact_23  contact_23_6
timestamp 1644951705
transform 1 0 38049 0 1 -24
box 0 0 1 1
use contact_22  contact_22_6
timestamp 1644951705
transform 1 0 38056 0 1 10
box 0 0 1 1
use contact_23  contact_23_7
timestamp 1644951705
transform 1 0 38049 0 1 808
box 0 0 1 1
use contact_22  contact_22_7
timestamp 1644951705
transform 1 0 38056 0 1 842
box 0 0 1 1
use contact_23  contact_23_8
timestamp 1644951705
transform 1 0 34937 0 1 -24
box 0 0 1 1
use contact_22  contact_22_8
timestamp 1644951705
transform 1 0 34944 0 1 10
box 0 0 1 1
use contact_23  contact_23_9
timestamp 1644951705
transform 1 0 34937 0 1 808
box 0 0 1 1
use contact_22  contact_22_9
timestamp 1644951705
transform 1 0 34944 0 1 842
box 0 0 1 1
use contact_23  contact_23_10
timestamp 1644951705
transform 1 0 31825 0 1 -24
box 0 0 1 1
use contact_22  contact_22_10
timestamp 1644951705
transform 1 0 31832 0 1 10
box 0 0 1 1
use contact_23  contact_23_11
timestamp 1644951705
transform 1 0 31825 0 1 808
box 0 0 1 1
use contact_22  contact_22_11
timestamp 1644951705
transform 1 0 31832 0 1 842
box 0 0 1 1
use contact_23  contact_23_12
timestamp 1644951705
transform 1 0 28713 0 1 -24
box 0 0 1 1
use contact_22  contact_22_12
timestamp 1644951705
transform 1 0 28720 0 1 10
box 0 0 1 1
use contact_23  contact_23_13
timestamp 1644951705
transform 1 0 28713 0 1 808
box 0 0 1 1
use contact_22  contact_22_13
timestamp 1644951705
transform 1 0 28720 0 1 842
box 0 0 1 1
use contact_23  contact_23_14
timestamp 1644951705
transform 1 0 25601 0 1 -24
box 0 0 1 1
use contact_22  contact_22_14
timestamp 1644951705
transform 1 0 25608 0 1 10
box 0 0 1 1
use contact_23  contact_23_15
timestamp 1644951705
transform 1 0 25601 0 1 808
box 0 0 1 1
use contact_22  contact_22_15
timestamp 1644951705
transform 1 0 25608 0 1 842
box 0 0 1 1
use contact_23  contact_23_16
timestamp 1644951705
transform 1 0 22489 0 1 -24
box 0 0 1 1
use contact_22  contact_22_16
timestamp 1644951705
transform 1 0 22496 0 1 10
box 0 0 1 1
use contact_23  contact_23_17
timestamp 1644951705
transform 1 0 22489 0 1 808
box 0 0 1 1
use contact_22  contact_22_17
timestamp 1644951705
transform 1 0 22496 0 1 842
box 0 0 1 1
use contact_23  contact_23_18
timestamp 1644951705
transform 1 0 19377 0 1 -24
box 0 0 1 1
use contact_22  contact_22_18
timestamp 1644951705
transform 1 0 19384 0 1 10
box 0 0 1 1
use contact_23  contact_23_19
timestamp 1644951705
transform 1 0 19377 0 1 808
box 0 0 1 1
use contact_22  contact_22_19
timestamp 1644951705
transform 1 0 19384 0 1 842
box 0 0 1 1
use contact_23  contact_23_20
timestamp 1644951705
transform 1 0 16265 0 1 -24
box 0 0 1 1
use contact_22  contact_22_20
timestamp 1644951705
transform 1 0 16272 0 1 10
box 0 0 1 1
use contact_23  contact_23_21
timestamp 1644951705
transform 1 0 16265 0 1 808
box 0 0 1 1
use contact_22  contact_22_21
timestamp 1644951705
transform 1 0 16272 0 1 842
box 0 0 1 1
use contact_23  contact_23_22
timestamp 1644951705
transform 1 0 13153 0 1 -24
box 0 0 1 1
use contact_22  contact_22_22
timestamp 1644951705
transform 1 0 13160 0 1 10
box 0 0 1 1
use contact_23  contact_23_23
timestamp 1644951705
transform 1 0 13153 0 1 808
box 0 0 1 1
use contact_22  contact_22_23
timestamp 1644951705
transform 1 0 13160 0 1 842
box 0 0 1 1
use contact_23  contact_23_24
timestamp 1644951705
transform 1 0 10041 0 1 -24
box 0 0 1 1
use contact_22  contact_22_24
timestamp 1644951705
transform 1 0 10048 0 1 10
box 0 0 1 1
use contact_23  contact_23_25
timestamp 1644951705
transform 1 0 10041 0 1 808
box 0 0 1 1
use contact_22  contact_22_25
timestamp 1644951705
transform 1 0 10048 0 1 842
box 0 0 1 1
use contact_23  contact_23_26
timestamp 1644951705
transform 1 0 6929 0 1 -24
box 0 0 1 1
use contact_22  contact_22_26
timestamp 1644951705
transform 1 0 6936 0 1 10
box 0 0 1 1
use contact_23  contact_23_27
timestamp 1644951705
transform 1 0 6929 0 1 808
box 0 0 1 1
use contact_22  contact_22_27
timestamp 1644951705
transform 1 0 6936 0 1 842
box 0 0 1 1
use contact_23  contact_23_28
timestamp 1644951705
transform 1 0 3817 0 1 -24
box 0 0 1 1
use contact_22  contact_22_28
timestamp 1644951705
transform 1 0 3824 0 1 10
box 0 0 1 1
use contact_23  contact_23_29
timestamp 1644951705
transform 1 0 3817 0 1 808
box 0 0 1 1
use contact_22  contact_22_29
timestamp 1644951705
transform 1 0 3824 0 1 842
box 0 0 1 1
use contact_23  contact_23_30
timestamp 1644951705
transform 1 0 705 0 1 -24
box 0 0 1 1
use contact_22  contact_22_30
timestamp 1644951705
transform 1 0 712 0 1 10
box 0 0 1 1
use contact_23  contact_23_31
timestamp 1644951705
transform 1 0 705 0 1 808
box 0 0 1 1
use contact_22  contact_22_31
timestamp 1644951705
transform 1 0 712 0 1 842
box 0 0 1 1
use write_driver_multiport  write_driver_multiport_0
timestamp 1644951705
transform 1 0 47069 0 1 0
box 0 0 698 952
use write_driver_multiport  write_driver_multiport_1
timestamp 1644951705
transform 1 0 43957 0 1 0
box 0 0 698 952
use write_driver_multiport  write_driver_multiport_2
timestamp 1644951705
transform 1 0 40845 0 1 0
box 0 0 698 952
use write_driver_multiport  write_driver_multiport_3
timestamp 1644951705
transform 1 0 37733 0 1 0
box 0 0 698 952
use write_driver_multiport  write_driver_multiport_4
timestamp 1644951705
transform 1 0 34621 0 1 0
box 0 0 698 952
use write_driver_multiport  write_driver_multiport_5
timestamp 1644951705
transform 1 0 31509 0 1 0
box 0 0 698 952
use write_driver_multiport  write_driver_multiport_6
timestamp 1644951705
transform 1 0 28397 0 1 0
box 0 0 698 952
use write_driver_multiport  write_driver_multiport_7
timestamp 1644951705
transform 1 0 25285 0 1 0
box 0 0 698 952
use write_driver_multiport  write_driver_multiport_8
timestamp 1644951705
transform 1 0 22173 0 1 0
box 0 0 698 952
use write_driver_multiport  write_driver_multiport_9
timestamp 1644951705
transform 1 0 19061 0 1 0
box 0 0 698 952
use write_driver_multiport  write_driver_multiport_10
timestamp 1644951705
transform 1 0 15949 0 1 0
box 0 0 698 952
use write_driver_multiport  write_driver_multiport_11
timestamp 1644951705
transform 1 0 12837 0 1 0
box 0 0 698 952
use write_driver_multiport  write_driver_multiport_12
timestamp 1644951705
transform 1 0 9725 0 1 0
box 0 0 698 952
use write_driver_multiport  write_driver_multiport_13
timestamp 1644951705
transform 1 0 6613 0 1 0
box 0 0 698 952
use write_driver_multiport  write_driver_multiport_14
timestamp 1644951705
transform 1 0 3501 0 1 0
box 0 0 698 952
use write_driver_multiport  write_driver_multiport_15
timestamp 1644951705
transform 1 0 389 0 1 0
box 0 0 698 952
<< labels >>
rlabel metal2 s 585 272 639 300 4 din_0
rlabel metal2 s 1019 322 1047 952 4 wbl0_0
rlabel metal3 s 41161 808 41227 940 4 vdd
rlabel metal3 s 47385 808 47451 940 4 vdd
rlabel metal3 s 705 808 771 940 4 vdd
rlabel metal3 s 10041 808 10107 940 4 vdd
rlabel metal3 s 13153 808 13219 940 4 vdd
rlabel metal3 s 6929 808 6995 940 4 vdd
rlabel metal3 s 16265 808 16331 940 4 vdd
rlabel metal3 s 28713 808 28779 940 4 vdd
rlabel metal3 s 19377 808 19443 940 4 vdd
rlabel metal3 s 25601 808 25667 940 4 vdd
rlabel metal3 s 38049 808 38115 940 4 vdd
rlabel metal3 s 44273 808 44339 940 4 vdd
rlabel metal3 s 34937 808 35003 940 4 vdd
rlabel metal3 s 22489 808 22555 940 4 vdd
rlabel metal3 s 31825 808 31891 940 4 vdd
rlabel metal3 s 3817 808 3883 940 4 vdd
rlabel metal3 s 6929 -24 6995 108 4 gnd
rlabel metal3 s 16265 -24 16331 108 4 gnd
rlabel metal3 s 3817 -24 3883 108 4 gnd
rlabel metal3 s 41161 -24 41227 108 4 gnd
rlabel metal3 s 28713 -24 28779 108 4 gnd
rlabel metal3 s 22489 -24 22555 108 4 gnd
rlabel metal3 s 31825 -24 31891 108 4 gnd
rlabel metal3 s 19377 -24 19443 108 4 gnd
rlabel metal3 s 34937 -24 35003 108 4 gnd
rlabel metal3 s 10041 -24 10107 108 4 gnd
rlabel metal3 s 705 -24 771 108 4 gnd
rlabel metal3 s 38049 -24 38115 108 4 gnd
rlabel metal3 s 44273 -24 44339 108 4 gnd
rlabel metal3 s 25601 -24 25667 108 4 gnd
rlabel metal3 s 13153 -24 13219 108 4 gnd
rlabel metal3 s 47385 -24 47451 108 4 gnd
rlabel metal2 s 3697 272 3751 300 4 din_1
rlabel metal2 s 4131 322 4159 952 4 wbl0_1
rlabel metal2 s 6809 272 6863 300 4 din_2
rlabel metal2 s 7243 322 7271 952 4 wbl0_2
rlabel metal2 s 9921 272 9975 300 4 din_3
rlabel metal2 s 10355 322 10383 952 4 wbl0_3
rlabel metal2 s 13033 272 13087 300 4 din_4
rlabel metal2 s 13467 322 13495 952 4 wbl0_4
rlabel metal2 s 16145 272 16199 300 4 din_5
rlabel metal2 s 16579 322 16607 952 4 wbl0_5
rlabel metal2 s 19257 272 19311 300 4 din_6
rlabel metal2 s 19691 322 19719 952 4 wbl0_6
rlabel metal2 s 22369 272 22423 300 4 din_7
rlabel metal2 s 22803 322 22831 952 4 wbl0_7
rlabel metal2 s 25481 272 25535 300 4 din_8
rlabel metal2 s 25915 322 25943 952 4 wbl0_8
rlabel metal2 s 28593 272 28647 300 4 din_9
rlabel metal2 s 29027 322 29055 952 4 wbl0_9
rlabel metal2 s 31705 272 31759 300 4 din_10
rlabel metal2 s 32139 322 32167 952 4 wbl0_10
rlabel metal2 s 34817 272 34871 300 4 din_11
rlabel metal2 s 35251 322 35279 952 4 wbl0_11
rlabel metal2 s 37929 272 37983 300 4 din_12
rlabel metal2 s 38363 322 38391 952 4 wbl0_12
rlabel metal2 s 41041 272 41095 300 4 din_13
rlabel metal2 s 41475 322 41503 952 4 wbl0_13
rlabel metal2 s 44153 272 44207 300 4 din_14
rlabel metal2 s 44587 322 44615 952 4 wbl0_14
rlabel metal2 s 47265 272 47319 300 4 din_15
rlabel metal2 s 47699 322 47727 952 4 wbl0_15
rlabel metal1 s 0 356 47767 384 4 en
<< properties >>
string FIXED_BBOX 47385 -24 47451 0
string GDS_FILE sram_0rw2r1w_16_128_sky130A.gds
string GDS_END 1512750
string GDS_START 1495014
<< end >>
