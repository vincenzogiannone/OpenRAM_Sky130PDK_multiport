magic
tech sky130A
magscale 1 2
timestamp 1644949024
<< checkpaint >>
rect -1296 -1277 3284 2155
<< nwell >>
rect -36 402 2024 895
<< pwell >>
rect 1878 51 1928 133
<< psubdiff >>
rect 1878 109 1928 133
rect 1878 75 1886 109
rect 1920 75 1928 109
rect 1878 51 1928 75
<< nsubdiff >>
rect 1878 763 1928 787
rect 1878 729 1886 763
rect 1920 729 1928 763
rect 1878 705 1928 729
<< psubdiffcont >>
rect 1886 75 1920 109
<< nsubdiffcont >>
rect 1886 729 1920 763
<< poly >>
rect 114 404 144 447
rect 48 388 144 404
rect 48 354 64 388
rect 98 354 144 388
rect 48 338 144 354
rect 114 201 144 338
<< polycont >>
rect 64 354 98 388
<< locali >>
rect 0 821 1988 855
rect 62 612 96 821
rect 274 612 308 821
rect 490 612 524 821
rect 706 612 740 821
rect 922 612 956 821
rect 1138 612 1172 821
rect 1354 612 1388 821
rect 1570 612 1604 821
rect 1782 612 1816 821
rect 1886 763 1920 821
rect 1886 713 1920 729
rect 48 388 114 404
rect 48 354 64 388
rect 98 354 114 388
rect 48 338 114 354
rect 922 388 956 578
rect 922 354 973 388
rect 922 165 956 354
rect 1886 109 1920 125
rect 62 17 96 65
rect 274 17 308 65
rect 490 17 524 65
rect 706 17 740 65
rect 922 17 956 65
rect 1138 17 1172 65
rect 1354 17 1388 65
rect 1570 17 1604 65
rect 1782 17 1816 65
rect 1886 17 1920 75
rect 0 -17 1988 17
use contact_12  contact_12_0
timestamp 1644949024
transform 1 0 48 0 1 338
box 0 0 1 1
use contact_11  contact_11_0
timestamp 1644949024
transform 1 0 1878 0 1 51
box 0 0 1 1
use contact_10  contact_10_0
timestamp 1644949024
transform 1 0 1878 0 1 705
box 0 0 1 1
use nmos_m16_w0_470_sli_dli_da_p  nmos_m16_w0_470_sli_dli_da_p_0
timestamp 1644949024
transform 1 0 54 0 1 51
box 0 -26 1770 150
use pmos_m16_w1_420_sli_dli_da_p  pmos_m16_w1_420_sli_dli_da_p_0
timestamp 1644949024
transform 1 0 54 0 1 503
box -59 -56 1829 338
<< labels >>
rlabel locali s 81 371 81 371 4 A
rlabel locali s 956 371 956 371 4 Z
rlabel locali s 994 0 994 0 4 gnd
rlabel locali s 994 838 994 838 4 vdd
<< properties >>
string FIXED_BBOX 0 0 1988 838
string GDS_FILE sram_0rw2r1w_4_16_sky130A.gds
string GDS_END 476638
string GDS_START 474122
<< end >>
