magic
tech sky130A
timestamp 1643153523
<< nwell >>
rect 0 488 602 808
<< nmos >>
rect 47 154 62 209
rect 95 154 110 209
rect 143 154 158 209
rect 191 154 206 209
rect 293 154 308 209
rect 341 154 356 209
rect 392 154 407 196
rect 492 154 507 196
rect 540 154 555 196
<< pmos >>
rect 47 506 62 548
rect 95 506 110 548
rect 143 506 158 548
rect 191 506 206 548
rect 293 506 308 548
rect 341 506 356 548
rect 392 506 407 641
rect 492 506 507 641
rect 540 506 555 641
<< ndiff >>
rect 18 191 47 209
rect 18 174 22 191
rect 39 174 47 191
rect 18 154 47 174
rect 62 154 95 209
rect 110 191 143 209
rect 110 174 118 191
rect 135 174 143 191
rect 110 154 143 174
rect 158 154 191 209
rect 206 191 235 209
rect 206 174 214 191
rect 231 174 235 191
rect 206 154 235 174
rect 264 191 293 209
rect 264 174 268 191
rect 285 174 293 191
rect 264 154 293 174
rect 308 154 341 209
rect 356 196 384 209
rect 356 191 392 196
rect 356 174 364 191
rect 381 174 392 191
rect 356 154 392 174
rect 407 184 436 196
rect 407 167 415 184
rect 432 167 436 184
rect 407 154 436 167
rect 463 184 492 196
rect 463 167 467 184
rect 484 167 492 184
rect 463 154 492 167
rect 507 184 540 196
rect 507 167 515 184
rect 532 167 540 184
rect 507 154 540 167
rect 555 184 584 196
rect 555 167 563 184
rect 580 167 584 184
rect 555 154 584 167
<< pdiff >>
rect 364 625 392 641
rect 364 608 368 625
rect 385 608 392 625
rect 364 583 392 608
rect 364 566 368 583
rect 385 566 392 583
rect 364 548 392 566
rect 18 535 47 548
rect 18 518 22 535
rect 39 518 47 535
rect 18 506 47 518
rect 62 535 95 548
rect 62 518 70 535
rect 87 518 95 535
rect 62 506 95 518
rect 110 535 143 548
rect 110 518 118 535
rect 135 518 143 535
rect 110 506 143 518
rect 158 535 191 548
rect 158 518 166 535
rect 183 518 191 535
rect 158 506 191 518
rect 206 535 235 548
rect 206 518 214 535
rect 231 518 235 535
rect 206 506 235 518
rect 264 535 293 548
rect 264 518 268 535
rect 285 518 293 535
rect 264 506 293 518
rect 308 534 341 548
rect 308 517 316 534
rect 333 517 341 534
rect 308 506 341 517
rect 356 534 392 548
rect 356 517 366 534
rect 383 517 392 534
rect 356 506 392 517
rect 407 625 436 641
rect 407 608 415 625
rect 432 608 436 625
rect 407 583 436 608
rect 407 566 415 583
rect 432 566 436 583
rect 407 540 436 566
rect 407 523 415 540
rect 432 523 436 540
rect 407 506 436 523
rect 463 625 492 641
rect 463 608 467 625
rect 484 608 492 625
rect 463 583 492 608
rect 463 566 467 583
rect 484 566 492 583
rect 463 540 492 566
rect 463 523 467 540
rect 484 523 492 540
rect 463 506 492 523
rect 507 625 540 641
rect 507 608 515 625
rect 532 608 540 625
rect 507 583 540 608
rect 507 566 515 583
rect 532 566 540 583
rect 507 540 540 566
rect 507 523 515 540
rect 532 523 540 540
rect 507 506 540 523
rect 555 625 584 641
rect 555 608 563 625
rect 580 608 584 625
rect 555 583 584 608
rect 555 566 563 583
rect 580 566 584 583
rect 555 540 584 566
rect 555 523 563 540
rect 580 523 584 540
rect 555 506 584 523
<< ndiffc >>
rect 22 174 39 191
rect 118 174 135 191
rect 214 174 231 191
rect 268 174 285 191
rect 364 174 381 191
rect 415 167 432 184
rect 467 167 484 184
rect 515 167 532 184
rect 563 167 580 184
<< pdiffc >>
rect 368 608 385 625
rect 368 566 385 583
rect 22 518 39 535
rect 70 518 87 535
rect 118 518 135 535
rect 166 518 183 535
rect 214 518 231 535
rect 268 518 285 535
rect 316 517 333 534
rect 366 517 383 534
rect 415 608 432 625
rect 415 566 432 583
rect 415 523 432 540
rect 467 608 484 625
rect 467 566 484 583
rect 467 523 484 540
rect 515 608 532 625
rect 515 566 532 583
rect 515 523 532 540
rect 563 608 580 625
rect 563 566 580 583
rect 563 523 580 540
<< psubdiff >>
rect 92 9 128 21
rect 92 -9 101 9
rect 119 -9 128 9
rect 92 -21 128 -9
rect 219 9 255 21
rect 219 -9 228 9
rect 246 -9 255 9
rect 219 -21 255 -9
rect 347 9 383 21
rect 347 -9 356 9
rect 374 -9 383 9
rect 347 -21 383 -9
rect 474 9 510 21
rect 474 -9 483 9
rect 500 -9 510 9
rect 474 -21 510 -9
<< nsubdiff >>
rect 92 778 128 790
rect 92 760 101 778
rect 119 760 128 778
rect 92 748 128 760
rect 219 778 255 790
rect 219 760 228 778
rect 246 760 255 778
rect 219 748 255 760
rect 347 778 383 790
rect 347 760 356 778
rect 374 760 383 778
rect 347 748 383 760
rect 474 778 510 790
rect 474 760 483 778
rect 501 760 510 778
rect 474 748 510 760
<< psubdiffcont >>
rect 101 -9 119 9
rect 228 -9 246 9
rect 356 -9 374 9
rect 483 -9 500 9
<< nsubdiffcont >>
rect 101 760 119 778
rect 228 760 246 778
rect 356 760 374 778
rect 483 760 501 778
<< poly >>
rect 392 641 407 654
rect 492 641 507 654
rect 540 641 555 654
rect 47 548 62 561
rect 95 548 110 561
rect 143 548 158 561
rect 191 548 206 561
rect 293 548 308 561
rect 341 548 356 561
rect 47 457 62 506
rect 35 449 62 457
rect 35 432 40 449
rect 57 432 62 449
rect 35 424 62 432
rect 95 429 110 506
rect 47 209 62 424
rect 83 421 110 429
rect 83 404 88 421
rect 105 404 110 421
rect 83 396 110 404
rect 143 401 158 506
rect 95 209 110 396
rect 131 393 158 401
rect 131 376 136 393
rect 153 376 158 393
rect 131 368 158 376
rect 191 373 206 506
rect 143 209 158 368
rect 179 365 206 373
rect 179 348 184 365
rect 201 348 206 365
rect 179 340 206 348
rect 191 209 206 340
rect 293 319 308 506
rect 281 311 308 319
rect 281 294 286 311
rect 303 294 308 311
rect 281 286 308 294
rect 341 291 356 506
rect 392 350 407 506
rect 380 342 407 350
rect 380 325 385 342
rect 402 325 407 342
rect 380 317 407 325
rect 293 209 308 286
rect 329 283 356 291
rect 329 266 334 283
rect 351 266 356 283
rect 329 258 356 266
rect 341 209 356 258
rect 392 196 407 317
rect 492 393 507 506
rect 540 457 555 506
rect 528 449 555 457
rect 528 432 533 449
rect 550 432 555 449
rect 528 424 555 432
rect 492 385 519 393
rect 492 368 497 385
rect 514 368 519 385
rect 492 360 519 368
rect 492 196 507 360
rect 540 196 555 424
rect 47 141 62 154
rect 95 141 110 154
rect 143 141 158 154
rect 191 141 206 154
rect 293 141 308 154
rect 341 141 356 154
rect 392 141 407 154
rect 492 141 507 154
rect 540 141 555 154
<< polycont >>
rect 40 432 57 449
rect 88 404 105 421
rect 136 376 153 393
rect 184 348 201 365
rect 286 294 303 311
rect 385 325 402 342
rect 334 266 351 283
rect 533 432 550 449
rect 497 368 514 385
<< locali >>
rect 22 778 580 786
rect 22 760 101 778
rect 119 760 228 778
rect 246 760 356 778
rect 374 760 483 778
rect 501 760 580 778
rect 22 752 580 760
rect 22 548 39 752
rect 118 548 135 752
rect 214 548 231 752
rect 268 548 285 752
rect 368 641 385 752
rect 515 641 532 752
rect 364 625 387 641
rect 364 608 368 625
rect 385 608 387 625
rect 364 583 387 608
rect 364 566 368 583
rect 385 566 387 583
rect 364 548 387 566
rect 18 535 42 548
rect 18 518 22 535
rect 39 518 42 535
rect 18 506 42 518
rect 67 535 90 548
rect 67 518 70 535
rect 87 518 90 535
rect 67 506 90 518
rect 115 535 138 548
rect 115 518 118 535
rect 135 518 138 535
rect 115 506 138 518
rect 163 535 186 548
rect 163 518 166 535
rect 183 518 186 535
rect 163 506 186 518
rect 211 535 235 548
rect 211 518 214 535
rect 231 518 235 535
rect 211 506 235 518
rect 264 535 288 548
rect 264 518 268 535
rect 285 518 288 535
rect 264 506 288 518
rect 313 534 336 548
rect 313 517 316 534
rect 333 517 336 534
rect 313 506 336 517
rect 361 534 387 548
rect 361 517 366 534
rect 383 517 387 534
rect 361 506 387 517
rect 412 625 436 641
rect 412 608 415 625
rect 432 608 436 625
rect 412 583 436 608
rect 412 566 415 583
rect 432 566 436 583
rect 412 540 436 566
rect 412 523 415 540
rect 432 523 436 540
rect 412 506 436 523
rect 40 449 57 457
rect 169 456 186 506
rect 169 439 255 456
rect 40 424 57 432
rect 88 421 105 429
rect 88 396 105 404
rect 136 393 153 401
rect 136 368 153 376
rect 184 365 201 373
rect 184 340 201 348
rect 218 323 235 392
rect 25 306 235 323
rect 25 209 42 306
rect 252 289 269 439
rect 316 376 333 506
rect 316 359 402 376
rect 380 342 402 359
rect 380 333 385 342
rect 218 272 269 289
rect 286 311 303 319
rect 385 317 402 325
rect 286 286 303 294
rect 419 298 436 506
rect 334 283 351 291
rect 218 209 235 272
rect 334 258 351 266
rect 18 191 42 209
rect 18 174 22 191
rect 39 174 42 191
rect 18 154 42 174
rect 115 191 138 209
rect 115 174 118 191
rect 135 174 138 191
rect 115 154 138 174
rect 211 191 235 209
rect 211 174 214 191
rect 231 174 235 191
rect 211 154 235 174
rect 264 191 288 209
rect 264 174 268 191
rect 285 174 288 191
rect 264 154 288 174
rect 361 191 384 209
rect 419 196 436 281
rect 361 174 364 191
rect 381 174 384 191
rect 361 154 384 174
rect 412 184 436 196
rect 412 167 415 184
rect 432 167 436 184
rect 412 154 436 167
rect 463 625 487 641
rect 463 608 467 625
rect 484 608 487 625
rect 463 583 487 608
rect 463 566 467 583
rect 484 566 487 583
rect 463 540 487 566
rect 463 523 467 540
rect 484 523 487 540
rect 463 506 487 523
rect 512 625 535 641
rect 512 608 515 625
rect 532 608 535 625
rect 512 583 535 608
rect 512 566 515 583
rect 532 566 535 583
rect 512 540 535 566
rect 512 523 515 540
rect 532 523 535 540
rect 512 506 535 523
rect 560 625 584 641
rect 560 608 563 625
rect 580 608 584 625
rect 560 583 584 608
rect 560 566 563 583
rect 580 566 584 583
rect 560 540 584 566
rect 560 523 563 540
rect 580 523 584 540
rect 560 506 584 523
rect 463 342 480 506
rect 533 449 550 457
rect 533 424 550 432
rect 567 439 584 506
rect 567 422 571 439
rect 497 385 514 393
rect 497 360 514 368
rect 463 196 480 325
rect 567 196 584 422
rect 463 184 487 196
rect 463 167 467 184
rect 484 167 487 184
rect 463 154 487 167
rect 512 184 535 196
rect 512 167 515 184
rect 532 167 535 184
rect 512 154 535 167
rect 560 184 584 196
rect 560 167 563 184
rect 580 167 584 184
rect 560 154 584 167
rect 118 17 135 154
rect 364 17 381 154
rect 515 17 532 154
rect 69 9 532 17
rect 69 -9 101 9
rect 119 -9 228 9
rect 246 -9 356 9
rect 374 -9 483 9
rect 500 -9 532 9
rect 69 -17 532 -9
<< viali >>
rect 101 760 119 778
rect 228 760 246 778
rect 356 760 374 778
rect 483 760 501 778
rect 70 518 87 535
rect 40 432 57 449
rect 255 439 272 456
rect 88 404 105 421
rect 136 376 153 393
rect 218 392 235 409
rect 184 348 201 365
rect 385 325 402 342
rect 286 294 303 311
rect 334 266 351 283
rect 419 281 436 298
rect 268 174 285 191
rect 533 432 550 449
rect 571 422 588 439
rect 497 368 514 385
rect 463 325 480 342
rect 101 -9 119 9
rect 228 -9 246 9
rect 356 -9 374 9
rect 483 -9 500 9
<< metal1 >>
rect 0 778 602 784
rect 0 760 101 778
rect 119 760 228 778
rect 246 760 356 778
rect 374 760 483 778
rect 501 760 602 778
rect 0 754 602 760
rect 67 535 90 541
rect 67 518 70 535
rect 87 526 90 535
rect 87 518 238 526
rect 67 512 238 518
rect 36 449 63 456
rect 36 439 40 449
rect 35 432 40 439
rect 57 432 63 449
rect 35 425 63 432
rect 84 421 111 428
rect 84 411 88 421
rect 83 404 88 411
rect 105 404 111 421
rect 224 415 238 512
rect 252 456 275 462
rect 252 439 255 456
rect 272 447 275 456
rect 529 449 553 455
rect 529 447 533 449
rect 272 439 533 447
rect 252 433 533 439
rect 529 432 533 433
rect 550 432 553 449
rect 529 425 553 432
rect 568 439 591 446
rect 568 422 571 439
rect 588 438 591 439
rect 588 424 602 438
rect 588 422 591 424
rect 568 415 591 422
rect 83 397 111 404
rect 215 409 238 415
rect 132 393 159 400
rect 132 383 136 393
rect 131 376 136 383
rect 153 376 159 393
rect 215 392 218 409
rect 235 400 238 409
rect 235 392 517 400
rect 215 386 517 392
rect 131 369 159 376
rect 494 385 517 386
rect 180 365 207 372
rect 180 355 184 365
rect 179 348 184 355
rect 201 348 207 365
rect 494 368 497 385
rect 514 368 517 385
rect 494 362 517 368
rect 556 351 602 365
rect 179 341 207 348
rect 371 342 406 349
rect 371 325 385 342
rect 402 325 406 342
rect 371 319 406 325
rect 460 343 483 348
rect 556 343 570 351
rect 460 342 570 343
rect 460 325 463 342
rect 480 329 570 342
rect 480 325 483 329
rect 460 319 483 325
rect 282 311 309 318
rect 282 301 286 311
rect 281 294 286 301
rect 303 294 309 311
rect 281 287 309 294
rect 330 283 357 290
rect 330 273 334 283
rect 329 266 334 273
rect 351 266 357 283
rect 329 259 357 266
rect 371 197 385 319
rect 416 298 602 304
rect 416 281 419 298
rect 436 290 602 298
rect 436 281 439 290
rect 416 275 439 281
rect 265 191 385 197
rect 265 174 268 191
rect 285 183 385 191
rect 285 174 288 183
rect 265 168 288 174
rect 0 9 602 15
rect 0 -9 101 9
rect 119 -9 228 9
rect 246 -9 356 9
rect 374 -9 483 9
rect 500 -9 602 9
rect 0 -15 602 -9
<< labels >>
flabel metal1 35 431 35 431 0 FreeSans 80 0 0 0 A0
port 0 nsew
flabel metal1 83 403 83 403 0 FreeSans 80 0 0 0 B0
port 1 nsew
flabel metal1 131 374 131 374 0 FreeSans 80 0 0 0 A1
port 3 nsew
flabel metal1 179 347 179 347 0 FreeSans 80 0 0 0 B1
port 4 nsew
flabel metal1 281 294 281 294 0 FreeSans 80 0 0 0 A2
port 5 nsew
flabel metal1 329 265 329 265 0 FreeSans 80 0 0 0 B2
port 6 nsew
flabel metal1 599 431 599 431 0 FreeSans 80 0 0 0 OUT1
port 7 nsew
flabel metal1 596 358 596 358 0 FreeSans 80 0 0 0 OUT0
port 8 nsew
flabel metal1 595 297 595 297 0 FreeSans 80 0 0 0 OUT2
port 9 nsew
flabel ndiff 78 178 78 178 0 FreeSans 80 0 0 0 net1
flabel metal1 229 478 229 478 0 FreeSans 80 0 0 0 net2
flabel ndiff 174 177 174 177 0 FreeSans 80 0 0 0 net3
flabel metal1 280 438 280 438 0 FreeSans 80 0 0 0 net4
flabel ndiff 326 174 326 174 0 FreeSans 80 0 0 0 net5
flabel metal1 378 281 378 281 0 FreeSans 80 0 0 0 net6
flabel metal1 298 764 298 764 0 FreeSans 80 0 0 0 vdd
port 10 nsew
flabel metal1 284 0 284 0 0 FreeSans 80 0 0 0 gnd
port 11 nsew
<< properties >>
string FIXED_BBOX 0 -21 602 769
<< end >>
