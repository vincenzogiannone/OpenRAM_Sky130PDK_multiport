magic
tech sky130A
magscale 1 2
timestamp 1643593061
<< checkpaint >>
rect -1296 -1277 2960 2155
<< nwell >>
rect -36 402 1700 895
<< pwell >>
rect 1554 51 1604 133
<< psubdiff >>
rect 1554 109 1604 133
rect 1554 75 1562 109
rect 1596 75 1604 109
rect 1554 51 1604 75
<< nsubdiff >>
rect 1554 763 1604 787
rect 1554 729 1562 763
rect 1596 729 1604 763
rect 1554 705 1604 729
<< psubdiffcont >>
rect 1562 75 1596 109
<< nsubdiffcont >>
rect 1562 729 1596 763
<< poly >>
rect 114 404 144 440
rect 48 388 144 404
rect 48 354 64 388
rect 98 354 144 388
rect 48 338 144 354
rect 114 204 144 338
<< polycont >>
rect 64 354 98 388
<< locali >>
rect 0 821 1664 855
rect 62 608 96 821
rect 274 608 308 821
rect 490 608 524 821
rect 706 608 740 821
rect 922 608 956 821
rect 1138 608 1172 821
rect 1354 608 1388 821
rect 1562 763 1596 821
rect 1562 713 1596 729
rect 48 388 114 404
rect 48 354 64 388
rect 98 354 114 388
rect 48 338 114 354
rect 812 388 846 574
rect 812 354 863 388
rect 812 167 846 354
rect 1562 109 1596 125
rect 62 17 96 67
rect 274 17 308 67
rect 490 17 524 67
rect 706 17 740 67
rect 922 17 956 67
rect 1138 17 1172 67
rect 1354 17 1388 67
rect 1562 17 1596 75
rect 0 -17 1664 17
use contact_12  contact_12_0
timestamp 1643593061
transform 1 0 48 0 1 338
box 0 0 1 1
use contact_11  contact_11_0
timestamp 1643593061
transform 1 0 1554 0 1 51
box 0 0 1 1
use contact_10  contact_10_0
timestamp 1643593061
transform 1 0 1554 0 1 705
box 0 0 1 1
use nmos_m13_w0_485_sli_dli_da_p  nmos_m13_w0_485_sli_dli_da_p_0
timestamp 1643593061
transform 1 0 54 0 1 51
box 0 -26 1446 153
use pmos_m13_w1_455_sli_dli_da_p  pmos_m13_w1_455_sli_dli_da_p_0
timestamp 1643593061
transform 1 0 54 0 1 496
box -59 -56 1505 345
<< labels >>
rlabel locali s 81 371 81 371 4 A
rlabel locali s 846 371 846 371 4 Z
rlabel locali s 832 0 832 0 4 gnd
rlabel locali s 832 838 832 838 4 vdd
<< properties >>
string FIXED_BBOX 0 0 1664 838
string GDS_FILE sram_0rw2r1w_2_16_sky130A.gds
string GDS_END 536556
string GDS_START 534296
<< end >>
