magic
tech sky130A
magscale 1 2
timestamp 1644951705
<< checkpaint >>
rect -1260 -1286 2382 1408
<< scnmos >>
rect 60 0 90 92
rect 168 0 198 92
rect 276 0 306 92
rect 384 0 414 92
rect 492 0 522 92
rect 600 0 630 92
rect 708 0 738 92
rect 816 0 846 92
rect 924 0 954 92
rect 1032 0 1062 92
<< ndiff >>
rect 0 63 60 92
rect 0 29 8 63
rect 42 29 60 63
rect 0 0 60 29
rect 90 63 168 92
rect 90 29 112 63
rect 146 29 168 63
rect 90 0 168 29
rect 198 63 276 92
rect 198 29 220 63
rect 254 29 276 63
rect 198 0 276 29
rect 306 63 384 92
rect 306 29 328 63
rect 362 29 384 63
rect 306 0 384 29
rect 414 63 492 92
rect 414 29 436 63
rect 470 29 492 63
rect 414 0 492 29
rect 522 63 600 92
rect 522 29 544 63
rect 578 29 600 63
rect 522 0 600 29
rect 630 63 708 92
rect 630 29 652 63
rect 686 29 708 63
rect 630 0 708 29
rect 738 63 816 92
rect 738 29 760 63
rect 794 29 816 63
rect 738 0 816 29
rect 846 63 924 92
rect 846 29 868 63
rect 902 29 924 63
rect 846 0 924 29
rect 954 63 1032 92
rect 954 29 976 63
rect 1010 29 1032 63
rect 954 0 1032 29
rect 1062 63 1122 92
rect 1062 29 1080 63
rect 1114 29 1122 63
rect 1062 0 1122 29
<< ndiffc >>
rect 8 29 42 63
rect 112 29 146 63
rect 220 29 254 63
rect 328 29 362 63
rect 436 29 470 63
rect 544 29 578 63
rect 652 29 686 63
rect 760 29 794 63
rect 868 29 902 63
rect 976 29 1010 63
rect 1080 29 1114 63
<< poly >>
rect 60 118 1062 148
rect 60 92 90 118
rect 168 92 198 118
rect 276 92 306 118
rect 384 92 414 118
rect 492 92 522 118
rect 600 92 630 118
rect 708 92 738 118
rect 816 92 846 118
rect 924 92 954 118
rect 1032 92 1062 118
rect 60 -26 90 0
rect 168 -26 198 0
rect 276 -26 306 0
rect 384 -26 414 0
rect 492 -26 522 0
rect 600 -26 630 0
rect 708 -26 738 0
rect 816 -26 846 0
rect 924 -26 954 0
rect 1032 -26 1062 0
<< locali >>
rect 112 113 1010 147
rect 8 63 42 79
rect 8 13 42 29
rect 112 63 146 113
rect 112 13 146 29
rect 220 63 254 79
rect 220 13 254 29
rect 328 63 362 113
rect 328 13 362 29
rect 436 63 470 79
rect 436 13 470 29
rect 544 63 578 113
rect 544 13 578 29
rect 652 63 686 79
rect 652 13 686 29
rect 760 63 794 113
rect 760 13 794 29
rect 868 63 902 79
rect 868 13 902 29
rect 976 63 1010 113
rect 976 13 1010 29
rect 1080 63 1114 79
rect 1080 13 1114 29
use contact_8  contact_8_0
timestamp 1644951705
transform 1 0 1072 0 1 5
box 0 0 1 1
use contact_8  contact_8_1
timestamp 1644951705
transform 1 0 968 0 1 5
box 0 0 1 1
use contact_8  contact_8_2
timestamp 1644951705
transform 1 0 860 0 1 5
box 0 0 1 1
use contact_8  contact_8_3
timestamp 1644951705
transform 1 0 752 0 1 5
box 0 0 1 1
use contact_8  contact_8_4
timestamp 1644951705
transform 1 0 644 0 1 5
box 0 0 1 1
use contact_8  contact_8_5
timestamp 1644951705
transform 1 0 536 0 1 5
box 0 0 1 1
use contact_8  contact_8_6
timestamp 1644951705
transform 1 0 428 0 1 5
box 0 0 1 1
use contact_8  contact_8_7
timestamp 1644951705
transform 1 0 320 0 1 5
box 0 0 1 1
use contact_8  contact_8_8
timestamp 1644951705
transform 1 0 212 0 1 5
box 0 0 1 1
use contact_8  contact_8_9
timestamp 1644951705
transform 1 0 104 0 1 5
box 0 0 1 1
use contact_8  contact_8_10
timestamp 1644951705
transform 1 0 0 0 1 5
box 0 0 1 1
<< labels >>
rlabel mvvaractor s 561 133 561 133 4 G
rlabel locali s 1097 46 1097 46 4 S
rlabel locali s 885 46 885 46 4 S
rlabel locali s 453 46 453 46 4 S
rlabel locali s 25 46 25 46 4 S
rlabel locali s 669 46 669 46 4 S
rlabel locali s 237 46 237 46 4 S
rlabel locali s 561 130 561 130 4 D
<< properties >>
string FIXED_BBOX -25 -26 1147 148
string GDS_FILE sram_0rw2r1w_16_128_sky130A.gds
string GDS_END 2040460
string GDS_START 2037840
<< end >>
