magic
tech sky130A
magscale 1 2
timestamp 1643678851
<< checkpaint >>
rect -1260 -1284 48638 2212
<< metal1 >>
rect 0 356 47378 384
<< via1 >>
rect 323 848 375 900
rect 3435 848 3487 900
rect 6547 848 6599 900
rect 9659 848 9711 900
rect 12771 848 12823 900
rect 15883 848 15935 900
rect 18995 848 19047 900
rect 22107 848 22159 900
rect 25219 848 25271 900
rect 28331 848 28383 900
rect 31443 848 31495 900
rect 34555 848 34607 900
rect 37667 848 37719 900
rect 40779 848 40831 900
rect 43891 848 43943 900
rect 47003 848 47055 900
rect 323 16 375 68
rect 3435 16 3487 68
rect 6547 16 6599 68
rect 9659 16 9711 68
rect 12771 16 12823 68
rect 15883 16 15935 68
rect 18995 16 19047 68
rect 22107 16 22159 68
rect 25219 16 25271 68
rect 28331 16 28383 68
rect 31443 16 31495 68
rect 34555 16 34607 68
rect 37667 16 37719 68
rect 40779 16 40831 68
rect 43891 16 43943 68
rect 47003 16 47055 68
<< metal2 >>
rect 329 902 369 908
rect 329 840 369 846
rect 630 322 658 952
rect 3441 902 3481 908
rect 3441 840 3481 846
rect 3742 322 3770 952
rect 6553 902 6593 908
rect 6553 840 6593 846
rect 6854 322 6882 952
rect 9665 902 9705 908
rect 9665 840 9705 846
rect 9966 322 9994 952
rect 12777 902 12817 908
rect 12777 840 12817 846
rect 13078 322 13106 952
rect 15889 902 15929 908
rect 15889 840 15929 846
rect 16190 322 16218 952
rect 19001 902 19041 908
rect 19001 840 19041 846
rect 19302 322 19330 952
rect 22113 902 22153 908
rect 22113 840 22153 846
rect 22414 322 22442 952
rect 25225 902 25265 908
rect 25225 840 25265 846
rect 25526 322 25554 952
rect 28337 902 28377 908
rect 28337 840 28377 846
rect 28638 322 28666 952
rect 31449 902 31489 908
rect 31449 840 31489 846
rect 31750 322 31778 952
rect 34561 902 34601 908
rect 34561 840 34601 846
rect 34862 322 34890 952
rect 37673 902 37713 908
rect 37673 840 37713 846
rect 37974 322 38002 952
rect 40785 902 40825 908
rect 40785 840 40825 846
rect 41086 322 41114 952
rect 43897 902 43937 908
rect 43897 840 43937 846
rect 44198 322 44226 952
rect 47009 902 47049 908
rect 47009 840 47049 846
rect 47310 322 47338 952
rect 196 272 250 300
rect 3308 272 3362 300
rect 6420 272 6474 300
rect 9532 272 9586 300
rect 12644 272 12698 300
rect 15756 272 15810 300
rect 18868 272 18922 300
rect 21980 272 22034 300
rect 25092 272 25146 300
rect 28204 272 28258 300
rect 31316 272 31370 300
rect 34428 272 34482 300
rect 37540 272 37594 300
rect 40652 272 40706 300
rect 43764 272 43818 300
rect 46876 272 46930 300
rect 329 70 369 76
rect 3441 70 3481 76
rect 6553 70 6593 76
rect 9665 70 9705 76
rect 12777 70 12817 76
rect 15889 70 15929 76
rect 19001 70 19041 76
rect 22113 70 22153 76
rect 25225 70 25265 76
rect 28337 70 28377 76
rect 31449 70 31489 76
rect 34561 70 34601 76
rect 37673 70 37713 76
rect 40785 70 40825 76
rect 43897 70 43937 76
rect 47009 70 47049 76
rect 329 8 369 14
rect 3441 8 3481 14
rect 6553 8 6593 14
rect 9665 8 9705 14
rect 12777 8 12817 14
rect 15889 8 15929 14
rect 19001 8 19041 14
rect 22113 8 22153 14
rect 25225 8 25265 14
rect 28337 8 28377 14
rect 31449 8 31489 14
rect 34561 8 34601 14
rect 37673 8 37713 14
rect 40785 8 40825 14
rect 43897 8 43937 14
rect 47009 8 47049 14
<< via2 >>
rect 321 900 377 902
rect 321 848 323 900
rect 323 848 375 900
rect 375 848 377 900
rect 321 846 377 848
rect 3433 900 3489 902
rect 3433 848 3435 900
rect 3435 848 3487 900
rect 3487 848 3489 900
rect 3433 846 3489 848
rect 6545 900 6601 902
rect 6545 848 6547 900
rect 6547 848 6599 900
rect 6599 848 6601 900
rect 6545 846 6601 848
rect 9657 900 9713 902
rect 9657 848 9659 900
rect 9659 848 9711 900
rect 9711 848 9713 900
rect 9657 846 9713 848
rect 12769 900 12825 902
rect 12769 848 12771 900
rect 12771 848 12823 900
rect 12823 848 12825 900
rect 12769 846 12825 848
rect 15881 900 15937 902
rect 15881 848 15883 900
rect 15883 848 15935 900
rect 15935 848 15937 900
rect 15881 846 15937 848
rect 18993 900 19049 902
rect 18993 848 18995 900
rect 18995 848 19047 900
rect 19047 848 19049 900
rect 18993 846 19049 848
rect 22105 900 22161 902
rect 22105 848 22107 900
rect 22107 848 22159 900
rect 22159 848 22161 900
rect 22105 846 22161 848
rect 25217 900 25273 902
rect 25217 848 25219 900
rect 25219 848 25271 900
rect 25271 848 25273 900
rect 25217 846 25273 848
rect 28329 900 28385 902
rect 28329 848 28331 900
rect 28331 848 28383 900
rect 28383 848 28385 900
rect 28329 846 28385 848
rect 31441 900 31497 902
rect 31441 848 31443 900
rect 31443 848 31495 900
rect 31495 848 31497 900
rect 31441 846 31497 848
rect 34553 900 34609 902
rect 34553 848 34555 900
rect 34555 848 34607 900
rect 34607 848 34609 900
rect 34553 846 34609 848
rect 37665 900 37721 902
rect 37665 848 37667 900
rect 37667 848 37719 900
rect 37719 848 37721 900
rect 37665 846 37721 848
rect 40777 900 40833 902
rect 40777 848 40779 900
rect 40779 848 40831 900
rect 40831 848 40833 900
rect 40777 846 40833 848
rect 43889 900 43945 902
rect 43889 848 43891 900
rect 43891 848 43943 900
rect 43943 848 43945 900
rect 43889 846 43945 848
rect 47001 900 47057 902
rect 47001 848 47003 900
rect 47003 848 47055 900
rect 47055 848 47057 900
rect 47001 846 47057 848
rect 321 68 377 70
rect 321 16 323 68
rect 323 16 375 68
rect 375 16 377 68
rect 321 14 377 16
rect 3433 68 3489 70
rect 3433 16 3435 68
rect 3435 16 3487 68
rect 3487 16 3489 68
rect 3433 14 3489 16
rect 6545 68 6601 70
rect 6545 16 6547 68
rect 6547 16 6599 68
rect 6599 16 6601 68
rect 6545 14 6601 16
rect 9657 68 9713 70
rect 9657 16 9659 68
rect 9659 16 9711 68
rect 9711 16 9713 68
rect 9657 14 9713 16
rect 12769 68 12825 70
rect 12769 16 12771 68
rect 12771 16 12823 68
rect 12823 16 12825 68
rect 12769 14 12825 16
rect 15881 68 15937 70
rect 15881 16 15883 68
rect 15883 16 15935 68
rect 15935 16 15937 68
rect 15881 14 15937 16
rect 18993 68 19049 70
rect 18993 16 18995 68
rect 18995 16 19047 68
rect 19047 16 19049 68
rect 18993 14 19049 16
rect 22105 68 22161 70
rect 22105 16 22107 68
rect 22107 16 22159 68
rect 22159 16 22161 68
rect 22105 14 22161 16
rect 25217 68 25273 70
rect 25217 16 25219 68
rect 25219 16 25271 68
rect 25271 16 25273 68
rect 25217 14 25273 16
rect 28329 68 28385 70
rect 28329 16 28331 68
rect 28331 16 28383 68
rect 28383 16 28385 68
rect 28329 14 28385 16
rect 31441 68 31497 70
rect 31441 16 31443 68
rect 31443 16 31495 68
rect 31495 16 31497 68
rect 31441 14 31497 16
rect 34553 68 34609 70
rect 34553 16 34555 68
rect 34555 16 34607 68
rect 34607 16 34609 68
rect 34553 14 34609 16
rect 37665 68 37721 70
rect 37665 16 37667 68
rect 37667 16 37719 68
rect 37719 16 37721 68
rect 37665 14 37721 16
rect 40777 68 40833 70
rect 40777 16 40779 68
rect 40779 16 40831 68
rect 40831 16 40833 68
rect 40777 14 40833 16
rect 43889 68 43945 70
rect 43889 16 43891 68
rect 43891 16 43943 68
rect 43943 16 43945 68
rect 43889 14 43945 16
rect 47001 68 47057 70
rect 47001 16 47003 68
rect 47003 16 47055 68
rect 47055 16 47057 68
rect 47001 14 47057 16
<< metal3 >>
rect 316 902 382 940
rect 316 846 321 902
rect 377 846 382 902
rect 316 808 382 846
rect 3428 902 3494 940
rect 3428 846 3433 902
rect 3489 846 3494 902
rect 3428 808 3494 846
rect 6540 902 6606 940
rect 6540 846 6545 902
rect 6601 846 6606 902
rect 6540 808 6606 846
rect 9652 902 9718 940
rect 9652 846 9657 902
rect 9713 846 9718 902
rect 9652 808 9718 846
rect 12764 902 12830 940
rect 12764 846 12769 902
rect 12825 846 12830 902
rect 12764 808 12830 846
rect 15876 902 15942 940
rect 15876 846 15881 902
rect 15937 846 15942 902
rect 15876 808 15942 846
rect 18988 902 19054 940
rect 18988 846 18993 902
rect 19049 846 19054 902
rect 18988 808 19054 846
rect 22100 902 22166 940
rect 22100 846 22105 902
rect 22161 846 22166 902
rect 22100 808 22166 846
rect 25212 902 25278 940
rect 25212 846 25217 902
rect 25273 846 25278 902
rect 25212 808 25278 846
rect 28324 902 28390 940
rect 28324 846 28329 902
rect 28385 846 28390 902
rect 28324 808 28390 846
rect 31436 902 31502 940
rect 31436 846 31441 902
rect 31497 846 31502 902
rect 31436 808 31502 846
rect 34548 902 34614 940
rect 34548 846 34553 902
rect 34609 846 34614 902
rect 34548 808 34614 846
rect 37660 902 37726 940
rect 37660 846 37665 902
rect 37721 846 37726 902
rect 37660 808 37726 846
rect 40772 902 40838 940
rect 40772 846 40777 902
rect 40833 846 40838 902
rect 40772 808 40838 846
rect 43884 902 43950 940
rect 43884 846 43889 902
rect 43945 846 43950 902
rect 43884 808 43950 846
rect 46996 902 47062 940
rect 46996 846 47001 902
rect 47057 846 47062 902
rect 46996 808 47062 846
rect 316 70 382 108
rect 316 14 321 70
rect 377 14 382 70
rect 316 -24 382 14
rect 3428 70 3494 108
rect 3428 14 3433 70
rect 3489 14 3494 70
rect 3428 -24 3494 14
rect 6540 70 6606 108
rect 6540 14 6545 70
rect 6601 14 6606 70
rect 6540 -24 6606 14
rect 9652 70 9718 108
rect 9652 14 9657 70
rect 9713 14 9718 70
rect 9652 -24 9718 14
rect 12764 70 12830 108
rect 12764 14 12769 70
rect 12825 14 12830 70
rect 12764 -24 12830 14
rect 15876 70 15942 108
rect 15876 14 15881 70
rect 15937 14 15942 70
rect 15876 -24 15942 14
rect 18988 70 19054 108
rect 18988 14 18993 70
rect 19049 14 19054 70
rect 18988 -24 19054 14
rect 22100 70 22166 108
rect 22100 14 22105 70
rect 22161 14 22166 70
rect 22100 -24 22166 14
rect 25212 70 25278 108
rect 25212 14 25217 70
rect 25273 14 25278 70
rect 25212 -24 25278 14
rect 28324 70 28390 108
rect 28324 14 28329 70
rect 28385 14 28390 70
rect 28324 -24 28390 14
rect 31436 70 31502 108
rect 31436 14 31441 70
rect 31497 14 31502 70
rect 31436 -24 31502 14
rect 34548 70 34614 108
rect 34548 14 34553 70
rect 34609 14 34614 70
rect 34548 -24 34614 14
rect 37660 70 37726 108
rect 37660 14 37665 70
rect 37721 14 37726 70
rect 37660 -24 37726 14
rect 40772 70 40838 108
rect 40772 14 40777 70
rect 40833 14 40838 70
rect 40772 -24 40838 14
rect 43884 70 43950 108
rect 43884 14 43889 70
rect 43945 14 43950 70
rect 43884 -24 43950 14
rect 46996 70 47062 108
rect 46996 14 47001 70
rect 47057 14 47062 70
rect 46996 -24 47062 14
use contact_23  contact_23_0
timestamp 1643678851
transform 1 0 46996 0 1 -24
box 0 0 1 1
use contact_22  contact_22_0
timestamp 1643678851
transform 1 0 47014 0 1 27
box 0 0 1 1
use contact_23  contact_23_1
timestamp 1643678851
transform 1 0 46996 0 1 808
box 0 0 1 1
use contact_22  contact_22_1
timestamp 1643678851
transform 1 0 47014 0 1 859
box 0 0 1 1
use contact_23  contact_23_2
timestamp 1643678851
transform 1 0 43884 0 1 -24
box 0 0 1 1
use contact_22  contact_22_2
timestamp 1643678851
transform 1 0 43902 0 1 27
box 0 0 1 1
use contact_23  contact_23_3
timestamp 1643678851
transform 1 0 43884 0 1 808
box 0 0 1 1
use contact_22  contact_22_3
timestamp 1643678851
transform 1 0 43902 0 1 859
box 0 0 1 1
use contact_23  contact_23_4
timestamp 1643678851
transform 1 0 40772 0 1 -24
box 0 0 1 1
use contact_22  contact_22_4
timestamp 1643678851
transform 1 0 40790 0 1 27
box 0 0 1 1
use contact_23  contact_23_5
timestamp 1643678851
transform 1 0 40772 0 1 808
box 0 0 1 1
use contact_22  contact_22_5
timestamp 1643678851
transform 1 0 40790 0 1 859
box 0 0 1 1
use contact_23  contact_23_6
timestamp 1643678851
transform 1 0 37660 0 1 -24
box 0 0 1 1
use contact_22  contact_22_6
timestamp 1643678851
transform 1 0 37678 0 1 27
box 0 0 1 1
use contact_23  contact_23_7
timestamp 1643678851
transform 1 0 37660 0 1 808
box 0 0 1 1
use contact_22  contact_22_7
timestamp 1643678851
transform 1 0 37678 0 1 859
box 0 0 1 1
use contact_23  contact_23_8
timestamp 1643678851
transform 1 0 34548 0 1 -24
box 0 0 1 1
use contact_22  contact_22_8
timestamp 1643678851
transform 1 0 34566 0 1 27
box 0 0 1 1
use contact_23  contact_23_9
timestamp 1643678851
transform 1 0 34548 0 1 808
box 0 0 1 1
use contact_22  contact_22_9
timestamp 1643678851
transform 1 0 34566 0 1 859
box 0 0 1 1
use contact_23  contact_23_10
timestamp 1643678851
transform 1 0 31436 0 1 -24
box 0 0 1 1
use contact_22  contact_22_10
timestamp 1643678851
transform 1 0 31454 0 1 27
box 0 0 1 1
use contact_23  contact_23_11
timestamp 1643678851
transform 1 0 31436 0 1 808
box 0 0 1 1
use contact_22  contact_22_11
timestamp 1643678851
transform 1 0 31454 0 1 859
box 0 0 1 1
use contact_23  contact_23_12
timestamp 1643678851
transform 1 0 28324 0 1 -24
box 0 0 1 1
use contact_22  contact_22_12
timestamp 1643678851
transform 1 0 28342 0 1 27
box 0 0 1 1
use contact_23  contact_23_13
timestamp 1643678851
transform 1 0 28324 0 1 808
box 0 0 1 1
use contact_22  contact_22_13
timestamp 1643678851
transform 1 0 28342 0 1 859
box 0 0 1 1
use contact_23  contact_23_14
timestamp 1643678851
transform 1 0 25212 0 1 -24
box 0 0 1 1
use contact_22  contact_22_14
timestamp 1643678851
transform 1 0 25230 0 1 27
box 0 0 1 1
use contact_23  contact_23_15
timestamp 1643678851
transform 1 0 25212 0 1 808
box 0 0 1 1
use contact_22  contact_22_15
timestamp 1643678851
transform 1 0 25230 0 1 859
box 0 0 1 1
use contact_23  contact_23_16
timestamp 1643678851
transform 1 0 22100 0 1 -24
box 0 0 1 1
use contact_22  contact_22_16
timestamp 1643678851
transform 1 0 22118 0 1 27
box 0 0 1 1
use contact_23  contact_23_17
timestamp 1643678851
transform 1 0 22100 0 1 808
box 0 0 1 1
use contact_22  contact_22_17
timestamp 1643678851
transform 1 0 22118 0 1 859
box 0 0 1 1
use contact_23  contact_23_18
timestamp 1643678851
transform 1 0 18988 0 1 -24
box 0 0 1 1
use contact_22  contact_22_18
timestamp 1643678851
transform 1 0 19006 0 1 27
box 0 0 1 1
use contact_23  contact_23_19
timestamp 1643678851
transform 1 0 18988 0 1 808
box 0 0 1 1
use contact_22  contact_22_19
timestamp 1643678851
transform 1 0 19006 0 1 859
box 0 0 1 1
use contact_23  contact_23_20
timestamp 1643678851
transform 1 0 15876 0 1 -24
box 0 0 1 1
use contact_22  contact_22_20
timestamp 1643678851
transform 1 0 15894 0 1 27
box 0 0 1 1
use contact_23  contact_23_21
timestamp 1643678851
transform 1 0 15876 0 1 808
box 0 0 1 1
use contact_22  contact_22_21
timestamp 1643678851
transform 1 0 15894 0 1 859
box 0 0 1 1
use contact_23  contact_23_22
timestamp 1643678851
transform 1 0 12764 0 1 -24
box 0 0 1 1
use contact_22  contact_22_22
timestamp 1643678851
transform 1 0 12782 0 1 27
box 0 0 1 1
use contact_23  contact_23_23
timestamp 1643678851
transform 1 0 12764 0 1 808
box 0 0 1 1
use contact_22  contact_22_23
timestamp 1643678851
transform 1 0 12782 0 1 859
box 0 0 1 1
use contact_23  contact_23_24
timestamp 1643678851
transform 1 0 9652 0 1 -24
box 0 0 1 1
use contact_22  contact_22_24
timestamp 1643678851
transform 1 0 9670 0 1 27
box 0 0 1 1
use contact_23  contact_23_25
timestamp 1643678851
transform 1 0 9652 0 1 808
box 0 0 1 1
use contact_22  contact_22_25
timestamp 1643678851
transform 1 0 9670 0 1 859
box 0 0 1 1
use contact_23  contact_23_26
timestamp 1643678851
transform 1 0 6540 0 1 -24
box 0 0 1 1
use contact_22  contact_22_26
timestamp 1643678851
transform 1 0 6558 0 1 27
box 0 0 1 1
use contact_23  contact_23_27
timestamp 1643678851
transform 1 0 6540 0 1 808
box 0 0 1 1
use contact_22  contact_22_27
timestamp 1643678851
transform 1 0 6558 0 1 859
box 0 0 1 1
use contact_23  contact_23_28
timestamp 1643678851
transform 1 0 3428 0 1 -24
box 0 0 1 1
use contact_22  contact_22_28
timestamp 1643678851
transform 1 0 3446 0 1 27
box 0 0 1 1
use contact_23  contact_23_29
timestamp 1643678851
transform 1 0 3428 0 1 808
box 0 0 1 1
use contact_22  contact_22_29
timestamp 1643678851
transform 1 0 3446 0 1 859
box 0 0 1 1
use contact_23  contact_23_30
timestamp 1643678851
transform 1 0 316 0 1 -24
box 0 0 1 1
use contact_22  contact_22_30
timestamp 1643678851
transform 1 0 334 0 1 27
box 0 0 1 1
use contact_23  contact_23_31
timestamp 1643678851
transform 1 0 316 0 1 808
box 0 0 1 1
use contact_22  contact_22_31
timestamp 1643678851
transform 1 0 334 0 1 859
box 0 0 1 1
use write_driver_multiport  write_driver_multiport_0
timestamp 1643678851
transform 1 0 46680 0 1 0
box 0 0 698 952
use write_driver_multiport  write_driver_multiport_1
timestamp 1643678851
transform 1 0 43568 0 1 0
box 0 0 698 952
use write_driver_multiport  write_driver_multiport_2
timestamp 1643678851
transform 1 0 40456 0 1 0
box 0 0 698 952
use write_driver_multiport  write_driver_multiport_3
timestamp 1643678851
transform 1 0 37344 0 1 0
box 0 0 698 952
use write_driver_multiport  write_driver_multiport_4
timestamp 1643678851
transform 1 0 34232 0 1 0
box 0 0 698 952
use write_driver_multiport  write_driver_multiport_5
timestamp 1643678851
transform 1 0 31120 0 1 0
box 0 0 698 952
use write_driver_multiport  write_driver_multiport_6
timestamp 1643678851
transform 1 0 28008 0 1 0
box 0 0 698 952
use write_driver_multiport  write_driver_multiport_7
timestamp 1643678851
transform 1 0 24896 0 1 0
box 0 0 698 952
use write_driver_multiport  write_driver_multiport_8
timestamp 1643678851
transform 1 0 21784 0 1 0
box 0 0 698 952
use write_driver_multiport  write_driver_multiport_9
timestamp 1643678851
transform 1 0 18672 0 1 0
box 0 0 698 952
use write_driver_multiport  write_driver_multiport_10
timestamp 1643678851
transform 1 0 15560 0 1 0
box 0 0 698 952
use write_driver_multiport  write_driver_multiport_11
timestamp 1643678851
transform 1 0 12448 0 1 0
box 0 0 698 952
use write_driver_multiport  write_driver_multiport_12
timestamp 1643678851
transform 1 0 9336 0 1 0
box 0 0 698 952
use write_driver_multiport  write_driver_multiport_13
timestamp 1643678851
transform 1 0 6224 0 1 0
box 0 0 698 952
use write_driver_multiport  write_driver_multiport_14
timestamp 1643678851
transform 1 0 3112 0 1 0
box 0 0 698 952
use write_driver_multiport  write_driver_multiport_15
timestamp 1643678851
transform 1 0 0 0 1 0
box 0 0 698 952
<< labels >>
rlabel metal2 s 196 272 250 300 4 din_0
rlabel metal2 s 630 322 658 952 4 wbl0_0
rlabel metal3 s 25212 808 25278 940 4 vdd
rlabel metal3 s 37660 808 37726 940 4 vdd
rlabel metal3 s 46996 808 47062 940 4 vdd
rlabel metal3 s 18988 808 19054 940 4 vdd
rlabel metal3 s 3428 808 3494 940 4 vdd
rlabel metal3 s 12764 808 12830 940 4 vdd
rlabel metal3 s 43884 808 43950 940 4 vdd
rlabel metal3 s 9652 808 9718 940 4 vdd
rlabel metal3 s 40772 808 40838 940 4 vdd
rlabel metal3 s 34548 808 34614 940 4 vdd
rlabel metal3 s 28324 808 28390 940 4 vdd
rlabel metal3 s 31436 808 31502 940 4 vdd
rlabel metal3 s 316 808 382 940 4 vdd
rlabel metal3 s 6540 808 6606 940 4 vdd
rlabel metal3 s 15876 808 15942 940 4 vdd
rlabel metal3 s 22100 808 22166 940 4 vdd
rlabel metal3 s 6540 -24 6606 108 4 gnd
rlabel metal3 s 40772 -24 40838 108 4 gnd
rlabel metal3 s 46996 -24 47062 108 4 gnd
rlabel metal3 s 28324 -24 28390 108 4 gnd
rlabel metal3 s 34548 -24 34614 108 4 gnd
rlabel metal3 s 43884 -24 43950 108 4 gnd
rlabel metal3 s 15876 -24 15942 108 4 gnd
rlabel metal3 s 37660 -24 37726 108 4 gnd
rlabel metal3 s 25212 -24 25278 108 4 gnd
rlabel metal3 s 12764 -24 12830 108 4 gnd
rlabel metal3 s 31436 -24 31502 108 4 gnd
rlabel metal3 s 9652 -24 9718 108 4 gnd
rlabel metal3 s 22100 -24 22166 108 4 gnd
rlabel metal3 s 18988 -24 19054 108 4 gnd
rlabel metal3 s 316 -24 382 108 4 gnd
rlabel metal3 s 3428 -24 3494 108 4 gnd
rlabel metal2 s 3308 272 3362 300 4 din_1
rlabel metal2 s 3742 322 3770 952 4 wbl0_1
rlabel metal2 s 6420 272 6474 300 4 din_2
rlabel metal2 s 6854 322 6882 952 4 wbl0_2
rlabel metal2 s 9532 272 9586 300 4 din_3
rlabel metal2 s 9966 322 9994 952 4 wbl0_3
rlabel metal2 s 12644 272 12698 300 4 din_4
rlabel metal2 s 13078 322 13106 952 4 wbl0_4
rlabel metal2 s 15756 272 15810 300 4 din_5
rlabel metal2 s 16190 322 16218 952 4 wbl0_5
rlabel metal2 s 18868 272 18922 300 4 din_6
rlabel metal2 s 19302 322 19330 952 4 wbl0_6
rlabel metal2 s 21980 272 22034 300 4 din_7
rlabel metal2 s 22414 322 22442 952 4 wbl0_7
rlabel metal2 s 25092 272 25146 300 4 din_8
rlabel metal2 s 25526 322 25554 952 4 wbl0_8
rlabel metal2 s 28204 272 28258 300 4 din_9
rlabel metal2 s 28638 322 28666 952 4 wbl0_9
rlabel metal2 s 31316 272 31370 300 4 din_10
rlabel metal2 s 31750 322 31778 952 4 wbl0_10
rlabel metal2 s 34428 272 34482 300 4 din_11
rlabel metal2 s 34862 322 34890 952 4 wbl0_11
rlabel metal2 s 37540 272 37594 300 4 din_12
rlabel metal2 s 37974 322 38002 952 4 wbl0_12
rlabel metal2 s 40652 272 40706 300 4 din_13
rlabel metal2 s 41086 322 41114 952 4 wbl0_13
rlabel metal2 s 43764 272 43818 300 4 din_14
rlabel metal2 s 44198 322 44226 952 4 wbl0_14
rlabel metal2 s 46876 272 46930 300 4 din_15
rlabel metal2 s 47310 322 47338 952 4 wbl0_15
rlabel metal1 s 0 356 47378 384 4 en
<< properties >>
string FIXED_BBOX 46996 -24 47062 0
string GDS_FILE sram_0rw2r1w_16_128_sky130A.gds
string GDS_END 1543614
string GDS_START 1525878
<< end >>
