magic
tech sky130A
magscale 1 2
timestamp 1643678851
<< checkpaint >>
rect -1260 -1228 51118 3174
<< poly >>
rect 374 221 404 434
rect 1152 279 1182 434
rect 1930 337 1960 434
rect 2708 395 2738 434
rect 2690 379 2756 395
rect 2690 345 2706 379
rect 2740 345 2756 379
rect 1912 321 1978 337
rect 2690 329 2756 345
rect 1912 287 1928 321
rect 1962 287 1978 321
rect 1134 263 1200 279
rect 1912 271 1978 287
rect 1134 229 1150 263
rect 1184 229 1200 263
rect 356 205 422 221
rect 1134 213 1200 229
rect 3486 221 3516 434
rect 4264 279 4294 434
rect 5042 337 5072 434
rect 5820 395 5850 434
rect 5802 379 5868 395
rect 5802 345 5818 379
rect 5852 345 5868 379
rect 5024 321 5090 337
rect 5802 329 5868 345
rect 5024 287 5040 321
rect 5074 287 5090 321
rect 4246 263 4312 279
rect 5024 271 5090 287
rect 4246 229 4262 263
rect 4296 229 4312 263
rect 356 171 372 205
rect 406 171 422 205
rect 356 155 422 171
rect 3468 205 3534 221
rect 4246 213 4312 229
rect 6598 221 6628 434
rect 7376 279 7406 434
rect 8154 337 8184 434
rect 8932 395 8962 434
rect 8914 379 8980 395
rect 8914 345 8930 379
rect 8964 345 8980 379
rect 8136 321 8202 337
rect 8914 329 8980 345
rect 8136 287 8152 321
rect 8186 287 8202 321
rect 7358 263 7424 279
rect 8136 271 8202 287
rect 7358 229 7374 263
rect 7408 229 7424 263
rect 3468 171 3484 205
rect 3518 171 3534 205
rect 3468 155 3534 171
rect 6580 205 6646 221
rect 7358 213 7424 229
rect 9710 221 9740 434
rect 10488 279 10518 434
rect 11266 337 11296 434
rect 12044 395 12074 434
rect 12026 379 12092 395
rect 12026 345 12042 379
rect 12076 345 12092 379
rect 11248 321 11314 337
rect 12026 329 12092 345
rect 11248 287 11264 321
rect 11298 287 11314 321
rect 10470 263 10536 279
rect 11248 271 11314 287
rect 10470 229 10486 263
rect 10520 229 10536 263
rect 6580 171 6596 205
rect 6630 171 6646 205
rect 6580 155 6646 171
rect 9692 205 9758 221
rect 10470 213 10536 229
rect 12822 221 12852 434
rect 13600 279 13630 434
rect 14378 337 14408 434
rect 15156 395 15186 434
rect 15138 379 15204 395
rect 15138 345 15154 379
rect 15188 345 15204 379
rect 14360 321 14426 337
rect 15138 329 15204 345
rect 14360 287 14376 321
rect 14410 287 14426 321
rect 13582 263 13648 279
rect 14360 271 14426 287
rect 13582 229 13598 263
rect 13632 229 13648 263
rect 9692 171 9708 205
rect 9742 171 9758 205
rect 9692 155 9758 171
rect 12804 205 12870 221
rect 13582 213 13648 229
rect 15934 221 15964 434
rect 16712 279 16742 434
rect 17490 337 17520 434
rect 18268 395 18298 434
rect 18250 379 18316 395
rect 18250 345 18266 379
rect 18300 345 18316 379
rect 17472 321 17538 337
rect 18250 329 18316 345
rect 17472 287 17488 321
rect 17522 287 17538 321
rect 16694 263 16760 279
rect 17472 271 17538 287
rect 16694 229 16710 263
rect 16744 229 16760 263
rect 12804 171 12820 205
rect 12854 171 12870 205
rect 12804 155 12870 171
rect 15916 205 15982 221
rect 16694 213 16760 229
rect 19046 221 19076 434
rect 19824 279 19854 434
rect 20602 337 20632 434
rect 21380 395 21410 434
rect 21362 379 21428 395
rect 21362 345 21378 379
rect 21412 345 21428 379
rect 20584 321 20650 337
rect 21362 329 21428 345
rect 20584 287 20600 321
rect 20634 287 20650 321
rect 19806 263 19872 279
rect 20584 271 20650 287
rect 19806 229 19822 263
rect 19856 229 19872 263
rect 15916 171 15932 205
rect 15966 171 15982 205
rect 15916 155 15982 171
rect 19028 205 19094 221
rect 19806 213 19872 229
rect 22158 221 22188 434
rect 22936 279 22966 434
rect 23714 337 23744 434
rect 24492 395 24522 434
rect 24474 379 24540 395
rect 24474 345 24490 379
rect 24524 345 24540 379
rect 23696 321 23762 337
rect 24474 329 24540 345
rect 23696 287 23712 321
rect 23746 287 23762 321
rect 22918 263 22984 279
rect 23696 271 23762 287
rect 22918 229 22934 263
rect 22968 229 22984 263
rect 19028 171 19044 205
rect 19078 171 19094 205
rect 19028 155 19094 171
rect 22140 205 22206 221
rect 22918 213 22984 229
rect 25270 221 25300 434
rect 26048 279 26078 434
rect 26826 337 26856 434
rect 27604 395 27634 434
rect 27586 379 27652 395
rect 27586 345 27602 379
rect 27636 345 27652 379
rect 26808 321 26874 337
rect 27586 329 27652 345
rect 26808 287 26824 321
rect 26858 287 26874 321
rect 26030 263 26096 279
rect 26808 271 26874 287
rect 26030 229 26046 263
rect 26080 229 26096 263
rect 22140 171 22156 205
rect 22190 171 22206 205
rect 22140 155 22206 171
rect 25252 205 25318 221
rect 26030 213 26096 229
rect 28382 221 28412 434
rect 29160 279 29190 434
rect 29938 337 29968 434
rect 30716 395 30746 434
rect 30698 379 30764 395
rect 30698 345 30714 379
rect 30748 345 30764 379
rect 29920 321 29986 337
rect 30698 329 30764 345
rect 29920 287 29936 321
rect 29970 287 29986 321
rect 29142 263 29208 279
rect 29920 271 29986 287
rect 29142 229 29158 263
rect 29192 229 29208 263
rect 25252 171 25268 205
rect 25302 171 25318 205
rect 25252 155 25318 171
rect 28364 205 28430 221
rect 29142 213 29208 229
rect 31494 221 31524 434
rect 32272 279 32302 434
rect 33050 337 33080 434
rect 33828 395 33858 434
rect 33810 379 33876 395
rect 33810 345 33826 379
rect 33860 345 33876 379
rect 33032 321 33098 337
rect 33810 329 33876 345
rect 33032 287 33048 321
rect 33082 287 33098 321
rect 32254 263 32320 279
rect 33032 271 33098 287
rect 32254 229 32270 263
rect 32304 229 32320 263
rect 28364 171 28380 205
rect 28414 171 28430 205
rect 28364 155 28430 171
rect 31476 205 31542 221
rect 32254 213 32320 229
rect 34606 221 34636 434
rect 35384 279 35414 434
rect 36162 337 36192 434
rect 36940 395 36970 434
rect 36922 379 36988 395
rect 36922 345 36938 379
rect 36972 345 36988 379
rect 36144 321 36210 337
rect 36922 329 36988 345
rect 36144 287 36160 321
rect 36194 287 36210 321
rect 35366 263 35432 279
rect 36144 271 36210 287
rect 35366 229 35382 263
rect 35416 229 35432 263
rect 31476 171 31492 205
rect 31526 171 31542 205
rect 31476 155 31542 171
rect 34588 205 34654 221
rect 35366 213 35432 229
rect 37718 221 37748 434
rect 38496 279 38526 434
rect 39274 337 39304 434
rect 40052 395 40082 434
rect 40034 379 40100 395
rect 40034 345 40050 379
rect 40084 345 40100 379
rect 39256 321 39322 337
rect 40034 329 40100 345
rect 39256 287 39272 321
rect 39306 287 39322 321
rect 38478 263 38544 279
rect 39256 271 39322 287
rect 38478 229 38494 263
rect 38528 229 38544 263
rect 34588 171 34604 205
rect 34638 171 34654 205
rect 34588 155 34654 171
rect 37700 205 37766 221
rect 38478 213 38544 229
rect 40830 221 40860 434
rect 41608 279 41638 434
rect 42386 337 42416 434
rect 43164 395 43194 434
rect 43146 379 43212 395
rect 43146 345 43162 379
rect 43196 345 43212 379
rect 42368 321 42434 337
rect 43146 329 43212 345
rect 42368 287 42384 321
rect 42418 287 42434 321
rect 41590 263 41656 279
rect 42368 271 42434 287
rect 41590 229 41606 263
rect 41640 229 41656 263
rect 37700 171 37716 205
rect 37750 171 37766 205
rect 37700 155 37766 171
rect 40812 205 40878 221
rect 41590 213 41656 229
rect 43942 221 43972 434
rect 44720 279 44750 434
rect 45498 337 45528 434
rect 46276 395 46306 434
rect 46258 379 46324 395
rect 46258 345 46274 379
rect 46308 345 46324 379
rect 45480 321 45546 337
rect 46258 329 46324 345
rect 45480 287 45496 321
rect 45530 287 45546 321
rect 44702 263 44768 279
rect 45480 271 45546 287
rect 44702 229 44718 263
rect 44752 229 44768 263
rect 40812 171 40828 205
rect 40862 171 40878 205
rect 40812 155 40878 171
rect 43924 205 43990 221
rect 44702 213 44768 229
rect 47054 221 47084 434
rect 47832 279 47862 434
rect 48610 337 48640 434
rect 49388 395 49418 434
rect 49370 379 49436 395
rect 49370 345 49386 379
rect 49420 345 49436 379
rect 48592 321 48658 337
rect 49370 329 49436 345
rect 48592 287 48608 321
rect 48642 287 48658 321
rect 47814 263 47880 279
rect 48592 271 48658 287
rect 47814 229 47830 263
rect 47864 229 47880 263
rect 43924 171 43940 205
rect 43974 171 43990 205
rect 43924 155 43990 171
rect 47036 205 47102 221
rect 47814 213 47880 229
rect 47036 171 47052 205
rect 47086 171 47102 205
rect 47036 155 47102 171
<< polycont >>
rect 2706 345 2740 379
rect 1928 287 1962 321
rect 1150 229 1184 263
rect 5818 345 5852 379
rect 5040 287 5074 321
rect 4262 229 4296 263
rect 372 171 406 205
rect 8930 345 8964 379
rect 8152 287 8186 321
rect 7374 229 7408 263
rect 3484 171 3518 205
rect 12042 345 12076 379
rect 11264 287 11298 321
rect 10486 229 10520 263
rect 6596 171 6630 205
rect 15154 345 15188 379
rect 14376 287 14410 321
rect 13598 229 13632 263
rect 9708 171 9742 205
rect 18266 345 18300 379
rect 17488 287 17522 321
rect 16710 229 16744 263
rect 12820 171 12854 205
rect 21378 345 21412 379
rect 20600 287 20634 321
rect 19822 229 19856 263
rect 15932 171 15966 205
rect 24490 345 24524 379
rect 23712 287 23746 321
rect 22934 229 22968 263
rect 19044 171 19078 205
rect 27602 345 27636 379
rect 26824 287 26858 321
rect 26046 229 26080 263
rect 22156 171 22190 205
rect 30714 345 30748 379
rect 29936 287 29970 321
rect 29158 229 29192 263
rect 25268 171 25302 205
rect 33826 345 33860 379
rect 33048 287 33082 321
rect 32270 229 32304 263
rect 28380 171 28414 205
rect 36938 345 36972 379
rect 36160 287 36194 321
rect 35382 229 35416 263
rect 31492 171 31526 205
rect 40050 345 40084 379
rect 39272 287 39306 321
rect 38494 229 38528 263
rect 34604 171 34638 205
rect 43162 345 43196 379
rect 42384 287 42418 321
rect 41606 229 41640 263
rect 37716 171 37750 205
rect 46274 345 46308 379
rect 45496 287 45530 321
rect 44718 229 44752 263
rect 40828 171 40862 205
rect 49386 345 49420 379
rect 48608 287 48642 321
rect 47830 229 47864 263
rect 43940 171 43974 205
rect 47052 171 47086 205
<< locali >>
rect 2690 379 2756 395
rect 2690 345 2706 379
rect 2740 345 2756 379
rect 1912 321 1978 337
rect 2690 329 2756 345
rect 5802 379 5868 395
rect 5802 345 5818 379
rect 5852 345 5868 379
rect 1912 287 1928 321
rect 1962 287 1978 321
rect 1134 263 1200 279
rect 1912 271 1978 287
rect 5024 321 5090 337
rect 5802 329 5868 345
rect 8914 379 8980 395
rect 8914 345 8930 379
rect 8964 345 8980 379
rect 5024 287 5040 321
rect 5074 287 5090 321
rect 1134 229 1150 263
rect 1184 229 1200 263
rect 356 205 422 221
rect 1134 213 1200 229
rect 4246 263 4312 279
rect 5024 271 5090 287
rect 8136 321 8202 337
rect 8914 329 8980 345
rect 12026 379 12092 395
rect 12026 345 12042 379
rect 12076 345 12092 379
rect 8136 287 8152 321
rect 8186 287 8202 321
rect 4246 229 4262 263
rect 4296 229 4312 263
rect 356 171 372 205
rect 406 171 422 205
rect 356 155 422 171
rect 3468 205 3534 221
rect 4246 213 4312 229
rect 7358 263 7424 279
rect 8136 271 8202 287
rect 11248 321 11314 337
rect 12026 329 12092 345
rect 15138 379 15204 395
rect 15138 345 15154 379
rect 15188 345 15204 379
rect 11248 287 11264 321
rect 11298 287 11314 321
rect 7358 229 7374 263
rect 7408 229 7424 263
rect 3468 171 3484 205
rect 3518 171 3534 205
rect 3468 155 3534 171
rect 6580 205 6646 221
rect 7358 213 7424 229
rect 10470 263 10536 279
rect 11248 271 11314 287
rect 14360 321 14426 337
rect 15138 329 15204 345
rect 18250 379 18316 395
rect 18250 345 18266 379
rect 18300 345 18316 379
rect 14360 287 14376 321
rect 14410 287 14426 321
rect 10470 229 10486 263
rect 10520 229 10536 263
rect 6580 171 6596 205
rect 6630 171 6646 205
rect 6580 155 6646 171
rect 9692 205 9758 221
rect 10470 213 10536 229
rect 13582 263 13648 279
rect 14360 271 14426 287
rect 17472 321 17538 337
rect 18250 329 18316 345
rect 21362 379 21428 395
rect 21362 345 21378 379
rect 21412 345 21428 379
rect 17472 287 17488 321
rect 17522 287 17538 321
rect 13582 229 13598 263
rect 13632 229 13648 263
rect 9692 171 9708 205
rect 9742 171 9758 205
rect 9692 155 9758 171
rect 12804 205 12870 221
rect 13582 213 13648 229
rect 16694 263 16760 279
rect 17472 271 17538 287
rect 20584 321 20650 337
rect 21362 329 21428 345
rect 24474 379 24540 395
rect 24474 345 24490 379
rect 24524 345 24540 379
rect 20584 287 20600 321
rect 20634 287 20650 321
rect 16694 229 16710 263
rect 16744 229 16760 263
rect 12804 171 12820 205
rect 12854 171 12870 205
rect 12804 155 12870 171
rect 15916 205 15982 221
rect 16694 213 16760 229
rect 19806 263 19872 279
rect 20584 271 20650 287
rect 23696 321 23762 337
rect 24474 329 24540 345
rect 27586 379 27652 395
rect 27586 345 27602 379
rect 27636 345 27652 379
rect 23696 287 23712 321
rect 23746 287 23762 321
rect 19806 229 19822 263
rect 19856 229 19872 263
rect 15916 171 15932 205
rect 15966 171 15982 205
rect 15916 155 15982 171
rect 19028 205 19094 221
rect 19806 213 19872 229
rect 22918 263 22984 279
rect 23696 271 23762 287
rect 26808 321 26874 337
rect 27586 329 27652 345
rect 30698 379 30764 395
rect 30698 345 30714 379
rect 30748 345 30764 379
rect 26808 287 26824 321
rect 26858 287 26874 321
rect 22918 229 22934 263
rect 22968 229 22984 263
rect 19028 171 19044 205
rect 19078 171 19094 205
rect 19028 155 19094 171
rect 22140 205 22206 221
rect 22918 213 22984 229
rect 26030 263 26096 279
rect 26808 271 26874 287
rect 29920 321 29986 337
rect 30698 329 30764 345
rect 33810 379 33876 395
rect 33810 345 33826 379
rect 33860 345 33876 379
rect 29920 287 29936 321
rect 29970 287 29986 321
rect 26030 229 26046 263
rect 26080 229 26096 263
rect 22140 171 22156 205
rect 22190 171 22206 205
rect 22140 155 22206 171
rect 25252 205 25318 221
rect 26030 213 26096 229
rect 29142 263 29208 279
rect 29920 271 29986 287
rect 33032 321 33098 337
rect 33810 329 33876 345
rect 36922 379 36988 395
rect 36922 345 36938 379
rect 36972 345 36988 379
rect 33032 287 33048 321
rect 33082 287 33098 321
rect 29142 229 29158 263
rect 29192 229 29208 263
rect 25252 171 25268 205
rect 25302 171 25318 205
rect 25252 155 25318 171
rect 28364 205 28430 221
rect 29142 213 29208 229
rect 32254 263 32320 279
rect 33032 271 33098 287
rect 36144 321 36210 337
rect 36922 329 36988 345
rect 40034 379 40100 395
rect 40034 345 40050 379
rect 40084 345 40100 379
rect 36144 287 36160 321
rect 36194 287 36210 321
rect 32254 229 32270 263
rect 32304 229 32320 263
rect 28364 171 28380 205
rect 28414 171 28430 205
rect 28364 155 28430 171
rect 31476 205 31542 221
rect 32254 213 32320 229
rect 35366 263 35432 279
rect 36144 271 36210 287
rect 39256 321 39322 337
rect 40034 329 40100 345
rect 43146 379 43212 395
rect 43146 345 43162 379
rect 43196 345 43212 379
rect 39256 287 39272 321
rect 39306 287 39322 321
rect 35366 229 35382 263
rect 35416 229 35432 263
rect 31476 171 31492 205
rect 31526 171 31542 205
rect 31476 155 31542 171
rect 34588 205 34654 221
rect 35366 213 35432 229
rect 38478 263 38544 279
rect 39256 271 39322 287
rect 42368 321 42434 337
rect 43146 329 43212 345
rect 46258 379 46324 395
rect 46258 345 46274 379
rect 46308 345 46324 379
rect 42368 287 42384 321
rect 42418 287 42434 321
rect 38478 229 38494 263
rect 38528 229 38544 263
rect 34588 171 34604 205
rect 34638 171 34654 205
rect 34588 155 34654 171
rect 37700 205 37766 221
rect 38478 213 38544 229
rect 41590 263 41656 279
rect 42368 271 42434 287
rect 45480 321 45546 337
rect 46258 329 46324 345
rect 49370 379 49436 395
rect 49370 345 49386 379
rect 49420 345 49436 379
rect 45480 287 45496 321
rect 45530 287 45546 321
rect 41590 229 41606 263
rect 41640 229 41656 263
rect 37700 171 37716 205
rect 37750 171 37766 205
rect 37700 155 37766 171
rect 40812 205 40878 221
rect 41590 213 41656 229
rect 44702 263 44768 279
rect 45480 271 45546 287
rect 48592 321 48658 337
rect 49370 329 49436 345
rect 48592 287 48608 321
rect 48642 287 48658 321
rect 44702 229 44718 263
rect 44752 229 44768 263
rect 40812 171 40828 205
rect 40862 171 40878 205
rect 40812 155 40878 171
rect 43924 205 43990 221
rect 44702 213 44768 229
rect 47814 263 47880 279
rect 48592 271 48658 287
rect 47814 229 47830 263
rect 47864 229 47880 263
rect 43924 171 43940 205
rect 43974 171 43990 205
rect 43924 155 43990 171
rect 47036 205 47102 221
rect 47814 213 47880 229
rect 47036 171 47052 205
rect 47086 171 47102 205
rect 47036 155 47102 171
<< viali >>
rect 2706 345 2740 379
rect 5818 345 5852 379
rect 1928 287 1962 321
rect 8930 345 8964 379
rect 5040 287 5074 321
rect 1150 229 1184 263
rect 12042 345 12076 379
rect 8152 287 8186 321
rect 4262 229 4296 263
rect 372 171 406 205
rect 15154 345 15188 379
rect 11264 287 11298 321
rect 7374 229 7408 263
rect 3484 171 3518 205
rect 18266 345 18300 379
rect 14376 287 14410 321
rect 10486 229 10520 263
rect 6596 171 6630 205
rect 21378 345 21412 379
rect 17488 287 17522 321
rect 13598 229 13632 263
rect 9708 171 9742 205
rect 24490 345 24524 379
rect 20600 287 20634 321
rect 16710 229 16744 263
rect 12820 171 12854 205
rect 27602 345 27636 379
rect 23712 287 23746 321
rect 19822 229 19856 263
rect 15932 171 15966 205
rect 30714 345 30748 379
rect 26824 287 26858 321
rect 22934 229 22968 263
rect 19044 171 19078 205
rect 33826 345 33860 379
rect 29936 287 29970 321
rect 26046 229 26080 263
rect 22156 171 22190 205
rect 36938 345 36972 379
rect 33048 287 33082 321
rect 29158 229 29192 263
rect 25268 171 25302 205
rect 40050 345 40084 379
rect 36160 287 36194 321
rect 32270 229 32304 263
rect 28380 171 28414 205
rect 43162 345 43196 379
rect 39272 287 39306 321
rect 35382 229 35416 263
rect 31492 171 31526 205
rect 46274 345 46308 379
rect 42384 287 42418 321
rect 38494 229 38528 263
rect 34604 171 34638 205
rect 49386 345 49420 379
rect 45496 287 45530 321
rect 41606 229 41640 263
rect 37716 171 37750 205
rect 48608 287 48642 321
rect 44718 229 44752 263
rect 40828 171 40862 205
rect 47830 229 47864 263
rect 43940 171 43974 205
rect 47052 171 47086 205
<< metal1 >>
rect 2694 379 2752 385
rect 2694 376 2706 379
rect 0 348 2706 376
rect 2694 345 2706 348
rect 2740 376 2752 379
rect 5806 379 5864 385
rect 5806 376 5818 379
rect 2740 348 5818 376
rect 2740 345 2752 348
rect 2694 339 2752 345
rect 5806 345 5818 348
rect 5852 376 5864 379
rect 8918 379 8976 385
rect 8918 376 8930 379
rect 5852 348 8930 376
rect 5852 345 5864 348
rect 5806 339 5864 345
rect 8918 345 8930 348
rect 8964 376 8976 379
rect 12030 379 12088 385
rect 12030 376 12042 379
rect 8964 348 12042 376
rect 8964 345 8976 348
rect 8918 339 8976 345
rect 12030 345 12042 348
rect 12076 376 12088 379
rect 15142 379 15200 385
rect 15142 376 15154 379
rect 12076 348 15154 376
rect 12076 345 12088 348
rect 12030 339 12088 345
rect 15142 345 15154 348
rect 15188 376 15200 379
rect 18254 379 18312 385
rect 18254 376 18266 379
rect 15188 348 18266 376
rect 15188 345 15200 348
rect 15142 339 15200 345
rect 18254 345 18266 348
rect 18300 376 18312 379
rect 21366 379 21424 385
rect 21366 376 21378 379
rect 18300 348 21378 376
rect 18300 345 18312 348
rect 18254 339 18312 345
rect 21366 345 21378 348
rect 21412 376 21424 379
rect 24478 379 24536 385
rect 24478 376 24490 379
rect 21412 348 24490 376
rect 21412 345 21424 348
rect 21366 339 21424 345
rect 24478 345 24490 348
rect 24524 376 24536 379
rect 27590 379 27648 385
rect 27590 376 27602 379
rect 24524 348 27602 376
rect 24524 345 24536 348
rect 24478 339 24536 345
rect 27590 345 27602 348
rect 27636 376 27648 379
rect 30702 379 30760 385
rect 30702 376 30714 379
rect 27636 348 30714 376
rect 27636 345 27648 348
rect 27590 339 27648 345
rect 30702 345 30714 348
rect 30748 376 30760 379
rect 33814 379 33872 385
rect 33814 376 33826 379
rect 30748 348 33826 376
rect 30748 345 30760 348
rect 30702 339 30760 345
rect 33814 345 33826 348
rect 33860 376 33872 379
rect 36926 379 36984 385
rect 36926 376 36938 379
rect 33860 348 36938 376
rect 33860 345 33872 348
rect 33814 339 33872 345
rect 36926 345 36938 348
rect 36972 376 36984 379
rect 40038 379 40096 385
rect 40038 376 40050 379
rect 36972 348 40050 376
rect 36972 345 36984 348
rect 36926 339 36984 345
rect 40038 345 40050 348
rect 40084 376 40096 379
rect 43150 379 43208 385
rect 43150 376 43162 379
rect 40084 348 43162 376
rect 40084 345 40096 348
rect 40038 339 40096 345
rect 43150 345 43162 348
rect 43196 376 43208 379
rect 46262 379 46320 385
rect 46262 376 46274 379
rect 43196 348 46274 376
rect 43196 345 43208 348
rect 43150 339 43208 345
rect 46262 345 46274 348
rect 46308 376 46320 379
rect 49374 379 49432 385
rect 49374 376 49386 379
rect 46308 348 49386 376
rect 46308 345 46320 348
rect 46262 339 46320 345
rect 49374 345 49386 348
rect 49420 376 49432 379
rect 49420 348 49792 376
rect 49420 345 49432 348
rect 49374 339 49432 345
rect 1916 321 1974 327
rect 1916 318 1928 321
rect 0 290 1928 318
rect 1916 287 1928 290
rect 1962 318 1974 321
rect 5028 321 5086 327
rect 5028 318 5040 321
rect 1962 290 5040 318
rect 1962 287 1974 290
rect 1916 281 1974 287
rect 5028 287 5040 290
rect 5074 318 5086 321
rect 8140 321 8198 327
rect 8140 318 8152 321
rect 5074 290 8152 318
rect 5074 287 5086 290
rect 5028 281 5086 287
rect 8140 287 8152 290
rect 8186 318 8198 321
rect 11252 321 11310 327
rect 11252 318 11264 321
rect 8186 290 11264 318
rect 8186 287 8198 290
rect 8140 281 8198 287
rect 11252 287 11264 290
rect 11298 318 11310 321
rect 14364 321 14422 327
rect 14364 318 14376 321
rect 11298 290 14376 318
rect 11298 287 11310 290
rect 11252 281 11310 287
rect 14364 287 14376 290
rect 14410 318 14422 321
rect 17476 321 17534 327
rect 17476 318 17488 321
rect 14410 290 17488 318
rect 14410 287 14422 290
rect 14364 281 14422 287
rect 17476 287 17488 290
rect 17522 318 17534 321
rect 20588 321 20646 327
rect 20588 318 20600 321
rect 17522 290 20600 318
rect 17522 287 17534 290
rect 17476 281 17534 287
rect 20588 287 20600 290
rect 20634 318 20646 321
rect 23700 321 23758 327
rect 23700 318 23712 321
rect 20634 290 23712 318
rect 20634 287 20646 290
rect 20588 281 20646 287
rect 23700 287 23712 290
rect 23746 318 23758 321
rect 26812 321 26870 327
rect 26812 318 26824 321
rect 23746 290 26824 318
rect 23746 287 23758 290
rect 23700 281 23758 287
rect 26812 287 26824 290
rect 26858 318 26870 321
rect 29924 321 29982 327
rect 29924 318 29936 321
rect 26858 290 29936 318
rect 26858 287 26870 290
rect 26812 281 26870 287
rect 29924 287 29936 290
rect 29970 318 29982 321
rect 33036 321 33094 327
rect 33036 318 33048 321
rect 29970 290 33048 318
rect 29970 287 29982 290
rect 29924 281 29982 287
rect 33036 287 33048 290
rect 33082 318 33094 321
rect 36148 321 36206 327
rect 36148 318 36160 321
rect 33082 290 36160 318
rect 33082 287 33094 290
rect 33036 281 33094 287
rect 36148 287 36160 290
rect 36194 318 36206 321
rect 39260 321 39318 327
rect 39260 318 39272 321
rect 36194 290 39272 318
rect 36194 287 36206 290
rect 36148 281 36206 287
rect 39260 287 39272 290
rect 39306 318 39318 321
rect 42372 321 42430 327
rect 42372 318 42384 321
rect 39306 290 42384 318
rect 39306 287 39318 290
rect 39260 281 39318 287
rect 42372 287 42384 290
rect 42418 318 42430 321
rect 45484 321 45542 327
rect 45484 318 45496 321
rect 42418 290 45496 318
rect 42418 287 42430 290
rect 42372 281 42430 287
rect 45484 287 45496 290
rect 45530 318 45542 321
rect 48596 321 48654 327
rect 48596 318 48608 321
rect 45530 290 48608 318
rect 45530 287 45542 290
rect 45484 281 45542 287
rect 48596 287 48608 290
rect 48642 318 48654 321
rect 48642 290 49792 318
rect 48642 287 48654 290
rect 48596 281 48654 287
rect 1138 263 1196 269
rect 1138 260 1150 263
rect 0 232 1150 260
rect 1138 229 1150 232
rect 1184 260 1196 263
rect 4250 263 4308 269
rect 4250 260 4262 263
rect 1184 232 4262 260
rect 1184 229 1196 232
rect 1138 223 1196 229
rect 4250 229 4262 232
rect 4296 260 4308 263
rect 7362 263 7420 269
rect 7362 260 7374 263
rect 4296 232 7374 260
rect 4296 229 4308 232
rect 4250 223 4308 229
rect 7362 229 7374 232
rect 7408 260 7420 263
rect 10474 263 10532 269
rect 10474 260 10486 263
rect 7408 232 10486 260
rect 7408 229 7420 232
rect 7362 223 7420 229
rect 10474 229 10486 232
rect 10520 260 10532 263
rect 13586 263 13644 269
rect 13586 260 13598 263
rect 10520 232 13598 260
rect 10520 229 10532 232
rect 10474 223 10532 229
rect 13586 229 13598 232
rect 13632 260 13644 263
rect 16698 263 16756 269
rect 16698 260 16710 263
rect 13632 232 16710 260
rect 13632 229 13644 232
rect 13586 223 13644 229
rect 16698 229 16710 232
rect 16744 260 16756 263
rect 19810 263 19868 269
rect 19810 260 19822 263
rect 16744 232 19822 260
rect 16744 229 16756 232
rect 16698 223 16756 229
rect 19810 229 19822 232
rect 19856 260 19868 263
rect 22922 263 22980 269
rect 22922 260 22934 263
rect 19856 232 22934 260
rect 19856 229 19868 232
rect 19810 223 19868 229
rect 22922 229 22934 232
rect 22968 260 22980 263
rect 26034 263 26092 269
rect 26034 260 26046 263
rect 22968 232 26046 260
rect 22968 229 22980 232
rect 22922 223 22980 229
rect 26034 229 26046 232
rect 26080 260 26092 263
rect 29146 263 29204 269
rect 29146 260 29158 263
rect 26080 232 29158 260
rect 26080 229 26092 232
rect 26034 223 26092 229
rect 29146 229 29158 232
rect 29192 260 29204 263
rect 32258 263 32316 269
rect 32258 260 32270 263
rect 29192 232 32270 260
rect 29192 229 29204 232
rect 29146 223 29204 229
rect 32258 229 32270 232
rect 32304 260 32316 263
rect 35370 263 35428 269
rect 35370 260 35382 263
rect 32304 232 35382 260
rect 32304 229 32316 232
rect 32258 223 32316 229
rect 35370 229 35382 232
rect 35416 260 35428 263
rect 38482 263 38540 269
rect 38482 260 38494 263
rect 35416 232 38494 260
rect 35416 229 35428 232
rect 35370 223 35428 229
rect 38482 229 38494 232
rect 38528 260 38540 263
rect 41594 263 41652 269
rect 41594 260 41606 263
rect 38528 232 41606 260
rect 38528 229 38540 232
rect 38482 223 38540 229
rect 41594 229 41606 232
rect 41640 260 41652 263
rect 44706 263 44764 269
rect 44706 260 44718 263
rect 41640 232 44718 260
rect 41640 229 41652 232
rect 41594 223 41652 229
rect 44706 229 44718 232
rect 44752 260 44764 263
rect 47818 263 47876 269
rect 47818 260 47830 263
rect 44752 232 47830 260
rect 44752 229 44764 232
rect 44706 223 44764 229
rect 47818 229 47830 232
rect 47864 260 47876 263
rect 47864 232 49792 260
rect 47864 229 47876 232
rect 47818 223 47876 229
rect 360 205 418 211
rect 360 202 372 205
rect 0 174 372 202
rect 360 171 372 174
rect 406 202 418 205
rect 3472 205 3530 211
rect 3472 202 3484 205
rect 406 174 3484 202
rect 406 171 418 174
rect 360 165 418 171
rect 3472 171 3484 174
rect 3518 202 3530 205
rect 6584 205 6642 211
rect 6584 202 6596 205
rect 3518 174 6596 202
rect 3518 171 3530 174
rect 3472 165 3530 171
rect 6584 171 6596 174
rect 6630 202 6642 205
rect 9696 205 9754 211
rect 9696 202 9708 205
rect 6630 174 9708 202
rect 6630 171 6642 174
rect 6584 165 6642 171
rect 9696 171 9708 174
rect 9742 202 9754 205
rect 12808 205 12866 211
rect 12808 202 12820 205
rect 9742 174 12820 202
rect 9742 171 9754 174
rect 9696 165 9754 171
rect 12808 171 12820 174
rect 12854 202 12866 205
rect 15920 205 15978 211
rect 15920 202 15932 205
rect 12854 174 15932 202
rect 12854 171 12866 174
rect 12808 165 12866 171
rect 15920 171 15932 174
rect 15966 202 15978 205
rect 19032 205 19090 211
rect 19032 202 19044 205
rect 15966 174 19044 202
rect 15966 171 15978 174
rect 15920 165 15978 171
rect 19032 171 19044 174
rect 19078 202 19090 205
rect 22144 205 22202 211
rect 22144 202 22156 205
rect 19078 174 22156 202
rect 19078 171 19090 174
rect 19032 165 19090 171
rect 22144 171 22156 174
rect 22190 202 22202 205
rect 25256 205 25314 211
rect 25256 202 25268 205
rect 22190 174 25268 202
rect 22190 171 22202 174
rect 22144 165 22202 171
rect 25256 171 25268 174
rect 25302 202 25314 205
rect 28368 205 28426 211
rect 28368 202 28380 205
rect 25302 174 28380 202
rect 25302 171 25314 174
rect 25256 165 25314 171
rect 28368 171 28380 174
rect 28414 202 28426 205
rect 31480 205 31538 211
rect 31480 202 31492 205
rect 28414 174 31492 202
rect 28414 171 28426 174
rect 28368 165 28426 171
rect 31480 171 31492 174
rect 31526 202 31538 205
rect 34592 205 34650 211
rect 34592 202 34604 205
rect 31526 174 34604 202
rect 31526 171 31538 174
rect 31480 165 31538 171
rect 34592 171 34604 174
rect 34638 202 34650 205
rect 37704 205 37762 211
rect 37704 202 37716 205
rect 34638 174 37716 202
rect 34638 171 34650 174
rect 34592 165 34650 171
rect 37704 171 37716 174
rect 37750 202 37762 205
rect 40816 205 40874 211
rect 40816 202 40828 205
rect 37750 174 40828 202
rect 37750 171 37762 174
rect 37704 165 37762 171
rect 40816 171 40828 174
rect 40862 202 40874 205
rect 43928 205 43986 211
rect 43928 202 43940 205
rect 40862 174 43940 202
rect 40862 171 40874 174
rect 40816 165 40874 171
rect 43928 171 43940 174
rect 43974 202 43986 205
rect 47040 205 47098 211
rect 47040 202 47052 205
rect 43974 174 47052 202
rect 43974 171 43986 174
rect 43928 165 43986 171
rect 47040 171 47052 174
rect 47086 202 47098 205
rect 47086 174 49792 202
rect 47086 171 47098 174
rect 47040 165 47098 171
rect 108 102 834 130
rect 886 102 1612 130
rect 1664 102 2390 130
rect 3220 102 3946 130
rect 3998 102 4724 130
rect 4776 102 5502 130
rect 6332 102 7058 130
rect 7110 102 7836 130
rect 7888 102 8614 130
rect 9444 102 10170 130
rect 10222 102 10948 130
rect 11000 102 11726 130
rect 12556 102 13282 130
rect 13334 102 14060 130
rect 14112 102 14838 130
rect 15668 102 16394 130
rect 16446 102 17172 130
rect 17224 102 17950 130
rect 18780 102 19506 130
rect 19558 102 20284 130
rect 20336 102 21062 130
rect 21892 102 22618 130
rect 22670 102 23396 130
rect 23448 102 24174 130
rect 25004 102 25730 130
rect 25782 102 26508 130
rect 26560 102 27286 130
rect 28116 102 28842 130
rect 28894 102 29620 130
rect 29672 102 30398 130
rect 31228 102 31954 130
rect 32006 102 32732 130
rect 32784 102 33510 130
rect 34340 102 35066 130
rect 35118 102 35844 130
rect 35896 102 36622 130
rect 37452 102 38178 130
rect 38230 102 38956 130
rect 39008 102 39734 130
rect 40564 102 41290 130
rect 41342 102 42068 130
rect 42120 102 42846 130
rect 43676 102 44402 130
rect 44454 102 45180 130
rect 45232 102 45958 130
rect 46788 102 47514 130
rect 47566 102 48292 130
rect 48344 102 49070 130
rect 750 44 1476 72
rect 1528 44 2254 72
rect 2306 44 3032 72
rect 3862 44 4588 72
rect 4640 44 5366 72
rect 5418 44 6144 72
rect 6974 44 7700 72
rect 7752 44 8478 72
rect 8530 44 9256 72
rect 10086 44 10812 72
rect 10864 44 11590 72
rect 11642 44 12368 72
rect 13198 44 13924 72
rect 13976 44 14702 72
rect 14754 44 15480 72
rect 16310 44 17036 72
rect 17088 44 17814 72
rect 17866 44 18592 72
rect 19422 44 20148 72
rect 20200 44 20926 72
rect 20978 44 21704 72
rect 22534 44 23260 72
rect 23312 44 24038 72
rect 24090 44 24816 72
rect 25646 44 26372 72
rect 26424 44 27150 72
rect 27202 44 27928 72
rect 28758 44 29484 72
rect 29536 44 30262 72
rect 30314 44 31040 72
rect 31870 44 32596 72
rect 32648 44 33374 72
rect 33426 44 34152 72
rect 34982 44 35708 72
rect 35760 44 36486 72
rect 36538 44 37264 72
rect 38094 44 38820 72
rect 38872 44 39598 72
rect 39650 44 40376 72
rect 41206 44 41932 72
rect 41984 44 42710 72
rect 42762 44 43488 72
rect 44318 44 45044 72
rect 45096 44 45822 72
rect 45874 44 46600 72
rect 47430 44 48156 72
rect 48208 44 48934 72
rect 48986 44 49712 72
<< via1 >>
rect 56 90 108 142
rect 834 90 886 142
rect 1612 90 1664 142
rect 2390 90 2442 142
rect 3168 90 3220 142
rect 3946 90 3998 142
rect 4724 90 4776 142
rect 5502 90 5554 142
rect 6280 90 6332 142
rect 7058 90 7110 142
rect 7836 90 7888 142
rect 8614 90 8666 142
rect 9392 90 9444 142
rect 10170 90 10222 142
rect 10948 90 11000 142
rect 11726 90 11778 142
rect 12504 90 12556 142
rect 13282 90 13334 142
rect 14060 90 14112 142
rect 14838 90 14890 142
rect 15616 90 15668 142
rect 16394 90 16446 142
rect 17172 90 17224 142
rect 17950 90 18002 142
rect 18728 90 18780 142
rect 19506 90 19558 142
rect 20284 90 20336 142
rect 21062 90 21114 142
rect 21840 90 21892 142
rect 22618 90 22670 142
rect 23396 90 23448 142
rect 24174 90 24226 142
rect 24952 90 25004 142
rect 25730 90 25782 142
rect 26508 90 26560 142
rect 27286 90 27338 142
rect 28064 90 28116 142
rect 28842 90 28894 142
rect 29620 90 29672 142
rect 30398 90 30450 142
rect 31176 90 31228 142
rect 31954 90 32006 142
rect 32732 90 32784 142
rect 33510 90 33562 142
rect 34288 90 34340 142
rect 35066 90 35118 142
rect 35844 90 35896 142
rect 36622 90 36674 142
rect 37400 90 37452 142
rect 38178 90 38230 142
rect 38956 90 39008 142
rect 39734 90 39786 142
rect 40512 90 40564 142
rect 41290 90 41342 142
rect 42068 90 42120 142
rect 42846 90 42898 142
rect 43624 90 43676 142
rect 44402 90 44454 142
rect 45180 90 45232 142
rect 45958 90 46010 142
rect 46736 90 46788 142
rect 47514 90 47566 142
rect 48292 90 48344 142
rect 49070 90 49122 142
rect 698 32 750 84
rect 1476 32 1528 84
rect 2254 32 2306 84
rect 3032 32 3084 84
rect 3810 32 3862 84
rect 4588 32 4640 84
rect 5366 32 5418 84
rect 6144 32 6196 84
rect 6922 32 6974 84
rect 7700 32 7752 84
rect 8478 32 8530 84
rect 9256 32 9308 84
rect 10034 32 10086 84
rect 10812 32 10864 84
rect 11590 32 11642 84
rect 12368 32 12420 84
rect 13146 32 13198 84
rect 13924 32 13976 84
rect 14702 32 14754 84
rect 15480 32 15532 84
rect 16258 32 16310 84
rect 17036 32 17088 84
rect 17814 32 17866 84
rect 18592 32 18644 84
rect 19370 32 19422 84
rect 20148 32 20200 84
rect 20926 32 20978 84
rect 21704 32 21756 84
rect 22482 32 22534 84
rect 23260 32 23312 84
rect 24038 32 24090 84
rect 24816 32 24868 84
rect 25594 32 25646 84
rect 26372 32 26424 84
rect 27150 32 27202 84
rect 27928 32 27980 84
rect 28706 32 28758 84
rect 29484 32 29536 84
rect 30262 32 30314 84
rect 31040 32 31092 84
rect 31818 32 31870 84
rect 32596 32 32648 84
rect 33374 32 33426 84
rect 34152 32 34204 84
rect 34930 32 34982 84
rect 35708 32 35760 84
rect 36486 32 36538 84
rect 37264 32 37316 84
rect 38042 32 38094 84
rect 38820 32 38872 84
rect 39598 32 39650 84
rect 40376 32 40428 84
rect 41154 32 41206 84
rect 41932 32 41984 84
rect 42710 32 42762 84
rect 43488 32 43540 84
rect 44266 32 44318 84
rect 45044 32 45096 84
rect 45822 32 45874 84
rect 46600 32 46652 84
rect 47378 32 47430 84
rect 48156 32 48208 84
rect 48934 32 48986 84
rect 49712 32 49764 84
<< metal2 >>
rect 68 1858 96 1914
rect 710 1858 738 1914
rect 846 1858 874 1914
rect 1488 1858 1516 1914
rect 1624 1858 1652 1914
rect 2266 1858 2294 1914
rect 2402 1858 2430 1914
rect 3044 1858 3072 1914
rect 3180 1858 3208 1914
rect 3822 1858 3850 1914
rect 3958 1858 3986 1914
rect 4600 1858 4628 1914
rect 4736 1858 4764 1914
rect 5378 1858 5406 1914
rect 5514 1858 5542 1914
rect 6156 1858 6184 1914
rect 6292 1858 6320 1914
rect 6934 1858 6962 1914
rect 7070 1858 7098 1914
rect 7712 1858 7740 1914
rect 7848 1858 7876 1914
rect 8490 1858 8518 1914
rect 8626 1858 8654 1914
rect 9268 1858 9296 1914
rect 9404 1858 9432 1914
rect 10046 1858 10074 1914
rect 10182 1858 10210 1914
rect 10824 1858 10852 1914
rect 10960 1858 10988 1914
rect 11602 1858 11630 1914
rect 11738 1858 11766 1914
rect 12380 1858 12408 1914
rect 12516 1858 12544 1914
rect 13158 1858 13186 1914
rect 13294 1858 13322 1914
rect 13936 1858 13964 1914
rect 14072 1858 14100 1914
rect 14714 1858 14742 1914
rect 14850 1858 14878 1914
rect 15492 1858 15520 1914
rect 15628 1858 15656 1914
rect 16270 1858 16298 1914
rect 16406 1858 16434 1914
rect 17048 1858 17076 1914
rect 17184 1858 17212 1914
rect 17826 1858 17854 1914
rect 17962 1858 17990 1914
rect 18604 1858 18632 1914
rect 18740 1858 18768 1914
rect 19382 1858 19410 1914
rect 19518 1858 19546 1914
rect 20160 1858 20188 1914
rect 20296 1858 20324 1914
rect 20938 1858 20966 1914
rect 21074 1858 21102 1914
rect 21716 1858 21744 1914
rect 21852 1858 21880 1914
rect 22494 1858 22522 1914
rect 22630 1858 22658 1914
rect 23272 1858 23300 1914
rect 23408 1858 23436 1914
rect 24050 1858 24078 1914
rect 24186 1858 24214 1914
rect 24828 1858 24856 1914
rect 24964 1858 24992 1914
rect 25606 1858 25634 1914
rect 25742 1858 25770 1914
rect 26384 1858 26412 1914
rect 26520 1858 26548 1914
rect 27162 1858 27190 1914
rect 27298 1858 27326 1914
rect 27940 1858 27968 1914
rect 28076 1858 28104 1914
rect 28718 1858 28746 1914
rect 28854 1858 28882 1914
rect 29496 1858 29524 1914
rect 29632 1858 29660 1914
rect 30274 1858 30302 1914
rect 30410 1858 30438 1914
rect 31052 1858 31080 1914
rect 31188 1858 31216 1914
rect 31830 1858 31858 1914
rect 31966 1858 31994 1914
rect 32608 1858 32636 1914
rect 32744 1858 32772 1914
rect 33386 1858 33414 1914
rect 33522 1858 33550 1914
rect 34164 1858 34192 1914
rect 34300 1858 34328 1914
rect 34942 1858 34970 1914
rect 35078 1858 35106 1914
rect 35720 1858 35748 1914
rect 35856 1858 35884 1914
rect 36498 1858 36526 1914
rect 36634 1858 36662 1914
rect 37276 1858 37304 1914
rect 37412 1858 37440 1914
rect 38054 1858 38082 1914
rect 38190 1858 38218 1914
rect 38832 1858 38860 1914
rect 38968 1858 38996 1914
rect 39610 1858 39638 1914
rect 39746 1858 39774 1914
rect 40388 1858 40416 1914
rect 40524 1858 40552 1914
rect 41166 1858 41194 1914
rect 41302 1858 41330 1914
rect 41944 1858 41972 1914
rect 42080 1858 42108 1914
rect 42722 1858 42750 1914
rect 42858 1858 42886 1914
rect 43500 1858 43528 1914
rect 43636 1858 43664 1914
rect 44278 1858 44306 1914
rect 44414 1858 44442 1914
rect 45056 1858 45084 1914
rect 45192 1858 45220 1914
rect 45834 1858 45862 1914
rect 45970 1858 45998 1914
rect 46612 1858 46640 1914
rect 46748 1858 46776 1914
rect 47390 1858 47418 1914
rect 47526 1858 47554 1914
rect 48168 1858 48196 1914
rect 48304 1858 48332 1914
rect 48946 1858 48974 1914
rect 49082 1858 49110 1914
rect 49724 1858 49752 1914
rect 68 142 96 406
rect 710 84 738 406
rect 846 142 874 406
rect 1488 84 1516 406
rect 1624 142 1652 406
rect 2266 84 2294 406
rect 2402 142 2430 406
rect 3044 84 3072 406
rect 3180 142 3208 406
rect 3822 84 3850 406
rect 3958 142 3986 406
rect 4600 84 4628 406
rect 4736 142 4764 406
rect 5378 84 5406 406
rect 5514 142 5542 406
rect 6156 84 6184 406
rect 6292 142 6320 406
rect 6934 84 6962 406
rect 7070 142 7098 406
rect 7712 84 7740 406
rect 7848 142 7876 406
rect 8490 84 8518 406
rect 8626 142 8654 406
rect 9268 84 9296 406
rect 9404 142 9432 406
rect 10046 84 10074 406
rect 10182 142 10210 406
rect 10824 84 10852 406
rect 10960 142 10988 406
rect 11602 84 11630 406
rect 11738 142 11766 406
rect 12380 84 12408 406
rect 12516 142 12544 406
rect 13158 84 13186 406
rect 13294 142 13322 406
rect 13936 84 13964 406
rect 14072 142 14100 406
rect 14714 84 14742 406
rect 14850 142 14878 406
rect 15492 84 15520 406
rect 15628 142 15656 406
rect 16270 84 16298 406
rect 16406 142 16434 406
rect 17048 84 17076 406
rect 17184 142 17212 406
rect 17826 84 17854 406
rect 17962 142 17990 406
rect 18604 84 18632 406
rect 18740 142 18768 406
rect 19382 84 19410 406
rect 19518 142 19546 406
rect 20160 84 20188 406
rect 20296 142 20324 406
rect 20938 84 20966 406
rect 21074 142 21102 406
rect 21716 84 21744 406
rect 21852 142 21880 406
rect 22494 84 22522 406
rect 22630 142 22658 406
rect 23272 84 23300 406
rect 23408 142 23436 406
rect 24050 84 24078 406
rect 24186 142 24214 406
rect 24828 84 24856 406
rect 24964 142 24992 406
rect 25606 84 25634 406
rect 25742 142 25770 406
rect 26384 84 26412 406
rect 26520 142 26548 406
rect 27162 84 27190 406
rect 27298 142 27326 406
rect 27940 84 27968 406
rect 28076 142 28104 406
rect 28718 84 28746 406
rect 28854 142 28882 406
rect 29496 84 29524 406
rect 29632 142 29660 406
rect 30274 84 30302 406
rect 30410 142 30438 406
rect 31052 84 31080 406
rect 31188 142 31216 406
rect 31830 84 31858 406
rect 31966 142 31994 406
rect 32608 84 32636 406
rect 32744 142 32772 406
rect 33386 84 33414 406
rect 33522 142 33550 406
rect 34164 84 34192 406
rect 34300 142 34328 406
rect 34942 84 34970 406
rect 35078 142 35106 406
rect 35720 84 35748 406
rect 35856 142 35884 406
rect 36498 84 36526 406
rect 36634 142 36662 406
rect 37276 84 37304 406
rect 37412 142 37440 406
rect 38054 84 38082 406
rect 38190 142 38218 406
rect 38832 84 38860 406
rect 38968 142 38996 406
rect 39610 84 39638 406
rect 39746 142 39774 406
rect 40388 84 40416 406
rect 40524 142 40552 406
rect 41166 84 41194 406
rect 41302 142 41330 406
rect 41944 84 41972 406
rect 42080 142 42108 406
rect 42722 84 42750 406
rect 42858 142 42886 406
rect 43500 84 43528 406
rect 43636 142 43664 406
rect 44278 84 44306 406
rect 44414 142 44442 406
rect 45056 84 45084 406
rect 45192 142 45220 406
rect 45834 84 45862 406
rect 45970 142 45998 406
rect 46612 84 46640 406
rect 46748 142 46776 406
rect 47390 84 47418 406
rect 47526 142 47554 406
rect 48168 84 48196 406
rect 48304 142 48332 406
rect 48946 84 48974 406
rect 49082 142 49110 406
rect 49724 84 49752 406
<< metal3 >>
rect 712 1132 844 1198
rect 1490 1132 1622 1198
rect 2268 1132 2400 1198
rect 3046 1132 3178 1198
rect 3824 1132 3956 1198
rect 4602 1132 4734 1198
rect 5380 1132 5512 1198
rect 6158 1132 6290 1198
rect 6936 1132 7068 1198
rect 7714 1132 7846 1198
rect 8492 1132 8624 1198
rect 9270 1132 9402 1198
rect 10048 1132 10180 1198
rect 10826 1132 10958 1198
rect 11604 1132 11736 1198
rect 12382 1132 12514 1198
rect 13160 1132 13292 1198
rect 13938 1132 14070 1198
rect 14716 1132 14848 1198
rect 15494 1132 15626 1198
rect 16272 1132 16404 1198
rect 17050 1132 17182 1198
rect 17828 1132 17960 1198
rect 18606 1132 18738 1198
rect 19384 1132 19516 1198
rect 20162 1132 20294 1198
rect 20940 1132 21072 1198
rect 21718 1132 21850 1198
rect 22496 1132 22628 1198
rect 23274 1132 23406 1198
rect 24052 1132 24184 1198
rect 24830 1132 24962 1198
rect 25608 1132 25740 1198
rect 26386 1132 26518 1198
rect 27164 1132 27296 1198
rect 27942 1132 28074 1198
rect 28720 1132 28852 1198
rect 29498 1132 29630 1198
rect 30276 1132 30408 1198
rect 31054 1132 31186 1198
rect 31832 1132 31964 1198
rect 32610 1132 32742 1198
rect 33388 1132 33520 1198
rect 34166 1132 34298 1198
rect 34944 1132 35076 1198
rect 35722 1132 35854 1198
rect 36500 1132 36632 1198
rect 37278 1132 37410 1198
rect 38056 1132 38188 1198
rect 38834 1132 38966 1198
rect 39612 1132 39744 1198
rect 40390 1132 40522 1198
rect 41168 1132 41300 1198
rect 41946 1132 42078 1198
rect 42724 1132 42856 1198
rect 43502 1132 43634 1198
rect 44280 1132 44412 1198
rect 45058 1132 45190 1198
rect 45836 1132 45968 1198
rect 46614 1132 46746 1198
rect 47392 1132 47524 1198
rect 48170 1132 48302 1198
rect 48948 1132 49080 1198
rect 49726 1132 49858 1198
use contact_14  contact_14_0
timestamp 1643678851
transform 1 0 49723 0 1 43
box 0 0 1 1
use contact_14  contact_14_1
timestamp 1643678851
transform 1 0 49081 0 1 101
box 0 0 1 1
use contact_14  contact_14_2
timestamp 1643678851
transform 1 0 48945 0 1 43
box 0 0 1 1
use contact_14  contact_14_3
timestamp 1643678851
transform 1 0 48303 0 1 101
box 0 0 1 1
use contact_14  contact_14_4
timestamp 1643678851
transform 1 0 48167 0 1 43
box 0 0 1 1
use contact_14  contact_14_5
timestamp 1643678851
transform 1 0 47525 0 1 101
box 0 0 1 1
use contact_14  contact_14_6
timestamp 1643678851
transform 1 0 47389 0 1 43
box 0 0 1 1
use contact_14  contact_14_7
timestamp 1643678851
transform 1 0 46747 0 1 101
box 0 0 1 1
use contact_14  contact_14_8
timestamp 1643678851
transform 1 0 46611 0 1 43
box 0 0 1 1
use contact_14  contact_14_9
timestamp 1643678851
transform 1 0 45969 0 1 101
box 0 0 1 1
use contact_14  contact_14_10
timestamp 1643678851
transform 1 0 45833 0 1 43
box 0 0 1 1
use contact_14  contact_14_11
timestamp 1643678851
transform 1 0 45191 0 1 101
box 0 0 1 1
use contact_14  contact_14_12
timestamp 1643678851
transform 1 0 45055 0 1 43
box 0 0 1 1
use contact_14  contact_14_13
timestamp 1643678851
transform 1 0 44413 0 1 101
box 0 0 1 1
use contact_14  contact_14_14
timestamp 1643678851
transform 1 0 44277 0 1 43
box 0 0 1 1
use contact_14  contact_14_15
timestamp 1643678851
transform 1 0 43635 0 1 101
box 0 0 1 1
use contact_14  contact_14_16
timestamp 1643678851
transform 1 0 43499 0 1 43
box 0 0 1 1
use contact_14  contact_14_17
timestamp 1643678851
transform 1 0 42857 0 1 101
box 0 0 1 1
use contact_14  contact_14_18
timestamp 1643678851
transform 1 0 42721 0 1 43
box 0 0 1 1
use contact_14  contact_14_19
timestamp 1643678851
transform 1 0 42079 0 1 101
box 0 0 1 1
use contact_14  contact_14_20
timestamp 1643678851
transform 1 0 41943 0 1 43
box 0 0 1 1
use contact_14  contact_14_21
timestamp 1643678851
transform 1 0 41301 0 1 101
box 0 0 1 1
use contact_14  contact_14_22
timestamp 1643678851
transform 1 0 41165 0 1 43
box 0 0 1 1
use contact_14  contact_14_23
timestamp 1643678851
transform 1 0 40523 0 1 101
box 0 0 1 1
use contact_14  contact_14_24
timestamp 1643678851
transform 1 0 40387 0 1 43
box 0 0 1 1
use contact_14  contact_14_25
timestamp 1643678851
transform 1 0 39745 0 1 101
box 0 0 1 1
use contact_14  contact_14_26
timestamp 1643678851
transform 1 0 39609 0 1 43
box 0 0 1 1
use contact_14  contact_14_27
timestamp 1643678851
transform 1 0 38967 0 1 101
box 0 0 1 1
use contact_14  contact_14_28
timestamp 1643678851
transform 1 0 38831 0 1 43
box 0 0 1 1
use contact_14  contact_14_29
timestamp 1643678851
transform 1 0 38189 0 1 101
box 0 0 1 1
use contact_14  contact_14_30
timestamp 1643678851
transform 1 0 38053 0 1 43
box 0 0 1 1
use contact_14  contact_14_31
timestamp 1643678851
transform 1 0 37411 0 1 101
box 0 0 1 1
use contact_14  contact_14_32
timestamp 1643678851
transform 1 0 37275 0 1 43
box 0 0 1 1
use contact_14  contact_14_33
timestamp 1643678851
transform 1 0 36633 0 1 101
box 0 0 1 1
use contact_14  contact_14_34
timestamp 1643678851
transform 1 0 36497 0 1 43
box 0 0 1 1
use contact_14  contact_14_35
timestamp 1643678851
transform 1 0 35855 0 1 101
box 0 0 1 1
use contact_14  contact_14_36
timestamp 1643678851
transform 1 0 35719 0 1 43
box 0 0 1 1
use contact_14  contact_14_37
timestamp 1643678851
transform 1 0 35077 0 1 101
box 0 0 1 1
use contact_14  contact_14_38
timestamp 1643678851
transform 1 0 34941 0 1 43
box 0 0 1 1
use contact_14  contact_14_39
timestamp 1643678851
transform 1 0 34299 0 1 101
box 0 0 1 1
use contact_14  contact_14_40
timestamp 1643678851
transform 1 0 34163 0 1 43
box 0 0 1 1
use contact_14  contact_14_41
timestamp 1643678851
transform 1 0 33521 0 1 101
box 0 0 1 1
use contact_14  contact_14_42
timestamp 1643678851
transform 1 0 33385 0 1 43
box 0 0 1 1
use contact_14  contact_14_43
timestamp 1643678851
transform 1 0 32743 0 1 101
box 0 0 1 1
use contact_14  contact_14_44
timestamp 1643678851
transform 1 0 32607 0 1 43
box 0 0 1 1
use contact_14  contact_14_45
timestamp 1643678851
transform 1 0 31965 0 1 101
box 0 0 1 1
use contact_14  contact_14_46
timestamp 1643678851
transform 1 0 31829 0 1 43
box 0 0 1 1
use contact_14  contact_14_47
timestamp 1643678851
transform 1 0 31187 0 1 101
box 0 0 1 1
use contact_14  contact_14_48
timestamp 1643678851
transform 1 0 31051 0 1 43
box 0 0 1 1
use contact_14  contact_14_49
timestamp 1643678851
transform 1 0 30409 0 1 101
box 0 0 1 1
use contact_14  contact_14_50
timestamp 1643678851
transform 1 0 30273 0 1 43
box 0 0 1 1
use contact_14  contact_14_51
timestamp 1643678851
transform 1 0 29631 0 1 101
box 0 0 1 1
use contact_14  contact_14_52
timestamp 1643678851
transform 1 0 29495 0 1 43
box 0 0 1 1
use contact_14  contact_14_53
timestamp 1643678851
transform 1 0 28853 0 1 101
box 0 0 1 1
use contact_14  contact_14_54
timestamp 1643678851
transform 1 0 28717 0 1 43
box 0 0 1 1
use contact_14  contact_14_55
timestamp 1643678851
transform 1 0 28075 0 1 101
box 0 0 1 1
use contact_14  contact_14_56
timestamp 1643678851
transform 1 0 27939 0 1 43
box 0 0 1 1
use contact_14  contact_14_57
timestamp 1643678851
transform 1 0 27297 0 1 101
box 0 0 1 1
use contact_14  contact_14_58
timestamp 1643678851
transform 1 0 27161 0 1 43
box 0 0 1 1
use contact_14  contact_14_59
timestamp 1643678851
transform 1 0 26519 0 1 101
box 0 0 1 1
use contact_14  contact_14_60
timestamp 1643678851
transform 1 0 26383 0 1 43
box 0 0 1 1
use contact_14  contact_14_61
timestamp 1643678851
transform 1 0 25741 0 1 101
box 0 0 1 1
use contact_14  contact_14_62
timestamp 1643678851
transform 1 0 25605 0 1 43
box 0 0 1 1
use contact_14  contact_14_63
timestamp 1643678851
transform 1 0 24963 0 1 101
box 0 0 1 1
use contact_14  contact_14_64
timestamp 1643678851
transform 1 0 24827 0 1 43
box 0 0 1 1
use contact_14  contact_14_65
timestamp 1643678851
transform 1 0 24185 0 1 101
box 0 0 1 1
use contact_14  contact_14_66
timestamp 1643678851
transform 1 0 24049 0 1 43
box 0 0 1 1
use contact_14  contact_14_67
timestamp 1643678851
transform 1 0 23407 0 1 101
box 0 0 1 1
use contact_14  contact_14_68
timestamp 1643678851
transform 1 0 23271 0 1 43
box 0 0 1 1
use contact_14  contact_14_69
timestamp 1643678851
transform 1 0 22629 0 1 101
box 0 0 1 1
use contact_14  contact_14_70
timestamp 1643678851
transform 1 0 22493 0 1 43
box 0 0 1 1
use contact_14  contact_14_71
timestamp 1643678851
transform 1 0 21851 0 1 101
box 0 0 1 1
use contact_14  contact_14_72
timestamp 1643678851
transform 1 0 21715 0 1 43
box 0 0 1 1
use contact_14  contact_14_73
timestamp 1643678851
transform 1 0 21073 0 1 101
box 0 0 1 1
use contact_14  contact_14_74
timestamp 1643678851
transform 1 0 20937 0 1 43
box 0 0 1 1
use contact_14  contact_14_75
timestamp 1643678851
transform 1 0 20295 0 1 101
box 0 0 1 1
use contact_14  contact_14_76
timestamp 1643678851
transform 1 0 20159 0 1 43
box 0 0 1 1
use contact_14  contact_14_77
timestamp 1643678851
transform 1 0 19517 0 1 101
box 0 0 1 1
use contact_14  contact_14_78
timestamp 1643678851
transform 1 0 19381 0 1 43
box 0 0 1 1
use contact_14  contact_14_79
timestamp 1643678851
transform 1 0 18739 0 1 101
box 0 0 1 1
use contact_14  contact_14_80
timestamp 1643678851
transform 1 0 18603 0 1 43
box 0 0 1 1
use contact_14  contact_14_81
timestamp 1643678851
transform 1 0 17961 0 1 101
box 0 0 1 1
use contact_14  contact_14_82
timestamp 1643678851
transform 1 0 17825 0 1 43
box 0 0 1 1
use contact_14  contact_14_83
timestamp 1643678851
transform 1 0 17183 0 1 101
box 0 0 1 1
use contact_14  contact_14_84
timestamp 1643678851
transform 1 0 17047 0 1 43
box 0 0 1 1
use contact_14  contact_14_85
timestamp 1643678851
transform 1 0 16405 0 1 101
box 0 0 1 1
use contact_14  contact_14_86
timestamp 1643678851
transform 1 0 16269 0 1 43
box 0 0 1 1
use contact_14  contact_14_87
timestamp 1643678851
transform 1 0 15627 0 1 101
box 0 0 1 1
use contact_14  contact_14_88
timestamp 1643678851
transform 1 0 15491 0 1 43
box 0 0 1 1
use contact_14  contact_14_89
timestamp 1643678851
transform 1 0 14849 0 1 101
box 0 0 1 1
use contact_14  contact_14_90
timestamp 1643678851
transform 1 0 14713 0 1 43
box 0 0 1 1
use contact_14  contact_14_91
timestamp 1643678851
transform 1 0 14071 0 1 101
box 0 0 1 1
use contact_14  contact_14_92
timestamp 1643678851
transform 1 0 13935 0 1 43
box 0 0 1 1
use contact_14  contact_14_93
timestamp 1643678851
transform 1 0 13293 0 1 101
box 0 0 1 1
use contact_14  contact_14_94
timestamp 1643678851
transform 1 0 13157 0 1 43
box 0 0 1 1
use contact_14  contact_14_95
timestamp 1643678851
transform 1 0 12515 0 1 101
box 0 0 1 1
use contact_14  contact_14_96
timestamp 1643678851
transform 1 0 12379 0 1 43
box 0 0 1 1
use contact_14  contact_14_97
timestamp 1643678851
transform 1 0 11737 0 1 101
box 0 0 1 1
use contact_14  contact_14_98
timestamp 1643678851
transform 1 0 11601 0 1 43
box 0 0 1 1
use contact_14  contact_14_99
timestamp 1643678851
transform 1 0 10959 0 1 101
box 0 0 1 1
use contact_14  contact_14_100
timestamp 1643678851
transform 1 0 10823 0 1 43
box 0 0 1 1
use contact_14  contact_14_101
timestamp 1643678851
transform 1 0 10181 0 1 101
box 0 0 1 1
use contact_14  contact_14_102
timestamp 1643678851
transform 1 0 10045 0 1 43
box 0 0 1 1
use contact_14  contact_14_103
timestamp 1643678851
transform 1 0 9403 0 1 101
box 0 0 1 1
use contact_14  contact_14_104
timestamp 1643678851
transform 1 0 9267 0 1 43
box 0 0 1 1
use contact_14  contact_14_105
timestamp 1643678851
transform 1 0 8625 0 1 101
box 0 0 1 1
use contact_14  contact_14_106
timestamp 1643678851
transform 1 0 8489 0 1 43
box 0 0 1 1
use contact_14  contact_14_107
timestamp 1643678851
transform 1 0 7847 0 1 101
box 0 0 1 1
use contact_14  contact_14_108
timestamp 1643678851
transform 1 0 7711 0 1 43
box 0 0 1 1
use contact_14  contact_14_109
timestamp 1643678851
transform 1 0 7069 0 1 101
box 0 0 1 1
use contact_14  contact_14_110
timestamp 1643678851
transform 1 0 6933 0 1 43
box 0 0 1 1
use contact_14  contact_14_111
timestamp 1643678851
transform 1 0 6291 0 1 101
box 0 0 1 1
use contact_14  contact_14_112
timestamp 1643678851
transform 1 0 6155 0 1 43
box 0 0 1 1
use contact_14  contact_14_113
timestamp 1643678851
transform 1 0 5513 0 1 101
box 0 0 1 1
use contact_14  contact_14_114
timestamp 1643678851
transform 1 0 5377 0 1 43
box 0 0 1 1
use contact_14  contact_14_115
timestamp 1643678851
transform 1 0 4735 0 1 101
box 0 0 1 1
use contact_14  contact_14_116
timestamp 1643678851
transform 1 0 4599 0 1 43
box 0 0 1 1
use contact_14  contact_14_117
timestamp 1643678851
transform 1 0 3957 0 1 101
box 0 0 1 1
use contact_14  contact_14_118
timestamp 1643678851
transform 1 0 3821 0 1 43
box 0 0 1 1
use contact_14  contact_14_119
timestamp 1643678851
transform 1 0 3179 0 1 101
box 0 0 1 1
use contact_14  contact_14_120
timestamp 1643678851
transform 1 0 3043 0 1 43
box 0 0 1 1
use contact_14  contact_14_121
timestamp 1643678851
transform 1 0 2401 0 1 101
box 0 0 1 1
use contact_14  contact_14_122
timestamp 1643678851
transform 1 0 2265 0 1 43
box 0 0 1 1
use contact_14  contact_14_123
timestamp 1643678851
transform 1 0 1623 0 1 101
box 0 0 1 1
use contact_14  contact_14_124
timestamp 1643678851
transform 1 0 1487 0 1 43
box 0 0 1 1
use contact_14  contact_14_125
timestamp 1643678851
transform 1 0 845 0 1 101
box 0 0 1 1
use contact_14  contact_14_126
timestamp 1643678851
transform 1 0 709 0 1 43
box 0 0 1 1
use contact_14  contact_14_127
timestamp 1643678851
transform 1 0 67 0 1 101
box 0 0 1 1
use contact_27  contact_27_0
timestamp 1643678851
transform 1 0 49374 0 1 339
box 0 0 1 1
use contact_26  contact_26_0
timestamp 1643678851
transform 1 0 49370 0 1 329
box 0 0 1 1
use contact_27  contact_27_1
timestamp 1643678851
transform 1 0 48596 0 1 281
box 0 0 1 1
use contact_26  contact_26_1
timestamp 1643678851
transform 1 0 48592 0 1 271
box 0 0 1 1
use contact_27  contact_27_2
timestamp 1643678851
transform 1 0 47818 0 1 223
box 0 0 1 1
use contact_26  contact_26_2
timestamp 1643678851
transform 1 0 47814 0 1 213
box 0 0 1 1
use contact_27  contact_27_3
timestamp 1643678851
transform 1 0 47040 0 1 165
box 0 0 1 1
use contact_26  contact_26_3
timestamp 1643678851
transform 1 0 47036 0 1 155
box 0 0 1 1
use contact_27  contact_27_4
timestamp 1643678851
transform 1 0 46262 0 1 339
box 0 0 1 1
use contact_26  contact_26_4
timestamp 1643678851
transform 1 0 46258 0 1 329
box 0 0 1 1
use contact_27  contact_27_5
timestamp 1643678851
transform 1 0 45484 0 1 281
box 0 0 1 1
use contact_26  contact_26_5
timestamp 1643678851
transform 1 0 45480 0 1 271
box 0 0 1 1
use contact_27  contact_27_6
timestamp 1643678851
transform 1 0 44706 0 1 223
box 0 0 1 1
use contact_26  contact_26_6
timestamp 1643678851
transform 1 0 44702 0 1 213
box 0 0 1 1
use contact_27  contact_27_7
timestamp 1643678851
transform 1 0 43928 0 1 165
box 0 0 1 1
use contact_26  contact_26_7
timestamp 1643678851
transform 1 0 43924 0 1 155
box 0 0 1 1
use contact_27  contact_27_8
timestamp 1643678851
transform 1 0 43150 0 1 339
box 0 0 1 1
use contact_26  contact_26_8
timestamp 1643678851
transform 1 0 43146 0 1 329
box 0 0 1 1
use contact_27  contact_27_9
timestamp 1643678851
transform 1 0 42372 0 1 281
box 0 0 1 1
use contact_26  contact_26_9
timestamp 1643678851
transform 1 0 42368 0 1 271
box 0 0 1 1
use contact_27  contact_27_10
timestamp 1643678851
transform 1 0 41594 0 1 223
box 0 0 1 1
use contact_26  contact_26_10
timestamp 1643678851
transform 1 0 41590 0 1 213
box 0 0 1 1
use contact_27  contact_27_11
timestamp 1643678851
transform 1 0 40816 0 1 165
box 0 0 1 1
use contact_26  contact_26_11
timestamp 1643678851
transform 1 0 40812 0 1 155
box 0 0 1 1
use contact_27  contact_27_12
timestamp 1643678851
transform 1 0 40038 0 1 339
box 0 0 1 1
use contact_26  contact_26_12
timestamp 1643678851
transform 1 0 40034 0 1 329
box 0 0 1 1
use contact_27  contact_27_13
timestamp 1643678851
transform 1 0 39260 0 1 281
box 0 0 1 1
use contact_26  contact_26_13
timestamp 1643678851
transform 1 0 39256 0 1 271
box 0 0 1 1
use contact_27  contact_27_14
timestamp 1643678851
transform 1 0 38482 0 1 223
box 0 0 1 1
use contact_26  contact_26_14
timestamp 1643678851
transform 1 0 38478 0 1 213
box 0 0 1 1
use contact_27  contact_27_15
timestamp 1643678851
transform 1 0 37704 0 1 165
box 0 0 1 1
use contact_26  contact_26_15
timestamp 1643678851
transform 1 0 37700 0 1 155
box 0 0 1 1
use contact_27  contact_27_16
timestamp 1643678851
transform 1 0 36926 0 1 339
box 0 0 1 1
use contact_26  contact_26_16
timestamp 1643678851
transform 1 0 36922 0 1 329
box 0 0 1 1
use contact_27  contact_27_17
timestamp 1643678851
transform 1 0 36148 0 1 281
box 0 0 1 1
use contact_26  contact_26_17
timestamp 1643678851
transform 1 0 36144 0 1 271
box 0 0 1 1
use contact_27  contact_27_18
timestamp 1643678851
transform 1 0 35370 0 1 223
box 0 0 1 1
use contact_26  contact_26_18
timestamp 1643678851
transform 1 0 35366 0 1 213
box 0 0 1 1
use contact_27  contact_27_19
timestamp 1643678851
transform 1 0 34592 0 1 165
box 0 0 1 1
use contact_26  contact_26_19
timestamp 1643678851
transform 1 0 34588 0 1 155
box 0 0 1 1
use contact_27  contact_27_20
timestamp 1643678851
transform 1 0 33814 0 1 339
box 0 0 1 1
use contact_26  contact_26_20
timestamp 1643678851
transform 1 0 33810 0 1 329
box 0 0 1 1
use contact_27  contact_27_21
timestamp 1643678851
transform 1 0 33036 0 1 281
box 0 0 1 1
use contact_26  contact_26_21
timestamp 1643678851
transform 1 0 33032 0 1 271
box 0 0 1 1
use contact_27  contact_27_22
timestamp 1643678851
transform 1 0 32258 0 1 223
box 0 0 1 1
use contact_26  contact_26_22
timestamp 1643678851
transform 1 0 32254 0 1 213
box 0 0 1 1
use contact_27  contact_27_23
timestamp 1643678851
transform 1 0 31480 0 1 165
box 0 0 1 1
use contact_26  contact_26_23
timestamp 1643678851
transform 1 0 31476 0 1 155
box 0 0 1 1
use contact_27  contact_27_24
timestamp 1643678851
transform 1 0 30702 0 1 339
box 0 0 1 1
use contact_26  contact_26_24
timestamp 1643678851
transform 1 0 30698 0 1 329
box 0 0 1 1
use contact_27  contact_27_25
timestamp 1643678851
transform 1 0 29924 0 1 281
box 0 0 1 1
use contact_26  contact_26_25
timestamp 1643678851
transform 1 0 29920 0 1 271
box 0 0 1 1
use contact_27  contact_27_26
timestamp 1643678851
transform 1 0 29146 0 1 223
box 0 0 1 1
use contact_26  contact_26_26
timestamp 1643678851
transform 1 0 29142 0 1 213
box 0 0 1 1
use contact_27  contact_27_27
timestamp 1643678851
transform 1 0 28368 0 1 165
box 0 0 1 1
use contact_26  contact_26_27
timestamp 1643678851
transform 1 0 28364 0 1 155
box 0 0 1 1
use contact_27  contact_27_28
timestamp 1643678851
transform 1 0 27590 0 1 339
box 0 0 1 1
use contact_26  contact_26_28
timestamp 1643678851
transform 1 0 27586 0 1 329
box 0 0 1 1
use contact_27  contact_27_29
timestamp 1643678851
transform 1 0 26812 0 1 281
box 0 0 1 1
use contact_26  contact_26_29
timestamp 1643678851
transform 1 0 26808 0 1 271
box 0 0 1 1
use contact_27  contact_27_30
timestamp 1643678851
transform 1 0 26034 0 1 223
box 0 0 1 1
use contact_26  contact_26_30
timestamp 1643678851
transform 1 0 26030 0 1 213
box 0 0 1 1
use contact_27  contact_27_31
timestamp 1643678851
transform 1 0 25256 0 1 165
box 0 0 1 1
use contact_26  contact_26_31
timestamp 1643678851
transform 1 0 25252 0 1 155
box 0 0 1 1
use contact_27  contact_27_32
timestamp 1643678851
transform 1 0 24478 0 1 339
box 0 0 1 1
use contact_26  contact_26_32
timestamp 1643678851
transform 1 0 24474 0 1 329
box 0 0 1 1
use contact_27  contact_27_33
timestamp 1643678851
transform 1 0 23700 0 1 281
box 0 0 1 1
use contact_26  contact_26_33
timestamp 1643678851
transform 1 0 23696 0 1 271
box 0 0 1 1
use contact_27  contact_27_34
timestamp 1643678851
transform 1 0 22922 0 1 223
box 0 0 1 1
use contact_26  contact_26_34
timestamp 1643678851
transform 1 0 22918 0 1 213
box 0 0 1 1
use contact_27  contact_27_35
timestamp 1643678851
transform 1 0 22144 0 1 165
box 0 0 1 1
use contact_26  contact_26_35
timestamp 1643678851
transform 1 0 22140 0 1 155
box 0 0 1 1
use contact_27  contact_27_36
timestamp 1643678851
transform 1 0 21366 0 1 339
box 0 0 1 1
use contact_26  contact_26_36
timestamp 1643678851
transform 1 0 21362 0 1 329
box 0 0 1 1
use contact_27  contact_27_37
timestamp 1643678851
transform 1 0 20588 0 1 281
box 0 0 1 1
use contact_26  contact_26_37
timestamp 1643678851
transform 1 0 20584 0 1 271
box 0 0 1 1
use contact_27  contact_27_38
timestamp 1643678851
transform 1 0 19810 0 1 223
box 0 0 1 1
use contact_26  contact_26_38
timestamp 1643678851
transform 1 0 19806 0 1 213
box 0 0 1 1
use contact_27  contact_27_39
timestamp 1643678851
transform 1 0 19032 0 1 165
box 0 0 1 1
use contact_26  contact_26_39
timestamp 1643678851
transform 1 0 19028 0 1 155
box 0 0 1 1
use contact_27  contact_27_40
timestamp 1643678851
transform 1 0 18254 0 1 339
box 0 0 1 1
use contact_26  contact_26_40
timestamp 1643678851
transform 1 0 18250 0 1 329
box 0 0 1 1
use contact_27  contact_27_41
timestamp 1643678851
transform 1 0 17476 0 1 281
box 0 0 1 1
use contact_26  contact_26_41
timestamp 1643678851
transform 1 0 17472 0 1 271
box 0 0 1 1
use contact_27  contact_27_42
timestamp 1643678851
transform 1 0 16698 0 1 223
box 0 0 1 1
use contact_26  contact_26_42
timestamp 1643678851
transform 1 0 16694 0 1 213
box 0 0 1 1
use contact_27  contact_27_43
timestamp 1643678851
transform 1 0 15920 0 1 165
box 0 0 1 1
use contact_26  contact_26_43
timestamp 1643678851
transform 1 0 15916 0 1 155
box 0 0 1 1
use contact_27  contact_27_44
timestamp 1643678851
transform 1 0 15142 0 1 339
box 0 0 1 1
use contact_26  contact_26_44
timestamp 1643678851
transform 1 0 15138 0 1 329
box 0 0 1 1
use contact_27  contact_27_45
timestamp 1643678851
transform 1 0 14364 0 1 281
box 0 0 1 1
use contact_26  contact_26_45
timestamp 1643678851
transform 1 0 14360 0 1 271
box 0 0 1 1
use contact_27  contact_27_46
timestamp 1643678851
transform 1 0 13586 0 1 223
box 0 0 1 1
use contact_26  contact_26_46
timestamp 1643678851
transform 1 0 13582 0 1 213
box 0 0 1 1
use contact_27  contact_27_47
timestamp 1643678851
transform 1 0 12808 0 1 165
box 0 0 1 1
use contact_26  contact_26_47
timestamp 1643678851
transform 1 0 12804 0 1 155
box 0 0 1 1
use contact_27  contact_27_48
timestamp 1643678851
transform 1 0 12030 0 1 339
box 0 0 1 1
use contact_26  contact_26_48
timestamp 1643678851
transform 1 0 12026 0 1 329
box 0 0 1 1
use contact_27  contact_27_49
timestamp 1643678851
transform 1 0 11252 0 1 281
box 0 0 1 1
use contact_26  contact_26_49
timestamp 1643678851
transform 1 0 11248 0 1 271
box 0 0 1 1
use contact_27  contact_27_50
timestamp 1643678851
transform 1 0 10474 0 1 223
box 0 0 1 1
use contact_26  contact_26_50
timestamp 1643678851
transform 1 0 10470 0 1 213
box 0 0 1 1
use contact_27  contact_27_51
timestamp 1643678851
transform 1 0 9696 0 1 165
box 0 0 1 1
use contact_26  contact_26_51
timestamp 1643678851
transform 1 0 9692 0 1 155
box 0 0 1 1
use contact_27  contact_27_52
timestamp 1643678851
transform 1 0 8918 0 1 339
box 0 0 1 1
use contact_26  contact_26_52
timestamp 1643678851
transform 1 0 8914 0 1 329
box 0 0 1 1
use contact_27  contact_27_53
timestamp 1643678851
transform 1 0 8140 0 1 281
box 0 0 1 1
use contact_26  contact_26_53
timestamp 1643678851
transform 1 0 8136 0 1 271
box 0 0 1 1
use contact_27  contact_27_54
timestamp 1643678851
transform 1 0 7362 0 1 223
box 0 0 1 1
use contact_26  contact_26_54
timestamp 1643678851
transform 1 0 7358 0 1 213
box 0 0 1 1
use contact_27  contact_27_55
timestamp 1643678851
transform 1 0 6584 0 1 165
box 0 0 1 1
use contact_26  contact_26_55
timestamp 1643678851
transform 1 0 6580 0 1 155
box 0 0 1 1
use contact_27  contact_27_56
timestamp 1643678851
transform 1 0 5806 0 1 339
box 0 0 1 1
use contact_26  contact_26_56
timestamp 1643678851
transform 1 0 5802 0 1 329
box 0 0 1 1
use contact_27  contact_27_57
timestamp 1643678851
transform 1 0 5028 0 1 281
box 0 0 1 1
use contact_26  contact_26_57
timestamp 1643678851
transform 1 0 5024 0 1 271
box 0 0 1 1
use contact_27  contact_27_58
timestamp 1643678851
transform 1 0 4250 0 1 223
box 0 0 1 1
use contact_26  contact_26_58
timestamp 1643678851
transform 1 0 4246 0 1 213
box 0 0 1 1
use contact_27  contact_27_59
timestamp 1643678851
transform 1 0 3472 0 1 165
box 0 0 1 1
use contact_26  contact_26_59
timestamp 1643678851
transform 1 0 3468 0 1 155
box 0 0 1 1
use contact_27  contact_27_60
timestamp 1643678851
transform 1 0 2694 0 1 339
box 0 0 1 1
use contact_26  contact_26_60
timestamp 1643678851
transform 1 0 2690 0 1 329
box 0 0 1 1
use contact_27  contact_27_61
timestamp 1643678851
transform 1 0 1916 0 1 281
box 0 0 1 1
use contact_26  contact_26_61
timestamp 1643678851
transform 1 0 1912 0 1 271
box 0 0 1 1
use contact_27  contact_27_62
timestamp 1643678851
transform 1 0 1138 0 1 223
box 0 0 1 1
use contact_26  contact_26_62
timestamp 1643678851
transform 1 0 1134 0 1 213
box 0 0 1 1
use contact_27  contact_27_63
timestamp 1643678851
transform 1 0 360 0 1 165
box 0 0 1 1
use contact_26  contact_26_63
timestamp 1643678851
transform 1 0 356 0 1 155
box 0 0 1 1
use column_mux_multiport  column_mux_multiport_0
timestamp 1643678851
transform 1 0 49014 0 1 406
box 33 0 844 1508
use column_mux_multiport  column_mux_multiport_1
timestamp 1643678851
transform 1 0 48236 0 1 406
box 33 0 844 1508
use column_mux_multiport  column_mux_multiport_2
timestamp 1643678851
transform 1 0 47458 0 1 406
box 33 0 844 1508
use column_mux_multiport  column_mux_multiport_3
timestamp 1643678851
transform 1 0 46680 0 1 406
box 33 0 844 1508
use column_mux_multiport  column_mux_multiport_4
timestamp 1643678851
transform 1 0 45902 0 1 406
box 33 0 844 1508
use column_mux_multiport  column_mux_multiport_5
timestamp 1643678851
transform 1 0 45124 0 1 406
box 33 0 844 1508
use column_mux_multiport  column_mux_multiport_6
timestamp 1643678851
transform 1 0 44346 0 1 406
box 33 0 844 1508
use column_mux_multiport  column_mux_multiport_7
timestamp 1643678851
transform 1 0 43568 0 1 406
box 33 0 844 1508
use column_mux_multiport  column_mux_multiport_8
timestamp 1643678851
transform 1 0 42790 0 1 406
box 33 0 844 1508
use column_mux_multiport  column_mux_multiport_9
timestamp 1643678851
transform 1 0 42012 0 1 406
box 33 0 844 1508
use column_mux_multiport  column_mux_multiport_10
timestamp 1643678851
transform 1 0 41234 0 1 406
box 33 0 844 1508
use column_mux_multiport  column_mux_multiport_11
timestamp 1643678851
transform 1 0 40456 0 1 406
box 33 0 844 1508
use column_mux_multiport  column_mux_multiport_12
timestamp 1643678851
transform 1 0 39678 0 1 406
box 33 0 844 1508
use column_mux_multiport  column_mux_multiport_13
timestamp 1643678851
transform 1 0 38900 0 1 406
box 33 0 844 1508
use column_mux_multiport  column_mux_multiport_14
timestamp 1643678851
transform 1 0 38122 0 1 406
box 33 0 844 1508
use column_mux_multiport  column_mux_multiport_15
timestamp 1643678851
transform 1 0 37344 0 1 406
box 33 0 844 1508
use column_mux_multiport  column_mux_multiport_16
timestamp 1643678851
transform 1 0 36566 0 1 406
box 33 0 844 1508
use column_mux_multiport  column_mux_multiport_17
timestamp 1643678851
transform 1 0 35788 0 1 406
box 33 0 844 1508
use column_mux_multiport  column_mux_multiport_18
timestamp 1643678851
transform 1 0 35010 0 1 406
box 33 0 844 1508
use column_mux_multiport  column_mux_multiport_19
timestamp 1643678851
transform 1 0 34232 0 1 406
box 33 0 844 1508
use column_mux_multiport  column_mux_multiport_20
timestamp 1643678851
transform 1 0 33454 0 1 406
box 33 0 844 1508
use column_mux_multiport  column_mux_multiport_21
timestamp 1643678851
transform 1 0 32676 0 1 406
box 33 0 844 1508
use column_mux_multiport  column_mux_multiport_22
timestamp 1643678851
transform 1 0 31898 0 1 406
box 33 0 844 1508
use column_mux_multiport  column_mux_multiport_23
timestamp 1643678851
transform 1 0 31120 0 1 406
box 33 0 844 1508
use column_mux_multiport  column_mux_multiport_24
timestamp 1643678851
transform 1 0 30342 0 1 406
box 33 0 844 1508
use column_mux_multiport  column_mux_multiport_25
timestamp 1643678851
transform 1 0 29564 0 1 406
box 33 0 844 1508
use column_mux_multiport  column_mux_multiport_26
timestamp 1643678851
transform 1 0 28786 0 1 406
box 33 0 844 1508
use column_mux_multiport  column_mux_multiport_27
timestamp 1643678851
transform 1 0 28008 0 1 406
box 33 0 844 1508
use column_mux_multiport  column_mux_multiport_28
timestamp 1643678851
transform 1 0 27230 0 1 406
box 33 0 844 1508
use column_mux_multiport  column_mux_multiport_29
timestamp 1643678851
transform 1 0 26452 0 1 406
box 33 0 844 1508
use column_mux_multiport  column_mux_multiport_30
timestamp 1643678851
transform 1 0 25674 0 1 406
box 33 0 844 1508
use column_mux_multiport  column_mux_multiport_31
timestamp 1643678851
transform 1 0 24896 0 1 406
box 33 0 844 1508
use column_mux_multiport  column_mux_multiport_32
timestamp 1643678851
transform 1 0 24118 0 1 406
box 33 0 844 1508
use column_mux_multiport  column_mux_multiport_33
timestamp 1643678851
transform 1 0 23340 0 1 406
box 33 0 844 1508
use column_mux_multiport  column_mux_multiport_34
timestamp 1643678851
transform 1 0 22562 0 1 406
box 33 0 844 1508
use column_mux_multiport  column_mux_multiport_35
timestamp 1643678851
transform 1 0 21784 0 1 406
box 33 0 844 1508
use column_mux_multiport  column_mux_multiport_36
timestamp 1643678851
transform 1 0 21006 0 1 406
box 33 0 844 1508
use column_mux_multiport  column_mux_multiport_37
timestamp 1643678851
transform 1 0 20228 0 1 406
box 33 0 844 1508
use column_mux_multiport  column_mux_multiport_38
timestamp 1643678851
transform 1 0 19450 0 1 406
box 33 0 844 1508
use column_mux_multiport  column_mux_multiport_39
timestamp 1643678851
transform 1 0 18672 0 1 406
box 33 0 844 1508
use column_mux_multiport  column_mux_multiport_40
timestamp 1643678851
transform 1 0 17894 0 1 406
box 33 0 844 1508
use column_mux_multiport  column_mux_multiport_41
timestamp 1643678851
transform 1 0 17116 0 1 406
box 33 0 844 1508
use column_mux_multiport  column_mux_multiport_42
timestamp 1643678851
transform 1 0 16338 0 1 406
box 33 0 844 1508
use column_mux_multiport  column_mux_multiport_43
timestamp 1643678851
transform 1 0 15560 0 1 406
box 33 0 844 1508
use column_mux_multiport  column_mux_multiport_44
timestamp 1643678851
transform 1 0 14782 0 1 406
box 33 0 844 1508
use column_mux_multiport  column_mux_multiport_45
timestamp 1643678851
transform 1 0 14004 0 1 406
box 33 0 844 1508
use column_mux_multiport  column_mux_multiport_46
timestamp 1643678851
transform 1 0 13226 0 1 406
box 33 0 844 1508
use column_mux_multiport  column_mux_multiport_47
timestamp 1643678851
transform 1 0 12448 0 1 406
box 33 0 844 1508
use column_mux_multiport  column_mux_multiport_48
timestamp 1643678851
transform 1 0 11670 0 1 406
box 33 0 844 1508
use column_mux_multiport  column_mux_multiport_49
timestamp 1643678851
transform 1 0 10892 0 1 406
box 33 0 844 1508
use column_mux_multiport  column_mux_multiport_50
timestamp 1643678851
transform 1 0 10114 0 1 406
box 33 0 844 1508
use column_mux_multiport  column_mux_multiport_51
timestamp 1643678851
transform 1 0 9336 0 1 406
box 33 0 844 1508
use column_mux_multiport  column_mux_multiport_52
timestamp 1643678851
transform 1 0 8558 0 1 406
box 33 0 844 1508
use column_mux_multiport  column_mux_multiport_53
timestamp 1643678851
transform 1 0 7780 0 1 406
box 33 0 844 1508
use column_mux_multiport  column_mux_multiport_54
timestamp 1643678851
transform 1 0 7002 0 1 406
box 33 0 844 1508
use column_mux_multiport  column_mux_multiport_55
timestamp 1643678851
transform 1 0 6224 0 1 406
box 33 0 844 1508
use column_mux_multiport  column_mux_multiport_56
timestamp 1643678851
transform 1 0 5446 0 1 406
box 33 0 844 1508
use column_mux_multiport  column_mux_multiport_57
timestamp 1643678851
transform 1 0 4668 0 1 406
box 33 0 844 1508
use column_mux_multiport  column_mux_multiport_58
timestamp 1643678851
transform 1 0 3890 0 1 406
box 33 0 844 1508
use column_mux_multiport  column_mux_multiport_59
timestamp 1643678851
transform 1 0 3112 0 1 406
box 33 0 844 1508
use column_mux_multiport  column_mux_multiport_60
timestamp 1643678851
transform 1 0 2334 0 1 406
box 33 0 844 1508
use column_mux_multiport  column_mux_multiport_61
timestamp 1643678851
transform 1 0 1556 0 1 406
box 33 0 844 1508
use column_mux_multiport  column_mux_multiport_62
timestamp 1643678851
transform 1 0 778 0 1 406
box 33 0 844 1508
use column_mux_multiport  column_mux_multiport_63
timestamp 1643678851
transform 1 0 0 0 1 406
box 33 0 844 1508
<< labels >>
rlabel metal1 s 0 174 49792 202 4 sel_0
rlabel metal1 s 0 232 49792 260 4 sel_1
rlabel metal1 s 0 290 49792 318 4 sel_2
rlabel metal1 s 0 348 49792 376 4 sel_3
rlabel metal2 s 68 116 96 406 4 rbl0_out_0
rlabel metal2 s 710 58 738 406 4 rbl1_out_0
rlabel metal2 s 3180 116 3208 406 4 rbl0_out_1
rlabel metal2 s 3822 58 3850 406 4 rbl1_out_1
rlabel metal2 s 6292 116 6320 406 4 rbl0_out_2
rlabel metal2 s 6934 58 6962 406 4 rbl1_out_2
rlabel metal2 s 9404 116 9432 406 4 rbl0_out_3
rlabel metal2 s 10046 58 10074 406 4 rbl1_out_3
rlabel metal2 s 12516 116 12544 406 4 rbl0_out_4
rlabel metal2 s 13158 58 13186 406 4 rbl1_out_4
rlabel metal2 s 15628 116 15656 406 4 rbl0_out_5
rlabel metal2 s 16270 58 16298 406 4 rbl1_out_5
rlabel metal2 s 18740 116 18768 406 4 rbl0_out_6
rlabel metal2 s 19382 58 19410 406 4 rbl1_out_6
rlabel metal2 s 21852 116 21880 406 4 rbl0_out_7
rlabel metal2 s 22494 58 22522 406 4 rbl1_out_7
rlabel metal2 s 24964 116 24992 406 4 rbl0_out_8
rlabel metal2 s 25606 58 25634 406 4 rbl1_out_8
rlabel metal2 s 28076 116 28104 406 4 rbl0_out_9
rlabel metal2 s 28718 58 28746 406 4 rbl1_out_9
rlabel metal2 s 31188 116 31216 406 4 rbl0_out_10
rlabel metal2 s 31830 58 31858 406 4 rbl1_out_10
rlabel metal2 s 34300 116 34328 406 4 rbl0_out_11
rlabel metal2 s 34942 58 34970 406 4 rbl1_out_11
rlabel metal2 s 37412 116 37440 406 4 rbl0_out_12
rlabel metal2 s 38054 58 38082 406 4 rbl1_out_12
rlabel metal2 s 40524 116 40552 406 4 rbl0_out_13
rlabel metal2 s 41166 58 41194 406 4 rbl1_out_13
rlabel metal2 s 43636 116 43664 406 4 rbl0_out_14
rlabel metal2 s 44278 58 44306 406 4 rbl1_out_14
rlabel metal2 s 46748 116 46776 406 4 rbl0_out_15
rlabel metal2 s 47390 58 47418 406 4 rbl1_out_15
rlabel metal2 s 68 1858 96 1914 4 rbl0_0
rlabel metal2 s 710 1858 738 1914 4 rbl1_0
rlabel metal2 s 846 1858 874 1914 4 rbl0_1
rlabel metal2 s 1488 1858 1516 1914 4 rbl1_1
rlabel metal2 s 1624 1858 1652 1914 4 rbl0_2
rlabel metal2 s 2266 1858 2294 1914 4 rbl1_2
rlabel metal2 s 2402 1858 2430 1914 4 rbl0_3
rlabel metal2 s 3044 1858 3072 1914 4 rbl1_3
rlabel metal2 s 3180 1858 3208 1914 4 rbl0_4
rlabel metal2 s 3822 1858 3850 1914 4 rbl1_4
rlabel metal2 s 3958 1858 3986 1914 4 rbl0_5
rlabel metal2 s 4600 1858 4628 1914 4 rbl1_5
rlabel metal2 s 4736 1858 4764 1914 4 rbl0_6
rlabel metal2 s 5378 1858 5406 1914 4 rbl1_6
rlabel metal2 s 5514 1858 5542 1914 4 rbl0_7
rlabel metal2 s 6156 1858 6184 1914 4 rbl1_7
rlabel metal2 s 6292 1858 6320 1914 4 rbl0_8
rlabel metal2 s 6934 1858 6962 1914 4 rbl1_8
rlabel metal2 s 7070 1858 7098 1914 4 rbl0_9
rlabel metal2 s 7712 1858 7740 1914 4 rbl1_9
rlabel metal2 s 7848 1858 7876 1914 4 rbl0_10
rlabel metal2 s 8490 1858 8518 1914 4 rbl1_10
rlabel metal2 s 8626 1858 8654 1914 4 rbl0_11
rlabel metal2 s 9268 1858 9296 1914 4 rbl1_11
rlabel metal2 s 9404 1858 9432 1914 4 rbl0_12
rlabel metal2 s 10046 1858 10074 1914 4 rbl1_12
rlabel metal2 s 10182 1858 10210 1914 4 rbl0_13
rlabel metal2 s 10824 1858 10852 1914 4 rbl1_13
rlabel metal2 s 10960 1858 10988 1914 4 rbl0_14
rlabel metal2 s 11602 1858 11630 1914 4 rbl1_14
rlabel metal2 s 11738 1858 11766 1914 4 rbl0_15
rlabel metal2 s 12380 1858 12408 1914 4 rbl1_15
rlabel metal2 s 12516 1858 12544 1914 4 rbl0_16
rlabel metal2 s 13158 1858 13186 1914 4 rbl1_16
rlabel metal2 s 13294 1858 13322 1914 4 rbl0_17
rlabel metal2 s 13936 1858 13964 1914 4 rbl1_17
rlabel metal2 s 14072 1858 14100 1914 4 rbl0_18
rlabel metal2 s 14714 1858 14742 1914 4 rbl1_18
rlabel metal2 s 14850 1858 14878 1914 4 rbl0_19
rlabel metal2 s 15492 1858 15520 1914 4 rbl1_19
rlabel metal2 s 15628 1858 15656 1914 4 rbl0_20
rlabel metal2 s 16270 1858 16298 1914 4 rbl1_20
rlabel metal2 s 16406 1858 16434 1914 4 rbl0_21
rlabel metal2 s 17048 1858 17076 1914 4 rbl1_21
rlabel metal2 s 17184 1858 17212 1914 4 rbl0_22
rlabel metal2 s 17826 1858 17854 1914 4 rbl1_22
rlabel metal2 s 17962 1858 17990 1914 4 rbl0_23
rlabel metal2 s 18604 1858 18632 1914 4 rbl1_23
rlabel metal2 s 18740 1858 18768 1914 4 rbl0_24
rlabel metal2 s 19382 1858 19410 1914 4 rbl1_24
rlabel metal2 s 19518 1858 19546 1914 4 rbl0_25
rlabel metal2 s 20160 1858 20188 1914 4 rbl1_25
rlabel metal2 s 20296 1858 20324 1914 4 rbl0_26
rlabel metal2 s 20938 1858 20966 1914 4 rbl1_26
rlabel metal2 s 21074 1858 21102 1914 4 rbl0_27
rlabel metal2 s 21716 1858 21744 1914 4 rbl1_27
rlabel metal2 s 21852 1858 21880 1914 4 rbl0_28
rlabel metal2 s 22494 1858 22522 1914 4 rbl1_28
rlabel metal2 s 22630 1858 22658 1914 4 rbl0_29
rlabel metal2 s 23272 1858 23300 1914 4 rbl1_29
rlabel metal2 s 23408 1858 23436 1914 4 rbl0_30
rlabel metal2 s 24050 1858 24078 1914 4 rbl1_30
rlabel metal2 s 24186 1858 24214 1914 4 rbl0_31
rlabel metal2 s 24828 1858 24856 1914 4 rbl1_31
rlabel metal2 s 24964 1858 24992 1914 4 rbl0_32
rlabel metal2 s 25606 1858 25634 1914 4 rbl1_32
rlabel metal2 s 25742 1858 25770 1914 4 rbl0_33
rlabel metal2 s 26384 1858 26412 1914 4 rbl1_33
rlabel metal2 s 26520 1858 26548 1914 4 rbl0_34
rlabel metal2 s 27162 1858 27190 1914 4 rbl1_34
rlabel metal2 s 27298 1858 27326 1914 4 rbl0_35
rlabel metal2 s 27940 1858 27968 1914 4 rbl1_35
rlabel metal2 s 28076 1858 28104 1914 4 rbl0_36
rlabel metal2 s 28718 1858 28746 1914 4 rbl1_36
rlabel metal2 s 28854 1858 28882 1914 4 rbl0_37
rlabel metal2 s 29496 1858 29524 1914 4 rbl1_37
rlabel metal2 s 29632 1858 29660 1914 4 rbl0_38
rlabel metal2 s 30274 1858 30302 1914 4 rbl1_38
rlabel metal2 s 30410 1858 30438 1914 4 rbl0_39
rlabel metal2 s 31052 1858 31080 1914 4 rbl1_39
rlabel metal2 s 31188 1858 31216 1914 4 rbl0_40
rlabel metal2 s 31830 1858 31858 1914 4 rbl1_40
rlabel metal2 s 31966 1858 31994 1914 4 rbl0_41
rlabel metal2 s 32608 1858 32636 1914 4 rbl1_41
rlabel metal2 s 32744 1858 32772 1914 4 rbl0_42
rlabel metal2 s 33386 1858 33414 1914 4 rbl1_42
rlabel metal2 s 33522 1858 33550 1914 4 rbl0_43
rlabel metal2 s 34164 1858 34192 1914 4 rbl1_43
rlabel metal2 s 34300 1858 34328 1914 4 rbl0_44
rlabel metal2 s 34942 1858 34970 1914 4 rbl1_44
rlabel metal2 s 35078 1858 35106 1914 4 rbl0_45
rlabel metal2 s 35720 1858 35748 1914 4 rbl1_45
rlabel metal2 s 35856 1858 35884 1914 4 rbl0_46
rlabel metal2 s 36498 1858 36526 1914 4 rbl1_46
rlabel metal2 s 36634 1858 36662 1914 4 rbl0_47
rlabel metal2 s 37276 1858 37304 1914 4 rbl1_47
rlabel metal2 s 37412 1858 37440 1914 4 rbl0_48
rlabel metal2 s 38054 1858 38082 1914 4 rbl1_48
rlabel metal2 s 38190 1858 38218 1914 4 rbl0_49
rlabel metal2 s 38832 1858 38860 1914 4 rbl1_49
rlabel metal2 s 38968 1858 38996 1914 4 rbl0_50
rlabel metal2 s 39610 1858 39638 1914 4 rbl1_50
rlabel metal2 s 39746 1858 39774 1914 4 rbl0_51
rlabel metal2 s 40388 1858 40416 1914 4 rbl1_51
rlabel metal2 s 40524 1858 40552 1914 4 rbl0_52
rlabel metal2 s 41166 1858 41194 1914 4 rbl1_52
rlabel metal2 s 41302 1858 41330 1914 4 rbl0_53
rlabel metal2 s 41944 1858 41972 1914 4 rbl1_53
rlabel metal2 s 42080 1858 42108 1914 4 rbl0_54
rlabel metal2 s 42722 1858 42750 1914 4 rbl1_54
rlabel metal2 s 42858 1858 42886 1914 4 rbl0_55
rlabel metal2 s 43500 1858 43528 1914 4 rbl1_55
rlabel metal2 s 43636 1858 43664 1914 4 rbl0_56
rlabel metal2 s 44278 1858 44306 1914 4 rbl1_56
rlabel metal2 s 44414 1858 44442 1914 4 rbl0_57
rlabel metal2 s 45056 1858 45084 1914 4 rbl1_57
rlabel metal2 s 45192 1858 45220 1914 4 rbl0_58
rlabel metal2 s 45834 1858 45862 1914 4 rbl1_58
rlabel metal2 s 45970 1858 45998 1914 4 rbl0_59
rlabel metal2 s 46612 1858 46640 1914 4 rbl1_59
rlabel metal2 s 46748 1858 46776 1914 4 rbl0_60
rlabel metal2 s 47390 1858 47418 1914 4 rbl1_60
rlabel metal2 s 47526 1858 47554 1914 4 rbl0_61
rlabel metal2 s 48168 1858 48196 1914 4 rbl1_61
rlabel metal2 s 48304 1858 48332 1914 4 rbl0_62
rlabel metal2 s 48946 1858 48974 1914 4 rbl1_62
rlabel metal2 s 49082 1858 49110 1914 4 rbl0_63
rlabel metal2 s 49724 1858 49752 1914 4 rbl1_63
rlabel metal3 s 3046 1132 3178 1198 4 gnd
rlabel metal3 s 5380 1132 5512 1198 4 gnd
rlabel metal3 s 11604 1132 11736 1198 4 gnd
rlabel metal3 s 20940 1132 21072 1198 4 gnd
rlabel metal3 s 24830 1132 24962 1198 4 gnd
rlabel metal3 s 37278 1132 37410 1198 4 gnd
rlabel metal3 s 41946 1132 42078 1198 4 gnd
rlabel metal3 s 20162 1132 20294 1198 4 gnd
rlabel metal3 s 13938 1132 14070 1198 4 gnd
rlabel metal3 s 21718 1132 21850 1198 4 gnd
rlabel metal3 s 36500 1132 36632 1198 4 gnd
rlabel metal3 s 22496 1132 22628 1198 4 gnd
rlabel metal3 s 25608 1132 25740 1198 4 gnd
rlabel metal3 s 45058 1132 45190 1198 4 gnd
rlabel metal3 s 31832 1132 31964 1198 4 gnd
rlabel metal3 s 17828 1132 17960 1198 4 gnd
rlabel metal3 s 18606 1132 18738 1198 4 gnd
rlabel metal3 s 1490 1132 1622 1198 4 gnd
rlabel metal3 s 10826 1132 10958 1198 4 gnd
rlabel metal3 s 17050 1132 17182 1198 4 gnd
rlabel metal3 s 4602 1132 4734 1198 4 gnd
rlabel metal3 s 14716 1132 14848 1198 4 gnd
rlabel metal3 s 29498 1132 29630 1198 4 gnd
rlabel metal3 s 6158 1132 6290 1198 4 gnd
rlabel metal3 s 26386 1132 26518 1198 4 gnd
rlabel metal3 s 32610 1132 32742 1198 4 gnd
rlabel metal3 s 45836 1132 45968 1198 4 gnd
rlabel metal3 s 28720 1132 28852 1198 4 gnd
rlabel metal3 s 47392 1132 47524 1198 4 gnd
rlabel metal3 s 42724 1132 42856 1198 4 gnd
rlabel metal3 s 39612 1132 39744 1198 4 gnd
rlabel metal3 s 12382 1132 12514 1198 4 gnd
rlabel metal3 s 15494 1132 15626 1198 4 gnd
rlabel metal3 s 38056 1132 38188 1198 4 gnd
rlabel metal3 s 712 1132 844 1198 4 gnd
rlabel metal3 s 38834 1132 38966 1198 4 gnd
rlabel metal3 s 46614 1132 46746 1198 4 gnd
rlabel metal3 s 10048 1132 10180 1198 4 gnd
rlabel metal3 s 34166 1132 34298 1198 4 gnd
rlabel metal3 s 33388 1132 33520 1198 4 gnd
rlabel metal3 s 8492 1132 8624 1198 4 gnd
rlabel metal3 s 30276 1132 30408 1198 4 gnd
rlabel metal3 s 44280 1132 44412 1198 4 gnd
rlabel metal3 s 3824 1132 3956 1198 4 gnd
rlabel metal3 s 9270 1132 9402 1198 4 gnd
rlabel metal3 s 27942 1132 28074 1198 4 gnd
rlabel metal3 s 34944 1132 35076 1198 4 gnd
rlabel metal3 s 16272 1132 16404 1198 4 gnd
rlabel metal3 s 41168 1132 41300 1198 4 gnd
rlabel metal3 s 31054 1132 31186 1198 4 gnd
rlabel metal3 s 6936 1132 7068 1198 4 gnd
rlabel metal3 s 24052 1132 24184 1198 4 gnd
rlabel metal3 s 48170 1132 48302 1198 4 gnd
rlabel metal3 s 7714 1132 7846 1198 4 gnd
rlabel metal3 s 19384 1132 19516 1198 4 gnd
rlabel metal3 s 2268 1132 2400 1198 4 gnd
rlabel metal3 s 13160 1132 13292 1198 4 gnd
rlabel metal3 s 23274 1132 23406 1198 4 gnd
rlabel metal3 s 49726 1132 49858 1198 4 gnd
rlabel metal3 s 48948 1132 49080 1198 4 gnd
rlabel metal3 s 27164 1132 27296 1198 4 gnd
rlabel metal3 s 43502 1132 43634 1198 4 gnd
rlabel metal3 s 40390 1132 40522 1198 4 gnd
rlabel metal3 s 35722 1132 35854 1198 4 gnd
<< properties >>
string FIXED_BBOX 0 0 49792 1914
string GDS_FILE sram_0rw2r1w_16_128_sky130A.gds
string GDS_END 1622846
string GDS_START 1553882
<< end >>
