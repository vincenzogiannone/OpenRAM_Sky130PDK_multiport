magic
tech sky130A
magscale 1 2
timestamp 1643671299
<< checkpaint >>
rect -1290 -1302 12496 7178
<< locali >>
rect 3833 4734 4035 4768
rect 4001 4550 4035 4734
rect 3807 2207 3983 2241
rect 3807 2154 3841 2207
rect 3682 2120 3841 2154
<< viali >>
rect 3550 5472 3584 5506
rect 5044 5472 5078 5506
rect 5929 4546 5963 4580
rect 3598 4463 3632 4497
rect 3598 3883 3632 3917
rect 5125 3802 5159 3836
rect 3698 3643 3732 3677
rect 3698 3027 3732 3061
rect 4585 2870 4619 2904
rect 3598 2787 3632 2821
rect 3550 2120 3584 2154
rect 4936 2124 4970 2158
rect 4049 1967 4083 2001
rect 3550 1198 3584 1232
rect 8988 1191 9022 1225
<< metal1 >>
rect 3538 5506 3596 5512
rect 3538 5503 3550 5506
rect 2982 5475 3550 5503
rect 3538 5472 3550 5475
rect 3584 5472 3596 5506
rect 5032 5504 5035 5512
rect 5006 5474 5035 5504
rect 3538 5466 3596 5472
rect 5032 5466 5035 5474
rect 5087 5504 5090 5512
rect 5087 5474 5117 5504
rect 5087 5466 5090 5474
rect 5917 4578 5920 4586
rect 5891 4548 5920 4578
rect 5917 4540 5920 4548
rect 5972 4578 5975 4586
rect 5972 4548 6002 4578
rect 5972 4540 5975 4548
rect 3586 4497 3644 4503
rect 3586 4494 3598 4497
rect 3050 4466 3598 4494
rect 3586 4463 3598 4466
rect 3632 4463 3644 4497
rect 3586 4457 3644 4463
rect 3586 3917 3644 3923
rect 3586 3914 3598 3917
rect 3118 3886 3598 3914
rect 3586 3883 3598 3886
rect 3632 3883 3644 3917
rect 3586 3877 3644 3883
rect 5113 3834 5116 3842
rect 5087 3804 5116 3834
rect 5113 3796 5116 3804
rect 5168 3834 5171 3842
rect 5168 3804 5198 3834
rect 5168 3796 5171 3804
rect 3686 3677 3744 3683
rect 3686 3674 3698 3677
rect 2982 3646 3698 3674
rect 3686 3643 3698 3646
rect 3732 3643 3744 3677
rect 3686 3637 3744 3643
rect 40 3280 3202 3308
rect 3686 3061 3744 3067
rect 3686 3058 3698 3061
rect 3322 3030 3698 3058
rect 3686 3027 3698 3030
rect 3732 3027 3744 3061
rect 3686 3021 3744 3027
rect 4573 2902 4576 2910
rect 4547 2872 4576 2902
rect 4573 2864 4576 2872
rect 4628 2902 4631 2910
rect 4628 2872 4658 2902
rect 4628 2864 4631 2872
rect 3586 2821 3644 2827
rect 3586 2818 3598 2821
rect 3254 2790 3598 2818
rect 3586 2787 3598 2790
rect 3632 2787 3644 2821
rect 3586 2781 3644 2787
rect 3538 2154 3596 2160
rect 4924 2156 4927 2164
rect 3538 2151 3550 2154
rect 3254 2123 3550 2151
rect 3538 2120 3550 2123
rect 3584 2120 3596 2154
rect 4898 2126 4927 2156
rect 3538 2114 3596 2120
rect 4924 2118 4927 2126
rect 4979 2156 4982 2164
rect 4979 2126 5009 2156
rect 4979 2118 4982 2126
rect 4037 1999 4040 2007
rect 4011 1969 4040 1999
rect 4037 1961 4040 1969
rect 4092 1999 4095 2007
rect 4092 1969 4122 1999
rect 4092 1961 4095 1969
rect 3538 1230 3541 1238
rect 3512 1200 3541 1230
rect 3538 1192 3541 1200
rect 3593 1230 3596 1238
rect 3593 1200 3623 1230
rect 8976 1223 8979 1231
rect 3593 1192 3596 1200
rect 8950 1193 8979 1223
rect 8976 1185 8979 1193
rect 9031 1223 9034 1231
rect 9031 1193 9061 1223
rect 9031 1185 9034 1193
<< via1 >>
rect 2930 5463 2982 5515
rect 5035 5506 5087 5515
rect 5035 5472 5044 5506
rect 5044 5472 5078 5506
rect 5078 5472 5087 5506
rect 5035 5463 5087 5472
rect 5920 4580 5972 4589
rect 5920 4546 5929 4580
rect 5929 4546 5963 4580
rect 5963 4546 5972 4580
rect 5920 4537 5972 4546
rect 2998 4454 3050 4506
rect 3066 3874 3118 3926
rect 5116 3836 5168 3845
rect 5116 3802 5125 3836
rect 5125 3802 5159 3836
rect 5159 3802 5168 3836
rect 5116 3793 5168 3802
rect 2930 3634 2982 3686
rect -12 3268 40 3320
rect 3202 3268 3254 3320
rect 3270 3018 3322 3070
rect 4576 2904 4628 2913
rect 4576 2870 4585 2904
rect 4585 2870 4619 2904
rect 4619 2870 4628 2904
rect 4576 2861 4628 2870
rect 3202 2778 3254 2830
rect 3202 2111 3254 2163
rect 4927 2158 4979 2167
rect 4927 2124 4936 2158
rect 4936 2124 4970 2158
rect 4970 2124 4979 2158
rect 4927 2115 4979 2124
rect 4040 2001 4092 2010
rect 4040 1967 4049 2001
rect 4049 1967 4083 2001
rect 4083 1967 4092 2001
rect 4040 1958 4092 1967
rect 3541 1232 3593 1241
rect 3541 1198 3550 1232
rect 3550 1198 3584 1232
rect 3584 1198 3593 1232
rect 8979 1225 9031 1234
rect 3541 1189 3593 1198
rect 8979 1191 8988 1225
rect 8988 1191 9022 1225
rect 9022 1191 9031 1225
rect 8979 1182 9031 1191
<< metal2 >>
rect 2942 5515 2970 5918
rect 2942 3686 2970 5463
rect 3010 4506 3038 5918
rect 0 1676 28 3268
rect 2942 1834 2970 3634
rect 3010 2915 3038 4454
rect 3078 3926 3106 5918
rect 180 1416 234 1444
rect 180 232 234 260
rect 2942 0 2970 1778
rect 3010 0 3038 2859
rect 3078 541 3106 3874
rect 3078 0 3106 485
rect 3146 269 3174 5918
rect 3214 3320 3242 5918
rect 3214 2830 3242 3268
rect 3282 3070 3310 5918
rect 3214 2163 3242 2778
rect 3214 901 3242 2111
rect 3282 2012 3310 3018
rect 3282 1191 3310 1956
rect 3350 1463 3378 5918
rect 5087 5475 11236 5503
rect 5972 4549 11236 4577
rect 5168 3805 11236 3833
rect 4582 2915 4622 2921
rect 4582 2853 4622 2859
rect 4046 2012 4086 2018
rect 4046 1950 4086 1956
rect 4939 1834 4967 2115
rect 3146 0 3174 213
rect 3214 0 3242 845
rect 3282 0 3310 1135
rect 3350 0 3378 1407
rect 9031 1194 11236 1222
rect 8991 901 9019 1182
<< via2 >>
rect 2996 2859 3052 2915
rect 2928 1778 2984 1834
rect 2615 1407 2671 1463
rect 2150 1135 2206 1191
rect 2150 485 2206 541
rect 2615 213 2671 269
rect 3064 485 3120 541
rect 3268 1956 3324 2012
rect 4574 2913 4630 2915
rect 4574 2861 4576 2913
rect 4576 2861 4628 2913
rect 4628 2861 4630 2913
rect 4574 2859 4630 2861
rect 4038 2010 4094 2012
rect 4038 1958 4040 2010
rect 4040 1958 4092 2010
rect 4092 1958 4094 2010
rect 4038 1956 4094 1958
rect 4925 1778 4981 1834
rect 3336 1407 3392 1463
rect 3268 1135 3324 1191
rect 3200 845 3256 901
rect 3132 213 3188 269
rect 8977 845 9033 901
<< metal3 >>
rect 2994 2915 4632 2917
rect 2994 2859 2996 2915
rect 3052 2859 4574 2915
rect 4630 2859 4632 2915
rect 2994 2857 4632 2859
rect 3266 2012 4096 2014
rect 3266 1956 3268 2012
rect 3324 1956 4038 2012
rect 4094 1956 4096 2012
rect 3266 1954 4096 1956
rect 2926 1834 4983 1836
rect 2926 1778 2928 1834
rect 2984 1778 4925 1834
rect 4981 1778 4983 1834
rect 2926 1776 4983 1778
rect -30 1646 30 1706
rect 2613 1463 3394 1465
rect 2613 1407 2615 1463
rect 2671 1407 3336 1463
rect 3392 1407 3394 1463
rect 2613 1405 3394 1407
rect 2148 1191 3326 1193
rect 2148 1135 2150 1191
rect 2206 1135 3268 1191
rect 3324 1135 3326 1191
rect 2148 1133 3326 1135
rect 3198 901 9035 903
rect -30 808 30 868
rect 3198 845 3200 901
rect 3256 845 8977 901
rect 9033 845 9035 901
rect 3198 843 9035 845
rect 2148 541 3122 543
rect 2148 485 2150 541
rect 2206 485 3064 541
rect 3120 485 3122 541
rect 2148 483 3122 485
rect 2613 269 3190 271
rect 2613 213 2615 269
rect 2671 213 3132 269
rect 3188 213 3190 269
rect 2613 211 3190 213
rect -30 -30 30 30
use contact_17  contact_17_0
timestamp 1643671299
transform 1 0 4587 0 1 2872
box 0 0 1 1
use contact_13  contact_13_0
timestamp 1643671299
transform 1 0 4573 0 1 2864
box 0 0 1 1
use contact_18  contact_18_0
timestamp 1643671299
transform 1 0 4572 0 1 2857
box 0 0 1 1
use contact_17  contact_17_1
timestamp 1643671299
transform 1 0 4587 0 1 2872
box 0 0 1 1
use contact_13  contact_13_1
timestamp 1643671299
transform 1 0 4573 0 1 2864
box 0 0 1 1
use contact_30  contact_30_0
timestamp 1643671299
transform 1 0 2994 0 1 2857
box 0 0 1 1
use contact_13  contact_13_2
timestamp 1643671299
transform 1 0 3686 0 1 3021
box 0 0 1 1
use contact_17  contact_17_2
timestamp 1643671299
transform 1 0 3281 0 1 3029
box 0 0 1 1
use contact_13  contact_13_3
timestamp 1643671299
transform 1 0 3586 0 1 2781
box 0 0 1 1
use contact_17  contact_17_3
timestamp 1643671299
transform 1 0 3213 0 1 2789
box 0 0 1 1
use contact_17  contact_17_4
timestamp 1643671299
transform 1 0 4938 0 1 2126
box 0 0 1 1
use contact_13  contact_13_4
timestamp 1643671299
transform 1 0 4924 0 1 2118
box 0 0 1 1
use contact_30  contact_30_1
timestamp 1643671299
transform 1 0 2926 0 1 1776
box 0 0 1 1
use contact_30  contact_30_2
timestamp 1643671299
transform 1 0 4923 0 1 1776
box 0 0 1 1
use contact_18  contact_18_1
timestamp 1643671299
transform 1 0 4036 0 1 1954
box 0 0 1 1
use contact_17  contact_17_5
timestamp 1643671299
transform 1 0 4051 0 1 1969
box 0 0 1 1
use contact_13  contact_13_5
timestamp 1643671299
transform 1 0 4037 0 1 1961
box 0 0 1 1
use contact_18  contact_18_2
timestamp 1643671299
transform 1 0 4036 0 1 1954
box 0 0 1 1
use contact_17  contact_17_6
timestamp 1643671299
transform 1 0 4051 0 1 1969
box 0 0 1 1
use contact_13  contact_13_6
timestamp 1643671299
transform 1 0 4037 0 1 1961
box 0 0 1 1
use contact_30  contact_30_3
timestamp 1643671299
transform 1 0 3266 0 1 1954
box 0 0 1 1
use contact_13  contact_13_7
timestamp 1643671299
transform 1 0 3538 0 1 2114
box 0 0 1 1
use contact_17  contact_17_7
timestamp 1643671299
transform 1 0 3213 0 1 2122
box 0 0 1 1
use contact_17  contact_17_8
timestamp 1643671299
transform 1 0 8990 0 1 1193
box 0 0 1 1
use contact_13  contact_13_8
timestamp 1643671299
transform 1 0 8976 0 1 1185
box 0 0 1 1
use contact_17  contact_17_9
timestamp 1643671299
transform 1 0 8990 0 1 1193
box 0 0 1 1
use contact_13  contact_13_9
timestamp 1643671299
transform 1 0 8976 0 1 1185
box 0 0 1 1
use contact_30  contact_30_4
timestamp 1643671299
transform 1 0 3198 0 1 843
box 0 0 1 1
use contact_30  contact_30_5
timestamp 1643671299
transform 1 0 8975 0 1 843
box 0 0 1 1
use contact_17  contact_17_10
timestamp 1643671299
transform 1 0 3552 0 1 1200
box 0 0 1 1
use contact_13  contact_13_10
timestamp 1643671299
transform 1 0 3538 0 1 1192
box 0 0 1 1
use contact_17  contact_17_11
timestamp 1643671299
transform 1 0 5931 0 1 4548
box 0 0 1 1
use contact_13  contact_13_11
timestamp 1643671299
transform 1 0 5917 0 1 4540
box 0 0 1 1
use contact_13  contact_13_12
timestamp 1643671299
transform 1 0 3586 0 1 4457
box 0 0 1 1
use contact_17  contact_17_12
timestamp 1643671299
transform 1 0 3009 0 1 4465
box 0 0 1 1
use contact_17  contact_17_13
timestamp 1643671299
transform 1 0 5127 0 1 3804
box 0 0 1 1
use contact_13  contact_13_13
timestamp 1643671299
transform 1 0 5113 0 1 3796
box 0 0 1 1
use contact_13  contact_13_14
timestamp 1643671299
transform 1 0 3686 0 1 3637
box 0 0 1 1
use contact_17  contact_17_14
timestamp 1643671299
transform 1 0 2941 0 1 3645
box 0 0 1 1
use contact_13  contact_13_15
timestamp 1643671299
transform 1 0 3586 0 1 3877
box 0 0 1 1
use contact_17  contact_17_15
timestamp 1643671299
transform 1 0 3077 0 1 3885
box 0 0 1 1
use contact_17  contact_17_16
timestamp 1643671299
transform 1 0 5046 0 1 5474
box 0 0 1 1
use contact_13  contact_13_16
timestamp 1643671299
transform 1 0 5032 0 1 5466
box 0 0 1 1
use contact_13  contact_13_17
timestamp 1643671299
transform 1 0 3538 0 1 5466
box 0 0 1 1
use contact_17  contact_17_17
timestamp 1643671299
transform 1 0 2941 0 1 5474
box 0 0 1 1
use contact_17  contact_17_18
timestamp 1643671299
transform 1 0 3213 0 1 3279
box 0 0 1 1
use contact_17  contact_17_19
timestamp 1643671299
transform 1 0 -1 0 1 3279
box 0 0 1 1
use contact_18  contact_18_3
timestamp 1643671299
transform 1 0 2613 0 1 1405
box 0 0 1 1
use contact_30  contact_30_6
timestamp 1643671299
transform 1 0 3334 0 1 1405
box 0 0 1 1
use contact_18  contact_18_4
timestamp 1643671299
transform 1 0 2148 0 1 1133
box 0 0 1 1
use contact_30  contact_30_7
timestamp 1643671299
transform 1 0 3266 0 1 1133
box 0 0 1 1
use contact_18  contact_18_5
timestamp 1643671299
transform 1 0 2613 0 1 211
box 0 0 1 1
use contact_30  contact_30_8
timestamp 1643671299
transform 1 0 3130 0 1 211
box 0 0 1 1
use contact_18  contact_18_6
timestamp 1643671299
transform 1 0 2148 0 1 483
box 0 0 1 1
use contact_30  contact_30_9
timestamp 1643671299
transform 1 0 3062 0 1 483
box 0 0 1 1
use pdriver_3  pdriver_3_0
timestamp 1643671299
transform 1 0 3937 0 1 4190
box -36 -17 2736 895
use pnand2_1  pnand2_1_0
timestamp 1643671299
transform 1 0 3486 0 1 4190
box -36 -17 487 895
use pand2_0  pand2_0_0
timestamp 1643671299
transform 1 0 3486 0 -1 4190
box -36 -17 2925 895
use pdriver_1  pdriver_1_0
timestamp 1643671299
transform 1 0 3486 0 -1 5866
box -36 -17 1980 895
use pand2  pand2_0
timestamp 1643671299
transform 1 0 3486 0 1 2514
box -36 -17 1845 895
use pand2  pand2_1
timestamp 1643671299
transform 1 0 3837 0 -1 2514
box -36 -17 1845 895
use pinv_0  pinv_0_0
timestamp 1643671299
transform 1 0 3486 0 -1 2514
box -36 -17 387 895
use pdriver_0  pdriver_0_0
timestamp 1643671299
transform 1 0 3486 0 1 838
box -36 -17 7650 895
use dff_buf_array  dff_buf_array_0
timestamp 1643671299
transform 1 0 0 0 1 0
box -30 -42 2978 1718
<< labels >>
rlabel metal2 s 180 1416 234 1444 4 csb
rlabel metal2 s 180 232 234 260 4 web
rlabel metal2 s 5061 5475 11236 5503 4 wl_en
rlabel metal2 s 5142 3805 11236 3833 4 w_en
rlabel metal2 s 5946 4549 11236 4577 4 p_en_bar
rlabel metal2 s 3553 1201 3581 1229 4 clk
rlabel metal2 s 9005 1194 11236 1222 4 clk_buf
rlabel metal3 s -30 1646 30 1706 4 gnd
rlabel metal3 s -30 -30 30 30 4 gnd
rlabel metal3 s -30 808 30 868 4 vdd
<< properties >>
string FIXED_BBOX 0 0 11236 116
string GDS_FILE sram_0rw2r1w_16_32_sky130A.gds
string GDS_END 1117480
string GDS_START 1108770
<< end >>
