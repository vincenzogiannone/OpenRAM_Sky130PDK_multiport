magic
tech sky130A
magscale 1 2
timestamp 1643678851
<< checkpaint >>
rect -1260 -1286 1410 1958
<< scnmos >>
rect 60 0 90 672
<< ndiff >>
rect 0 353 60 672
rect 0 319 8 353
rect 42 319 60 353
rect 0 0 60 319
rect 90 353 150 672
rect 90 319 108 353
rect 142 319 150 353
rect 90 0 150 319
<< ndiffc >>
rect 8 319 42 353
rect 108 319 142 353
<< poly >>
rect 60 672 90 698
rect 60 -26 90 0
<< locali >>
rect 8 353 42 369
rect 8 303 42 319
rect 108 353 142 369
rect 108 303 142 319
use contact_8  contact_8_0
timestamp 1643678851
transform 1 0 100 0 1 295
box 0 0 1 1
use contact_8  contact_8_1
timestamp 1643678851
transform 1 0 0 0 1 295
box 0 0 1 1
<< labels >>
rlabel mvvaractor s 75 336 75 336 4 G
rlabel locali s 25 336 25 336 4 S
rlabel locali s 125 336 125 336 4 D
<< properties >>
string FIXED_BBOX -25 -26 175 698
string GDS_FILE sram_0rw2r1w_16_128_sky130A.gds
string GDS_END 1626692
string GDS_START 1625928
<< end >>
