magic
tech sky130A
magscale 1 2
timestamp 1644951705
<< checkpaint >>
rect -1299 -1302 4224 2176
<< metal1 >>
rect 709 812 715 864
rect 767 812 773 864
rect 2191 812 2197 864
rect 2249 812 2255 864
rect 709 -26 715 26
rect 767 -26 773 26
rect 2191 -26 2197 26
rect 2249 -26 2255 26
<< via1 >>
rect 715 812 767 864
rect 2197 812 2249 864
rect 715 -26 767 26
rect 2197 -26 2249 26
<< metal2 >>
rect 713 866 769 875
rect 0 345 28 838
rect 2195 866 2251 875
rect 713 801 769 810
rect 1482 345 1510 838
rect 2195 801 2251 810
rect -1 336 55 345
rect -1 271 55 280
rect 1481 336 1537 345
rect 1481 271 1537 280
rect 0 0 28 271
rect 180 232 234 260
rect 1260 228 1314 256
rect 713 28 769 37
rect 1482 0 1510 271
rect 1662 232 1716 260
rect 2742 228 2796 256
rect 2195 28 2251 37
rect 713 -37 769 -28
rect 2195 -37 2251 -28
<< via2 >>
rect 713 864 769 866
rect 713 812 715 864
rect 715 812 767 864
rect 767 812 769 864
rect 2195 864 2251 866
rect 713 810 769 812
rect 2195 812 2197 864
rect 2197 812 2249 864
rect 2249 812 2251 864
rect 2195 810 2251 812
rect -1 280 55 336
rect 1481 280 1537 336
rect 713 26 769 28
rect 713 -26 715 26
rect 715 -26 767 26
rect 767 -26 769 26
rect 2195 26 2251 28
rect 713 -28 769 -26
rect 2195 -26 2197 26
rect 2197 -26 2249 26
rect 2249 -26 2251 26
rect 2195 -28 2251 -26
<< metal3 >>
rect 675 866 807 875
rect 675 810 713 866
rect 769 810 807 866
rect 675 801 807 810
rect 2157 866 2289 875
rect 2157 810 2195 866
rect 2251 810 2289 866
rect 2157 801 2289 810
rect -39 338 93 341
rect 1443 338 1575 341
rect -39 336 2964 338
rect -39 280 -1 336
rect 55 280 1481 336
rect 1537 280 2964 336
rect -39 278 2964 280
rect -39 275 93 278
rect 1443 275 1575 278
rect 675 28 807 37
rect 675 -28 713 28
rect 769 -28 807 28
rect 675 -37 807 -28
rect 2157 28 2289 37
rect 2157 -28 2195 28
rect 2251 -28 2289 28
rect 2157 -37 2289 -28
use contact_18  contact_18_0
timestamp 1644951705
transform 1 0 1443 0 1 271
box 0 0 1 1
use contact_18  contact_18_1
timestamp 1644951705
transform 1 0 -39 0 1 271
box 0 0 1 1
use contact_18  contact_18_2
timestamp 1644951705
transform 1 0 2157 0 1 -37
box 0 0 1 1
use contact_17  contact_17_0
timestamp 1644951705
transform 1 0 2191 0 1 -32
box 0 0 1 1
use contact_18  contact_18_3
timestamp 1644951705
transform 1 0 2157 0 1 801
box 0 0 1 1
use contact_17  contact_17_1
timestamp 1644951705
transform 1 0 2191 0 1 806
box 0 0 1 1
use contact_18  contact_18_4
timestamp 1644951705
transform 1 0 675 0 1 -37
box 0 0 1 1
use contact_17  contact_17_2
timestamp 1644951705
transform 1 0 709 0 1 -32
box 0 0 1 1
use contact_18  contact_18_5
timestamp 1644951705
transform 1 0 675 0 1 801
box 0 0 1 1
use contact_17  contact_17_3
timestamp 1644951705
transform 1 0 709 0 1 806
box 0 0 1 1
use dff  dff_0
timestamp 1644951705
transform 1 0 1482 0 1 0
box 0 -42 1482 916
use dff  dff_1
timestamp 1644951705
transform 1 0 0 0 1 0
box 0 -42 1482 916
<< labels >>
rlabel metal3 s 2157 801 2289 875 4 vdd
rlabel metal3 s 675 801 807 875 4 vdd
rlabel metal3 s 675 -37 807 37 4 gnd
rlabel metal3 s 2157 -37 2289 37 4 gnd
rlabel metal2 s 180 232 234 260 4 din_0
rlabel metal2 s 1260 228 1314 256 4 dout_0
rlabel metal2 s 1662 232 1716 260 4 din_1
rlabel metal2 s 2742 228 2796 256 4 dout_1
rlabel metal3 s 0 278 2964 338 4 clk
<< properties >>
string FIXED_BBOX 2157 -37 2289 0
string GDS_FILE sram_0rw2r1w_16_128_sky130A.gds
string GDS_END 2088022
string GDS_START 2085356
<< end >>
