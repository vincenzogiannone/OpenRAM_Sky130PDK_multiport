magic
tech sky130A
magscale 1 2
timestamp 1643671299
<< checkpaint >>
rect -1319 -1316 5249 1608
<< nwell >>
rect -54 231 3984 348
rect -59 63 3989 231
rect -54 -54 3984 63
<< scpmos >>
rect 60 0 90 294
rect 168 0 198 294
rect 276 0 306 294
rect 384 0 414 294
rect 492 0 522 294
rect 600 0 630 294
rect 708 0 738 294
rect 816 0 846 294
rect 924 0 954 294
rect 1032 0 1062 294
rect 1140 0 1170 294
rect 1248 0 1278 294
rect 1356 0 1386 294
rect 1464 0 1494 294
rect 1572 0 1602 294
rect 1680 0 1710 294
rect 1788 0 1818 294
rect 1896 0 1926 294
rect 2004 0 2034 294
rect 2112 0 2142 294
rect 2220 0 2250 294
rect 2328 0 2358 294
rect 2436 0 2466 294
rect 2544 0 2574 294
rect 2652 0 2682 294
rect 2760 0 2790 294
rect 2868 0 2898 294
rect 2976 0 3006 294
rect 3084 0 3114 294
rect 3192 0 3222 294
rect 3300 0 3330 294
rect 3408 0 3438 294
rect 3516 0 3546 294
rect 3624 0 3654 294
rect 3732 0 3762 294
rect 3840 0 3870 294
<< pdiff >>
rect 0 164 60 294
rect 0 130 8 164
rect 42 130 60 164
rect 0 0 60 130
rect 90 164 168 294
rect 90 130 112 164
rect 146 130 168 164
rect 90 0 168 130
rect 198 164 276 294
rect 198 130 220 164
rect 254 130 276 164
rect 198 0 276 130
rect 306 164 384 294
rect 306 130 328 164
rect 362 130 384 164
rect 306 0 384 130
rect 414 164 492 294
rect 414 130 436 164
rect 470 130 492 164
rect 414 0 492 130
rect 522 164 600 294
rect 522 130 544 164
rect 578 130 600 164
rect 522 0 600 130
rect 630 164 708 294
rect 630 130 652 164
rect 686 130 708 164
rect 630 0 708 130
rect 738 164 816 294
rect 738 130 760 164
rect 794 130 816 164
rect 738 0 816 130
rect 846 164 924 294
rect 846 130 868 164
rect 902 130 924 164
rect 846 0 924 130
rect 954 164 1032 294
rect 954 130 976 164
rect 1010 130 1032 164
rect 954 0 1032 130
rect 1062 164 1140 294
rect 1062 130 1084 164
rect 1118 130 1140 164
rect 1062 0 1140 130
rect 1170 164 1248 294
rect 1170 130 1192 164
rect 1226 130 1248 164
rect 1170 0 1248 130
rect 1278 164 1356 294
rect 1278 130 1300 164
rect 1334 130 1356 164
rect 1278 0 1356 130
rect 1386 164 1464 294
rect 1386 130 1408 164
rect 1442 130 1464 164
rect 1386 0 1464 130
rect 1494 164 1572 294
rect 1494 130 1516 164
rect 1550 130 1572 164
rect 1494 0 1572 130
rect 1602 164 1680 294
rect 1602 130 1624 164
rect 1658 130 1680 164
rect 1602 0 1680 130
rect 1710 164 1788 294
rect 1710 130 1732 164
rect 1766 130 1788 164
rect 1710 0 1788 130
rect 1818 164 1896 294
rect 1818 130 1840 164
rect 1874 130 1896 164
rect 1818 0 1896 130
rect 1926 164 2004 294
rect 1926 130 1948 164
rect 1982 130 2004 164
rect 1926 0 2004 130
rect 2034 164 2112 294
rect 2034 130 2056 164
rect 2090 130 2112 164
rect 2034 0 2112 130
rect 2142 164 2220 294
rect 2142 130 2164 164
rect 2198 130 2220 164
rect 2142 0 2220 130
rect 2250 164 2328 294
rect 2250 130 2272 164
rect 2306 130 2328 164
rect 2250 0 2328 130
rect 2358 164 2436 294
rect 2358 130 2380 164
rect 2414 130 2436 164
rect 2358 0 2436 130
rect 2466 164 2544 294
rect 2466 130 2488 164
rect 2522 130 2544 164
rect 2466 0 2544 130
rect 2574 164 2652 294
rect 2574 130 2596 164
rect 2630 130 2652 164
rect 2574 0 2652 130
rect 2682 164 2760 294
rect 2682 130 2704 164
rect 2738 130 2760 164
rect 2682 0 2760 130
rect 2790 164 2868 294
rect 2790 130 2812 164
rect 2846 130 2868 164
rect 2790 0 2868 130
rect 2898 164 2976 294
rect 2898 130 2920 164
rect 2954 130 2976 164
rect 2898 0 2976 130
rect 3006 164 3084 294
rect 3006 130 3028 164
rect 3062 130 3084 164
rect 3006 0 3084 130
rect 3114 164 3192 294
rect 3114 130 3136 164
rect 3170 130 3192 164
rect 3114 0 3192 130
rect 3222 164 3300 294
rect 3222 130 3244 164
rect 3278 130 3300 164
rect 3222 0 3300 130
rect 3330 164 3408 294
rect 3330 130 3352 164
rect 3386 130 3408 164
rect 3330 0 3408 130
rect 3438 164 3516 294
rect 3438 130 3460 164
rect 3494 130 3516 164
rect 3438 0 3516 130
rect 3546 164 3624 294
rect 3546 130 3568 164
rect 3602 130 3624 164
rect 3546 0 3624 130
rect 3654 164 3732 294
rect 3654 130 3676 164
rect 3710 130 3732 164
rect 3654 0 3732 130
rect 3762 164 3840 294
rect 3762 130 3784 164
rect 3818 130 3840 164
rect 3762 0 3840 130
rect 3870 164 3930 294
rect 3870 130 3888 164
rect 3922 130 3930 164
rect 3870 0 3930 130
<< pdiffc >>
rect 8 130 42 164
rect 112 130 146 164
rect 220 130 254 164
rect 328 130 362 164
rect 436 130 470 164
rect 544 130 578 164
rect 652 130 686 164
rect 760 130 794 164
rect 868 130 902 164
rect 976 130 1010 164
rect 1084 130 1118 164
rect 1192 130 1226 164
rect 1300 130 1334 164
rect 1408 130 1442 164
rect 1516 130 1550 164
rect 1624 130 1658 164
rect 1732 130 1766 164
rect 1840 130 1874 164
rect 1948 130 1982 164
rect 2056 130 2090 164
rect 2164 130 2198 164
rect 2272 130 2306 164
rect 2380 130 2414 164
rect 2488 130 2522 164
rect 2596 130 2630 164
rect 2704 130 2738 164
rect 2812 130 2846 164
rect 2920 130 2954 164
rect 3028 130 3062 164
rect 3136 130 3170 164
rect 3244 130 3278 164
rect 3352 130 3386 164
rect 3460 130 3494 164
rect 3568 130 3602 164
rect 3676 130 3710 164
rect 3784 130 3818 164
rect 3888 130 3922 164
<< poly >>
rect 60 294 90 320
rect 168 294 198 320
rect 276 294 306 320
rect 384 294 414 320
rect 492 294 522 320
rect 600 294 630 320
rect 708 294 738 320
rect 816 294 846 320
rect 924 294 954 320
rect 1032 294 1062 320
rect 1140 294 1170 320
rect 1248 294 1278 320
rect 1356 294 1386 320
rect 1464 294 1494 320
rect 1572 294 1602 320
rect 1680 294 1710 320
rect 1788 294 1818 320
rect 1896 294 1926 320
rect 2004 294 2034 320
rect 2112 294 2142 320
rect 2220 294 2250 320
rect 2328 294 2358 320
rect 2436 294 2466 320
rect 2544 294 2574 320
rect 2652 294 2682 320
rect 2760 294 2790 320
rect 2868 294 2898 320
rect 2976 294 3006 320
rect 3084 294 3114 320
rect 3192 294 3222 320
rect 3300 294 3330 320
rect 3408 294 3438 320
rect 3516 294 3546 320
rect 3624 294 3654 320
rect 3732 294 3762 320
rect 3840 294 3870 320
rect 60 -26 90 0
rect 168 -26 198 0
rect 276 -26 306 0
rect 384 -26 414 0
rect 492 -26 522 0
rect 600 -26 630 0
rect 708 -26 738 0
rect 816 -26 846 0
rect 924 -26 954 0
rect 1032 -26 1062 0
rect 1140 -26 1170 0
rect 1248 -26 1278 0
rect 1356 -26 1386 0
rect 1464 -26 1494 0
rect 1572 -26 1602 0
rect 1680 -26 1710 0
rect 1788 -26 1818 0
rect 1896 -26 1926 0
rect 2004 -26 2034 0
rect 2112 -26 2142 0
rect 2220 -26 2250 0
rect 2328 -26 2358 0
rect 2436 -26 2466 0
rect 2544 -26 2574 0
rect 2652 -26 2682 0
rect 2760 -26 2790 0
rect 2868 -26 2898 0
rect 2976 -26 3006 0
rect 3084 -26 3114 0
rect 3192 -26 3222 0
rect 3300 -26 3330 0
rect 3408 -26 3438 0
rect 3516 -26 3546 0
rect 3624 -26 3654 0
rect 3732 -26 3762 0
rect 3840 -26 3870 0
rect 60 -56 3870 -26
<< locali >>
rect 8 164 42 180
rect 8 114 42 130
rect 112 164 146 180
rect 112 80 146 130
rect 220 164 254 180
rect 220 114 254 130
rect 328 164 362 180
rect 328 80 362 130
rect 436 164 470 180
rect 436 114 470 130
rect 544 164 578 180
rect 544 80 578 130
rect 652 164 686 180
rect 652 114 686 130
rect 760 164 794 180
rect 760 80 794 130
rect 868 164 902 180
rect 868 114 902 130
rect 976 164 1010 180
rect 976 80 1010 130
rect 1084 164 1118 180
rect 1084 114 1118 130
rect 1192 164 1226 180
rect 1192 80 1226 130
rect 1300 164 1334 180
rect 1300 114 1334 130
rect 1408 164 1442 180
rect 1408 80 1442 130
rect 1516 164 1550 180
rect 1516 114 1550 130
rect 1624 164 1658 180
rect 1624 80 1658 130
rect 1732 164 1766 180
rect 1732 114 1766 130
rect 1840 164 1874 180
rect 1840 80 1874 130
rect 1948 164 1982 180
rect 1948 114 1982 130
rect 2056 164 2090 180
rect 2056 80 2090 130
rect 2164 164 2198 180
rect 2164 114 2198 130
rect 2272 164 2306 180
rect 2272 80 2306 130
rect 2380 164 2414 180
rect 2380 114 2414 130
rect 2488 164 2522 180
rect 2488 80 2522 130
rect 2596 164 2630 180
rect 2596 114 2630 130
rect 2704 164 2738 180
rect 2704 80 2738 130
rect 2812 164 2846 180
rect 2812 114 2846 130
rect 2920 164 2954 180
rect 2920 80 2954 130
rect 3028 164 3062 180
rect 3028 114 3062 130
rect 3136 164 3170 180
rect 3136 80 3170 130
rect 3244 164 3278 180
rect 3244 114 3278 130
rect 3352 164 3386 180
rect 3352 80 3386 130
rect 3460 164 3494 180
rect 3460 114 3494 130
rect 3568 164 3602 180
rect 3568 80 3602 130
rect 3676 164 3710 180
rect 3676 114 3710 130
rect 3784 164 3818 180
rect 3784 80 3818 130
rect 3888 164 3922 180
rect 3888 114 3922 130
rect 112 46 3818 80
use contact_9  contact_9_0
timestamp 1643671299
transform 1 0 3880 0 1 106
box 0 0 2 2
use contact_9  contact_9_1
timestamp 1643671299
transform 1 0 3776 0 1 106
box 0 0 2 2
use contact_9  contact_9_2
timestamp 1643671299
transform 1 0 3668 0 1 106
box 0 0 2 2
use contact_9  contact_9_3
timestamp 1643671299
transform 1 0 3560 0 1 106
box 0 0 2 2
use contact_9  contact_9_4
timestamp 1643671299
transform 1 0 3452 0 1 106
box 0 0 2 2
use contact_9  contact_9_5
timestamp 1643671299
transform 1 0 3344 0 1 106
box 0 0 2 2
use contact_9  contact_9_6
timestamp 1643671299
transform 1 0 3236 0 1 106
box 0 0 2 2
use contact_9  contact_9_7
timestamp 1643671299
transform 1 0 3128 0 1 106
box 0 0 2 2
use contact_9  contact_9_8
timestamp 1643671299
transform 1 0 3020 0 1 106
box 0 0 2 2
use contact_9  contact_9_9
timestamp 1643671299
transform 1 0 2912 0 1 106
box 0 0 2 2
use contact_9  contact_9_10
timestamp 1643671299
transform 1 0 2804 0 1 106
box 0 0 2 2
use contact_9  contact_9_11
timestamp 1643671299
transform 1 0 2696 0 1 106
box 0 0 2 2
use contact_9  contact_9_12
timestamp 1643671299
transform 1 0 2588 0 1 106
box 0 0 2 2
use contact_9  contact_9_13
timestamp 1643671299
transform 1 0 2480 0 1 106
box 0 0 2 2
use contact_9  contact_9_14
timestamp 1643671299
transform 1 0 2372 0 1 106
box 0 0 2 2
use contact_9  contact_9_15
timestamp 1643671299
transform 1 0 2264 0 1 106
box 0 0 2 2
use contact_9  contact_9_16
timestamp 1643671299
transform 1 0 2156 0 1 106
box 0 0 2 2
use contact_9  contact_9_17
timestamp 1643671299
transform 1 0 2048 0 1 106
box 0 0 2 2
use contact_9  contact_9_18
timestamp 1643671299
transform 1 0 1940 0 1 106
box 0 0 2 2
use contact_9  contact_9_19
timestamp 1643671299
transform 1 0 1832 0 1 106
box 0 0 2 2
use contact_9  contact_9_20
timestamp 1643671299
transform 1 0 1724 0 1 106
box 0 0 2 2
use contact_9  contact_9_21
timestamp 1643671299
transform 1 0 1616 0 1 106
box 0 0 2 2
use contact_9  contact_9_22
timestamp 1643671299
transform 1 0 1508 0 1 106
box 0 0 2 2
use contact_9  contact_9_23
timestamp 1643671299
transform 1 0 1400 0 1 106
box 0 0 2 2
use contact_9  contact_9_24
timestamp 1643671299
transform 1 0 1292 0 1 106
box 0 0 2 2
use contact_9  contact_9_25
timestamp 1643671299
transform 1 0 1184 0 1 106
box 0 0 2 2
use contact_9  contact_9_26
timestamp 1643671299
transform 1 0 1076 0 1 106
box 0 0 2 2
use contact_9  contact_9_27
timestamp 1643671299
transform 1 0 968 0 1 106
box 0 0 2 2
use contact_9  contact_9_28
timestamp 1643671299
transform 1 0 860 0 1 106
box 0 0 2 2
use contact_9  contact_9_29
timestamp 1643671299
transform 1 0 752 0 1 106
box 0 0 2 2
use contact_9  contact_9_30
timestamp 1643671299
transform 1 0 644 0 1 106
box 0 0 2 2
use contact_9  contact_9_31
timestamp 1643671299
transform 1 0 536 0 1 106
box 0 0 2 2
use contact_9  contact_9_32
timestamp 1643671299
transform 1 0 428 0 1 106
box 0 0 2 2
use contact_9  contact_9_33
timestamp 1643671299
transform 1 0 320 0 1 106
box 0 0 2 2
use contact_9  contact_9_34
timestamp 1643671299
transform 1 0 212 0 1 106
box 0 0 2 2
use contact_9  contact_9_35
timestamp 1643671299
transform 1 0 104 0 1 106
box 0 0 2 2
use contact_9  contact_9_36
timestamp 1643671299
transform 1 0 0 0 1 106
box 0 0 2 2
<< labels >>
rlabel mvvaractor s 1965 -41 1965 -41 4 G
rlabel locali s 885 147 885 147 4 S
rlabel locali s 1101 147 1101 147 4 S
rlabel locali s 237 147 237 147 4 S
rlabel locali s 2397 147 2397 147 4 S
rlabel locali s 1965 147 1965 147 4 S
rlabel locali s 669 147 669 147 4 S
rlabel locali s 453 147 453 147 4 S
rlabel locali s 1533 147 1533 147 4 S
rlabel locali s 1317 147 1317 147 4 S
rlabel locali s 1749 147 1749 147 4 S
rlabel locali s 2181 147 2181 147 4 S
rlabel locali s 3477 147 3477 147 4 S
rlabel locali s 2613 147 2613 147 4 S
rlabel locali s 3905 147 3905 147 4 S
rlabel locali s 3693 147 3693 147 4 S
rlabel locali s 3045 147 3045 147 4 S
rlabel locali s 3261 147 3261 147 4 S
rlabel locali s 25 147 25 147 4 S
rlabel locali s 2829 147 2829 147 4 S
rlabel locali s 1965 63 1965 63 4 D
<< properties >>
string FIXED_BBOX -54 -56 3984 63
string GDS_FILE sram_0rw2r1w_16_32_sky130A.gds
string GDS_END 1174530
string GDS_START 1166750
<< end >>
