magic
tech sky130A
timestamp 1643678851
<< checkpaint >>
rect -630 -651 25526 25291
<< metal1 >>
rect 0 24625 24896 24656
rect 0 24304 24896 24318
rect 0 24241 24896 24255
rect 0 24128 24896 24142
rect 0 23854 24896 23886
rect 0 23598 24896 23612
rect 0 23485 24896 23499
rect 0 23422 24896 23436
rect 0 23084 24896 23116
rect 0 22764 24896 22778
rect 0 22701 24896 22715
rect 0 22588 24896 22602
rect 0 22314 24896 22346
rect 0 22058 24896 22072
rect 0 21945 24896 21959
rect 0 21882 24896 21896
rect 0 21544 24896 21576
rect 0 21224 24896 21238
rect 0 21161 24896 21175
rect 0 21048 24896 21062
rect 0 20774 24896 20806
rect 0 20518 24896 20532
rect 0 20405 24896 20419
rect 0 20342 24896 20356
rect 0 20004 24896 20036
rect 0 19684 24896 19698
rect 0 19621 24896 19635
rect 0 19508 24896 19522
rect 0 19234 24896 19266
rect 0 18978 24896 18992
rect 0 18865 24896 18879
rect 0 18802 24896 18816
rect 0 18464 24896 18496
rect 0 18144 24896 18158
rect 0 18081 24896 18095
rect 0 17968 24896 17982
rect 0 17694 24896 17726
rect 0 17438 24896 17452
rect 0 17325 24896 17339
rect 0 17262 24896 17276
rect 0 16924 24896 16956
rect 0 16604 24896 16618
rect 0 16541 24896 16555
rect 0 16428 24896 16442
rect 0 16154 24896 16186
rect 0 15898 24896 15912
rect 0 15785 24896 15799
rect 0 15722 24896 15736
rect 0 15384 24896 15416
rect 0 15064 24896 15078
rect 0 15001 24896 15015
rect 0 14888 24896 14902
rect 0 14614 24896 14646
rect 0 14358 24896 14372
rect 0 14245 24896 14259
rect 0 14182 24896 14196
rect 0 13844 24896 13876
rect 0 13524 24896 13538
rect 0 13461 24896 13475
rect 0 13348 24896 13362
rect 0 13074 24896 13106
rect 0 12818 24896 12832
rect 0 12705 24896 12719
rect 0 12642 24896 12656
rect 0 12304 24896 12336
rect 0 11984 24896 11998
rect 0 11921 24896 11935
rect 0 11808 24896 11822
rect 0 11534 24896 11566
rect 0 11278 24896 11292
rect 0 11165 24896 11179
rect 0 11102 24896 11116
rect 0 10764 24896 10796
rect 0 10444 24896 10458
rect 0 10381 24896 10395
rect 0 10268 24896 10282
rect 0 9994 24896 10026
rect 0 9738 24896 9752
rect 0 9625 24896 9639
rect 0 9562 24896 9576
rect 0 9224 24896 9256
rect 0 8904 24896 8918
rect 0 8841 24896 8855
rect 0 8728 24896 8742
rect 0 8454 24896 8486
rect 0 8198 24896 8212
rect 0 8085 24896 8099
rect 0 8022 24896 8036
rect 0 7684 24896 7716
rect 0 7364 24896 7378
rect 0 7301 24896 7315
rect 0 7188 24896 7202
rect 0 6914 24896 6946
rect 0 6658 24896 6672
rect 0 6545 24896 6559
rect 0 6482 24896 6496
rect 0 6144 24896 6176
rect 0 5824 24896 5838
rect 0 5761 24896 5775
rect 0 5648 24896 5662
rect 0 5374 24896 5406
rect 0 5118 24896 5132
rect 0 5005 24896 5019
rect 0 4942 24896 4956
rect 0 4604 24896 4636
rect 0 4284 24896 4298
rect 0 4221 24896 4235
rect 0 4108 24896 4122
rect 0 3834 24896 3866
rect 0 3578 24896 3592
rect 0 3465 24896 3479
rect 0 3402 24896 3416
rect 0 3064 24896 3096
rect 0 2744 24896 2758
rect 0 2681 24896 2695
rect 0 2568 24896 2582
rect 0 2294 24896 2326
rect 0 2038 24896 2052
rect 0 1925 24896 1939
rect 0 1862 24896 1876
rect 0 1524 24896 1556
rect 0 1204 24896 1218
rect 0 1141 24896 1155
rect 0 1028 24896 1042
rect 0 754 24896 786
rect 0 498 24896 512
rect 0 385 24896 399
rect 0 322 24896 336
rect 0 -16 24896 15
<< metal2 >>
rect 96 0 110 24640
rect 222 0 236 24640
rect 313 0 327 24640
rect 485 0 499 24640
rect 611 0 625 24640
rect 702 0 716 24640
rect 874 0 888 24640
rect 1000 0 1014 24640
rect 1091 0 1105 24640
rect 1263 0 1277 24640
rect 1389 0 1403 24640
rect 1480 0 1494 24640
rect 1652 0 1666 24640
rect 1778 0 1792 24640
rect 1869 0 1883 24640
rect 2041 0 2055 24640
rect 2167 0 2181 24640
rect 2258 0 2272 24640
rect 2430 0 2444 24640
rect 2556 0 2570 24640
rect 2647 0 2661 24640
rect 2819 0 2833 24640
rect 2945 0 2959 24640
rect 3036 0 3050 24640
rect 3208 0 3222 24640
rect 3334 0 3348 24640
rect 3425 0 3439 24640
rect 3597 0 3611 24640
rect 3723 0 3737 24640
rect 3814 0 3828 24640
rect 3986 0 4000 24640
rect 4112 0 4126 24640
rect 4203 0 4217 24640
rect 4375 0 4389 24640
rect 4501 0 4515 24640
rect 4592 0 4606 24640
rect 4764 0 4778 24640
rect 4890 0 4904 24640
rect 4981 0 4995 24640
rect 5153 0 5167 24640
rect 5279 0 5293 24640
rect 5370 0 5384 24640
rect 5542 0 5556 24640
rect 5668 0 5682 24640
rect 5759 0 5773 24640
rect 5931 0 5945 24640
rect 6057 0 6071 24640
rect 6148 0 6162 24640
rect 6320 0 6334 24640
rect 6446 0 6460 24640
rect 6537 0 6551 24640
rect 6709 0 6723 24640
rect 6835 0 6849 24640
rect 6926 0 6940 24640
rect 7098 0 7112 24640
rect 7224 0 7238 24640
rect 7315 0 7329 24640
rect 7487 0 7501 24640
rect 7613 0 7627 24640
rect 7704 0 7718 24640
rect 7876 0 7890 24640
rect 8002 0 8016 24640
rect 8093 0 8107 24640
rect 8265 0 8279 24640
rect 8391 0 8405 24640
rect 8482 0 8496 24640
rect 8654 0 8668 24640
rect 8780 0 8794 24640
rect 8871 0 8885 24640
rect 9043 0 9057 24640
rect 9169 0 9183 24640
rect 9260 0 9274 24640
rect 9432 0 9446 24640
rect 9558 0 9572 24640
rect 9649 0 9663 24640
rect 9821 0 9835 24640
rect 9947 0 9961 24640
rect 10038 0 10052 24640
rect 10210 0 10224 24640
rect 10336 0 10350 24640
rect 10427 0 10441 24640
rect 10599 0 10613 24640
rect 10725 0 10739 24640
rect 10816 0 10830 24640
rect 10988 0 11002 24640
rect 11114 0 11128 24640
rect 11205 0 11219 24640
rect 11377 0 11391 24640
rect 11503 0 11517 24640
rect 11594 0 11608 24640
rect 11766 0 11780 24640
rect 11892 0 11906 24640
rect 11983 0 11997 24640
rect 12155 0 12169 24640
rect 12281 0 12295 24640
rect 12372 0 12386 24640
rect 12544 0 12558 24640
rect 12670 0 12684 24640
rect 12761 0 12775 24640
rect 12933 0 12947 24640
rect 13059 0 13073 24640
rect 13150 0 13164 24640
rect 13322 0 13336 24640
rect 13448 0 13462 24640
rect 13539 0 13553 24640
rect 13711 0 13725 24640
rect 13837 0 13851 24640
rect 13928 0 13942 24640
rect 14100 0 14114 24640
rect 14226 0 14240 24640
rect 14317 0 14331 24640
rect 14489 0 14503 24640
rect 14615 0 14629 24640
rect 14706 0 14720 24640
rect 14878 0 14892 24640
rect 15004 0 15018 24640
rect 15095 0 15109 24640
rect 15267 0 15281 24640
rect 15393 0 15407 24640
rect 15484 0 15498 24640
rect 15656 0 15670 24640
rect 15782 0 15796 24640
rect 15873 0 15887 24640
rect 16045 0 16059 24640
rect 16171 0 16185 24640
rect 16262 0 16276 24640
rect 16434 0 16448 24640
rect 16560 0 16574 24640
rect 16651 0 16665 24640
rect 16823 0 16837 24640
rect 16949 0 16963 24640
rect 17040 0 17054 24640
rect 17212 0 17226 24640
rect 17338 0 17352 24640
rect 17429 0 17443 24640
rect 17601 0 17615 24640
rect 17727 0 17741 24640
rect 17818 0 17832 24640
rect 17990 0 18004 24640
rect 18116 0 18130 24640
rect 18207 0 18221 24640
rect 18379 0 18393 24640
rect 18505 0 18519 24640
rect 18596 0 18610 24640
rect 18768 0 18782 24640
rect 18894 0 18908 24640
rect 18985 0 18999 24640
rect 19157 0 19171 24640
rect 19283 0 19297 24640
rect 19374 0 19388 24640
rect 19546 0 19560 24640
rect 19672 0 19686 24640
rect 19763 0 19777 24640
rect 19935 0 19949 24640
rect 20061 0 20075 24640
rect 20152 0 20166 24640
rect 20324 0 20338 24640
rect 20450 0 20464 24640
rect 20541 0 20555 24640
rect 20713 0 20727 24640
rect 20839 0 20853 24640
rect 20930 0 20944 24640
rect 21102 0 21116 24640
rect 21228 0 21242 24640
rect 21319 0 21333 24640
rect 21491 0 21505 24640
rect 21617 0 21631 24640
rect 21708 0 21722 24640
rect 21880 0 21894 24640
rect 22006 0 22020 24640
rect 22097 0 22111 24640
rect 22269 0 22283 24640
rect 22395 0 22409 24640
rect 22486 0 22500 24640
rect 22658 0 22672 24640
rect 22784 0 22798 24640
rect 22875 0 22889 24640
rect 23047 0 23061 24640
rect 23173 0 23187 24640
rect 23264 0 23278 24640
rect 23436 0 23450 24640
rect 23562 0 23576 24640
rect 23653 0 23667 24640
rect 23825 0 23839 24640
rect 23951 0 23965 24640
rect 24042 0 24056 24640
rect 24214 0 24228 24640
rect 24340 0 24354 24640
rect 24431 0 24445 24640
rect 24603 0 24617 24640
rect 24729 0 24743 24640
rect 24820 0 24834 24640
use cell_2r1w  cell_2r1w_0
timestamp 1643678851
transform 1 0 24507 0 -1 24640
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1
timestamp 1643678851
transform 1 0 24507 0 1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_2
timestamp 1643678851
transform 1 0 24507 0 -1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_3
timestamp 1643678851
transform 1 0 24507 0 1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_4
timestamp 1643678851
transform 1 0 24507 0 -1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_5
timestamp 1643678851
transform 1 0 24507 0 1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_6
timestamp 1643678851
transform 1 0 24507 0 -1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_7
timestamp 1643678851
transform 1 0 24507 0 1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_8
timestamp 1643678851
transform 1 0 24507 0 -1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_9
timestamp 1643678851
transform 1 0 24507 0 1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_10
timestamp 1643678851
transform 1 0 24507 0 -1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_11
timestamp 1643678851
transform 1 0 24507 0 1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_12
timestamp 1643678851
transform 1 0 24507 0 -1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_13
timestamp 1643678851
transform 1 0 24507 0 1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_14
timestamp 1643678851
transform 1 0 24507 0 -1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_15
timestamp 1643678851
transform 1 0 24507 0 1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_16
timestamp 1643678851
transform 1 0 24507 0 -1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_17
timestamp 1643678851
transform 1 0 24507 0 1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_18
timestamp 1643678851
transform 1 0 24507 0 -1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_19
timestamp 1643678851
transform 1 0 24507 0 1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_20
timestamp 1643678851
transform 1 0 24507 0 -1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_21
timestamp 1643678851
transform 1 0 24507 0 1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_22
timestamp 1643678851
transform 1 0 24507 0 -1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_23
timestamp 1643678851
transform 1 0 24507 0 1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_24
timestamp 1643678851
transform 1 0 24507 0 -1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_25
timestamp 1643678851
transform 1 0 24507 0 1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_26
timestamp 1643678851
transform 1 0 24507 0 -1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_27
timestamp 1643678851
transform 1 0 24507 0 1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_28
timestamp 1643678851
transform 1 0 24507 0 -1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_29
timestamp 1643678851
transform 1 0 24507 0 1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_30
timestamp 1643678851
transform 1 0 24507 0 -1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_31
timestamp 1643678851
transform 1 0 24507 0 1 0
box 0 -21 389 808
use cell_2r1w  cell_2r1w_32
timestamp 1643678851
transform 1 0 24118 0 -1 24640
box 0 -21 389 808
use cell_2r1w  cell_2r1w_33
timestamp 1643678851
transform 1 0 24118 0 1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_34
timestamp 1643678851
transform 1 0 24118 0 -1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_35
timestamp 1643678851
transform 1 0 24118 0 1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_36
timestamp 1643678851
transform 1 0 24118 0 -1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_37
timestamp 1643678851
transform 1 0 24118 0 1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_38
timestamp 1643678851
transform 1 0 24118 0 -1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_39
timestamp 1643678851
transform 1 0 24118 0 1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_40
timestamp 1643678851
transform 1 0 24118 0 -1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_41
timestamp 1643678851
transform 1 0 24118 0 1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_42
timestamp 1643678851
transform 1 0 24118 0 -1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_43
timestamp 1643678851
transform 1 0 24118 0 1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_44
timestamp 1643678851
transform 1 0 24118 0 -1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_45
timestamp 1643678851
transform 1 0 24118 0 1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_46
timestamp 1643678851
transform 1 0 24118 0 -1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_47
timestamp 1643678851
transform 1 0 24118 0 1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_48
timestamp 1643678851
transform 1 0 24118 0 -1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_49
timestamp 1643678851
transform 1 0 24118 0 1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_50
timestamp 1643678851
transform 1 0 24118 0 -1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_51
timestamp 1643678851
transform 1 0 24118 0 1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_52
timestamp 1643678851
transform 1 0 24118 0 -1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_53
timestamp 1643678851
transform 1 0 24118 0 1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_54
timestamp 1643678851
transform 1 0 24118 0 -1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_55
timestamp 1643678851
transform 1 0 24118 0 1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_56
timestamp 1643678851
transform 1 0 24118 0 -1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_57
timestamp 1643678851
transform 1 0 24118 0 1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_58
timestamp 1643678851
transform 1 0 24118 0 -1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_59
timestamp 1643678851
transform 1 0 24118 0 1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_60
timestamp 1643678851
transform 1 0 24118 0 -1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_61
timestamp 1643678851
transform 1 0 24118 0 1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_62
timestamp 1643678851
transform 1 0 24118 0 -1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_63
timestamp 1643678851
transform 1 0 24118 0 1 0
box 0 -21 389 808
use cell_2r1w  cell_2r1w_64
timestamp 1643678851
transform 1 0 23729 0 -1 24640
box 0 -21 389 808
use cell_2r1w  cell_2r1w_65
timestamp 1643678851
transform 1 0 23729 0 1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_66
timestamp 1643678851
transform 1 0 23729 0 -1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_67
timestamp 1643678851
transform 1 0 23729 0 1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_68
timestamp 1643678851
transform 1 0 23729 0 -1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_69
timestamp 1643678851
transform 1 0 23729 0 1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_70
timestamp 1643678851
transform 1 0 23729 0 -1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_71
timestamp 1643678851
transform 1 0 23729 0 1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_72
timestamp 1643678851
transform 1 0 23729 0 -1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_73
timestamp 1643678851
transform 1 0 23729 0 1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_74
timestamp 1643678851
transform 1 0 23729 0 -1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_75
timestamp 1643678851
transform 1 0 23729 0 1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_76
timestamp 1643678851
transform 1 0 23729 0 -1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_77
timestamp 1643678851
transform 1 0 23729 0 1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_78
timestamp 1643678851
transform 1 0 23729 0 -1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_79
timestamp 1643678851
transform 1 0 23729 0 1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_80
timestamp 1643678851
transform 1 0 23729 0 -1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_81
timestamp 1643678851
transform 1 0 23729 0 1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_82
timestamp 1643678851
transform 1 0 23729 0 -1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_83
timestamp 1643678851
transform 1 0 23729 0 1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_84
timestamp 1643678851
transform 1 0 23729 0 -1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_85
timestamp 1643678851
transform 1 0 23729 0 1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_86
timestamp 1643678851
transform 1 0 23729 0 -1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_87
timestamp 1643678851
transform 1 0 23729 0 1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_88
timestamp 1643678851
transform 1 0 23729 0 -1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_89
timestamp 1643678851
transform 1 0 23729 0 1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_90
timestamp 1643678851
transform 1 0 23729 0 -1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_91
timestamp 1643678851
transform 1 0 23729 0 1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_92
timestamp 1643678851
transform 1 0 23729 0 -1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_93
timestamp 1643678851
transform 1 0 23729 0 1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_94
timestamp 1643678851
transform 1 0 23729 0 -1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_95
timestamp 1643678851
transform 1 0 23729 0 1 0
box 0 -21 389 808
use cell_2r1w  cell_2r1w_96
timestamp 1643678851
transform 1 0 23340 0 -1 24640
box 0 -21 389 808
use cell_2r1w  cell_2r1w_97
timestamp 1643678851
transform 1 0 23340 0 1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_98
timestamp 1643678851
transform 1 0 23340 0 -1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_99
timestamp 1643678851
transform 1 0 23340 0 1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_100
timestamp 1643678851
transform 1 0 23340 0 -1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_101
timestamp 1643678851
transform 1 0 23340 0 1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_102
timestamp 1643678851
transform 1 0 23340 0 -1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_103
timestamp 1643678851
transform 1 0 23340 0 1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_104
timestamp 1643678851
transform 1 0 23340 0 -1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_105
timestamp 1643678851
transform 1 0 23340 0 1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_106
timestamp 1643678851
transform 1 0 23340 0 -1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_107
timestamp 1643678851
transform 1 0 23340 0 1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_108
timestamp 1643678851
transform 1 0 23340 0 -1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_109
timestamp 1643678851
transform 1 0 23340 0 1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_110
timestamp 1643678851
transform 1 0 23340 0 -1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_111
timestamp 1643678851
transform 1 0 23340 0 1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_112
timestamp 1643678851
transform 1 0 23340 0 -1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_113
timestamp 1643678851
transform 1 0 23340 0 1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_114
timestamp 1643678851
transform 1 0 23340 0 -1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_115
timestamp 1643678851
transform 1 0 23340 0 1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_116
timestamp 1643678851
transform 1 0 23340 0 -1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_117
timestamp 1643678851
transform 1 0 23340 0 1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_118
timestamp 1643678851
transform 1 0 23340 0 -1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_119
timestamp 1643678851
transform 1 0 23340 0 1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_120
timestamp 1643678851
transform 1 0 23340 0 -1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_121
timestamp 1643678851
transform 1 0 23340 0 1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_122
timestamp 1643678851
transform 1 0 23340 0 -1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_123
timestamp 1643678851
transform 1 0 23340 0 1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_124
timestamp 1643678851
transform 1 0 23340 0 -1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_125
timestamp 1643678851
transform 1 0 23340 0 1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_126
timestamp 1643678851
transform 1 0 23340 0 -1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_127
timestamp 1643678851
transform 1 0 23340 0 1 0
box 0 -21 389 808
use cell_2r1w  cell_2r1w_128
timestamp 1643678851
transform 1 0 22951 0 -1 24640
box 0 -21 389 808
use cell_2r1w  cell_2r1w_129
timestamp 1643678851
transform 1 0 22951 0 1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_130
timestamp 1643678851
transform 1 0 22951 0 -1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_131
timestamp 1643678851
transform 1 0 22951 0 1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_132
timestamp 1643678851
transform 1 0 22951 0 -1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_133
timestamp 1643678851
transform 1 0 22951 0 1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_134
timestamp 1643678851
transform 1 0 22951 0 -1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_135
timestamp 1643678851
transform 1 0 22951 0 1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_136
timestamp 1643678851
transform 1 0 22951 0 -1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_137
timestamp 1643678851
transform 1 0 22951 0 1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_138
timestamp 1643678851
transform 1 0 22951 0 -1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_139
timestamp 1643678851
transform 1 0 22951 0 1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_140
timestamp 1643678851
transform 1 0 22951 0 -1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_141
timestamp 1643678851
transform 1 0 22951 0 1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_142
timestamp 1643678851
transform 1 0 22951 0 -1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_143
timestamp 1643678851
transform 1 0 22951 0 1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_144
timestamp 1643678851
transform 1 0 22951 0 -1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_145
timestamp 1643678851
transform 1 0 22951 0 1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_146
timestamp 1643678851
transform 1 0 22951 0 -1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_147
timestamp 1643678851
transform 1 0 22951 0 1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_148
timestamp 1643678851
transform 1 0 22951 0 -1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_149
timestamp 1643678851
transform 1 0 22951 0 1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_150
timestamp 1643678851
transform 1 0 22951 0 -1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_151
timestamp 1643678851
transform 1 0 22951 0 1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_152
timestamp 1643678851
transform 1 0 22951 0 -1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_153
timestamp 1643678851
transform 1 0 22951 0 1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_154
timestamp 1643678851
transform 1 0 22951 0 -1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_155
timestamp 1643678851
transform 1 0 22951 0 1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_156
timestamp 1643678851
transform 1 0 22951 0 -1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_157
timestamp 1643678851
transform 1 0 22951 0 1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_158
timestamp 1643678851
transform 1 0 22951 0 -1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_159
timestamp 1643678851
transform 1 0 22951 0 1 0
box 0 -21 389 808
use cell_2r1w  cell_2r1w_160
timestamp 1643678851
transform 1 0 22562 0 -1 24640
box 0 -21 389 808
use cell_2r1w  cell_2r1w_161
timestamp 1643678851
transform 1 0 22562 0 1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_162
timestamp 1643678851
transform 1 0 22562 0 -1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_163
timestamp 1643678851
transform 1 0 22562 0 1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_164
timestamp 1643678851
transform 1 0 22562 0 -1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_165
timestamp 1643678851
transform 1 0 22562 0 1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_166
timestamp 1643678851
transform 1 0 22562 0 -1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_167
timestamp 1643678851
transform 1 0 22562 0 1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_168
timestamp 1643678851
transform 1 0 22562 0 -1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_169
timestamp 1643678851
transform 1 0 22562 0 1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_170
timestamp 1643678851
transform 1 0 22562 0 -1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_171
timestamp 1643678851
transform 1 0 22562 0 1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_172
timestamp 1643678851
transform 1 0 22562 0 -1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_173
timestamp 1643678851
transform 1 0 22562 0 1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_174
timestamp 1643678851
transform 1 0 22562 0 -1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_175
timestamp 1643678851
transform 1 0 22562 0 1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_176
timestamp 1643678851
transform 1 0 22562 0 -1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_177
timestamp 1643678851
transform 1 0 22562 0 1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_178
timestamp 1643678851
transform 1 0 22562 0 -1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_179
timestamp 1643678851
transform 1 0 22562 0 1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_180
timestamp 1643678851
transform 1 0 22562 0 -1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_181
timestamp 1643678851
transform 1 0 22562 0 1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_182
timestamp 1643678851
transform 1 0 22562 0 -1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_183
timestamp 1643678851
transform 1 0 22562 0 1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_184
timestamp 1643678851
transform 1 0 22562 0 -1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_185
timestamp 1643678851
transform 1 0 22562 0 1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_186
timestamp 1643678851
transform 1 0 22562 0 -1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_187
timestamp 1643678851
transform 1 0 22562 0 1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_188
timestamp 1643678851
transform 1 0 22562 0 -1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_189
timestamp 1643678851
transform 1 0 22562 0 1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_190
timestamp 1643678851
transform 1 0 22562 0 -1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_191
timestamp 1643678851
transform 1 0 22562 0 1 0
box 0 -21 389 808
use cell_2r1w  cell_2r1w_192
timestamp 1643678851
transform 1 0 22173 0 -1 24640
box 0 -21 389 808
use cell_2r1w  cell_2r1w_193
timestamp 1643678851
transform 1 0 22173 0 1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_194
timestamp 1643678851
transform 1 0 22173 0 -1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_195
timestamp 1643678851
transform 1 0 22173 0 1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_196
timestamp 1643678851
transform 1 0 22173 0 -1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_197
timestamp 1643678851
transform 1 0 22173 0 1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_198
timestamp 1643678851
transform 1 0 22173 0 -1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_199
timestamp 1643678851
transform 1 0 22173 0 1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_200
timestamp 1643678851
transform 1 0 22173 0 -1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_201
timestamp 1643678851
transform 1 0 22173 0 1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_202
timestamp 1643678851
transform 1 0 22173 0 -1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_203
timestamp 1643678851
transform 1 0 22173 0 1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_204
timestamp 1643678851
transform 1 0 22173 0 -1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_205
timestamp 1643678851
transform 1 0 22173 0 1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_206
timestamp 1643678851
transform 1 0 22173 0 -1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_207
timestamp 1643678851
transform 1 0 22173 0 1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_208
timestamp 1643678851
transform 1 0 22173 0 -1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_209
timestamp 1643678851
transform 1 0 22173 0 1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_210
timestamp 1643678851
transform 1 0 22173 0 -1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_211
timestamp 1643678851
transform 1 0 22173 0 1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_212
timestamp 1643678851
transform 1 0 22173 0 -1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_213
timestamp 1643678851
transform 1 0 22173 0 1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_214
timestamp 1643678851
transform 1 0 22173 0 -1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_215
timestamp 1643678851
transform 1 0 22173 0 1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_216
timestamp 1643678851
transform 1 0 22173 0 -1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_217
timestamp 1643678851
transform 1 0 22173 0 1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_218
timestamp 1643678851
transform 1 0 22173 0 -1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_219
timestamp 1643678851
transform 1 0 22173 0 1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_220
timestamp 1643678851
transform 1 0 22173 0 -1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_221
timestamp 1643678851
transform 1 0 22173 0 1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_222
timestamp 1643678851
transform 1 0 22173 0 -1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_223
timestamp 1643678851
transform 1 0 22173 0 1 0
box 0 -21 389 808
use cell_2r1w  cell_2r1w_224
timestamp 1643678851
transform 1 0 21784 0 -1 24640
box 0 -21 389 808
use cell_2r1w  cell_2r1w_225
timestamp 1643678851
transform 1 0 21784 0 1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_226
timestamp 1643678851
transform 1 0 21784 0 -1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_227
timestamp 1643678851
transform 1 0 21784 0 1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_228
timestamp 1643678851
transform 1 0 21784 0 -1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_229
timestamp 1643678851
transform 1 0 21784 0 1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_230
timestamp 1643678851
transform 1 0 21784 0 -1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_231
timestamp 1643678851
transform 1 0 21784 0 1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_232
timestamp 1643678851
transform 1 0 21784 0 -1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_233
timestamp 1643678851
transform 1 0 21784 0 1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_234
timestamp 1643678851
transform 1 0 21784 0 -1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_235
timestamp 1643678851
transform 1 0 21784 0 1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_236
timestamp 1643678851
transform 1 0 21784 0 -1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_237
timestamp 1643678851
transform 1 0 21784 0 1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_238
timestamp 1643678851
transform 1 0 21784 0 -1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_239
timestamp 1643678851
transform 1 0 21784 0 1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_240
timestamp 1643678851
transform 1 0 21784 0 -1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_241
timestamp 1643678851
transform 1 0 21784 0 1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_242
timestamp 1643678851
transform 1 0 21784 0 -1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_243
timestamp 1643678851
transform 1 0 21784 0 1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_244
timestamp 1643678851
transform 1 0 21784 0 -1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_245
timestamp 1643678851
transform 1 0 21784 0 1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_246
timestamp 1643678851
transform 1 0 21784 0 -1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_247
timestamp 1643678851
transform 1 0 21784 0 1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_248
timestamp 1643678851
transform 1 0 21784 0 -1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_249
timestamp 1643678851
transform 1 0 21784 0 1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_250
timestamp 1643678851
transform 1 0 21784 0 -1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_251
timestamp 1643678851
transform 1 0 21784 0 1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_252
timestamp 1643678851
transform 1 0 21784 0 -1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_253
timestamp 1643678851
transform 1 0 21784 0 1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_254
timestamp 1643678851
transform 1 0 21784 0 -1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_255
timestamp 1643678851
transform 1 0 21784 0 1 0
box 0 -21 389 808
use cell_2r1w  cell_2r1w_256
timestamp 1643678851
transform 1 0 21395 0 -1 24640
box 0 -21 389 808
use cell_2r1w  cell_2r1w_257
timestamp 1643678851
transform 1 0 21395 0 1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_258
timestamp 1643678851
transform 1 0 21395 0 -1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_259
timestamp 1643678851
transform 1 0 21395 0 1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_260
timestamp 1643678851
transform 1 0 21395 0 -1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_261
timestamp 1643678851
transform 1 0 21395 0 1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_262
timestamp 1643678851
transform 1 0 21395 0 -1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_263
timestamp 1643678851
transform 1 0 21395 0 1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_264
timestamp 1643678851
transform 1 0 21395 0 -1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_265
timestamp 1643678851
transform 1 0 21395 0 1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_266
timestamp 1643678851
transform 1 0 21395 0 -1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_267
timestamp 1643678851
transform 1 0 21395 0 1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_268
timestamp 1643678851
transform 1 0 21395 0 -1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_269
timestamp 1643678851
transform 1 0 21395 0 1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_270
timestamp 1643678851
transform 1 0 21395 0 -1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_271
timestamp 1643678851
transform 1 0 21395 0 1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_272
timestamp 1643678851
transform 1 0 21395 0 -1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_273
timestamp 1643678851
transform 1 0 21395 0 1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_274
timestamp 1643678851
transform 1 0 21395 0 -1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_275
timestamp 1643678851
transform 1 0 21395 0 1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_276
timestamp 1643678851
transform 1 0 21395 0 -1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_277
timestamp 1643678851
transform 1 0 21395 0 1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_278
timestamp 1643678851
transform 1 0 21395 0 -1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_279
timestamp 1643678851
transform 1 0 21395 0 1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_280
timestamp 1643678851
transform 1 0 21395 0 -1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_281
timestamp 1643678851
transform 1 0 21395 0 1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_282
timestamp 1643678851
transform 1 0 21395 0 -1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_283
timestamp 1643678851
transform 1 0 21395 0 1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_284
timestamp 1643678851
transform 1 0 21395 0 -1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_285
timestamp 1643678851
transform 1 0 21395 0 1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_286
timestamp 1643678851
transform 1 0 21395 0 -1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_287
timestamp 1643678851
transform 1 0 21395 0 1 0
box 0 -21 389 808
use cell_2r1w  cell_2r1w_288
timestamp 1643678851
transform 1 0 21006 0 -1 24640
box 0 -21 389 808
use cell_2r1w  cell_2r1w_289
timestamp 1643678851
transform 1 0 21006 0 1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_290
timestamp 1643678851
transform 1 0 21006 0 -1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_291
timestamp 1643678851
transform 1 0 21006 0 1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_292
timestamp 1643678851
transform 1 0 21006 0 -1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_293
timestamp 1643678851
transform 1 0 21006 0 1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_294
timestamp 1643678851
transform 1 0 21006 0 -1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_295
timestamp 1643678851
transform 1 0 21006 0 1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_296
timestamp 1643678851
transform 1 0 21006 0 -1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_297
timestamp 1643678851
transform 1 0 21006 0 1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_298
timestamp 1643678851
transform 1 0 21006 0 -1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_299
timestamp 1643678851
transform 1 0 21006 0 1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_300
timestamp 1643678851
transform 1 0 21006 0 -1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_301
timestamp 1643678851
transform 1 0 21006 0 1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_302
timestamp 1643678851
transform 1 0 21006 0 -1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_303
timestamp 1643678851
transform 1 0 21006 0 1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_304
timestamp 1643678851
transform 1 0 21006 0 -1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_305
timestamp 1643678851
transform 1 0 21006 0 1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_306
timestamp 1643678851
transform 1 0 21006 0 -1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_307
timestamp 1643678851
transform 1 0 21006 0 1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_308
timestamp 1643678851
transform 1 0 21006 0 -1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_309
timestamp 1643678851
transform 1 0 21006 0 1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_310
timestamp 1643678851
transform 1 0 21006 0 -1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_311
timestamp 1643678851
transform 1 0 21006 0 1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_312
timestamp 1643678851
transform 1 0 21006 0 -1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_313
timestamp 1643678851
transform 1 0 21006 0 1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_314
timestamp 1643678851
transform 1 0 21006 0 -1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_315
timestamp 1643678851
transform 1 0 21006 0 1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_316
timestamp 1643678851
transform 1 0 21006 0 -1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_317
timestamp 1643678851
transform 1 0 21006 0 1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_318
timestamp 1643678851
transform 1 0 21006 0 -1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_319
timestamp 1643678851
transform 1 0 21006 0 1 0
box 0 -21 389 808
use cell_2r1w  cell_2r1w_320
timestamp 1643678851
transform 1 0 20617 0 -1 24640
box 0 -21 389 808
use cell_2r1w  cell_2r1w_321
timestamp 1643678851
transform 1 0 20617 0 1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_322
timestamp 1643678851
transform 1 0 20617 0 -1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_323
timestamp 1643678851
transform 1 0 20617 0 1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_324
timestamp 1643678851
transform 1 0 20617 0 -1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_325
timestamp 1643678851
transform 1 0 20617 0 1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_326
timestamp 1643678851
transform 1 0 20617 0 -1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_327
timestamp 1643678851
transform 1 0 20617 0 1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_328
timestamp 1643678851
transform 1 0 20617 0 -1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_329
timestamp 1643678851
transform 1 0 20617 0 1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_330
timestamp 1643678851
transform 1 0 20617 0 -1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_331
timestamp 1643678851
transform 1 0 20617 0 1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_332
timestamp 1643678851
transform 1 0 20617 0 -1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_333
timestamp 1643678851
transform 1 0 20617 0 1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_334
timestamp 1643678851
transform 1 0 20617 0 -1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_335
timestamp 1643678851
transform 1 0 20617 0 1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_336
timestamp 1643678851
transform 1 0 20617 0 -1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_337
timestamp 1643678851
transform 1 0 20617 0 1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_338
timestamp 1643678851
transform 1 0 20617 0 -1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_339
timestamp 1643678851
transform 1 0 20617 0 1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_340
timestamp 1643678851
transform 1 0 20617 0 -1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_341
timestamp 1643678851
transform 1 0 20617 0 1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_342
timestamp 1643678851
transform 1 0 20617 0 -1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_343
timestamp 1643678851
transform 1 0 20617 0 1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_344
timestamp 1643678851
transform 1 0 20617 0 -1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_345
timestamp 1643678851
transform 1 0 20617 0 1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_346
timestamp 1643678851
transform 1 0 20617 0 -1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_347
timestamp 1643678851
transform 1 0 20617 0 1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_348
timestamp 1643678851
transform 1 0 20617 0 -1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_349
timestamp 1643678851
transform 1 0 20617 0 1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_350
timestamp 1643678851
transform 1 0 20617 0 -1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_351
timestamp 1643678851
transform 1 0 20617 0 1 0
box 0 -21 389 808
use cell_2r1w  cell_2r1w_352
timestamp 1643678851
transform 1 0 20228 0 -1 24640
box 0 -21 389 808
use cell_2r1w  cell_2r1w_353
timestamp 1643678851
transform 1 0 20228 0 1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_354
timestamp 1643678851
transform 1 0 20228 0 -1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_355
timestamp 1643678851
transform 1 0 20228 0 1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_356
timestamp 1643678851
transform 1 0 20228 0 -1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_357
timestamp 1643678851
transform 1 0 20228 0 1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_358
timestamp 1643678851
transform 1 0 20228 0 -1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_359
timestamp 1643678851
transform 1 0 20228 0 1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_360
timestamp 1643678851
transform 1 0 20228 0 -1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_361
timestamp 1643678851
transform 1 0 20228 0 1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_362
timestamp 1643678851
transform 1 0 20228 0 -1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_363
timestamp 1643678851
transform 1 0 20228 0 1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_364
timestamp 1643678851
transform 1 0 20228 0 -1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_365
timestamp 1643678851
transform 1 0 20228 0 1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_366
timestamp 1643678851
transform 1 0 20228 0 -1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_367
timestamp 1643678851
transform 1 0 20228 0 1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_368
timestamp 1643678851
transform 1 0 20228 0 -1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_369
timestamp 1643678851
transform 1 0 20228 0 1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_370
timestamp 1643678851
transform 1 0 20228 0 -1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_371
timestamp 1643678851
transform 1 0 20228 0 1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_372
timestamp 1643678851
transform 1 0 20228 0 -1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_373
timestamp 1643678851
transform 1 0 20228 0 1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_374
timestamp 1643678851
transform 1 0 20228 0 -1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_375
timestamp 1643678851
transform 1 0 20228 0 1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_376
timestamp 1643678851
transform 1 0 20228 0 -1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_377
timestamp 1643678851
transform 1 0 20228 0 1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_378
timestamp 1643678851
transform 1 0 20228 0 -1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_379
timestamp 1643678851
transform 1 0 20228 0 1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_380
timestamp 1643678851
transform 1 0 20228 0 -1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_381
timestamp 1643678851
transform 1 0 20228 0 1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_382
timestamp 1643678851
transform 1 0 20228 0 -1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_383
timestamp 1643678851
transform 1 0 20228 0 1 0
box 0 -21 389 808
use cell_2r1w  cell_2r1w_384
timestamp 1643678851
transform 1 0 19839 0 -1 24640
box 0 -21 389 808
use cell_2r1w  cell_2r1w_385
timestamp 1643678851
transform 1 0 19839 0 1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_386
timestamp 1643678851
transform 1 0 19839 0 -1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_387
timestamp 1643678851
transform 1 0 19839 0 1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_388
timestamp 1643678851
transform 1 0 19839 0 -1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_389
timestamp 1643678851
transform 1 0 19839 0 1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_390
timestamp 1643678851
transform 1 0 19839 0 -1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_391
timestamp 1643678851
transform 1 0 19839 0 1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_392
timestamp 1643678851
transform 1 0 19839 0 -1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_393
timestamp 1643678851
transform 1 0 19839 0 1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_394
timestamp 1643678851
transform 1 0 19839 0 -1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_395
timestamp 1643678851
transform 1 0 19839 0 1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_396
timestamp 1643678851
transform 1 0 19839 0 -1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_397
timestamp 1643678851
transform 1 0 19839 0 1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_398
timestamp 1643678851
transform 1 0 19839 0 -1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_399
timestamp 1643678851
transform 1 0 19839 0 1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_400
timestamp 1643678851
transform 1 0 19839 0 -1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_401
timestamp 1643678851
transform 1 0 19839 0 1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_402
timestamp 1643678851
transform 1 0 19839 0 -1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_403
timestamp 1643678851
transform 1 0 19839 0 1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_404
timestamp 1643678851
transform 1 0 19839 0 -1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_405
timestamp 1643678851
transform 1 0 19839 0 1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_406
timestamp 1643678851
transform 1 0 19839 0 -1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_407
timestamp 1643678851
transform 1 0 19839 0 1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_408
timestamp 1643678851
transform 1 0 19839 0 -1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_409
timestamp 1643678851
transform 1 0 19839 0 1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_410
timestamp 1643678851
transform 1 0 19839 0 -1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_411
timestamp 1643678851
transform 1 0 19839 0 1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_412
timestamp 1643678851
transform 1 0 19839 0 -1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_413
timestamp 1643678851
transform 1 0 19839 0 1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_414
timestamp 1643678851
transform 1 0 19839 0 -1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_415
timestamp 1643678851
transform 1 0 19839 0 1 0
box 0 -21 389 808
use cell_2r1w  cell_2r1w_416
timestamp 1643678851
transform 1 0 19450 0 -1 24640
box 0 -21 389 808
use cell_2r1w  cell_2r1w_417
timestamp 1643678851
transform 1 0 19450 0 1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_418
timestamp 1643678851
transform 1 0 19450 0 -1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_419
timestamp 1643678851
transform 1 0 19450 0 1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_420
timestamp 1643678851
transform 1 0 19450 0 -1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_421
timestamp 1643678851
transform 1 0 19450 0 1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_422
timestamp 1643678851
transform 1 0 19450 0 -1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_423
timestamp 1643678851
transform 1 0 19450 0 1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_424
timestamp 1643678851
transform 1 0 19450 0 -1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_425
timestamp 1643678851
transform 1 0 19450 0 1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_426
timestamp 1643678851
transform 1 0 19450 0 -1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_427
timestamp 1643678851
transform 1 0 19450 0 1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_428
timestamp 1643678851
transform 1 0 19450 0 -1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_429
timestamp 1643678851
transform 1 0 19450 0 1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_430
timestamp 1643678851
transform 1 0 19450 0 -1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_431
timestamp 1643678851
transform 1 0 19450 0 1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_432
timestamp 1643678851
transform 1 0 19450 0 -1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_433
timestamp 1643678851
transform 1 0 19450 0 1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_434
timestamp 1643678851
transform 1 0 19450 0 -1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_435
timestamp 1643678851
transform 1 0 19450 0 1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_436
timestamp 1643678851
transform 1 0 19450 0 -1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_437
timestamp 1643678851
transform 1 0 19450 0 1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_438
timestamp 1643678851
transform 1 0 19450 0 -1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_439
timestamp 1643678851
transform 1 0 19450 0 1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_440
timestamp 1643678851
transform 1 0 19450 0 -1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_441
timestamp 1643678851
transform 1 0 19450 0 1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_442
timestamp 1643678851
transform 1 0 19450 0 -1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_443
timestamp 1643678851
transform 1 0 19450 0 1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_444
timestamp 1643678851
transform 1 0 19450 0 -1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_445
timestamp 1643678851
transform 1 0 19450 0 1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_446
timestamp 1643678851
transform 1 0 19450 0 -1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_447
timestamp 1643678851
transform 1 0 19450 0 1 0
box 0 -21 389 808
use cell_2r1w  cell_2r1w_448
timestamp 1643678851
transform 1 0 19061 0 -1 24640
box 0 -21 389 808
use cell_2r1w  cell_2r1w_449
timestamp 1643678851
transform 1 0 19061 0 1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_450
timestamp 1643678851
transform 1 0 19061 0 -1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_451
timestamp 1643678851
transform 1 0 19061 0 1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_452
timestamp 1643678851
transform 1 0 19061 0 -1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_453
timestamp 1643678851
transform 1 0 19061 0 1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_454
timestamp 1643678851
transform 1 0 19061 0 -1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_455
timestamp 1643678851
transform 1 0 19061 0 1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_456
timestamp 1643678851
transform 1 0 19061 0 -1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_457
timestamp 1643678851
transform 1 0 19061 0 1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_458
timestamp 1643678851
transform 1 0 19061 0 -1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_459
timestamp 1643678851
transform 1 0 19061 0 1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_460
timestamp 1643678851
transform 1 0 19061 0 -1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_461
timestamp 1643678851
transform 1 0 19061 0 1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_462
timestamp 1643678851
transform 1 0 19061 0 -1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_463
timestamp 1643678851
transform 1 0 19061 0 1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_464
timestamp 1643678851
transform 1 0 19061 0 -1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_465
timestamp 1643678851
transform 1 0 19061 0 1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_466
timestamp 1643678851
transform 1 0 19061 0 -1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_467
timestamp 1643678851
transform 1 0 19061 0 1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_468
timestamp 1643678851
transform 1 0 19061 0 -1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_469
timestamp 1643678851
transform 1 0 19061 0 1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_470
timestamp 1643678851
transform 1 0 19061 0 -1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_471
timestamp 1643678851
transform 1 0 19061 0 1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_472
timestamp 1643678851
transform 1 0 19061 0 -1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_473
timestamp 1643678851
transform 1 0 19061 0 1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_474
timestamp 1643678851
transform 1 0 19061 0 -1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_475
timestamp 1643678851
transform 1 0 19061 0 1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_476
timestamp 1643678851
transform 1 0 19061 0 -1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_477
timestamp 1643678851
transform 1 0 19061 0 1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_478
timestamp 1643678851
transform 1 0 19061 0 -1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_479
timestamp 1643678851
transform 1 0 19061 0 1 0
box 0 -21 389 808
use cell_2r1w  cell_2r1w_480
timestamp 1643678851
transform 1 0 18672 0 -1 24640
box 0 -21 389 808
use cell_2r1w  cell_2r1w_481
timestamp 1643678851
transform 1 0 18672 0 1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_482
timestamp 1643678851
transform 1 0 18672 0 -1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_483
timestamp 1643678851
transform 1 0 18672 0 1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_484
timestamp 1643678851
transform 1 0 18672 0 -1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_485
timestamp 1643678851
transform 1 0 18672 0 1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_486
timestamp 1643678851
transform 1 0 18672 0 -1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_487
timestamp 1643678851
transform 1 0 18672 0 1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_488
timestamp 1643678851
transform 1 0 18672 0 -1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_489
timestamp 1643678851
transform 1 0 18672 0 1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_490
timestamp 1643678851
transform 1 0 18672 0 -1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_491
timestamp 1643678851
transform 1 0 18672 0 1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_492
timestamp 1643678851
transform 1 0 18672 0 -1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_493
timestamp 1643678851
transform 1 0 18672 0 1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_494
timestamp 1643678851
transform 1 0 18672 0 -1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_495
timestamp 1643678851
transform 1 0 18672 0 1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_496
timestamp 1643678851
transform 1 0 18672 0 -1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_497
timestamp 1643678851
transform 1 0 18672 0 1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_498
timestamp 1643678851
transform 1 0 18672 0 -1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_499
timestamp 1643678851
transform 1 0 18672 0 1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_500
timestamp 1643678851
transform 1 0 18672 0 -1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_501
timestamp 1643678851
transform 1 0 18672 0 1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_502
timestamp 1643678851
transform 1 0 18672 0 -1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_503
timestamp 1643678851
transform 1 0 18672 0 1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_504
timestamp 1643678851
transform 1 0 18672 0 -1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_505
timestamp 1643678851
transform 1 0 18672 0 1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_506
timestamp 1643678851
transform 1 0 18672 0 -1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_507
timestamp 1643678851
transform 1 0 18672 0 1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_508
timestamp 1643678851
transform 1 0 18672 0 -1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_509
timestamp 1643678851
transform 1 0 18672 0 1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_510
timestamp 1643678851
transform 1 0 18672 0 -1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_511
timestamp 1643678851
transform 1 0 18672 0 1 0
box 0 -21 389 808
use cell_2r1w  cell_2r1w_512
timestamp 1643678851
transform 1 0 18283 0 -1 24640
box 0 -21 389 808
use cell_2r1w  cell_2r1w_513
timestamp 1643678851
transform 1 0 18283 0 1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_514
timestamp 1643678851
transform 1 0 18283 0 -1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_515
timestamp 1643678851
transform 1 0 18283 0 1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_516
timestamp 1643678851
transform 1 0 18283 0 -1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_517
timestamp 1643678851
transform 1 0 18283 0 1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_518
timestamp 1643678851
transform 1 0 18283 0 -1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_519
timestamp 1643678851
transform 1 0 18283 0 1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_520
timestamp 1643678851
transform 1 0 18283 0 -1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_521
timestamp 1643678851
transform 1 0 18283 0 1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_522
timestamp 1643678851
transform 1 0 18283 0 -1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_523
timestamp 1643678851
transform 1 0 18283 0 1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_524
timestamp 1643678851
transform 1 0 18283 0 -1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_525
timestamp 1643678851
transform 1 0 18283 0 1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_526
timestamp 1643678851
transform 1 0 18283 0 -1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_527
timestamp 1643678851
transform 1 0 18283 0 1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_528
timestamp 1643678851
transform 1 0 18283 0 -1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_529
timestamp 1643678851
transform 1 0 18283 0 1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_530
timestamp 1643678851
transform 1 0 18283 0 -1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_531
timestamp 1643678851
transform 1 0 18283 0 1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_532
timestamp 1643678851
transform 1 0 18283 0 -1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_533
timestamp 1643678851
transform 1 0 18283 0 1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_534
timestamp 1643678851
transform 1 0 18283 0 -1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_535
timestamp 1643678851
transform 1 0 18283 0 1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_536
timestamp 1643678851
transform 1 0 18283 0 -1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_537
timestamp 1643678851
transform 1 0 18283 0 1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_538
timestamp 1643678851
transform 1 0 18283 0 -1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_539
timestamp 1643678851
transform 1 0 18283 0 1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_540
timestamp 1643678851
transform 1 0 18283 0 -1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_541
timestamp 1643678851
transform 1 0 18283 0 1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_542
timestamp 1643678851
transform 1 0 18283 0 -1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_543
timestamp 1643678851
transform 1 0 18283 0 1 0
box 0 -21 389 808
use cell_2r1w  cell_2r1w_544
timestamp 1643678851
transform 1 0 17894 0 -1 24640
box 0 -21 389 808
use cell_2r1w  cell_2r1w_545
timestamp 1643678851
transform 1 0 17894 0 1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_546
timestamp 1643678851
transform 1 0 17894 0 -1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_547
timestamp 1643678851
transform 1 0 17894 0 1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_548
timestamp 1643678851
transform 1 0 17894 0 -1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_549
timestamp 1643678851
transform 1 0 17894 0 1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_550
timestamp 1643678851
transform 1 0 17894 0 -1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_551
timestamp 1643678851
transform 1 0 17894 0 1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_552
timestamp 1643678851
transform 1 0 17894 0 -1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_553
timestamp 1643678851
transform 1 0 17894 0 1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_554
timestamp 1643678851
transform 1 0 17894 0 -1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_555
timestamp 1643678851
transform 1 0 17894 0 1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_556
timestamp 1643678851
transform 1 0 17894 0 -1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_557
timestamp 1643678851
transform 1 0 17894 0 1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_558
timestamp 1643678851
transform 1 0 17894 0 -1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_559
timestamp 1643678851
transform 1 0 17894 0 1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_560
timestamp 1643678851
transform 1 0 17894 0 -1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_561
timestamp 1643678851
transform 1 0 17894 0 1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_562
timestamp 1643678851
transform 1 0 17894 0 -1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_563
timestamp 1643678851
transform 1 0 17894 0 1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_564
timestamp 1643678851
transform 1 0 17894 0 -1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_565
timestamp 1643678851
transform 1 0 17894 0 1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_566
timestamp 1643678851
transform 1 0 17894 0 -1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_567
timestamp 1643678851
transform 1 0 17894 0 1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_568
timestamp 1643678851
transform 1 0 17894 0 -1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_569
timestamp 1643678851
transform 1 0 17894 0 1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_570
timestamp 1643678851
transform 1 0 17894 0 -1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_571
timestamp 1643678851
transform 1 0 17894 0 1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_572
timestamp 1643678851
transform 1 0 17894 0 -1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_573
timestamp 1643678851
transform 1 0 17894 0 1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_574
timestamp 1643678851
transform 1 0 17894 0 -1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_575
timestamp 1643678851
transform 1 0 17894 0 1 0
box 0 -21 389 808
use cell_2r1w  cell_2r1w_576
timestamp 1643678851
transform 1 0 17505 0 -1 24640
box 0 -21 389 808
use cell_2r1w  cell_2r1w_577
timestamp 1643678851
transform 1 0 17505 0 1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_578
timestamp 1643678851
transform 1 0 17505 0 -1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_579
timestamp 1643678851
transform 1 0 17505 0 1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_580
timestamp 1643678851
transform 1 0 17505 0 -1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_581
timestamp 1643678851
transform 1 0 17505 0 1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_582
timestamp 1643678851
transform 1 0 17505 0 -1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_583
timestamp 1643678851
transform 1 0 17505 0 1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_584
timestamp 1643678851
transform 1 0 17505 0 -1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_585
timestamp 1643678851
transform 1 0 17505 0 1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_586
timestamp 1643678851
transform 1 0 17505 0 -1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_587
timestamp 1643678851
transform 1 0 17505 0 1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_588
timestamp 1643678851
transform 1 0 17505 0 -1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_589
timestamp 1643678851
transform 1 0 17505 0 1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_590
timestamp 1643678851
transform 1 0 17505 0 -1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_591
timestamp 1643678851
transform 1 0 17505 0 1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_592
timestamp 1643678851
transform 1 0 17505 0 -1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_593
timestamp 1643678851
transform 1 0 17505 0 1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_594
timestamp 1643678851
transform 1 0 17505 0 -1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_595
timestamp 1643678851
transform 1 0 17505 0 1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_596
timestamp 1643678851
transform 1 0 17505 0 -1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_597
timestamp 1643678851
transform 1 0 17505 0 1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_598
timestamp 1643678851
transform 1 0 17505 0 -1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_599
timestamp 1643678851
transform 1 0 17505 0 1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_600
timestamp 1643678851
transform 1 0 17505 0 -1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_601
timestamp 1643678851
transform 1 0 17505 0 1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_602
timestamp 1643678851
transform 1 0 17505 0 -1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_603
timestamp 1643678851
transform 1 0 17505 0 1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_604
timestamp 1643678851
transform 1 0 17505 0 -1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_605
timestamp 1643678851
transform 1 0 17505 0 1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_606
timestamp 1643678851
transform 1 0 17505 0 -1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_607
timestamp 1643678851
transform 1 0 17505 0 1 0
box 0 -21 389 808
use cell_2r1w  cell_2r1w_608
timestamp 1643678851
transform 1 0 17116 0 -1 24640
box 0 -21 389 808
use cell_2r1w  cell_2r1w_609
timestamp 1643678851
transform 1 0 17116 0 1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_610
timestamp 1643678851
transform 1 0 17116 0 -1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_611
timestamp 1643678851
transform 1 0 17116 0 1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_612
timestamp 1643678851
transform 1 0 17116 0 -1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_613
timestamp 1643678851
transform 1 0 17116 0 1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_614
timestamp 1643678851
transform 1 0 17116 0 -1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_615
timestamp 1643678851
transform 1 0 17116 0 1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_616
timestamp 1643678851
transform 1 0 17116 0 -1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_617
timestamp 1643678851
transform 1 0 17116 0 1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_618
timestamp 1643678851
transform 1 0 17116 0 -1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_619
timestamp 1643678851
transform 1 0 17116 0 1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_620
timestamp 1643678851
transform 1 0 17116 0 -1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_621
timestamp 1643678851
transform 1 0 17116 0 1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_622
timestamp 1643678851
transform 1 0 17116 0 -1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_623
timestamp 1643678851
transform 1 0 17116 0 1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_624
timestamp 1643678851
transform 1 0 17116 0 -1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_625
timestamp 1643678851
transform 1 0 17116 0 1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_626
timestamp 1643678851
transform 1 0 17116 0 -1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_627
timestamp 1643678851
transform 1 0 17116 0 1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_628
timestamp 1643678851
transform 1 0 17116 0 -1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_629
timestamp 1643678851
transform 1 0 17116 0 1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_630
timestamp 1643678851
transform 1 0 17116 0 -1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_631
timestamp 1643678851
transform 1 0 17116 0 1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_632
timestamp 1643678851
transform 1 0 17116 0 -1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_633
timestamp 1643678851
transform 1 0 17116 0 1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_634
timestamp 1643678851
transform 1 0 17116 0 -1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_635
timestamp 1643678851
transform 1 0 17116 0 1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_636
timestamp 1643678851
transform 1 0 17116 0 -1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_637
timestamp 1643678851
transform 1 0 17116 0 1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_638
timestamp 1643678851
transform 1 0 17116 0 -1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_639
timestamp 1643678851
transform 1 0 17116 0 1 0
box 0 -21 389 808
use cell_2r1w  cell_2r1w_640
timestamp 1643678851
transform 1 0 16727 0 -1 24640
box 0 -21 389 808
use cell_2r1w  cell_2r1w_641
timestamp 1643678851
transform 1 0 16727 0 1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_642
timestamp 1643678851
transform 1 0 16727 0 -1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_643
timestamp 1643678851
transform 1 0 16727 0 1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_644
timestamp 1643678851
transform 1 0 16727 0 -1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_645
timestamp 1643678851
transform 1 0 16727 0 1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_646
timestamp 1643678851
transform 1 0 16727 0 -1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_647
timestamp 1643678851
transform 1 0 16727 0 1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_648
timestamp 1643678851
transform 1 0 16727 0 -1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_649
timestamp 1643678851
transform 1 0 16727 0 1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_650
timestamp 1643678851
transform 1 0 16727 0 -1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_651
timestamp 1643678851
transform 1 0 16727 0 1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_652
timestamp 1643678851
transform 1 0 16727 0 -1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_653
timestamp 1643678851
transform 1 0 16727 0 1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_654
timestamp 1643678851
transform 1 0 16727 0 -1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_655
timestamp 1643678851
transform 1 0 16727 0 1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_656
timestamp 1643678851
transform 1 0 16727 0 -1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_657
timestamp 1643678851
transform 1 0 16727 0 1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_658
timestamp 1643678851
transform 1 0 16727 0 -1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_659
timestamp 1643678851
transform 1 0 16727 0 1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_660
timestamp 1643678851
transform 1 0 16727 0 -1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_661
timestamp 1643678851
transform 1 0 16727 0 1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_662
timestamp 1643678851
transform 1 0 16727 0 -1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_663
timestamp 1643678851
transform 1 0 16727 0 1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_664
timestamp 1643678851
transform 1 0 16727 0 -1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_665
timestamp 1643678851
transform 1 0 16727 0 1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_666
timestamp 1643678851
transform 1 0 16727 0 -1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_667
timestamp 1643678851
transform 1 0 16727 0 1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_668
timestamp 1643678851
transform 1 0 16727 0 -1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_669
timestamp 1643678851
transform 1 0 16727 0 1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_670
timestamp 1643678851
transform 1 0 16727 0 -1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_671
timestamp 1643678851
transform 1 0 16727 0 1 0
box 0 -21 389 808
use cell_2r1w  cell_2r1w_672
timestamp 1643678851
transform 1 0 16338 0 -1 24640
box 0 -21 389 808
use cell_2r1w  cell_2r1w_673
timestamp 1643678851
transform 1 0 16338 0 1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_674
timestamp 1643678851
transform 1 0 16338 0 -1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_675
timestamp 1643678851
transform 1 0 16338 0 1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_676
timestamp 1643678851
transform 1 0 16338 0 -1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_677
timestamp 1643678851
transform 1 0 16338 0 1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_678
timestamp 1643678851
transform 1 0 16338 0 -1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_679
timestamp 1643678851
transform 1 0 16338 0 1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_680
timestamp 1643678851
transform 1 0 16338 0 -1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_681
timestamp 1643678851
transform 1 0 16338 0 1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_682
timestamp 1643678851
transform 1 0 16338 0 -1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_683
timestamp 1643678851
transform 1 0 16338 0 1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_684
timestamp 1643678851
transform 1 0 16338 0 -1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_685
timestamp 1643678851
transform 1 0 16338 0 1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_686
timestamp 1643678851
transform 1 0 16338 0 -1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_687
timestamp 1643678851
transform 1 0 16338 0 1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_688
timestamp 1643678851
transform 1 0 16338 0 -1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_689
timestamp 1643678851
transform 1 0 16338 0 1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_690
timestamp 1643678851
transform 1 0 16338 0 -1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_691
timestamp 1643678851
transform 1 0 16338 0 1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_692
timestamp 1643678851
transform 1 0 16338 0 -1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_693
timestamp 1643678851
transform 1 0 16338 0 1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_694
timestamp 1643678851
transform 1 0 16338 0 -1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_695
timestamp 1643678851
transform 1 0 16338 0 1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_696
timestamp 1643678851
transform 1 0 16338 0 -1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_697
timestamp 1643678851
transform 1 0 16338 0 1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_698
timestamp 1643678851
transform 1 0 16338 0 -1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_699
timestamp 1643678851
transform 1 0 16338 0 1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_700
timestamp 1643678851
transform 1 0 16338 0 -1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_701
timestamp 1643678851
transform 1 0 16338 0 1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_702
timestamp 1643678851
transform 1 0 16338 0 -1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_703
timestamp 1643678851
transform 1 0 16338 0 1 0
box 0 -21 389 808
use cell_2r1w  cell_2r1w_704
timestamp 1643678851
transform 1 0 15949 0 -1 24640
box 0 -21 389 808
use cell_2r1w  cell_2r1w_705
timestamp 1643678851
transform 1 0 15949 0 1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_706
timestamp 1643678851
transform 1 0 15949 0 -1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_707
timestamp 1643678851
transform 1 0 15949 0 1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_708
timestamp 1643678851
transform 1 0 15949 0 -1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_709
timestamp 1643678851
transform 1 0 15949 0 1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_710
timestamp 1643678851
transform 1 0 15949 0 -1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_711
timestamp 1643678851
transform 1 0 15949 0 1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_712
timestamp 1643678851
transform 1 0 15949 0 -1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_713
timestamp 1643678851
transform 1 0 15949 0 1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_714
timestamp 1643678851
transform 1 0 15949 0 -1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_715
timestamp 1643678851
transform 1 0 15949 0 1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_716
timestamp 1643678851
transform 1 0 15949 0 -1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_717
timestamp 1643678851
transform 1 0 15949 0 1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_718
timestamp 1643678851
transform 1 0 15949 0 -1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_719
timestamp 1643678851
transform 1 0 15949 0 1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_720
timestamp 1643678851
transform 1 0 15949 0 -1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_721
timestamp 1643678851
transform 1 0 15949 0 1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_722
timestamp 1643678851
transform 1 0 15949 0 -1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_723
timestamp 1643678851
transform 1 0 15949 0 1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_724
timestamp 1643678851
transform 1 0 15949 0 -1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_725
timestamp 1643678851
transform 1 0 15949 0 1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_726
timestamp 1643678851
transform 1 0 15949 0 -1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_727
timestamp 1643678851
transform 1 0 15949 0 1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_728
timestamp 1643678851
transform 1 0 15949 0 -1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_729
timestamp 1643678851
transform 1 0 15949 0 1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_730
timestamp 1643678851
transform 1 0 15949 0 -1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_731
timestamp 1643678851
transform 1 0 15949 0 1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_732
timestamp 1643678851
transform 1 0 15949 0 -1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_733
timestamp 1643678851
transform 1 0 15949 0 1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_734
timestamp 1643678851
transform 1 0 15949 0 -1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_735
timestamp 1643678851
transform 1 0 15949 0 1 0
box 0 -21 389 808
use cell_2r1w  cell_2r1w_736
timestamp 1643678851
transform 1 0 15560 0 -1 24640
box 0 -21 389 808
use cell_2r1w  cell_2r1w_737
timestamp 1643678851
transform 1 0 15560 0 1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_738
timestamp 1643678851
transform 1 0 15560 0 -1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_739
timestamp 1643678851
transform 1 0 15560 0 1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_740
timestamp 1643678851
transform 1 0 15560 0 -1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_741
timestamp 1643678851
transform 1 0 15560 0 1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_742
timestamp 1643678851
transform 1 0 15560 0 -1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_743
timestamp 1643678851
transform 1 0 15560 0 1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_744
timestamp 1643678851
transform 1 0 15560 0 -1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_745
timestamp 1643678851
transform 1 0 15560 0 1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_746
timestamp 1643678851
transform 1 0 15560 0 -1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_747
timestamp 1643678851
transform 1 0 15560 0 1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_748
timestamp 1643678851
transform 1 0 15560 0 -1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_749
timestamp 1643678851
transform 1 0 15560 0 1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_750
timestamp 1643678851
transform 1 0 15560 0 -1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_751
timestamp 1643678851
transform 1 0 15560 0 1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_752
timestamp 1643678851
transform 1 0 15560 0 -1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_753
timestamp 1643678851
transform 1 0 15560 0 1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_754
timestamp 1643678851
transform 1 0 15560 0 -1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_755
timestamp 1643678851
transform 1 0 15560 0 1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_756
timestamp 1643678851
transform 1 0 15560 0 -1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_757
timestamp 1643678851
transform 1 0 15560 0 1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_758
timestamp 1643678851
transform 1 0 15560 0 -1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_759
timestamp 1643678851
transform 1 0 15560 0 1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_760
timestamp 1643678851
transform 1 0 15560 0 -1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_761
timestamp 1643678851
transform 1 0 15560 0 1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_762
timestamp 1643678851
transform 1 0 15560 0 -1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_763
timestamp 1643678851
transform 1 0 15560 0 1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_764
timestamp 1643678851
transform 1 0 15560 0 -1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_765
timestamp 1643678851
transform 1 0 15560 0 1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_766
timestamp 1643678851
transform 1 0 15560 0 -1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_767
timestamp 1643678851
transform 1 0 15560 0 1 0
box 0 -21 389 808
use cell_2r1w  cell_2r1w_768
timestamp 1643678851
transform 1 0 15171 0 -1 24640
box 0 -21 389 808
use cell_2r1w  cell_2r1w_769
timestamp 1643678851
transform 1 0 15171 0 1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_770
timestamp 1643678851
transform 1 0 15171 0 -1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_771
timestamp 1643678851
transform 1 0 15171 0 1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_772
timestamp 1643678851
transform 1 0 15171 0 -1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_773
timestamp 1643678851
transform 1 0 15171 0 1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_774
timestamp 1643678851
transform 1 0 15171 0 -1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_775
timestamp 1643678851
transform 1 0 15171 0 1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_776
timestamp 1643678851
transform 1 0 15171 0 -1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_777
timestamp 1643678851
transform 1 0 15171 0 1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_778
timestamp 1643678851
transform 1 0 15171 0 -1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_779
timestamp 1643678851
transform 1 0 15171 0 1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_780
timestamp 1643678851
transform 1 0 15171 0 -1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_781
timestamp 1643678851
transform 1 0 15171 0 1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_782
timestamp 1643678851
transform 1 0 15171 0 -1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_783
timestamp 1643678851
transform 1 0 15171 0 1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_784
timestamp 1643678851
transform 1 0 15171 0 -1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_785
timestamp 1643678851
transform 1 0 15171 0 1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_786
timestamp 1643678851
transform 1 0 15171 0 -1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_787
timestamp 1643678851
transform 1 0 15171 0 1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_788
timestamp 1643678851
transform 1 0 15171 0 -1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_789
timestamp 1643678851
transform 1 0 15171 0 1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_790
timestamp 1643678851
transform 1 0 15171 0 -1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_791
timestamp 1643678851
transform 1 0 15171 0 1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_792
timestamp 1643678851
transform 1 0 15171 0 -1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_793
timestamp 1643678851
transform 1 0 15171 0 1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_794
timestamp 1643678851
transform 1 0 15171 0 -1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_795
timestamp 1643678851
transform 1 0 15171 0 1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_796
timestamp 1643678851
transform 1 0 15171 0 -1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_797
timestamp 1643678851
transform 1 0 15171 0 1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_798
timestamp 1643678851
transform 1 0 15171 0 -1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_799
timestamp 1643678851
transform 1 0 15171 0 1 0
box 0 -21 389 808
use cell_2r1w  cell_2r1w_800
timestamp 1643678851
transform 1 0 14782 0 -1 24640
box 0 -21 389 808
use cell_2r1w  cell_2r1w_801
timestamp 1643678851
transform 1 0 14782 0 1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_802
timestamp 1643678851
transform 1 0 14782 0 -1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_803
timestamp 1643678851
transform 1 0 14782 0 1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_804
timestamp 1643678851
transform 1 0 14782 0 -1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_805
timestamp 1643678851
transform 1 0 14782 0 1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_806
timestamp 1643678851
transform 1 0 14782 0 -1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_807
timestamp 1643678851
transform 1 0 14782 0 1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_808
timestamp 1643678851
transform 1 0 14782 0 -1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_809
timestamp 1643678851
transform 1 0 14782 0 1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_810
timestamp 1643678851
transform 1 0 14782 0 -1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_811
timestamp 1643678851
transform 1 0 14782 0 1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_812
timestamp 1643678851
transform 1 0 14782 0 -1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_813
timestamp 1643678851
transform 1 0 14782 0 1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_814
timestamp 1643678851
transform 1 0 14782 0 -1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_815
timestamp 1643678851
transform 1 0 14782 0 1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_816
timestamp 1643678851
transform 1 0 14782 0 -1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_817
timestamp 1643678851
transform 1 0 14782 0 1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_818
timestamp 1643678851
transform 1 0 14782 0 -1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_819
timestamp 1643678851
transform 1 0 14782 0 1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_820
timestamp 1643678851
transform 1 0 14782 0 -1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_821
timestamp 1643678851
transform 1 0 14782 0 1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_822
timestamp 1643678851
transform 1 0 14782 0 -1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_823
timestamp 1643678851
transform 1 0 14782 0 1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_824
timestamp 1643678851
transform 1 0 14782 0 -1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_825
timestamp 1643678851
transform 1 0 14782 0 1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_826
timestamp 1643678851
transform 1 0 14782 0 -1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_827
timestamp 1643678851
transform 1 0 14782 0 1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_828
timestamp 1643678851
transform 1 0 14782 0 -1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_829
timestamp 1643678851
transform 1 0 14782 0 1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_830
timestamp 1643678851
transform 1 0 14782 0 -1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_831
timestamp 1643678851
transform 1 0 14782 0 1 0
box 0 -21 389 808
use cell_2r1w  cell_2r1w_832
timestamp 1643678851
transform 1 0 14393 0 -1 24640
box 0 -21 389 808
use cell_2r1w  cell_2r1w_833
timestamp 1643678851
transform 1 0 14393 0 1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_834
timestamp 1643678851
transform 1 0 14393 0 -1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_835
timestamp 1643678851
transform 1 0 14393 0 1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_836
timestamp 1643678851
transform 1 0 14393 0 -1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_837
timestamp 1643678851
transform 1 0 14393 0 1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_838
timestamp 1643678851
transform 1 0 14393 0 -1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_839
timestamp 1643678851
transform 1 0 14393 0 1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_840
timestamp 1643678851
transform 1 0 14393 0 -1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_841
timestamp 1643678851
transform 1 0 14393 0 1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_842
timestamp 1643678851
transform 1 0 14393 0 -1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_843
timestamp 1643678851
transform 1 0 14393 0 1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_844
timestamp 1643678851
transform 1 0 14393 0 -1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_845
timestamp 1643678851
transform 1 0 14393 0 1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_846
timestamp 1643678851
transform 1 0 14393 0 -1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_847
timestamp 1643678851
transform 1 0 14393 0 1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_848
timestamp 1643678851
transform 1 0 14393 0 -1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_849
timestamp 1643678851
transform 1 0 14393 0 1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_850
timestamp 1643678851
transform 1 0 14393 0 -1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_851
timestamp 1643678851
transform 1 0 14393 0 1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_852
timestamp 1643678851
transform 1 0 14393 0 -1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_853
timestamp 1643678851
transform 1 0 14393 0 1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_854
timestamp 1643678851
transform 1 0 14393 0 -1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_855
timestamp 1643678851
transform 1 0 14393 0 1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_856
timestamp 1643678851
transform 1 0 14393 0 -1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_857
timestamp 1643678851
transform 1 0 14393 0 1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_858
timestamp 1643678851
transform 1 0 14393 0 -1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_859
timestamp 1643678851
transform 1 0 14393 0 1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_860
timestamp 1643678851
transform 1 0 14393 0 -1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_861
timestamp 1643678851
transform 1 0 14393 0 1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_862
timestamp 1643678851
transform 1 0 14393 0 -1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_863
timestamp 1643678851
transform 1 0 14393 0 1 0
box 0 -21 389 808
use cell_2r1w  cell_2r1w_864
timestamp 1643678851
transform 1 0 14004 0 -1 24640
box 0 -21 389 808
use cell_2r1w  cell_2r1w_865
timestamp 1643678851
transform 1 0 14004 0 1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_866
timestamp 1643678851
transform 1 0 14004 0 -1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_867
timestamp 1643678851
transform 1 0 14004 0 1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_868
timestamp 1643678851
transform 1 0 14004 0 -1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_869
timestamp 1643678851
transform 1 0 14004 0 1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_870
timestamp 1643678851
transform 1 0 14004 0 -1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_871
timestamp 1643678851
transform 1 0 14004 0 1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_872
timestamp 1643678851
transform 1 0 14004 0 -1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_873
timestamp 1643678851
transform 1 0 14004 0 1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_874
timestamp 1643678851
transform 1 0 14004 0 -1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_875
timestamp 1643678851
transform 1 0 14004 0 1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_876
timestamp 1643678851
transform 1 0 14004 0 -1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_877
timestamp 1643678851
transform 1 0 14004 0 1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_878
timestamp 1643678851
transform 1 0 14004 0 -1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_879
timestamp 1643678851
transform 1 0 14004 0 1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_880
timestamp 1643678851
transform 1 0 14004 0 -1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_881
timestamp 1643678851
transform 1 0 14004 0 1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_882
timestamp 1643678851
transform 1 0 14004 0 -1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_883
timestamp 1643678851
transform 1 0 14004 0 1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_884
timestamp 1643678851
transform 1 0 14004 0 -1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_885
timestamp 1643678851
transform 1 0 14004 0 1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_886
timestamp 1643678851
transform 1 0 14004 0 -1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_887
timestamp 1643678851
transform 1 0 14004 0 1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_888
timestamp 1643678851
transform 1 0 14004 0 -1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_889
timestamp 1643678851
transform 1 0 14004 0 1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_890
timestamp 1643678851
transform 1 0 14004 0 -1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_891
timestamp 1643678851
transform 1 0 14004 0 1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_892
timestamp 1643678851
transform 1 0 14004 0 -1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_893
timestamp 1643678851
transform 1 0 14004 0 1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_894
timestamp 1643678851
transform 1 0 14004 0 -1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_895
timestamp 1643678851
transform 1 0 14004 0 1 0
box 0 -21 389 808
use cell_2r1w  cell_2r1w_896
timestamp 1643678851
transform 1 0 13615 0 -1 24640
box 0 -21 389 808
use cell_2r1w  cell_2r1w_897
timestamp 1643678851
transform 1 0 13615 0 1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_898
timestamp 1643678851
transform 1 0 13615 0 -1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_899
timestamp 1643678851
transform 1 0 13615 0 1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_900
timestamp 1643678851
transform 1 0 13615 0 -1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_901
timestamp 1643678851
transform 1 0 13615 0 1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_902
timestamp 1643678851
transform 1 0 13615 0 -1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_903
timestamp 1643678851
transform 1 0 13615 0 1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_904
timestamp 1643678851
transform 1 0 13615 0 -1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_905
timestamp 1643678851
transform 1 0 13615 0 1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_906
timestamp 1643678851
transform 1 0 13615 0 -1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_907
timestamp 1643678851
transform 1 0 13615 0 1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_908
timestamp 1643678851
transform 1 0 13615 0 -1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_909
timestamp 1643678851
transform 1 0 13615 0 1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_910
timestamp 1643678851
transform 1 0 13615 0 -1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_911
timestamp 1643678851
transform 1 0 13615 0 1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_912
timestamp 1643678851
transform 1 0 13615 0 -1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_913
timestamp 1643678851
transform 1 0 13615 0 1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_914
timestamp 1643678851
transform 1 0 13615 0 -1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_915
timestamp 1643678851
transform 1 0 13615 0 1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_916
timestamp 1643678851
transform 1 0 13615 0 -1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_917
timestamp 1643678851
transform 1 0 13615 0 1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_918
timestamp 1643678851
transform 1 0 13615 0 -1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_919
timestamp 1643678851
transform 1 0 13615 0 1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_920
timestamp 1643678851
transform 1 0 13615 0 -1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_921
timestamp 1643678851
transform 1 0 13615 0 1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_922
timestamp 1643678851
transform 1 0 13615 0 -1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_923
timestamp 1643678851
transform 1 0 13615 0 1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_924
timestamp 1643678851
transform 1 0 13615 0 -1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_925
timestamp 1643678851
transform 1 0 13615 0 1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_926
timestamp 1643678851
transform 1 0 13615 0 -1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_927
timestamp 1643678851
transform 1 0 13615 0 1 0
box 0 -21 389 808
use cell_2r1w  cell_2r1w_928
timestamp 1643678851
transform 1 0 13226 0 -1 24640
box 0 -21 389 808
use cell_2r1w  cell_2r1w_929
timestamp 1643678851
transform 1 0 13226 0 1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_930
timestamp 1643678851
transform 1 0 13226 0 -1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_931
timestamp 1643678851
transform 1 0 13226 0 1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_932
timestamp 1643678851
transform 1 0 13226 0 -1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_933
timestamp 1643678851
transform 1 0 13226 0 1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_934
timestamp 1643678851
transform 1 0 13226 0 -1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_935
timestamp 1643678851
transform 1 0 13226 0 1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_936
timestamp 1643678851
transform 1 0 13226 0 -1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_937
timestamp 1643678851
transform 1 0 13226 0 1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_938
timestamp 1643678851
transform 1 0 13226 0 -1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_939
timestamp 1643678851
transform 1 0 13226 0 1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_940
timestamp 1643678851
transform 1 0 13226 0 -1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_941
timestamp 1643678851
transform 1 0 13226 0 1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_942
timestamp 1643678851
transform 1 0 13226 0 -1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_943
timestamp 1643678851
transform 1 0 13226 0 1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_944
timestamp 1643678851
transform 1 0 13226 0 -1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_945
timestamp 1643678851
transform 1 0 13226 0 1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_946
timestamp 1643678851
transform 1 0 13226 0 -1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_947
timestamp 1643678851
transform 1 0 13226 0 1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_948
timestamp 1643678851
transform 1 0 13226 0 -1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_949
timestamp 1643678851
transform 1 0 13226 0 1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_950
timestamp 1643678851
transform 1 0 13226 0 -1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_951
timestamp 1643678851
transform 1 0 13226 0 1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_952
timestamp 1643678851
transform 1 0 13226 0 -1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_953
timestamp 1643678851
transform 1 0 13226 0 1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_954
timestamp 1643678851
transform 1 0 13226 0 -1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_955
timestamp 1643678851
transform 1 0 13226 0 1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_956
timestamp 1643678851
transform 1 0 13226 0 -1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_957
timestamp 1643678851
transform 1 0 13226 0 1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_958
timestamp 1643678851
transform 1 0 13226 0 -1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_959
timestamp 1643678851
transform 1 0 13226 0 1 0
box 0 -21 389 808
use cell_2r1w  cell_2r1w_960
timestamp 1643678851
transform 1 0 12837 0 -1 24640
box 0 -21 389 808
use cell_2r1w  cell_2r1w_961
timestamp 1643678851
transform 1 0 12837 0 1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_962
timestamp 1643678851
transform 1 0 12837 0 -1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_963
timestamp 1643678851
transform 1 0 12837 0 1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_964
timestamp 1643678851
transform 1 0 12837 0 -1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_965
timestamp 1643678851
transform 1 0 12837 0 1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_966
timestamp 1643678851
transform 1 0 12837 0 -1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_967
timestamp 1643678851
transform 1 0 12837 0 1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_968
timestamp 1643678851
transform 1 0 12837 0 -1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_969
timestamp 1643678851
transform 1 0 12837 0 1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_970
timestamp 1643678851
transform 1 0 12837 0 -1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_971
timestamp 1643678851
transform 1 0 12837 0 1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_972
timestamp 1643678851
transform 1 0 12837 0 -1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_973
timestamp 1643678851
transform 1 0 12837 0 1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_974
timestamp 1643678851
transform 1 0 12837 0 -1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_975
timestamp 1643678851
transform 1 0 12837 0 1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_976
timestamp 1643678851
transform 1 0 12837 0 -1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_977
timestamp 1643678851
transform 1 0 12837 0 1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_978
timestamp 1643678851
transform 1 0 12837 0 -1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_979
timestamp 1643678851
transform 1 0 12837 0 1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_980
timestamp 1643678851
transform 1 0 12837 0 -1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_981
timestamp 1643678851
transform 1 0 12837 0 1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_982
timestamp 1643678851
transform 1 0 12837 0 -1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_983
timestamp 1643678851
transform 1 0 12837 0 1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_984
timestamp 1643678851
transform 1 0 12837 0 -1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_985
timestamp 1643678851
transform 1 0 12837 0 1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_986
timestamp 1643678851
transform 1 0 12837 0 -1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_987
timestamp 1643678851
transform 1 0 12837 0 1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_988
timestamp 1643678851
transform 1 0 12837 0 -1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_989
timestamp 1643678851
transform 1 0 12837 0 1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_990
timestamp 1643678851
transform 1 0 12837 0 -1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_991
timestamp 1643678851
transform 1 0 12837 0 1 0
box 0 -21 389 808
use cell_2r1w  cell_2r1w_992
timestamp 1643678851
transform 1 0 12448 0 -1 24640
box 0 -21 389 808
use cell_2r1w  cell_2r1w_993
timestamp 1643678851
transform 1 0 12448 0 1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_994
timestamp 1643678851
transform 1 0 12448 0 -1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_995
timestamp 1643678851
transform 1 0 12448 0 1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_996
timestamp 1643678851
transform 1 0 12448 0 -1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_997
timestamp 1643678851
transform 1 0 12448 0 1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_998
timestamp 1643678851
transform 1 0 12448 0 -1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_999
timestamp 1643678851
transform 1 0 12448 0 1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1000
timestamp 1643678851
transform 1 0 12448 0 -1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1001
timestamp 1643678851
transform 1 0 12448 0 1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1002
timestamp 1643678851
transform 1 0 12448 0 -1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1003
timestamp 1643678851
transform 1 0 12448 0 1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1004
timestamp 1643678851
transform 1 0 12448 0 -1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1005
timestamp 1643678851
transform 1 0 12448 0 1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1006
timestamp 1643678851
transform 1 0 12448 0 -1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1007
timestamp 1643678851
transform 1 0 12448 0 1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1008
timestamp 1643678851
transform 1 0 12448 0 -1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1009
timestamp 1643678851
transform 1 0 12448 0 1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1010
timestamp 1643678851
transform 1 0 12448 0 -1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1011
timestamp 1643678851
transform 1 0 12448 0 1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1012
timestamp 1643678851
transform 1 0 12448 0 -1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1013
timestamp 1643678851
transform 1 0 12448 0 1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1014
timestamp 1643678851
transform 1 0 12448 0 -1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1015
timestamp 1643678851
transform 1 0 12448 0 1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1016
timestamp 1643678851
transform 1 0 12448 0 -1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1017
timestamp 1643678851
transform 1 0 12448 0 1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1018
timestamp 1643678851
transform 1 0 12448 0 -1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1019
timestamp 1643678851
transform 1 0 12448 0 1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1020
timestamp 1643678851
transform 1 0 12448 0 -1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1021
timestamp 1643678851
transform 1 0 12448 0 1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1022
timestamp 1643678851
transform 1 0 12448 0 -1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1023
timestamp 1643678851
transform 1 0 12448 0 1 0
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1024
timestamp 1643678851
transform 1 0 12059 0 -1 24640
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1025
timestamp 1643678851
transform 1 0 12059 0 1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1026
timestamp 1643678851
transform 1 0 12059 0 -1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1027
timestamp 1643678851
transform 1 0 12059 0 1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1028
timestamp 1643678851
transform 1 0 12059 0 -1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1029
timestamp 1643678851
transform 1 0 12059 0 1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1030
timestamp 1643678851
transform 1 0 12059 0 -1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1031
timestamp 1643678851
transform 1 0 12059 0 1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1032
timestamp 1643678851
transform 1 0 12059 0 -1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1033
timestamp 1643678851
transform 1 0 12059 0 1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1034
timestamp 1643678851
transform 1 0 12059 0 -1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1035
timestamp 1643678851
transform 1 0 12059 0 1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1036
timestamp 1643678851
transform 1 0 12059 0 -1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1037
timestamp 1643678851
transform 1 0 12059 0 1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1038
timestamp 1643678851
transform 1 0 12059 0 -1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1039
timestamp 1643678851
transform 1 0 12059 0 1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1040
timestamp 1643678851
transform 1 0 12059 0 -1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1041
timestamp 1643678851
transform 1 0 12059 0 1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1042
timestamp 1643678851
transform 1 0 12059 0 -1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1043
timestamp 1643678851
transform 1 0 12059 0 1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1044
timestamp 1643678851
transform 1 0 12059 0 -1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1045
timestamp 1643678851
transform 1 0 12059 0 1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1046
timestamp 1643678851
transform 1 0 12059 0 -1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1047
timestamp 1643678851
transform 1 0 12059 0 1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1048
timestamp 1643678851
transform 1 0 12059 0 -1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1049
timestamp 1643678851
transform 1 0 12059 0 1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1050
timestamp 1643678851
transform 1 0 12059 0 -1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1051
timestamp 1643678851
transform 1 0 12059 0 1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1052
timestamp 1643678851
transform 1 0 12059 0 -1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1053
timestamp 1643678851
transform 1 0 12059 0 1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1054
timestamp 1643678851
transform 1 0 12059 0 -1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1055
timestamp 1643678851
transform 1 0 12059 0 1 0
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1056
timestamp 1643678851
transform 1 0 11670 0 -1 24640
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1057
timestamp 1643678851
transform 1 0 11670 0 1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1058
timestamp 1643678851
transform 1 0 11670 0 -1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1059
timestamp 1643678851
transform 1 0 11670 0 1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1060
timestamp 1643678851
transform 1 0 11670 0 -1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1061
timestamp 1643678851
transform 1 0 11670 0 1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1062
timestamp 1643678851
transform 1 0 11670 0 -1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1063
timestamp 1643678851
transform 1 0 11670 0 1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1064
timestamp 1643678851
transform 1 0 11670 0 -1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1065
timestamp 1643678851
transform 1 0 11670 0 1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1066
timestamp 1643678851
transform 1 0 11670 0 -1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1067
timestamp 1643678851
transform 1 0 11670 0 1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1068
timestamp 1643678851
transform 1 0 11670 0 -1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1069
timestamp 1643678851
transform 1 0 11670 0 1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1070
timestamp 1643678851
transform 1 0 11670 0 -1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1071
timestamp 1643678851
transform 1 0 11670 0 1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1072
timestamp 1643678851
transform 1 0 11670 0 -1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1073
timestamp 1643678851
transform 1 0 11670 0 1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1074
timestamp 1643678851
transform 1 0 11670 0 -1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1075
timestamp 1643678851
transform 1 0 11670 0 1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1076
timestamp 1643678851
transform 1 0 11670 0 -1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1077
timestamp 1643678851
transform 1 0 11670 0 1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1078
timestamp 1643678851
transform 1 0 11670 0 -1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1079
timestamp 1643678851
transform 1 0 11670 0 1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1080
timestamp 1643678851
transform 1 0 11670 0 -1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1081
timestamp 1643678851
transform 1 0 11670 0 1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1082
timestamp 1643678851
transform 1 0 11670 0 -1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1083
timestamp 1643678851
transform 1 0 11670 0 1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1084
timestamp 1643678851
transform 1 0 11670 0 -1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1085
timestamp 1643678851
transform 1 0 11670 0 1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1086
timestamp 1643678851
transform 1 0 11670 0 -1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1087
timestamp 1643678851
transform 1 0 11670 0 1 0
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1088
timestamp 1643678851
transform 1 0 11281 0 -1 24640
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1089
timestamp 1643678851
transform 1 0 11281 0 1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1090
timestamp 1643678851
transform 1 0 11281 0 -1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1091
timestamp 1643678851
transform 1 0 11281 0 1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1092
timestamp 1643678851
transform 1 0 11281 0 -1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1093
timestamp 1643678851
transform 1 0 11281 0 1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1094
timestamp 1643678851
transform 1 0 11281 0 -1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1095
timestamp 1643678851
transform 1 0 11281 0 1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1096
timestamp 1643678851
transform 1 0 11281 0 -1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1097
timestamp 1643678851
transform 1 0 11281 0 1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1098
timestamp 1643678851
transform 1 0 11281 0 -1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1099
timestamp 1643678851
transform 1 0 11281 0 1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1100
timestamp 1643678851
transform 1 0 11281 0 -1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1101
timestamp 1643678851
transform 1 0 11281 0 1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1102
timestamp 1643678851
transform 1 0 11281 0 -1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1103
timestamp 1643678851
transform 1 0 11281 0 1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1104
timestamp 1643678851
transform 1 0 11281 0 -1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1105
timestamp 1643678851
transform 1 0 11281 0 1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1106
timestamp 1643678851
transform 1 0 11281 0 -1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1107
timestamp 1643678851
transform 1 0 11281 0 1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1108
timestamp 1643678851
transform 1 0 11281 0 -1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1109
timestamp 1643678851
transform 1 0 11281 0 1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1110
timestamp 1643678851
transform 1 0 11281 0 -1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1111
timestamp 1643678851
transform 1 0 11281 0 1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1112
timestamp 1643678851
transform 1 0 11281 0 -1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1113
timestamp 1643678851
transform 1 0 11281 0 1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1114
timestamp 1643678851
transform 1 0 11281 0 -1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1115
timestamp 1643678851
transform 1 0 11281 0 1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1116
timestamp 1643678851
transform 1 0 11281 0 -1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1117
timestamp 1643678851
transform 1 0 11281 0 1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1118
timestamp 1643678851
transform 1 0 11281 0 -1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1119
timestamp 1643678851
transform 1 0 11281 0 1 0
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1120
timestamp 1643678851
transform 1 0 10892 0 -1 24640
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1121
timestamp 1643678851
transform 1 0 10892 0 1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1122
timestamp 1643678851
transform 1 0 10892 0 -1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1123
timestamp 1643678851
transform 1 0 10892 0 1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1124
timestamp 1643678851
transform 1 0 10892 0 -1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1125
timestamp 1643678851
transform 1 0 10892 0 1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1126
timestamp 1643678851
transform 1 0 10892 0 -1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1127
timestamp 1643678851
transform 1 0 10892 0 1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1128
timestamp 1643678851
transform 1 0 10892 0 -1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1129
timestamp 1643678851
transform 1 0 10892 0 1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1130
timestamp 1643678851
transform 1 0 10892 0 -1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1131
timestamp 1643678851
transform 1 0 10892 0 1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1132
timestamp 1643678851
transform 1 0 10892 0 -1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1133
timestamp 1643678851
transform 1 0 10892 0 1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1134
timestamp 1643678851
transform 1 0 10892 0 -1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1135
timestamp 1643678851
transform 1 0 10892 0 1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1136
timestamp 1643678851
transform 1 0 10892 0 -1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1137
timestamp 1643678851
transform 1 0 10892 0 1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1138
timestamp 1643678851
transform 1 0 10892 0 -1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1139
timestamp 1643678851
transform 1 0 10892 0 1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1140
timestamp 1643678851
transform 1 0 10892 0 -1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1141
timestamp 1643678851
transform 1 0 10892 0 1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1142
timestamp 1643678851
transform 1 0 10892 0 -1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1143
timestamp 1643678851
transform 1 0 10892 0 1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1144
timestamp 1643678851
transform 1 0 10892 0 -1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1145
timestamp 1643678851
transform 1 0 10892 0 1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1146
timestamp 1643678851
transform 1 0 10892 0 -1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1147
timestamp 1643678851
transform 1 0 10892 0 1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1148
timestamp 1643678851
transform 1 0 10892 0 -1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1149
timestamp 1643678851
transform 1 0 10892 0 1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1150
timestamp 1643678851
transform 1 0 10892 0 -1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1151
timestamp 1643678851
transform 1 0 10892 0 1 0
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1152
timestamp 1643678851
transform 1 0 10503 0 -1 24640
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1153
timestamp 1643678851
transform 1 0 10503 0 1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1154
timestamp 1643678851
transform 1 0 10503 0 -1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1155
timestamp 1643678851
transform 1 0 10503 0 1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1156
timestamp 1643678851
transform 1 0 10503 0 -1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1157
timestamp 1643678851
transform 1 0 10503 0 1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1158
timestamp 1643678851
transform 1 0 10503 0 -1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1159
timestamp 1643678851
transform 1 0 10503 0 1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1160
timestamp 1643678851
transform 1 0 10503 0 -1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1161
timestamp 1643678851
transform 1 0 10503 0 1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1162
timestamp 1643678851
transform 1 0 10503 0 -1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1163
timestamp 1643678851
transform 1 0 10503 0 1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1164
timestamp 1643678851
transform 1 0 10503 0 -1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1165
timestamp 1643678851
transform 1 0 10503 0 1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1166
timestamp 1643678851
transform 1 0 10503 0 -1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1167
timestamp 1643678851
transform 1 0 10503 0 1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1168
timestamp 1643678851
transform 1 0 10503 0 -1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1169
timestamp 1643678851
transform 1 0 10503 0 1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1170
timestamp 1643678851
transform 1 0 10503 0 -1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1171
timestamp 1643678851
transform 1 0 10503 0 1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1172
timestamp 1643678851
transform 1 0 10503 0 -1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1173
timestamp 1643678851
transform 1 0 10503 0 1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1174
timestamp 1643678851
transform 1 0 10503 0 -1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1175
timestamp 1643678851
transform 1 0 10503 0 1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1176
timestamp 1643678851
transform 1 0 10503 0 -1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1177
timestamp 1643678851
transform 1 0 10503 0 1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1178
timestamp 1643678851
transform 1 0 10503 0 -1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1179
timestamp 1643678851
transform 1 0 10503 0 1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1180
timestamp 1643678851
transform 1 0 10503 0 -1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1181
timestamp 1643678851
transform 1 0 10503 0 1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1182
timestamp 1643678851
transform 1 0 10503 0 -1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1183
timestamp 1643678851
transform 1 0 10503 0 1 0
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1184
timestamp 1643678851
transform 1 0 10114 0 -1 24640
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1185
timestamp 1643678851
transform 1 0 10114 0 1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1186
timestamp 1643678851
transform 1 0 10114 0 -1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1187
timestamp 1643678851
transform 1 0 10114 0 1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1188
timestamp 1643678851
transform 1 0 10114 0 -1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1189
timestamp 1643678851
transform 1 0 10114 0 1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1190
timestamp 1643678851
transform 1 0 10114 0 -1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1191
timestamp 1643678851
transform 1 0 10114 0 1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1192
timestamp 1643678851
transform 1 0 10114 0 -1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1193
timestamp 1643678851
transform 1 0 10114 0 1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1194
timestamp 1643678851
transform 1 0 10114 0 -1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1195
timestamp 1643678851
transform 1 0 10114 0 1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1196
timestamp 1643678851
transform 1 0 10114 0 -1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1197
timestamp 1643678851
transform 1 0 10114 0 1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1198
timestamp 1643678851
transform 1 0 10114 0 -1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1199
timestamp 1643678851
transform 1 0 10114 0 1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1200
timestamp 1643678851
transform 1 0 10114 0 -1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1201
timestamp 1643678851
transform 1 0 10114 0 1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1202
timestamp 1643678851
transform 1 0 10114 0 -1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1203
timestamp 1643678851
transform 1 0 10114 0 1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1204
timestamp 1643678851
transform 1 0 10114 0 -1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1205
timestamp 1643678851
transform 1 0 10114 0 1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1206
timestamp 1643678851
transform 1 0 10114 0 -1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1207
timestamp 1643678851
transform 1 0 10114 0 1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1208
timestamp 1643678851
transform 1 0 10114 0 -1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1209
timestamp 1643678851
transform 1 0 10114 0 1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1210
timestamp 1643678851
transform 1 0 10114 0 -1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1211
timestamp 1643678851
transform 1 0 10114 0 1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1212
timestamp 1643678851
transform 1 0 10114 0 -1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1213
timestamp 1643678851
transform 1 0 10114 0 1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1214
timestamp 1643678851
transform 1 0 10114 0 -1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1215
timestamp 1643678851
transform 1 0 10114 0 1 0
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1216
timestamp 1643678851
transform 1 0 9725 0 -1 24640
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1217
timestamp 1643678851
transform 1 0 9725 0 1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1218
timestamp 1643678851
transform 1 0 9725 0 -1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1219
timestamp 1643678851
transform 1 0 9725 0 1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1220
timestamp 1643678851
transform 1 0 9725 0 -1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1221
timestamp 1643678851
transform 1 0 9725 0 1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1222
timestamp 1643678851
transform 1 0 9725 0 -1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1223
timestamp 1643678851
transform 1 0 9725 0 1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1224
timestamp 1643678851
transform 1 0 9725 0 -1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1225
timestamp 1643678851
transform 1 0 9725 0 1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1226
timestamp 1643678851
transform 1 0 9725 0 -1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1227
timestamp 1643678851
transform 1 0 9725 0 1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1228
timestamp 1643678851
transform 1 0 9725 0 -1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1229
timestamp 1643678851
transform 1 0 9725 0 1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1230
timestamp 1643678851
transform 1 0 9725 0 -1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1231
timestamp 1643678851
transform 1 0 9725 0 1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1232
timestamp 1643678851
transform 1 0 9725 0 -1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1233
timestamp 1643678851
transform 1 0 9725 0 1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1234
timestamp 1643678851
transform 1 0 9725 0 -1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1235
timestamp 1643678851
transform 1 0 9725 0 1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1236
timestamp 1643678851
transform 1 0 9725 0 -1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1237
timestamp 1643678851
transform 1 0 9725 0 1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1238
timestamp 1643678851
transform 1 0 9725 0 -1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1239
timestamp 1643678851
transform 1 0 9725 0 1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1240
timestamp 1643678851
transform 1 0 9725 0 -1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1241
timestamp 1643678851
transform 1 0 9725 0 1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1242
timestamp 1643678851
transform 1 0 9725 0 -1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1243
timestamp 1643678851
transform 1 0 9725 0 1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1244
timestamp 1643678851
transform 1 0 9725 0 -1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1245
timestamp 1643678851
transform 1 0 9725 0 1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1246
timestamp 1643678851
transform 1 0 9725 0 -1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1247
timestamp 1643678851
transform 1 0 9725 0 1 0
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1248
timestamp 1643678851
transform 1 0 9336 0 -1 24640
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1249
timestamp 1643678851
transform 1 0 9336 0 1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1250
timestamp 1643678851
transform 1 0 9336 0 -1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1251
timestamp 1643678851
transform 1 0 9336 0 1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1252
timestamp 1643678851
transform 1 0 9336 0 -1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1253
timestamp 1643678851
transform 1 0 9336 0 1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1254
timestamp 1643678851
transform 1 0 9336 0 -1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1255
timestamp 1643678851
transform 1 0 9336 0 1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1256
timestamp 1643678851
transform 1 0 9336 0 -1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1257
timestamp 1643678851
transform 1 0 9336 0 1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1258
timestamp 1643678851
transform 1 0 9336 0 -1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1259
timestamp 1643678851
transform 1 0 9336 0 1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1260
timestamp 1643678851
transform 1 0 9336 0 -1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1261
timestamp 1643678851
transform 1 0 9336 0 1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1262
timestamp 1643678851
transform 1 0 9336 0 -1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1263
timestamp 1643678851
transform 1 0 9336 0 1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1264
timestamp 1643678851
transform 1 0 9336 0 -1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1265
timestamp 1643678851
transform 1 0 9336 0 1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1266
timestamp 1643678851
transform 1 0 9336 0 -1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1267
timestamp 1643678851
transform 1 0 9336 0 1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1268
timestamp 1643678851
transform 1 0 9336 0 -1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1269
timestamp 1643678851
transform 1 0 9336 0 1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1270
timestamp 1643678851
transform 1 0 9336 0 -1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1271
timestamp 1643678851
transform 1 0 9336 0 1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1272
timestamp 1643678851
transform 1 0 9336 0 -1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1273
timestamp 1643678851
transform 1 0 9336 0 1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1274
timestamp 1643678851
transform 1 0 9336 0 -1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1275
timestamp 1643678851
transform 1 0 9336 0 1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1276
timestamp 1643678851
transform 1 0 9336 0 -1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1277
timestamp 1643678851
transform 1 0 9336 0 1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1278
timestamp 1643678851
transform 1 0 9336 0 -1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1279
timestamp 1643678851
transform 1 0 9336 0 1 0
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1280
timestamp 1643678851
transform 1 0 8947 0 -1 24640
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1281
timestamp 1643678851
transform 1 0 8947 0 1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1282
timestamp 1643678851
transform 1 0 8947 0 -1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1283
timestamp 1643678851
transform 1 0 8947 0 1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1284
timestamp 1643678851
transform 1 0 8947 0 -1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1285
timestamp 1643678851
transform 1 0 8947 0 1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1286
timestamp 1643678851
transform 1 0 8947 0 -1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1287
timestamp 1643678851
transform 1 0 8947 0 1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1288
timestamp 1643678851
transform 1 0 8947 0 -1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1289
timestamp 1643678851
transform 1 0 8947 0 1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1290
timestamp 1643678851
transform 1 0 8947 0 -1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1291
timestamp 1643678851
transform 1 0 8947 0 1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1292
timestamp 1643678851
transform 1 0 8947 0 -1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1293
timestamp 1643678851
transform 1 0 8947 0 1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1294
timestamp 1643678851
transform 1 0 8947 0 -1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1295
timestamp 1643678851
transform 1 0 8947 0 1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1296
timestamp 1643678851
transform 1 0 8947 0 -1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1297
timestamp 1643678851
transform 1 0 8947 0 1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1298
timestamp 1643678851
transform 1 0 8947 0 -1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1299
timestamp 1643678851
transform 1 0 8947 0 1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1300
timestamp 1643678851
transform 1 0 8947 0 -1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1301
timestamp 1643678851
transform 1 0 8947 0 1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1302
timestamp 1643678851
transform 1 0 8947 0 -1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1303
timestamp 1643678851
transform 1 0 8947 0 1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1304
timestamp 1643678851
transform 1 0 8947 0 -1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1305
timestamp 1643678851
transform 1 0 8947 0 1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1306
timestamp 1643678851
transform 1 0 8947 0 -1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1307
timestamp 1643678851
transform 1 0 8947 0 1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1308
timestamp 1643678851
transform 1 0 8947 0 -1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1309
timestamp 1643678851
transform 1 0 8947 0 1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1310
timestamp 1643678851
transform 1 0 8947 0 -1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1311
timestamp 1643678851
transform 1 0 8947 0 1 0
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1312
timestamp 1643678851
transform 1 0 8558 0 -1 24640
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1313
timestamp 1643678851
transform 1 0 8558 0 1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1314
timestamp 1643678851
transform 1 0 8558 0 -1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1315
timestamp 1643678851
transform 1 0 8558 0 1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1316
timestamp 1643678851
transform 1 0 8558 0 -1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1317
timestamp 1643678851
transform 1 0 8558 0 1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1318
timestamp 1643678851
transform 1 0 8558 0 -1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1319
timestamp 1643678851
transform 1 0 8558 0 1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1320
timestamp 1643678851
transform 1 0 8558 0 -1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1321
timestamp 1643678851
transform 1 0 8558 0 1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1322
timestamp 1643678851
transform 1 0 8558 0 -1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1323
timestamp 1643678851
transform 1 0 8558 0 1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1324
timestamp 1643678851
transform 1 0 8558 0 -1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1325
timestamp 1643678851
transform 1 0 8558 0 1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1326
timestamp 1643678851
transform 1 0 8558 0 -1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1327
timestamp 1643678851
transform 1 0 8558 0 1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1328
timestamp 1643678851
transform 1 0 8558 0 -1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1329
timestamp 1643678851
transform 1 0 8558 0 1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1330
timestamp 1643678851
transform 1 0 8558 0 -1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1331
timestamp 1643678851
transform 1 0 8558 0 1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1332
timestamp 1643678851
transform 1 0 8558 0 -1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1333
timestamp 1643678851
transform 1 0 8558 0 1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1334
timestamp 1643678851
transform 1 0 8558 0 -1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1335
timestamp 1643678851
transform 1 0 8558 0 1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1336
timestamp 1643678851
transform 1 0 8558 0 -1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1337
timestamp 1643678851
transform 1 0 8558 0 1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1338
timestamp 1643678851
transform 1 0 8558 0 -1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1339
timestamp 1643678851
transform 1 0 8558 0 1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1340
timestamp 1643678851
transform 1 0 8558 0 -1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1341
timestamp 1643678851
transform 1 0 8558 0 1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1342
timestamp 1643678851
transform 1 0 8558 0 -1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1343
timestamp 1643678851
transform 1 0 8558 0 1 0
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1344
timestamp 1643678851
transform 1 0 8169 0 -1 24640
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1345
timestamp 1643678851
transform 1 0 8169 0 1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1346
timestamp 1643678851
transform 1 0 8169 0 -1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1347
timestamp 1643678851
transform 1 0 8169 0 1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1348
timestamp 1643678851
transform 1 0 8169 0 -1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1349
timestamp 1643678851
transform 1 0 8169 0 1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1350
timestamp 1643678851
transform 1 0 8169 0 -1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1351
timestamp 1643678851
transform 1 0 8169 0 1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1352
timestamp 1643678851
transform 1 0 8169 0 -1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1353
timestamp 1643678851
transform 1 0 8169 0 1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1354
timestamp 1643678851
transform 1 0 8169 0 -1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1355
timestamp 1643678851
transform 1 0 8169 0 1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1356
timestamp 1643678851
transform 1 0 8169 0 -1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1357
timestamp 1643678851
transform 1 0 8169 0 1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1358
timestamp 1643678851
transform 1 0 8169 0 -1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1359
timestamp 1643678851
transform 1 0 8169 0 1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1360
timestamp 1643678851
transform 1 0 8169 0 -1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1361
timestamp 1643678851
transform 1 0 8169 0 1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1362
timestamp 1643678851
transform 1 0 8169 0 -1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1363
timestamp 1643678851
transform 1 0 8169 0 1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1364
timestamp 1643678851
transform 1 0 8169 0 -1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1365
timestamp 1643678851
transform 1 0 8169 0 1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1366
timestamp 1643678851
transform 1 0 8169 0 -1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1367
timestamp 1643678851
transform 1 0 8169 0 1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1368
timestamp 1643678851
transform 1 0 8169 0 -1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1369
timestamp 1643678851
transform 1 0 8169 0 1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1370
timestamp 1643678851
transform 1 0 8169 0 -1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1371
timestamp 1643678851
transform 1 0 8169 0 1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1372
timestamp 1643678851
transform 1 0 8169 0 -1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1373
timestamp 1643678851
transform 1 0 8169 0 1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1374
timestamp 1643678851
transform 1 0 8169 0 -1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1375
timestamp 1643678851
transform 1 0 8169 0 1 0
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1376
timestamp 1643678851
transform 1 0 7780 0 -1 24640
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1377
timestamp 1643678851
transform 1 0 7780 0 1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1378
timestamp 1643678851
transform 1 0 7780 0 -1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1379
timestamp 1643678851
transform 1 0 7780 0 1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1380
timestamp 1643678851
transform 1 0 7780 0 -1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1381
timestamp 1643678851
transform 1 0 7780 0 1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1382
timestamp 1643678851
transform 1 0 7780 0 -1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1383
timestamp 1643678851
transform 1 0 7780 0 1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1384
timestamp 1643678851
transform 1 0 7780 0 -1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1385
timestamp 1643678851
transform 1 0 7780 0 1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1386
timestamp 1643678851
transform 1 0 7780 0 -1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1387
timestamp 1643678851
transform 1 0 7780 0 1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1388
timestamp 1643678851
transform 1 0 7780 0 -1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1389
timestamp 1643678851
transform 1 0 7780 0 1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1390
timestamp 1643678851
transform 1 0 7780 0 -1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1391
timestamp 1643678851
transform 1 0 7780 0 1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1392
timestamp 1643678851
transform 1 0 7780 0 -1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1393
timestamp 1643678851
transform 1 0 7780 0 1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1394
timestamp 1643678851
transform 1 0 7780 0 -1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1395
timestamp 1643678851
transform 1 0 7780 0 1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1396
timestamp 1643678851
transform 1 0 7780 0 -1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1397
timestamp 1643678851
transform 1 0 7780 0 1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1398
timestamp 1643678851
transform 1 0 7780 0 -1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1399
timestamp 1643678851
transform 1 0 7780 0 1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1400
timestamp 1643678851
transform 1 0 7780 0 -1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1401
timestamp 1643678851
transform 1 0 7780 0 1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1402
timestamp 1643678851
transform 1 0 7780 0 -1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1403
timestamp 1643678851
transform 1 0 7780 0 1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1404
timestamp 1643678851
transform 1 0 7780 0 -1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1405
timestamp 1643678851
transform 1 0 7780 0 1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1406
timestamp 1643678851
transform 1 0 7780 0 -1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1407
timestamp 1643678851
transform 1 0 7780 0 1 0
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1408
timestamp 1643678851
transform 1 0 7391 0 -1 24640
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1409
timestamp 1643678851
transform 1 0 7391 0 1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1410
timestamp 1643678851
transform 1 0 7391 0 -1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1411
timestamp 1643678851
transform 1 0 7391 0 1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1412
timestamp 1643678851
transform 1 0 7391 0 -1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1413
timestamp 1643678851
transform 1 0 7391 0 1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1414
timestamp 1643678851
transform 1 0 7391 0 -1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1415
timestamp 1643678851
transform 1 0 7391 0 1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1416
timestamp 1643678851
transform 1 0 7391 0 -1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1417
timestamp 1643678851
transform 1 0 7391 0 1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1418
timestamp 1643678851
transform 1 0 7391 0 -1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1419
timestamp 1643678851
transform 1 0 7391 0 1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1420
timestamp 1643678851
transform 1 0 7391 0 -1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1421
timestamp 1643678851
transform 1 0 7391 0 1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1422
timestamp 1643678851
transform 1 0 7391 0 -1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1423
timestamp 1643678851
transform 1 0 7391 0 1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1424
timestamp 1643678851
transform 1 0 7391 0 -1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1425
timestamp 1643678851
transform 1 0 7391 0 1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1426
timestamp 1643678851
transform 1 0 7391 0 -1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1427
timestamp 1643678851
transform 1 0 7391 0 1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1428
timestamp 1643678851
transform 1 0 7391 0 -1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1429
timestamp 1643678851
transform 1 0 7391 0 1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1430
timestamp 1643678851
transform 1 0 7391 0 -1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1431
timestamp 1643678851
transform 1 0 7391 0 1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1432
timestamp 1643678851
transform 1 0 7391 0 -1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1433
timestamp 1643678851
transform 1 0 7391 0 1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1434
timestamp 1643678851
transform 1 0 7391 0 -1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1435
timestamp 1643678851
transform 1 0 7391 0 1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1436
timestamp 1643678851
transform 1 0 7391 0 -1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1437
timestamp 1643678851
transform 1 0 7391 0 1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1438
timestamp 1643678851
transform 1 0 7391 0 -1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1439
timestamp 1643678851
transform 1 0 7391 0 1 0
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1440
timestamp 1643678851
transform 1 0 7002 0 -1 24640
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1441
timestamp 1643678851
transform 1 0 7002 0 1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1442
timestamp 1643678851
transform 1 0 7002 0 -1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1443
timestamp 1643678851
transform 1 0 7002 0 1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1444
timestamp 1643678851
transform 1 0 7002 0 -1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1445
timestamp 1643678851
transform 1 0 7002 0 1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1446
timestamp 1643678851
transform 1 0 7002 0 -1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1447
timestamp 1643678851
transform 1 0 7002 0 1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1448
timestamp 1643678851
transform 1 0 7002 0 -1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1449
timestamp 1643678851
transform 1 0 7002 0 1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1450
timestamp 1643678851
transform 1 0 7002 0 -1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1451
timestamp 1643678851
transform 1 0 7002 0 1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1452
timestamp 1643678851
transform 1 0 7002 0 -1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1453
timestamp 1643678851
transform 1 0 7002 0 1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1454
timestamp 1643678851
transform 1 0 7002 0 -1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1455
timestamp 1643678851
transform 1 0 7002 0 1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1456
timestamp 1643678851
transform 1 0 7002 0 -1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1457
timestamp 1643678851
transform 1 0 7002 0 1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1458
timestamp 1643678851
transform 1 0 7002 0 -1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1459
timestamp 1643678851
transform 1 0 7002 0 1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1460
timestamp 1643678851
transform 1 0 7002 0 -1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1461
timestamp 1643678851
transform 1 0 7002 0 1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1462
timestamp 1643678851
transform 1 0 7002 0 -1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1463
timestamp 1643678851
transform 1 0 7002 0 1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1464
timestamp 1643678851
transform 1 0 7002 0 -1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1465
timestamp 1643678851
transform 1 0 7002 0 1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1466
timestamp 1643678851
transform 1 0 7002 0 -1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1467
timestamp 1643678851
transform 1 0 7002 0 1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1468
timestamp 1643678851
transform 1 0 7002 0 -1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1469
timestamp 1643678851
transform 1 0 7002 0 1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1470
timestamp 1643678851
transform 1 0 7002 0 -1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1471
timestamp 1643678851
transform 1 0 7002 0 1 0
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1472
timestamp 1643678851
transform 1 0 6613 0 -1 24640
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1473
timestamp 1643678851
transform 1 0 6613 0 1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1474
timestamp 1643678851
transform 1 0 6613 0 -1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1475
timestamp 1643678851
transform 1 0 6613 0 1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1476
timestamp 1643678851
transform 1 0 6613 0 -1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1477
timestamp 1643678851
transform 1 0 6613 0 1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1478
timestamp 1643678851
transform 1 0 6613 0 -1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1479
timestamp 1643678851
transform 1 0 6613 0 1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1480
timestamp 1643678851
transform 1 0 6613 0 -1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1481
timestamp 1643678851
transform 1 0 6613 0 1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1482
timestamp 1643678851
transform 1 0 6613 0 -1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1483
timestamp 1643678851
transform 1 0 6613 0 1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1484
timestamp 1643678851
transform 1 0 6613 0 -1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1485
timestamp 1643678851
transform 1 0 6613 0 1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1486
timestamp 1643678851
transform 1 0 6613 0 -1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1487
timestamp 1643678851
transform 1 0 6613 0 1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1488
timestamp 1643678851
transform 1 0 6613 0 -1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1489
timestamp 1643678851
transform 1 0 6613 0 1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1490
timestamp 1643678851
transform 1 0 6613 0 -1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1491
timestamp 1643678851
transform 1 0 6613 0 1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1492
timestamp 1643678851
transform 1 0 6613 0 -1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1493
timestamp 1643678851
transform 1 0 6613 0 1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1494
timestamp 1643678851
transform 1 0 6613 0 -1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1495
timestamp 1643678851
transform 1 0 6613 0 1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1496
timestamp 1643678851
transform 1 0 6613 0 -1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1497
timestamp 1643678851
transform 1 0 6613 0 1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1498
timestamp 1643678851
transform 1 0 6613 0 -1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1499
timestamp 1643678851
transform 1 0 6613 0 1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1500
timestamp 1643678851
transform 1 0 6613 0 -1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1501
timestamp 1643678851
transform 1 0 6613 0 1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1502
timestamp 1643678851
transform 1 0 6613 0 -1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1503
timestamp 1643678851
transform 1 0 6613 0 1 0
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1504
timestamp 1643678851
transform 1 0 6224 0 -1 24640
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1505
timestamp 1643678851
transform 1 0 6224 0 1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1506
timestamp 1643678851
transform 1 0 6224 0 -1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1507
timestamp 1643678851
transform 1 0 6224 0 1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1508
timestamp 1643678851
transform 1 0 6224 0 -1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1509
timestamp 1643678851
transform 1 0 6224 0 1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1510
timestamp 1643678851
transform 1 0 6224 0 -1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1511
timestamp 1643678851
transform 1 0 6224 0 1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1512
timestamp 1643678851
transform 1 0 6224 0 -1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1513
timestamp 1643678851
transform 1 0 6224 0 1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1514
timestamp 1643678851
transform 1 0 6224 0 -1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1515
timestamp 1643678851
transform 1 0 6224 0 1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1516
timestamp 1643678851
transform 1 0 6224 0 -1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1517
timestamp 1643678851
transform 1 0 6224 0 1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1518
timestamp 1643678851
transform 1 0 6224 0 -1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1519
timestamp 1643678851
transform 1 0 6224 0 1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1520
timestamp 1643678851
transform 1 0 6224 0 -1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1521
timestamp 1643678851
transform 1 0 6224 0 1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1522
timestamp 1643678851
transform 1 0 6224 0 -1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1523
timestamp 1643678851
transform 1 0 6224 0 1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1524
timestamp 1643678851
transform 1 0 6224 0 -1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1525
timestamp 1643678851
transform 1 0 6224 0 1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1526
timestamp 1643678851
transform 1 0 6224 0 -1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1527
timestamp 1643678851
transform 1 0 6224 0 1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1528
timestamp 1643678851
transform 1 0 6224 0 -1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1529
timestamp 1643678851
transform 1 0 6224 0 1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1530
timestamp 1643678851
transform 1 0 6224 0 -1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1531
timestamp 1643678851
transform 1 0 6224 0 1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1532
timestamp 1643678851
transform 1 0 6224 0 -1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1533
timestamp 1643678851
transform 1 0 6224 0 1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1534
timestamp 1643678851
transform 1 0 6224 0 -1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1535
timestamp 1643678851
transform 1 0 6224 0 1 0
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1536
timestamp 1643678851
transform 1 0 5835 0 -1 24640
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1537
timestamp 1643678851
transform 1 0 5835 0 1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1538
timestamp 1643678851
transform 1 0 5835 0 -1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1539
timestamp 1643678851
transform 1 0 5835 0 1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1540
timestamp 1643678851
transform 1 0 5835 0 -1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1541
timestamp 1643678851
transform 1 0 5835 0 1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1542
timestamp 1643678851
transform 1 0 5835 0 -1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1543
timestamp 1643678851
transform 1 0 5835 0 1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1544
timestamp 1643678851
transform 1 0 5835 0 -1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1545
timestamp 1643678851
transform 1 0 5835 0 1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1546
timestamp 1643678851
transform 1 0 5835 0 -1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1547
timestamp 1643678851
transform 1 0 5835 0 1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1548
timestamp 1643678851
transform 1 0 5835 0 -1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1549
timestamp 1643678851
transform 1 0 5835 0 1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1550
timestamp 1643678851
transform 1 0 5835 0 -1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1551
timestamp 1643678851
transform 1 0 5835 0 1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1552
timestamp 1643678851
transform 1 0 5835 0 -1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1553
timestamp 1643678851
transform 1 0 5835 0 1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1554
timestamp 1643678851
transform 1 0 5835 0 -1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1555
timestamp 1643678851
transform 1 0 5835 0 1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1556
timestamp 1643678851
transform 1 0 5835 0 -1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1557
timestamp 1643678851
transform 1 0 5835 0 1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1558
timestamp 1643678851
transform 1 0 5835 0 -1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1559
timestamp 1643678851
transform 1 0 5835 0 1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1560
timestamp 1643678851
transform 1 0 5835 0 -1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1561
timestamp 1643678851
transform 1 0 5835 0 1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1562
timestamp 1643678851
transform 1 0 5835 0 -1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1563
timestamp 1643678851
transform 1 0 5835 0 1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1564
timestamp 1643678851
transform 1 0 5835 0 -1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1565
timestamp 1643678851
transform 1 0 5835 0 1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1566
timestamp 1643678851
transform 1 0 5835 0 -1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1567
timestamp 1643678851
transform 1 0 5835 0 1 0
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1568
timestamp 1643678851
transform 1 0 5446 0 -1 24640
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1569
timestamp 1643678851
transform 1 0 5446 0 1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1570
timestamp 1643678851
transform 1 0 5446 0 -1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1571
timestamp 1643678851
transform 1 0 5446 0 1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1572
timestamp 1643678851
transform 1 0 5446 0 -1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1573
timestamp 1643678851
transform 1 0 5446 0 1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1574
timestamp 1643678851
transform 1 0 5446 0 -1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1575
timestamp 1643678851
transform 1 0 5446 0 1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1576
timestamp 1643678851
transform 1 0 5446 0 -1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1577
timestamp 1643678851
transform 1 0 5446 0 1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1578
timestamp 1643678851
transform 1 0 5446 0 -1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1579
timestamp 1643678851
transform 1 0 5446 0 1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1580
timestamp 1643678851
transform 1 0 5446 0 -1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1581
timestamp 1643678851
transform 1 0 5446 0 1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1582
timestamp 1643678851
transform 1 0 5446 0 -1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1583
timestamp 1643678851
transform 1 0 5446 0 1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1584
timestamp 1643678851
transform 1 0 5446 0 -1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1585
timestamp 1643678851
transform 1 0 5446 0 1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1586
timestamp 1643678851
transform 1 0 5446 0 -1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1587
timestamp 1643678851
transform 1 0 5446 0 1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1588
timestamp 1643678851
transform 1 0 5446 0 -1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1589
timestamp 1643678851
transform 1 0 5446 0 1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1590
timestamp 1643678851
transform 1 0 5446 0 -1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1591
timestamp 1643678851
transform 1 0 5446 0 1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1592
timestamp 1643678851
transform 1 0 5446 0 -1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1593
timestamp 1643678851
transform 1 0 5446 0 1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1594
timestamp 1643678851
transform 1 0 5446 0 -1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1595
timestamp 1643678851
transform 1 0 5446 0 1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1596
timestamp 1643678851
transform 1 0 5446 0 -1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1597
timestamp 1643678851
transform 1 0 5446 0 1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1598
timestamp 1643678851
transform 1 0 5446 0 -1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1599
timestamp 1643678851
transform 1 0 5446 0 1 0
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1600
timestamp 1643678851
transform 1 0 5057 0 -1 24640
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1601
timestamp 1643678851
transform 1 0 5057 0 1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1602
timestamp 1643678851
transform 1 0 5057 0 -1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1603
timestamp 1643678851
transform 1 0 5057 0 1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1604
timestamp 1643678851
transform 1 0 5057 0 -1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1605
timestamp 1643678851
transform 1 0 5057 0 1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1606
timestamp 1643678851
transform 1 0 5057 0 -1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1607
timestamp 1643678851
transform 1 0 5057 0 1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1608
timestamp 1643678851
transform 1 0 5057 0 -1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1609
timestamp 1643678851
transform 1 0 5057 0 1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1610
timestamp 1643678851
transform 1 0 5057 0 -1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1611
timestamp 1643678851
transform 1 0 5057 0 1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1612
timestamp 1643678851
transform 1 0 5057 0 -1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1613
timestamp 1643678851
transform 1 0 5057 0 1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1614
timestamp 1643678851
transform 1 0 5057 0 -1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1615
timestamp 1643678851
transform 1 0 5057 0 1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1616
timestamp 1643678851
transform 1 0 5057 0 -1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1617
timestamp 1643678851
transform 1 0 5057 0 1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1618
timestamp 1643678851
transform 1 0 5057 0 -1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1619
timestamp 1643678851
transform 1 0 5057 0 1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1620
timestamp 1643678851
transform 1 0 5057 0 -1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1621
timestamp 1643678851
transform 1 0 5057 0 1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1622
timestamp 1643678851
transform 1 0 5057 0 -1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1623
timestamp 1643678851
transform 1 0 5057 0 1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1624
timestamp 1643678851
transform 1 0 5057 0 -1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1625
timestamp 1643678851
transform 1 0 5057 0 1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1626
timestamp 1643678851
transform 1 0 5057 0 -1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1627
timestamp 1643678851
transform 1 0 5057 0 1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1628
timestamp 1643678851
transform 1 0 5057 0 -1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1629
timestamp 1643678851
transform 1 0 5057 0 1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1630
timestamp 1643678851
transform 1 0 5057 0 -1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1631
timestamp 1643678851
transform 1 0 5057 0 1 0
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1632
timestamp 1643678851
transform 1 0 4668 0 -1 24640
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1633
timestamp 1643678851
transform 1 0 4668 0 1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1634
timestamp 1643678851
transform 1 0 4668 0 -1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1635
timestamp 1643678851
transform 1 0 4668 0 1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1636
timestamp 1643678851
transform 1 0 4668 0 -1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1637
timestamp 1643678851
transform 1 0 4668 0 1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1638
timestamp 1643678851
transform 1 0 4668 0 -1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1639
timestamp 1643678851
transform 1 0 4668 0 1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1640
timestamp 1643678851
transform 1 0 4668 0 -1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1641
timestamp 1643678851
transform 1 0 4668 0 1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1642
timestamp 1643678851
transform 1 0 4668 0 -1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1643
timestamp 1643678851
transform 1 0 4668 0 1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1644
timestamp 1643678851
transform 1 0 4668 0 -1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1645
timestamp 1643678851
transform 1 0 4668 0 1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1646
timestamp 1643678851
transform 1 0 4668 0 -1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1647
timestamp 1643678851
transform 1 0 4668 0 1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1648
timestamp 1643678851
transform 1 0 4668 0 -1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1649
timestamp 1643678851
transform 1 0 4668 0 1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1650
timestamp 1643678851
transform 1 0 4668 0 -1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1651
timestamp 1643678851
transform 1 0 4668 0 1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1652
timestamp 1643678851
transform 1 0 4668 0 -1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1653
timestamp 1643678851
transform 1 0 4668 0 1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1654
timestamp 1643678851
transform 1 0 4668 0 -1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1655
timestamp 1643678851
transform 1 0 4668 0 1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1656
timestamp 1643678851
transform 1 0 4668 0 -1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1657
timestamp 1643678851
transform 1 0 4668 0 1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1658
timestamp 1643678851
transform 1 0 4668 0 -1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1659
timestamp 1643678851
transform 1 0 4668 0 1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1660
timestamp 1643678851
transform 1 0 4668 0 -1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1661
timestamp 1643678851
transform 1 0 4668 0 1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1662
timestamp 1643678851
transform 1 0 4668 0 -1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1663
timestamp 1643678851
transform 1 0 4668 0 1 0
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1664
timestamp 1643678851
transform 1 0 4279 0 -1 24640
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1665
timestamp 1643678851
transform 1 0 4279 0 1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1666
timestamp 1643678851
transform 1 0 4279 0 -1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1667
timestamp 1643678851
transform 1 0 4279 0 1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1668
timestamp 1643678851
transform 1 0 4279 0 -1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1669
timestamp 1643678851
transform 1 0 4279 0 1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1670
timestamp 1643678851
transform 1 0 4279 0 -1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1671
timestamp 1643678851
transform 1 0 4279 0 1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1672
timestamp 1643678851
transform 1 0 4279 0 -1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1673
timestamp 1643678851
transform 1 0 4279 0 1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1674
timestamp 1643678851
transform 1 0 4279 0 -1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1675
timestamp 1643678851
transform 1 0 4279 0 1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1676
timestamp 1643678851
transform 1 0 4279 0 -1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1677
timestamp 1643678851
transform 1 0 4279 0 1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1678
timestamp 1643678851
transform 1 0 4279 0 -1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1679
timestamp 1643678851
transform 1 0 4279 0 1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1680
timestamp 1643678851
transform 1 0 4279 0 -1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1681
timestamp 1643678851
transform 1 0 4279 0 1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1682
timestamp 1643678851
transform 1 0 4279 0 -1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1683
timestamp 1643678851
transform 1 0 4279 0 1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1684
timestamp 1643678851
transform 1 0 4279 0 -1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1685
timestamp 1643678851
transform 1 0 4279 0 1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1686
timestamp 1643678851
transform 1 0 4279 0 -1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1687
timestamp 1643678851
transform 1 0 4279 0 1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1688
timestamp 1643678851
transform 1 0 4279 0 -1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1689
timestamp 1643678851
transform 1 0 4279 0 1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1690
timestamp 1643678851
transform 1 0 4279 0 -1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1691
timestamp 1643678851
transform 1 0 4279 0 1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1692
timestamp 1643678851
transform 1 0 4279 0 -1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1693
timestamp 1643678851
transform 1 0 4279 0 1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1694
timestamp 1643678851
transform 1 0 4279 0 -1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1695
timestamp 1643678851
transform 1 0 4279 0 1 0
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1696
timestamp 1643678851
transform 1 0 3890 0 -1 24640
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1697
timestamp 1643678851
transform 1 0 3890 0 1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1698
timestamp 1643678851
transform 1 0 3890 0 -1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1699
timestamp 1643678851
transform 1 0 3890 0 1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1700
timestamp 1643678851
transform 1 0 3890 0 -1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1701
timestamp 1643678851
transform 1 0 3890 0 1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1702
timestamp 1643678851
transform 1 0 3890 0 -1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1703
timestamp 1643678851
transform 1 0 3890 0 1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1704
timestamp 1643678851
transform 1 0 3890 0 -1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1705
timestamp 1643678851
transform 1 0 3890 0 1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1706
timestamp 1643678851
transform 1 0 3890 0 -1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1707
timestamp 1643678851
transform 1 0 3890 0 1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1708
timestamp 1643678851
transform 1 0 3890 0 -1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1709
timestamp 1643678851
transform 1 0 3890 0 1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1710
timestamp 1643678851
transform 1 0 3890 0 -1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1711
timestamp 1643678851
transform 1 0 3890 0 1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1712
timestamp 1643678851
transform 1 0 3890 0 -1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1713
timestamp 1643678851
transform 1 0 3890 0 1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1714
timestamp 1643678851
transform 1 0 3890 0 -1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1715
timestamp 1643678851
transform 1 0 3890 0 1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1716
timestamp 1643678851
transform 1 0 3890 0 -1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1717
timestamp 1643678851
transform 1 0 3890 0 1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1718
timestamp 1643678851
transform 1 0 3890 0 -1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1719
timestamp 1643678851
transform 1 0 3890 0 1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1720
timestamp 1643678851
transform 1 0 3890 0 -1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1721
timestamp 1643678851
transform 1 0 3890 0 1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1722
timestamp 1643678851
transform 1 0 3890 0 -1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1723
timestamp 1643678851
transform 1 0 3890 0 1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1724
timestamp 1643678851
transform 1 0 3890 0 -1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1725
timestamp 1643678851
transform 1 0 3890 0 1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1726
timestamp 1643678851
transform 1 0 3890 0 -1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1727
timestamp 1643678851
transform 1 0 3890 0 1 0
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1728
timestamp 1643678851
transform 1 0 3501 0 -1 24640
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1729
timestamp 1643678851
transform 1 0 3501 0 1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1730
timestamp 1643678851
transform 1 0 3501 0 -1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1731
timestamp 1643678851
transform 1 0 3501 0 1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1732
timestamp 1643678851
transform 1 0 3501 0 -1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1733
timestamp 1643678851
transform 1 0 3501 0 1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1734
timestamp 1643678851
transform 1 0 3501 0 -1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1735
timestamp 1643678851
transform 1 0 3501 0 1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1736
timestamp 1643678851
transform 1 0 3501 0 -1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1737
timestamp 1643678851
transform 1 0 3501 0 1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1738
timestamp 1643678851
transform 1 0 3501 0 -1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1739
timestamp 1643678851
transform 1 0 3501 0 1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1740
timestamp 1643678851
transform 1 0 3501 0 -1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1741
timestamp 1643678851
transform 1 0 3501 0 1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1742
timestamp 1643678851
transform 1 0 3501 0 -1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1743
timestamp 1643678851
transform 1 0 3501 0 1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1744
timestamp 1643678851
transform 1 0 3501 0 -1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1745
timestamp 1643678851
transform 1 0 3501 0 1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1746
timestamp 1643678851
transform 1 0 3501 0 -1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1747
timestamp 1643678851
transform 1 0 3501 0 1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1748
timestamp 1643678851
transform 1 0 3501 0 -1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1749
timestamp 1643678851
transform 1 0 3501 0 1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1750
timestamp 1643678851
transform 1 0 3501 0 -1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1751
timestamp 1643678851
transform 1 0 3501 0 1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1752
timestamp 1643678851
transform 1 0 3501 0 -1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1753
timestamp 1643678851
transform 1 0 3501 0 1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1754
timestamp 1643678851
transform 1 0 3501 0 -1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1755
timestamp 1643678851
transform 1 0 3501 0 1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1756
timestamp 1643678851
transform 1 0 3501 0 -1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1757
timestamp 1643678851
transform 1 0 3501 0 1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1758
timestamp 1643678851
transform 1 0 3501 0 -1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1759
timestamp 1643678851
transform 1 0 3501 0 1 0
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1760
timestamp 1643678851
transform 1 0 3112 0 -1 24640
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1761
timestamp 1643678851
transform 1 0 3112 0 1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1762
timestamp 1643678851
transform 1 0 3112 0 -1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1763
timestamp 1643678851
transform 1 0 3112 0 1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1764
timestamp 1643678851
transform 1 0 3112 0 -1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1765
timestamp 1643678851
transform 1 0 3112 0 1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1766
timestamp 1643678851
transform 1 0 3112 0 -1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1767
timestamp 1643678851
transform 1 0 3112 0 1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1768
timestamp 1643678851
transform 1 0 3112 0 -1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1769
timestamp 1643678851
transform 1 0 3112 0 1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1770
timestamp 1643678851
transform 1 0 3112 0 -1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1771
timestamp 1643678851
transform 1 0 3112 0 1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1772
timestamp 1643678851
transform 1 0 3112 0 -1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1773
timestamp 1643678851
transform 1 0 3112 0 1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1774
timestamp 1643678851
transform 1 0 3112 0 -1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1775
timestamp 1643678851
transform 1 0 3112 0 1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1776
timestamp 1643678851
transform 1 0 3112 0 -1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1777
timestamp 1643678851
transform 1 0 3112 0 1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1778
timestamp 1643678851
transform 1 0 3112 0 -1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1779
timestamp 1643678851
transform 1 0 3112 0 1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1780
timestamp 1643678851
transform 1 0 3112 0 -1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1781
timestamp 1643678851
transform 1 0 3112 0 1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1782
timestamp 1643678851
transform 1 0 3112 0 -1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1783
timestamp 1643678851
transform 1 0 3112 0 1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1784
timestamp 1643678851
transform 1 0 3112 0 -1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1785
timestamp 1643678851
transform 1 0 3112 0 1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1786
timestamp 1643678851
transform 1 0 3112 0 -1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1787
timestamp 1643678851
transform 1 0 3112 0 1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1788
timestamp 1643678851
transform 1 0 3112 0 -1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1789
timestamp 1643678851
transform 1 0 3112 0 1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1790
timestamp 1643678851
transform 1 0 3112 0 -1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1791
timestamp 1643678851
transform 1 0 3112 0 1 0
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1792
timestamp 1643678851
transform 1 0 2723 0 -1 24640
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1793
timestamp 1643678851
transform 1 0 2723 0 1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1794
timestamp 1643678851
transform 1 0 2723 0 -1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1795
timestamp 1643678851
transform 1 0 2723 0 1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1796
timestamp 1643678851
transform 1 0 2723 0 -1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1797
timestamp 1643678851
transform 1 0 2723 0 1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1798
timestamp 1643678851
transform 1 0 2723 0 -1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1799
timestamp 1643678851
transform 1 0 2723 0 1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1800
timestamp 1643678851
transform 1 0 2723 0 -1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1801
timestamp 1643678851
transform 1 0 2723 0 1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1802
timestamp 1643678851
transform 1 0 2723 0 -1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1803
timestamp 1643678851
transform 1 0 2723 0 1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1804
timestamp 1643678851
transform 1 0 2723 0 -1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1805
timestamp 1643678851
transform 1 0 2723 0 1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1806
timestamp 1643678851
transform 1 0 2723 0 -1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1807
timestamp 1643678851
transform 1 0 2723 0 1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1808
timestamp 1643678851
transform 1 0 2723 0 -1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1809
timestamp 1643678851
transform 1 0 2723 0 1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1810
timestamp 1643678851
transform 1 0 2723 0 -1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1811
timestamp 1643678851
transform 1 0 2723 0 1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1812
timestamp 1643678851
transform 1 0 2723 0 -1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1813
timestamp 1643678851
transform 1 0 2723 0 1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1814
timestamp 1643678851
transform 1 0 2723 0 -1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1815
timestamp 1643678851
transform 1 0 2723 0 1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1816
timestamp 1643678851
transform 1 0 2723 0 -1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1817
timestamp 1643678851
transform 1 0 2723 0 1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1818
timestamp 1643678851
transform 1 0 2723 0 -1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1819
timestamp 1643678851
transform 1 0 2723 0 1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1820
timestamp 1643678851
transform 1 0 2723 0 -1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1821
timestamp 1643678851
transform 1 0 2723 0 1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1822
timestamp 1643678851
transform 1 0 2723 0 -1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1823
timestamp 1643678851
transform 1 0 2723 0 1 0
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1824
timestamp 1643678851
transform 1 0 2334 0 -1 24640
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1825
timestamp 1643678851
transform 1 0 2334 0 1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1826
timestamp 1643678851
transform 1 0 2334 0 -1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1827
timestamp 1643678851
transform 1 0 2334 0 1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1828
timestamp 1643678851
transform 1 0 2334 0 -1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1829
timestamp 1643678851
transform 1 0 2334 0 1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1830
timestamp 1643678851
transform 1 0 2334 0 -1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1831
timestamp 1643678851
transform 1 0 2334 0 1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1832
timestamp 1643678851
transform 1 0 2334 0 -1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1833
timestamp 1643678851
transform 1 0 2334 0 1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1834
timestamp 1643678851
transform 1 0 2334 0 -1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1835
timestamp 1643678851
transform 1 0 2334 0 1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1836
timestamp 1643678851
transform 1 0 2334 0 -1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1837
timestamp 1643678851
transform 1 0 2334 0 1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1838
timestamp 1643678851
transform 1 0 2334 0 -1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1839
timestamp 1643678851
transform 1 0 2334 0 1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1840
timestamp 1643678851
transform 1 0 2334 0 -1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1841
timestamp 1643678851
transform 1 0 2334 0 1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1842
timestamp 1643678851
transform 1 0 2334 0 -1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1843
timestamp 1643678851
transform 1 0 2334 0 1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1844
timestamp 1643678851
transform 1 0 2334 0 -1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1845
timestamp 1643678851
transform 1 0 2334 0 1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1846
timestamp 1643678851
transform 1 0 2334 0 -1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1847
timestamp 1643678851
transform 1 0 2334 0 1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1848
timestamp 1643678851
transform 1 0 2334 0 -1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1849
timestamp 1643678851
transform 1 0 2334 0 1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1850
timestamp 1643678851
transform 1 0 2334 0 -1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1851
timestamp 1643678851
transform 1 0 2334 0 1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1852
timestamp 1643678851
transform 1 0 2334 0 -1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1853
timestamp 1643678851
transform 1 0 2334 0 1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1854
timestamp 1643678851
transform 1 0 2334 0 -1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1855
timestamp 1643678851
transform 1 0 2334 0 1 0
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1856
timestamp 1643678851
transform 1 0 1945 0 -1 24640
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1857
timestamp 1643678851
transform 1 0 1945 0 1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1858
timestamp 1643678851
transform 1 0 1945 0 -1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1859
timestamp 1643678851
transform 1 0 1945 0 1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1860
timestamp 1643678851
transform 1 0 1945 0 -1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1861
timestamp 1643678851
transform 1 0 1945 0 1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1862
timestamp 1643678851
transform 1 0 1945 0 -1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1863
timestamp 1643678851
transform 1 0 1945 0 1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1864
timestamp 1643678851
transform 1 0 1945 0 -1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1865
timestamp 1643678851
transform 1 0 1945 0 1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1866
timestamp 1643678851
transform 1 0 1945 0 -1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1867
timestamp 1643678851
transform 1 0 1945 0 1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1868
timestamp 1643678851
transform 1 0 1945 0 -1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1869
timestamp 1643678851
transform 1 0 1945 0 1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1870
timestamp 1643678851
transform 1 0 1945 0 -1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1871
timestamp 1643678851
transform 1 0 1945 0 1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1872
timestamp 1643678851
transform 1 0 1945 0 -1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1873
timestamp 1643678851
transform 1 0 1945 0 1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1874
timestamp 1643678851
transform 1 0 1945 0 -1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1875
timestamp 1643678851
transform 1 0 1945 0 1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1876
timestamp 1643678851
transform 1 0 1945 0 -1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1877
timestamp 1643678851
transform 1 0 1945 0 1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1878
timestamp 1643678851
transform 1 0 1945 0 -1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1879
timestamp 1643678851
transform 1 0 1945 0 1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1880
timestamp 1643678851
transform 1 0 1945 0 -1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1881
timestamp 1643678851
transform 1 0 1945 0 1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1882
timestamp 1643678851
transform 1 0 1945 0 -1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1883
timestamp 1643678851
transform 1 0 1945 0 1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1884
timestamp 1643678851
transform 1 0 1945 0 -1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1885
timestamp 1643678851
transform 1 0 1945 0 1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1886
timestamp 1643678851
transform 1 0 1945 0 -1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1887
timestamp 1643678851
transform 1 0 1945 0 1 0
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1888
timestamp 1643678851
transform 1 0 1556 0 -1 24640
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1889
timestamp 1643678851
transform 1 0 1556 0 1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1890
timestamp 1643678851
transform 1 0 1556 0 -1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1891
timestamp 1643678851
transform 1 0 1556 0 1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1892
timestamp 1643678851
transform 1 0 1556 0 -1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1893
timestamp 1643678851
transform 1 0 1556 0 1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1894
timestamp 1643678851
transform 1 0 1556 0 -1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1895
timestamp 1643678851
transform 1 0 1556 0 1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1896
timestamp 1643678851
transform 1 0 1556 0 -1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1897
timestamp 1643678851
transform 1 0 1556 0 1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1898
timestamp 1643678851
transform 1 0 1556 0 -1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1899
timestamp 1643678851
transform 1 0 1556 0 1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1900
timestamp 1643678851
transform 1 0 1556 0 -1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1901
timestamp 1643678851
transform 1 0 1556 0 1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1902
timestamp 1643678851
transform 1 0 1556 0 -1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1903
timestamp 1643678851
transform 1 0 1556 0 1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1904
timestamp 1643678851
transform 1 0 1556 0 -1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1905
timestamp 1643678851
transform 1 0 1556 0 1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1906
timestamp 1643678851
transform 1 0 1556 0 -1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1907
timestamp 1643678851
transform 1 0 1556 0 1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1908
timestamp 1643678851
transform 1 0 1556 0 -1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1909
timestamp 1643678851
transform 1 0 1556 0 1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1910
timestamp 1643678851
transform 1 0 1556 0 -1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1911
timestamp 1643678851
transform 1 0 1556 0 1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1912
timestamp 1643678851
transform 1 0 1556 0 -1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1913
timestamp 1643678851
transform 1 0 1556 0 1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1914
timestamp 1643678851
transform 1 0 1556 0 -1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1915
timestamp 1643678851
transform 1 0 1556 0 1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1916
timestamp 1643678851
transform 1 0 1556 0 -1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1917
timestamp 1643678851
transform 1 0 1556 0 1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1918
timestamp 1643678851
transform 1 0 1556 0 -1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1919
timestamp 1643678851
transform 1 0 1556 0 1 0
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1920
timestamp 1643678851
transform 1 0 1167 0 -1 24640
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1921
timestamp 1643678851
transform 1 0 1167 0 1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1922
timestamp 1643678851
transform 1 0 1167 0 -1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1923
timestamp 1643678851
transform 1 0 1167 0 1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1924
timestamp 1643678851
transform 1 0 1167 0 -1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1925
timestamp 1643678851
transform 1 0 1167 0 1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1926
timestamp 1643678851
transform 1 0 1167 0 -1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1927
timestamp 1643678851
transform 1 0 1167 0 1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1928
timestamp 1643678851
transform 1 0 1167 0 -1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1929
timestamp 1643678851
transform 1 0 1167 0 1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1930
timestamp 1643678851
transform 1 0 1167 0 -1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1931
timestamp 1643678851
transform 1 0 1167 0 1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1932
timestamp 1643678851
transform 1 0 1167 0 -1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1933
timestamp 1643678851
transform 1 0 1167 0 1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1934
timestamp 1643678851
transform 1 0 1167 0 -1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1935
timestamp 1643678851
transform 1 0 1167 0 1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1936
timestamp 1643678851
transform 1 0 1167 0 -1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1937
timestamp 1643678851
transform 1 0 1167 0 1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1938
timestamp 1643678851
transform 1 0 1167 0 -1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1939
timestamp 1643678851
transform 1 0 1167 0 1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1940
timestamp 1643678851
transform 1 0 1167 0 -1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1941
timestamp 1643678851
transform 1 0 1167 0 1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1942
timestamp 1643678851
transform 1 0 1167 0 -1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1943
timestamp 1643678851
transform 1 0 1167 0 1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1944
timestamp 1643678851
transform 1 0 1167 0 -1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1945
timestamp 1643678851
transform 1 0 1167 0 1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1946
timestamp 1643678851
transform 1 0 1167 0 -1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1947
timestamp 1643678851
transform 1 0 1167 0 1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1948
timestamp 1643678851
transform 1 0 1167 0 -1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1949
timestamp 1643678851
transform 1 0 1167 0 1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1950
timestamp 1643678851
transform 1 0 1167 0 -1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1951
timestamp 1643678851
transform 1 0 1167 0 1 0
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1952
timestamp 1643678851
transform 1 0 778 0 -1 24640
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1953
timestamp 1643678851
transform 1 0 778 0 1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1954
timestamp 1643678851
transform 1 0 778 0 -1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1955
timestamp 1643678851
transform 1 0 778 0 1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1956
timestamp 1643678851
transform 1 0 778 0 -1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1957
timestamp 1643678851
transform 1 0 778 0 1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1958
timestamp 1643678851
transform 1 0 778 0 -1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1959
timestamp 1643678851
transform 1 0 778 0 1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1960
timestamp 1643678851
transform 1 0 778 0 -1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1961
timestamp 1643678851
transform 1 0 778 0 1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1962
timestamp 1643678851
transform 1 0 778 0 -1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1963
timestamp 1643678851
transform 1 0 778 0 1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1964
timestamp 1643678851
transform 1 0 778 0 -1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1965
timestamp 1643678851
transform 1 0 778 0 1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1966
timestamp 1643678851
transform 1 0 778 0 -1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1967
timestamp 1643678851
transform 1 0 778 0 1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1968
timestamp 1643678851
transform 1 0 778 0 -1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1969
timestamp 1643678851
transform 1 0 778 0 1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1970
timestamp 1643678851
transform 1 0 778 0 -1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1971
timestamp 1643678851
transform 1 0 778 0 1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1972
timestamp 1643678851
transform 1 0 778 0 -1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1973
timestamp 1643678851
transform 1 0 778 0 1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1974
timestamp 1643678851
transform 1 0 778 0 -1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1975
timestamp 1643678851
transform 1 0 778 0 1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1976
timestamp 1643678851
transform 1 0 778 0 -1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1977
timestamp 1643678851
transform 1 0 778 0 1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1978
timestamp 1643678851
transform 1 0 778 0 -1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1979
timestamp 1643678851
transform 1 0 778 0 1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1980
timestamp 1643678851
transform 1 0 778 0 -1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1981
timestamp 1643678851
transform 1 0 778 0 1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1982
timestamp 1643678851
transform 1 0 778 0 -1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1983
timestamp 1643678851
transform 1 0 778 0 1 0
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1984
timestamp 1643678851
transform 1 0 389 0 -1 24640
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1985
timestamp 1643678851
transform 1 0 389 0 1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1986
timestamp 1643678851
transform 1 0 389 0 -1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1987
timestamp 1643678851
transform 1 0 389 0 1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1988
timestamp 1643678851
transform 1 0 389 0 -1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1989
timestamp 1643678851
transform 1 0 389 0 1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1990
timestamp 1643678851
transform 1 0 389 0 -1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1991
timestamp 1643678851
transform 1 0 389 0 1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1992
timestamp 1643678851
transform 1 0 389 0 -1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1993
timestamp 1643678851
transform 1 0 389 0 1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1994
timestamp 1643678851
transform 1 0 389 0 -1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1995
timestamp 1643678851
transform 1 0 389 0 1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1996
timestamp 1643678851
transform 1 0 389 0 -1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1997
timestamp 1643678851
transform 1 0 389 0 1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1998
timestamp 1643678851
transform 1 0 389 0 -1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_1999
timestamp 1643678851
transform 1 0 389 0 1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_2000
timestamp 1643678851
transform 1 0 389 0 -1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_2001
timestamp 1643678851
transform 1 0 389 0 1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_2002
timestamp 1643678851
transform 1 0 389 0 -1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_2003
timestamp 1643678851
transform 1 0 389 0 1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_2004
timestamp 1643678851
transform 1 0 389 0 -1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_2005
timestamp 1643678851
transform 1 0 389 0 1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_2006
timestamp 1643678851
transform 1 0 389 0 -1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_2007
timestamp 1643678851
transform 1 0 389 0 1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_2008
timestamp 1643678851
transform 1 0 389 0 -1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_2009
timestamp 1643678851
transform 1 0 389 0 1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_2010
timestamp 1643678851
transform 1 0 389 0 -1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_2011
timestamp 1643678851
transform 1 0 389 0 1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_2012
timestamp 1643678851
transform 1 0 389 0 -1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_2013
timestamp 1643678851
transform 1 0 389 0 1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_2014
timestamp 1643678851
transform 1 0 389 0 -1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_2015
timestamp 1643678851
transform 1 0 389 0 1 0
box 0 -21 389 808
use cell_2r1w  cell_2r1w_2016
timestamp 1643678851
transform 1 0 0 0 -1 24640
box 0 -21 389 808
use cell_2r1w  cell_2r1w_2017
timestamp 1643678851
transform 1 0 0 0 1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_2018
timestamp 1643678851
transform 1 0 0 0 -1 23100
box 0 -21 389 808
use cell_2r1w  cell_2r1w_2019
timestamp 1643678851
transform 1 0 0 0 1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_2020
timestamp 1643678851
transform 1 0 0 0 -1 21560
box 0 -21 389 808
use cell_2r1w  cell_2r1w_2021
timestamp 1643678851
transform 1 0 0 0 1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_2022
timestamp 1643678851
transform 1 0 0 0 -1 20020
box 0 -21 389 808
use cell_2r1w  cell_2r1w_2023
timestamp 1643678851
transform 1 0 0 0 1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_2024
timestamp 1643678851
transform 1 0 0 0 -1 18480
box 0 -21 389 808
use cell_2r1w  cell_2r1w_2025
timestamp 1643678851
transform 1 0 0 0 1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_2026
timestamp 1643678851
transform 1 0 0 0 -1 16940
box 0 -21 389 808
use cell_2r1w  cell_2r1w_2027
timestamp 1643678851
transform 1 0 0 0 1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_2028
timestamp 1643678851
transform 1 0 0 0 -1 15400
box 0 -21 389 808
use cell_2r1w  cell_2r1w_2029
timestamp 1643678851
transform 1 0 0 0 1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_2030
timestamp 1643678851
transform 1 0 0 0 -1 13860
box 0 -21 389 808
use cell_2r1w  cell_2r1w_2031
timestamp 1643678851
transform 1 0 0 0 1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_2032
timestamp 1643678851
transform 1 0 0 0 -1 12320
box 0 -21 389 808
use cell_2r1w  cell_2r1w_2033
timestamp 1643678851
transform 1 0 0 0 1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_2034
timestamp 1643678851
transform 1 0 0 0 -1 10780
box 0 -21 389 808
use cell_2r1w  cell_2r1w_2035
timestamp 1643678851
transform 1 0 0 0 1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_2036
timestamp 1643678851
transform 1 0 0 0 -1 9240
box 0 -21 389 808
use cell_2r1w  cell_2r1w_2037
timestamp 1643678851
transform 1 0 0 0 1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_2038
timestamp 1643678851
transform 1 0 0 0 -1 7700
box 0 -21 389 808
use cell_2r1w  cell_2r1w_2039
timestamp 1643678851
transform 1 0 0 0 1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_2040
timestamp 1643678851
transform 1 0 0 0 -1 6160
box 0 -21 389 808
use cell_2r1w  cell_2r1w_2041
timestamp 1643678851
transform 1 0 0 0 1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_2042
timestamp 1643678851
transform 1 0 0 0 -1 4620
box 0 -21 389 808
use cell_2r1w  cell_2r1w_2043
timestamp 1643678851
transform 1 0 0 0 1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_2044
timestamp 1643678851
transform 1 0 0 0 -1 3080
box 0 -21 389 808
use cell_2r1w  cell_2r1w_2045
timestamp 1643678851
transform 1 0 0 0 1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_2046
timestamp 1643678851
transform 1 0 0 0 -1 1540
box 0 -21 389 808
use cell_2r1w  cell_2r1w_2047
timestamp 1643678851
transform 1 0 0 0 1 0
box 0 -21 389 808
<< labels >>
rlabel metal2 s 96 0 110 24640 4 read_bl_0_0
rlabel metal2 s 222 0 236 24640 4 read_bl_1_0
rlabel metal2 s 313 0 327 24640 4 write_bl_0_0
rlabel metal2 s 485 0 499 24640 4 read_bl_0_1
rlabel metal2 s 611 0 625 24640 4 read_bl_1_1
rlabel metal2 s 702 0 716 24640 4 write_bl_0_1
rlabel metal2 s 874 0 888 24640 4 read_bl_0_2
rlabel metal2 s 1000 0 1014 24640 4 read_bl_1_2
rlabel metal2 s 1091 0 1105 24640 4 write_bl_0_2
rlabel metal2 s 1263 0 1277 24640 4 read_bl_0_3
rlabel metal2 s 1389 0 1403 24640 4 read_bl_1_3
rlabel metal2 s 1480 0 1494 24640 4 write_bl_0_3
rlabel metal2 s 1652 0 1666 24640 4 read_bl_0_4
rlabel metal2 s 1778 0 1792 24640 4 read_bl_1_4
rlabel metal2 s 1869 0 1883 24640 4 write_bl_0_4
rlabel metal2 s 2041 0 2055 24640 4 read_bl_0_5
rlabel metal2 s 2167 0 2181 24640 4 read_bl_1_5
rlabel metal2 s 2258 0 2272 24640 4 write_bl_0_5
rlabel metal2 s 2430 0 2444 24640 4 read_bl_0_6
rlabel metal2 s 2556 0 2570 24640 4 read_bl_1_6
rlabel metal2 s 2647 0 2661 24640 4 write_bl_0_6
rlabel metal2 s 2819 0 2833 24640 4 read_bl_0_7
rlabel metal2 s 2945 0 2959 24640 4 read_bl_1_7
rlabel metal2 s 3036 0 3050 24640 4 write_bl_0_7
rlabel metal2 s 3208 0 3222 24640 4 read_bl_0_8
rlabel metal2 s 3334 0 3348 24640 4 read_bl_1_8
rlabel metal2 s 3425 0 3439 24640 4 write_bl_0_8
rlabel metal2 s 3597 0 3611 24640 4 read_bl_0_9
rlabel metal2 s 3723 0 3737 24640 4 read_bl_1_9
rlabel metal2 s 3814 0 3828 24640 4 write_bl_0_9
rlabel metal2 s 3986 0 4000 24640 4 read_bl_0_10
rlabel metal2 s 4112 0 4126 24640 4 read_bl_1_10
rlabel metal2 s 4203 0 4217 24640 4 write_bl_0_10
rlabel metal2 s 4375 0 4389 24640 4 read_bl_0_11
rlabel metal2 s 4501 0 4515 24640 4 read_bl_1_11
rlabel metal2 s 4592 0 4606 24640 4 write_bl_0_11
rlabel metal2 s 4764 0 4778 24640 4 read_bl_0_12
rlabel metal2 s 4890 0 4904 24640 4 read_bl_1_12
rlabel metal2 s 4981 0 4995 24640 4 write_bl_0_12
rlabel metal2 s 5153 0 5167 24640 4 read_bl_0_13
rlabel metal2 s 5279 0 5293 24640 4 read_bl_1_13
rlabel metal2 s 5370 0 5384 24640 4 write_bl_0_13
rlabel metal2 s 5542 0 5556 24640 4 read_bl_0_14
rlabel metal2 s 5668 0 5682 24640 4 read_bl_1_14
rlabel metal2 s 5759 0 5773 24640 4 write_bl_0_14
rlabel metal2 s 5931 0 5945 24640 4 read_bl_0_15
rlabel metal2 s 6057 0 6071 24640 4 read_bl_1_15
rlabel metal2 s 6148 0 6162 24640 4 write_bl_0_15
rlabel metal2 s 6320 0 6334 24640 4 read_bl_0_16
rlabel metal2 s 6446 0 6460 24640 4 read_bl_1_16
rlabel metal2 s 6537 0 6551 24640 4 write_bl_0_16
rlabel metal2 s 6709 0 6723 24640 4 read_bl_0_17
rlabel metal2 s 6835 0 6849 24640 4 read_bl_1_17
rlabel metal2 s 6926 0 6940 24640 4 write_bl_0_17
rlabel metal2 s 7098 0 7112 24640 4 read_bl_0_18
rlabel metal2 s 7224 0 7238 24640 4 read_bl_1_18
rlabel metal2 s 7315 0 7329 24640 4 write_bl_0_18
rlabel metal2 s 7487 0 7501 24640 4 read_bl_0_19
rlabel metal2 s 7613 0 7627 24640 4 read_bl_1_19
rlabel metal2 s 7704 0 7718 24640 4 write_bl_0_19
rlabel metal2 s 7876 0 7890 24640 4 read_bl_0_20
rlabel metal2 s 8002 0 8016 24640 4 read_bl_1_20
rlabel metal2 s 8093 0 8107 24640 4 write_bl_0_20
rlabel metal2 s 8265 0 8279 24640 4 read_bl_0_21
rlabel metal2 s 8391 0 8405 24640 4 read_bl_1_21
rlabel metal2 s 8482 0 8496 24640 4 write_bl_0_21
rlabel metal2 s 8654 0 8668 24640 4 read_bl_0_22
rlabel metal2 s 8780 0 8794 24640 4 read_bl_1_22
rlabel metal2 s 8871 0 8885 24640 4 write_bl_0_22
rlabel metal2 s 9043 0 9057 24640 4 read_bl_0_23
rlabel metal2 s 9169 0 9183 24640 4 read_bl_1_23
rlabel metal2 s 9260 0 9274 24640 4 write_bl_0_23
rlabel metal2 s 9432 0 9446 24640 4 read_bl_0_24
rlabel metal2 s 9558 0 9572 24640 4 read_bl_1_24
rlabel metal2 s 9649 0 9663 24640 4 write_bl_0_24
rlabel metal2 s 9821 0 9835 24640 4 read_bl_0_25
rlabel metal2 s 9947 0 9961 24640 4 read_bl_1_25
rlabel metal2 s 10038 0 10052 24640 4 write_bl_0_25
rlabel metal2 s 10210 0 10224 24640 4 read_bl_0_26
rlabel metal2 s 10336 0 10350 24640 4 read_bl_1_26
rlabel metal2 s 10427 0 10441 24640 4 write_bl_0_26
rlabel metal2 s 10599 0 10613 24640 4 read_bl_0_27
rlabel metal2 s 10725 0 10739 24640 4 read_bl_1_27
rlabel metal2 s 10816 0 10830 24640 4 write_bl_0_27
rlabel metal2 s 10988 0 11002 24640 4 read_bl_0_28
rlabel metal2 s 11114 0 11128 24640 4 read_bl_1_28
rlabel metal2 s 11205 0 11219 24640 4 write_bl_0_28
rlabel metal2 s 11377 0 11391 24640 4 read_bl_0_29
rlabel metal2 s 11503 0 11517 24640 4 read_bl_1_29
rlabel metal2 s 11594 0 11608 24640 4 write_bl_0_29
rlabel metal2 s 11766 0 11780 24640 4 read_bl_0_30
rlabel metal2 s 11892 0 11906 24640 4 read_bl_1_30
rlabel metal2 s 11983 0 11997 24640 4 write_bl_0_30
rlabel metal2 s 12155 0 12169 24640 4 read_bl_0_31
rlabel metal2 s 12281 0 12295 24640 4 read_bl_1_31
rlabel metal2 s 12372 0 12386 24640 4 write_bl_0_31
rlabel metal2 s 12544 0 12558 24640 4 read_bl_0_32
rlabel metal2 s 12670 0 12684 24640 4 read_bl_1_32
rlabel metal2 s 12761 0 12775 24640 4 write_bl_0_32
rlabel metal2 s 12933 0 12947 24640 4 read_bl_0_33
rlabel metal2 s 13059 0 13073 24640 4 read_bl_1_33
rlabel metal2 s 13150 0 13164 24640 4 write_bl_0_33
rlabel metal2 s 13322 0 13336 24640 4 read_bl_0_34
rlabel metal2 s 13448 0 13462 24640 4 read_bl_1_34
rlabel metal2 s 13539 0 13553 24640 4 write_bl_0_34
rlabel metal2 s 13711 0 13725 24640 4 read_bl_0_35
rlabel metal2 s 13837 0 13851 24640 4 read_bl_1_35
rlabel metal2 s 13928 0 13942 24640 4 write_bl_0_35
rlabel metal2 s 14100 0 14114 24640 4 read_bl_0_36
rlabel metal2 s 14226 0 14240 24640 4 read_bl_1_36
rlabel metal2 s 14317 0 14331 24640 4 write_bl_0_36
rlabel metal2 s 14489 0 14503 24640 4 read_bl_0_37
rlabel metal2 s 14615 0 14629 24640 4 read_bl_1_37
rlabel metal2 s 14706 0 14720 24640 4 write_bl_0_37
rlabel metal2 s 14878 0 14892 24640 4 read_bl_0_38
rlabel metal2 s 15004 0 15018 24640 4 read_bl_1_38
rlabel metal2 s 15095 0 15109 24640 4 write_bl_0_38
rlabel metal2 s 15267 0 15281 24640 4 read_bl_0_39
rlabel metal2 s 15393 0 15407 24640 4 read_bl_1_39
rlabel metal2 s 15484 0 15498 24640 4 write_bl_0_39
rlabel metal2 s 15656 0 15670 24640 4 read_bl_0_40
rlabel metal2 s 15782 0 15796 24640 4 read_bl_1_40
rlabel metal2 s 15873 0 15887 24640 4 write_bl_0_40
rlabel metal2 s 16045 0 16059 24640 4 read_bl_0_41
rlabel metal2 s 16171 0 16185 24640 4 read_bl_1_41
rlabel metal2 s 16262 0 16276 24640 4 write_bl_0_41
rlabel metal2 s 16434 0 16448 24640 4 read_bl_0_42
rlabel metal2 s 16560 0 16574 24640 4 read_bl_1_42
rlabel metal2 s 16651 0 16665 24640 4 write_bl_0_42
rlabel metal2 s 16823 0 16837 24640 4 read_bl_0_43
rlabel metal2 s 16949 0 16963 24640 4 read_bl_1_43
rlabel metal2 s 17040 0 17054 24640 4 write_bl_0_43
rlabel metal2 s 17212 0 17226 24640 4 read_bl_0_44
rlabel metal2 s 17338 0 17352 24640 4 read_bl_1_44
rlabel metal2 s 17429 0 17443 24640 4 write_bl_0_44
rlabel metal2 s 17601 0 17615 24640 4 read_bl_0_45
rlabel metal2 s 17727 0 17741 24640 4 read_bl_1_45
rlabel metal2 s 17818 0 17832 24640 4 write_bl_0_45
rlabel metal2 s 17990 0 18004 24640 4 read_bl_0_46
rlabel metal2 s 18116 0 18130 24640 4 read_bl_1_46
rlabel metal2 s 18207 0 18221 24640 4 write_bl_0_46
rlabel metal2 s 18379 0 18393 24640 4 read_bl_0_47
rlabel metal2 s 18505 0 18519 24640 4 read_bl_1_47
rlabel metal2 s 18596 0 18610 24640 4 write_bl_0_47
rlabel metal2 s 18768 0 18782 24640 4 read_bl_0_48
rlabel metal2 s 18894 0 18908 24640 4 read_bl_1_48
rlabel metal2 s 18985 0 18999 24640 4 write_bl_0_48
rlabel metal2 s 19157 0 19171 24640 4 read_bl_0_49
rlabel metal2 s 19283 0 19297 24640 4 read_bl_1_49
rlabel metal2 s 19374 0 19388 24640 4 write_bl_0_49
rlabel metal2 s 19546 0 19560 24640 4 read_bl_0_50
rlabel metal2 s 19672 0 19686 24640 4 read_bl_1_50
rlabel metal2 s 19763 0 19777 24640 4 write_bl_0_50
rlabel metal2 s 19935 0 19949 24640 4 read_bl_0_51
rlabel metal2 s 20061 0 20075 24640 4 read_bl_1_51
rlabel metal2 s 20152 0 20166 24640 4 write_bl_0_51
rlabel metal2 s 20324 0 20338 24640 4 read_bl_0_52
rlabel metal2 s 20450 0 20464 24640 4 read_bl_1_52
rlabel metal2 s 20541 0 20555 24640 4 write_bl_0_52
rlabel metal2 s 20713 0 20727 24640 4 read_bl_0_53
rlabel metal2 s 20839 0 20853 24640 4 read_bl_1_53
rlabel metal2 s 20930 0 20944 24640 4 write_bl_0_53
rlabel metal2 s 21102 0 21116 24640 4 read_bl_0_54
rlabel metal2 s 21228 0 21242 24640 4 read_bl_1_54
rlabel metal2 s 21319 0 21333 24640 4 write_bl_0_54
rlabel metal2 s 21491 0 21505 24640 4 read_bl_0_55
rlabel metal2 s 21617 0 21631 24640 4 read_bl_1_55
rlabel metal2 s 21708 0 21722 24640 4 write_bl_0_55
rlabel metal2 s 21880 0 21894 24640 4 read_bl_0_56
rlabel metal2 s 22006 0 22020 24640 4 read_bl_1_56
rlabel metal2 s 22097 0 22111 24640 4 write_bl_0_56
rlabel metal2 s 22269 0 22283 24640 4 read_bl_0_57
rlabel metal2 s 22395 0 22409 24640 4 read_bl_1_57
rlabel metal2 s 22486 0 22500 24640 4 write_bl_0_57
rlabel metal2 s 22658 0 22672 24640 4 read_bl_0_58
rlabel metal2 s 22784 0 22798 24640 4 read_bl_1_58
rlabel metal2 s 22875 0 22889 24640 4 write_bl_0_58
rlabel metal2 s 23047 0 23061 24640 4 read_bl_0_59
rlabel metal2 s 23173 0 23187 24640 4 read_bl_1_59
rlabel metal2 s 23264 0 23278 24640 4 write_bl_0_59
rlabel metal2 s 23436 0 23450 24640 4 read_bl_0_60
rlabel metal2 s 23562 0 23576 24640 4 read_bl_1_60
rlabel metal2 s 23653 0 23667 24640 4 write_bl_0_60
rlabel metal2 s 23825 0 23839 24640 4 read_bl_0_61
rlabel metal2 s 23951 0 23965 24640 4 read_bl_1_61
rlabel metal2 s 24042 0 24056 24640 4 write_bl_0_61
rlabel metal2 s 24214 0 24228 24640 4 read_bl_0_62
rlabel metal2 s 24340 0 24354 24640 4 read_bl_1_62
rlabel metal2 s 24431 0 24445 24640 4 write_bl_0_62
rlabel metal2 s 24603 0 24617 24640 4 read_bl_0_63
rlabel metal2 s 24729 0 24743 24640 4 read_bl_1_63
rlabel metal2 s 24820 0 24834 24640 4 write_bl_0_63
rlabel metal1 s 0 385 24896 399 4 rwl_0_0
rlabel metal1 s 0 498 24896 512 4 rwl_1_0
rlabel metal1 s 0 322 24896 336 4 wwl_0_0
rlabel metal1 s 0 1141 24896 1155 4 rwl_0_1
rlabel metal1 s 0 1028 24896 1042 4 rwl_1_1
rlabel metal1 s 0 1204 24896 1218 4 wwl_0_1
rlabel metal1 s 0 1925 24896 1939 4 rwl_0_2
rlabel metal1 s 0 2038 24896 2052 4 rwl_1_2
rlabel metal1 s 0 1862 24896 1876 4 wwl_0_2
rlabel metal1 s 0 2681 24896 2695 4 rwl_0_3
rlabel metal1 s 0 2568 24896 2582 4 rwl_1_3
rlabel metal1 s 0 2744 24896 2758 4 wwl_0_3
rlabel metal1 s 0 3465 24896 3479 4 rwl_0_4
rlabel metal1 s 0 3578 24896 3592 4 rwl_1_4
rlabel metal1 s 0 3402 24896 3416 4 wwl_0_4
rlabel metal1 s 0 4221 24896 4235 4 rwl_0_5
rlabel metal1 s 0 4108 24896 4122 4 rwl_1_5
rlabel metal1 s 0 4284 24896 4298 4 wwl_0_5
rlabel metal1 s 0 5005 24896 5019 4 rwl_0_6
rlabel metal1 s 0 5118 24896 5132 4 rwl_1_6
rlabel metal1 s 0 4942 24896 4956 4 wwl_0_6
rlabel metal1 s 0 5761 24896 5775 4 rwl_0_7
rlabel metal1 s 0 5648 24896 5662 4 rwl_1_7
rlabel metal1 s 0 5824 24896 5838 4 wwl_0_7
rlabel metal1 s 0 6545 24896 6559 4 rwl_0_8
rlabel metal1 s 0 6658 24896 6672 4 rwl_1_8
rlabel metal1 s 0 6482 24896 6496 4 wwl_0_8
rlabel metal1 s 0 7301 24896 7315 4 rwl_0_9
rlabel metal1 s 0 7188 24896 7202 4 rwl_1_9
rlabel metal1 s 0 7364 24896 7378 4 wwl_0_9
rlabel metal1 s 0 8085 24896 8099 4 rwl_0_10
rlabel metal1 s 0 8198 24896 8212 4 rwl_1_10
rlabel metal1 s 0 8022 24896 8036 4 wwl_0_10
rlabel metal1 s 0 8841 24896 8855 4 rwl_0_11
rlabel metal1 s 0 8728 24896 8742 4 rwl_1_11
rlabel metal1 s 0 8904 24896 8918 4 wwl_0_11
rlabel metal1 s 0 9625 24896 9639 4 rwl_0_12
rlabel metal1 s 0 9738 24896 9752 4 rwl_1_12
rlabel metal1 s 0 9562 24896 9576 4 wwl_0_12
rlabel metal1 s 0 10381 24896 10395 4 rwl_0_13
rlabel metal1 s 0 10268 24896 10282 4 rwl_1_13
rlabel metal1 s 0 10444 24896 10458 4 wwl_0_13
rlabel metal1 s 0 11165 24896 11179 4 rwl_0_14
rlabel metal1 s 0 11278 24896 11292 4 rwl_1_14
rlabel metal1 s 0 11102 24896 11116 4 wwl_0_14
rlabel metal1 s 0 11921 24896 11935 4 rwl_0_15
rlabel metal1 s 0 11808 24896 11822 4 rwl_1_15
rlabel metal1 s 0 11984 24896 11998 4 wwl_0_15
rlabel metal1 s 0 12705 24896 12719 4 rwl_0_16
rlabel metal1 s 0 12818 24896 12832 4 rwl_1_16
rlabel metal1 s 0 12642 24896 12656 4 wwl_0_16
rlabel metal1 s 0 13461 24896 13475 4 rwl_0_17
rlabel metal1 s 0 13348 24896 13362 4 rwl_1_17
rlabel metal1 s 0 13524 24896 13538 4 wwl_0_17
rlabel metal1 s 0 14245 24896 14259 4 rwl_0_18
rlabel metal1 s 0 14358 24896 14372 4 rwl_1_18
rlabel metal1 s 0 14182 24896 14196 4 wwl_0_18
rlabel metal1 s 0 15001 24896 15015 4 rwl_0_19
rlabel metal1 s 0 14888 24896 14902 4 rwl_1_19
rlabel metal1 s 0 15064 24896 15078 4 wwl_0_19
rlabel metal1 s 0 15785 24896 15799 4 rwl_0_20
rlabel metal1 s 0 15898 24896 15912 4 rwl_1_20
rlabel metal1 s 0 15722 24896 15736 4 wwl_0_20
rlabel metal1 s 0 16541 24896 16555 4 rwl_0_21
rlabel metal1 s 0 16428 24896 16442 4 rwl_1_21
rlabel metal1 s 0 16604 24896 16618 4 wwl_0_21
rlabel metal1 s 0 17325 24896 17339 4 rwl_0_22
rlabel metal1 s 0 17438 24896 17452 4 rwl_1_22
rlabel metal1 s 0 17262 24896 17276 4 wwl_0_22
rlabel metal1 s 0 18081 24896 18095 4 rwl_0_23
rlabel metal1 s 0 17968 24896 17982 4 rwl_1_23
rlabel metal1 s 0 18144 24896 18158 4 wwl_0_23
rlabel metal1 s 0 18865 24896 18879 4 rwl_0_24
rlabel metal1 s 0 18978 24896 18992 4 rwl_1_24
rlabel metal1 s 0 18802 24896 18816 4 wwl_0_24
rlabel metal1 s 0 19621 24896 19635 4 rwl_0_25
rlabel metal1 s 0 19508 24896 19522 4 rwl_1_25
rlabel metal1 s 0 19684 24896 19698 4 wwl_0_25
rlabel metal1 s 0 20405 24896 20419 4 rwl_0_26
rlabel metal1 s 0 20518 24896 20532 4 rwl_1_26
rlabel metal1 s 0 20342 24896 20356 4 wwl_0_26
rlabel metal1 s 0 21161 24896 21175 4 rwl_0_27
rlabel metal1 s 0 21048 24896 21062 4 rwl_1_27
rlabel metal1 s 0 21224 24896 21238 4 wwl_0_27
rlabel metal1 s 0 21945 24896 21959 4 rwl_0_28
rlabel metal1 s 0 22058 24896 22072 4 rwl_1_28
rlabel metal1 s 0 21882 24896 21896 4 wwl_0_28
rlabel metal1 s 0 22701 24896 22715 4 rwl_0_29
rlabel metal1 s 0 22588 24896 22602 4 rwl_1_29
rlabel metal1 s 0 22764 24896 22778 4 wwl_0_29
rlabel metal1 s 0 23485 24896 23499 4 rwl_0_30
rlabel metal1 s 0 23598 24896 23612 4 rwl_1_30
rlabel metal1 s 0 23422 24896 23436 4 wwl_0_30
rlabel metal1 s 0 24241 24896 24255 4 rwl_0_31
rlabel metal1 s 0 24128 24896 24142 4 rwl_1_31
rlabel metal1 s 0 24304 24896 24318 4 wwl_0_31
rlabel metal1 s 1556 755 1945 786 4 vdd
rlabel metal1 s 10114 23855 10503 23886 4 vdd
rlabel metal1 s 22951 23855 23340 23886 4 vdd
rlabel metal1 s 11281 2295 11670 2326 4 vdd
rlabel metal1 s 18283 20775 18672 20806 4 vdd
rlabel metal1 s 2723 3835 3112 3866 4 vdd
rlabel metal1 s 17116 6914 17505 6945 4 vdd
rlabel metal1 s 22951 23854 23340 23885 4 vdd
rlabel metal1 s 24118 2295 24507 2326 4 vdd
rlabel metal1 s 7391 20775 7780 20806 4 vdd
rlabel metal1 s 1945 17694 2334 17725 4 vdd
rlabel metal1 s 1556 3835 1945 3866 4 vdd
rlabel metal1 s 0 19235 389 19266 4 vdd
rlabel metal1 s 20228 8454 20617 8485 4 vdd
rlabel metal1 s 1945 2294 2334 2325 4 vdd
rlabel metal1 s 22173 16154 22562 16185 4 vdd
rlabel metal1 s 19061 20775 19450 20806 4 vdd
rlabel metal1 s 2723 22315 3112 22346 4 vdd
rlabel metal1 s 13226 23854 13615 23885 4 vdd
rlabel metal1 s 7780 23855 8169 23886 4 vdd
rlabel metal1 s 21395 11534 21784 11565 4 vdd
rlabel metal1 s 16727 19234 17116 19265 4 vdd
rlabel metal1 s 6613 11534 7002 11565 4 vdd
rlabel metal1 s 15949 5374 16338 5405 4 vdd
rlabel metal1 s 2334 6914 2723 6945 4 vdd
rlabel metal1 s 7391 755 7780 786 4 vdd
rlabel metal1 s 18283 14614 18672 14645 4 vdd
rlabel metal1 s 20228 19235 20617 19266 4 vdd
rlabel metal1 s 14782 8455 15171 8486 4 vdd
rlabel metal1 s 24118 22315 24507 22346 4 vdd
rlabel metal1 s 17894 5374 18283 5405 4 vdd
rlabel metal1 s 21784 6914 22173 6945 4 vdd
rlabel metal1 s 1556 2295 1945 2326 4 vdd
rlabel metal1 s 24507 23854 24896 23885 4 vdd
rlabel metal1 s 9336 8454 9725 8485 4 vdd
rlabel metal1 s 24118 6915 24507 6946 4 vdd
rlabel metal1 s 3890 13074 4279 13105 4 vdd
rlabel metal1 s 10114 17695 10503 17726 4 vdd
rlabel metal1 s 19450 23855 19839 23886 4 vdd
rlabel metal1 s 4668 22315 5057 22346 4 vdd
rlabel metal1 s 9725 13075 10114 13106 4 vdd
rlabel metal1 s 20228 20774 20617 20805 4 vdd
rlabel metal1 s 19839 19234 20228 19265 4 vdd
rlabel metal1 s 18672 20775 19061 20806 4 vdd
rlabel metal1 s 7780 19234 8169 19265 4 vdd
rlabel metal1 s 17505 17694 17894 17725 4 vdd
rlabel metal1 s 23340 13074 23729 13105 4 vdd
rlabel metal1 s 9336 3835 9725 3866 4 vdd
rlabel metal1 s 2723 20775 3112 20806 4 vdd
rlabel metal1 s 14393 14615 14782 14646 4 vdd
rlabel metal1 s 16727 23854 17116 23885 4 vdd
rlabel metal1 s 1167 20774 1556 20805 4 vdd
rlabel metal1 s 1945 23854 2334 23885 4 vdd
rlabel metal1 s 10503 3834 10892 3865 4 vdd
rlabel metal1 s 16727 6914 17116 6945 4 vdd
rlabel metal1 s 15949 13074 16338 13105 4 vdd
rlabel metal1 s 1556 14614 1945 14645 4 vdd
rlabel metal1 s 17116 22314 17505 22345 4 vdd
rlabel metal1 s 23729 23855 24118 23886 4 vdd
rlabel metal1 s 8947 17694 9336 17725 4 vdd
rlabel metal1 s 20617 20775 21006 20806 4 vdd
rlabel metal1 s 22951 13075 23340 13106 4 vdd
rlabel metal1 s 23729 754 24118 785 4 vdd
rlabel metal1 s 17894 16154 18283 16185 4 vdd
rlabel metal1 s 5057 3834 5446 3865 4 vdd
rlabel metal1 s 8558 23855 8947 23886 4 vdd
rlabel metal1 s 9725 14614 10114 14645 4 vdd
rlabel metal1 s 16338 6914 16727 6945 4 vdd
rlabel metal1 s 0 8455 389 8486 4 vdd
rlabel metal1 s 22173 3835 22562 3866 4 vdd
rlabel metal1 s 20617 755 21006 786 4 vdd
rlabel metal1 s 16727 754 17116 785 4 vdd
rlabel metal1 s 18672 16155 19061 16186 4 vdd
rlabel metal1 s 11281 6915 11670 6946 4 vdd
rlabel metal1 s 22951 20775 23340 20806 4 vdd
rlabel metal1 s 16338 14614 16727 14645 4 vdd
rlabel metal1 s 21784 755 22173 786 4 vdd
rlabel metal1 s 17894 11535 18283 11566 4 vdd
rlabel metal1 s 8169 755 8558 786 4 vdd
rlabel metal1 s 23340 20774 23729 20805 4 vdd
rlabel metal1 s 16338 20775 16727 20806 4 vdd
rlabel metal1 s 17505 3835 17894 3866 4 vdd
rlabel metal1 s 5835 754 6224 785 4 vdd
rlabel metal1 s 8947 3835 9336 3866 4 vdd
rlabel metal1 s 18283 754 18672 785 4 vdd
rlabel metal1 s 17894 11534 18283 11565 4 vdd
rlabel metal1 s 17116 20775 17505 20806 4 vdd
rlabel metal1 s 12059 11535 12448 11566 4 vdd
rlabel metal1 s 5057 11534 5446 11565 4 vdd
rlabel metal1 s 22562 23855 22951 23886 4 vdd
rlabel metal1 s 23729 20775 24118 20806 4 vdd
rlabel metal1 s 19061 13074 19450 13105 4 vdd
rlabel metal1 s 2334 2295 2723 2326 4 vdd
rlabel metal1 s 15171 2295 15560 2326 4 vdd
rlabel metal1 s 15560 8454 15949 8485 4 vdd
rlabel metal1 s 15171 11535 15560 11566 4 vdd
rlabel metal1 s 24118 6914 24507 6945 4 vdd
rlabel metal1 s 4668 3835 5057 3866 4 vdd
rlabel metal1 s 16338 2295 16727 2326 4 vdd
rlabel metal1 s 11281 9994 11670 10025 4 vdd
rlabel metal1 s 8947 2294 9336 2325 4 vdd
rlabel metal1 s 7780 22315 8169 22346 4 vdd
rlabel metal1 s 19061 6915 19450 6946 4 vdd
rlabel metal1 s 23729 13075 24118 13106 4 vdd
rlabel metal1 s 1167 3835 1556 3866 4 vdd
rlabel metal1 s 14004 3835 14393 3866 4 vdd
rlabel metal1 s 14782 754 15171 785 4 vdd
rlabel metal1 s 3890 17694 4279 17725 4 vdd
rlabel metal1 s 5446 16155 5835 16186 4 vdd
rlabel metal1 s 10503 11534 10892 11565 4 vdd
rlabel metal1 s 7002 2294 7391 2325 4 vdd
rlabel metal1 s 4279 20775 4668 20806 4 vdd
rlabel metal1 s 12448 14615 12837 14646 4 vdd
rlabel metal1 s 23729 19235 24118 19266 4 vdd
rlabel metal1 s 8169 11535 8558 11566 4 vdd
rlabel metal1 s 14782 20774 15171 20805 4 vdd
rlabel metal1 s 12448 16154 12837 16185 4 vdd
rlabel metal1 s 13226 20775 13615 20806 4 vdd
rlabel metal1 s 8947 6914 9336 6945 4 vdd
rlabel metal1 s 9725 9994 10114 10025 4 vdd
rlabel metal1 s 2334 22315 2723 22346 4 vdd
rlabel metal1 s 1556 20774 1945 20805 4 vdd
rlabel metal1 s 7780 19235 8169 19266 4 vdd
rlabel metal1 s 4668 20775 5057 20806 4 vdd
rlabel metal1 s 7002 14614 7391 14645 4 vdd
rlabel metal1 s 8947 19234 9336 19265 4 vdd
rlabel metal1 s 19061 19235 19450 19266 4 vdd
rlabel metal1 s 4668 16155 5057 16186 4 vdd
rlabel metal1 s 0 11535 389 11566 4 vdd
rlabel metal1 s 9336 6915 9725 6946 4 vdd
rlabel metal1 s 24118 3835 24507 3866 4 vdd
rlabel metal1 s 20228 16154 20617 16185 4 vdd
rlabel metal1 s 1556 22315 1945 22346 4 vdd
rlabel metal1 s 8558 6915 8947 6946 4 vdd
rlabel metal1 s 10503 17694 10892 17725 4 vdd
rlabel metal1 s 10114 16154 10503 16185 4 vdd
rlabel metal1 s 21395 5374 21784 5405 4 vdd
rlabel metal1 s 5446 17695 5835 17726 4 vdd
rlabel metal1 s 12837 2295 13226 2326 4 vdd
rlabel metal1 s 9336 755 9725 786 4 vdd
rlabel metal1 s 6613 9994 7002 10025 4 vdd
rlabel metal1 s 389 5375 778 5406 4 vdd
rlabel metal1 s 17894 14614 18283 14645 4 vdd
rlabel metal1 s 4279 13074 4668 13105 4 vdd
rlabel metal1 s 6613 11535 7002 11566 4 vdd
rlabel metal1 s 7391 17694 7780 17725 4 vdd
rlabel metal1 s 8169 6915 8558 6946 4 vdd
rlabel metal1 s 20228 5375 20617 5406 4 vdd
rlabel metal1 s 21006 8455 21395 8486 4 vdd
rlabel metal1 s 16727 13075 17116 13106 4 vdd
rlabel metal1 s 24118 8455 24507 8486 4 vdd
rlabel metal1 s 18672 22315 19061 22346 4 vdd
rlabel metal1 s 14393 22315 14782 22346 4 vdd
rlabel metal1 s 24118 22314 24507 22345 4 vdd
rlabel metal1 s 778 16154 1167 16185 4 vdd
rlabel metal1 s 10892 754 11281 785 4 vdd
rlabel metal1 s 3501 8454 3890 8485 4 vdd
rlabel metal1 s 9725 19235 10114 19266 4 vdd
rlabel metal1 s 5835 8455 6224 8486 4 vdd
rlabel metal1 s 5835 14614 6224 14645 4 vdd
rlabel metal1 s 8169 23854 8558 23885 4 vdd
rlabel metal1 s 14393 6915 14782 6946 4 vdd
rlabel metal1 s 12448 9995 12837 10026 4 vdd
rlabel metal1 s 16727 22314 17116 22345 4 vdd
rlabel metal1 s 8947 9995 9336 10026 4 vdd
rlabel metal1 s 5057 11535 5446 11566 4 vdd
rlabel metal1 s 12837 755 13226 786 4 vdd
rlabel metal1 s 24118 16154 24507 16185 4 vdd
rlabel metal1 s 16727 2295 17116 2326 4 vdd
rlabel metal1 s 17116 11534 17505 11565 4 vdd
rlabel metal1 s 8169 9995 8558 10026 4 vdd
rlabel metal1 s 3112 3835 3501 3866 4 vdd
rlabel metal1 s 5446 14615 5835 14646 4 vdd
rlabel metal1 s 20617 22314 21006 22345 4 vdd
rlabel metal1 s 16338 11535 16727 11566 4 vdd
rlabel metal1 s 0 22314 389 22345 4 vdd
rlabel metal1 s 389 2294 778 2325 4 vdd
rlabel metal1 s 12448 5375 12837 5406 4 vdd
rlabel metal1 s 12837 14614 13226 14645 4 vdd
rlabel metal1 s 10503 8455 10892 8486 4 vdd
rlabel metal1 s 11670 23854 12059 23885 4 vdd
rlabel metal1 s 2723 16155 3112 16186 4 vdd
rlabel metal1 s 10892 9995 11281 10026 4 vdd
rlabel metal1 s 16338 755 16727 786 4 vdd
rlabel metal1 s 389 755 778 786 4 vdd
rlabel metal1 s 8947 14615 9336 14646 4 vdd
rlabel metal1 s 8169 2295 8558 2326 4 vdd
rlabel metal1 s 20228 3834 20617 3865 4 vdd
rlabel metal1 s 8169 3835 8558 3866 4 vdd
rlabel metal1 s 778 20774 1167 20805 4 vdd
rlabel metal1 s 8947 5374 9336 5405 4 vdd
rlabel metal1 s 17894 23854 18283 23885 4 vdd
rlabel metal1 s 4668 6915 5057 6946 4 vdd
rlabel metal1 s 18283 11534 18672 11565 4 vdd
rlabel metal1 s 15560 3834 15949 3865 4 vdd
rlabel metal1 s 18283 14615 18672 14646 4 vdd
rlabel metal1 s 1945 6914 2334 6945 4 vdd
rlabel metal1 s 13226 6914 13615 6945 4 vdd
rlabel metal1 s 4668 9995 5057 10026 4 vdd
rlabel metal1 s 12059 17695 12448 17726 4 vdd
rlabel metal1 s 6613 14615 7002 14646 4 vdd
rlabel metal1 s 18283 22315 18672 22346 4 vdd
rlabel metal1 s 20617 14614 21006 14645 4 vdd
rlabel metal1 s 12059 3835 12448 3866 4 vdd
rlabel metal1 s 9336 8455 9725 8486 4 vdd
rlabel metal1 s 2334 17694 2723 17725 4 vdd
rlabel metal1 s 8558 20775 8947 20806 4 vdd
rlabel metal1 s 11281 20775 11670 20806 4 vdd
rlabel metal1 s 23729 22315 24118 22346 4 vdd
rlabel metal1 s 7002 3834 7391 3865 4 vdd
rlabel metal1 s 8169 23855 8558 23886 4 vdd
rlabel metal1 s 7391 3834 7780 3865 4 vdd
rlabel metal1 s 12837 5375 13226 5406 4 vdd
rlabel metal1 s 4668 17695 5057 17726 4 vdd
rlabel metal1 s 1945 22315 2334 22346 4 vdd
rlabel metal1 s 22562 19235 22951 19266 4 vdd
rlabel metal1 s 21395 3834 21784 3865 4 vdd
rlabel metal1 s 13226 8455 13615 8486 4 vdd
rlabel metal1 s 3890 19235 4279 19266 4 vdd
rlabel metal1 s 23340 23854 23729 23885 4 vdd
rlabel metal1 s 15949 5375 16338 5406 4 vdd
rlabel metal1 s 0 20774 389 20805 4 vdd
rlabel metal1 s 10114 6914 10503 6945 4 vdd
rlabel metal1 s 15171 23854 15560 23885 4 vdd
rlabel metal1 s 13226 2295 13615 2326 4 vdd
rlabel metal1 s 16338 8455 16727 8486 4 vdd
rlabel metal1 s 10503 22315 10892 22346 4 vdd
rlabel metal1 s 17505 23854 17894 23885 4 vdd
rlabel metal1 s 9725 8455 10114 8486 4 vdd
rlabel metal1 s 21784 13074 22173 13105 4 vdd
rlabel metal1 s 23340 3834 23729 3865 4 vdd
rlabel metal1 s 17116 23855 17505 23886 4 vdd
rlabel metal1 s 14782 8454 15171 8485 4 vdd
rlabel metal1 s 19450 17695 19839 17726 4 vdd
rlabel metal1 s 3501 20775 3890 20806 4 vdd
rlabel metal1 s 23340 9995 23729 10026 4 vdd
rlabel metal1 s 14393 5374 14782 5405 4 vdd
rlabel metal1 s 13615 2295 14004 2326 4 vdd
rlabel metal1 s 8947 14614 9336 14645 4 vdd
rlabel metal1 s 10114 14615 10503 14646 4 vdd
rlabel metal1 s 3112 17694 3501 17725 4 vdd
rlabel metal1 s 1556 11534 1945 11565 4 vdd
rlabel metal1 s 5057 20774 5446 20805 4 vdd
rlabel metal1 s 15560 2295 15949 2326 4 vdd
rlabel metal1 s 5057 9994 5446 10025 4 vdd
rlabel metal1 s 23729 20774 24118 20805 4 vdd
rlabel metal1 s 6613 8455 7002 8486 4 vdd
rlabel metal1 s 7391 754 7780 785 4 vdd
rlabel metal1 s 9336 5374 9725 5405 4 vdd
rlabel metal1 s 7002 22315 7391 22346 4 vdd
rlabel metal1 s 24507 23855 24896 23886 4 vdd
rlabel metal1 s 5446 20774 5835 20805 4 vdd
rlabel metal1 s 20228 23854 20617 23885 4 vdd
rlabel metal1 s 0 2295 389 2326 4 vdd
rlabel metal1 s 19450 23854 19839 23885 4 vdd
rlabel metal1 s 5446 19235 5835 19266 4 vdd
rlabel metal1 s 10114 6915 10503 6946 4 vdd
rlabel metal1 s 1945 5374 2334 5405 4 vdd
rlabel metal1 s 24118 2294 24507 2325 4 vdd
rlabel metal1 s 2334 754 2723 785 4 vdd
rlabel metal1 s 21006 16155 21395 16186 4 vdd
rlabel metal1 s 15949 23854 16338 23885 4 vdd
rlabel metal1 s 2334 13074 2723 13105 4 vdd
rlabel metal1 s 1945 8455 2334 8486 4 vdd
rlabel metal1 s 24507 20774 24896 20805 4 vdd
rlabel metal1 s 14782 16155 15171 16186 4 vdd
rlabel metal1 s 5835 22315 6224 22346 4 vdd
rlabel metal1 s 6224 9995 6613 10026 4 vdd
rlabel metal1 s 3501 13074 3890 13105 4 vdd
rlabel metal1 s 5835 22314 6224 22345 4 vdd
rlabel metal1 s 8947 8455 9336 8486 4 vdd
rlabel metal1 s 19450 9994 19839 10025 4 vdd
rlabel metal1 s 7002 6914 7391 6945 4 vdd
rlabel metal1 s 21784 3835 22173 3866 4 vdd
rlabel metal1 s 8169 14615 8558 14646 4 vdd
rlabel metal1 s 3112 20774 3501 20805 4 vdd
rlabel metal1 s 2723 23855 3112 23886 4 vdd
rlabel metal1 s 20228 6914 20617 6945 4 vdd
rlabel metal1 s 14004 9995 14393 10026 4 vdd
rlabel metal1 s 15171 16155 15560 16186 4 vdd
rlabel metal1 s 22173 754 22562 785 4 vdd
rlabel metal1 s 8558 16155 8947 16186 4 vdd
rlabel metal1 s 12448 23855 12837 23886 4 vdd
rlabel metal1 s 17505 17695 17894 17726 4 vdd
rlabel metal1 s 3501 23855 3890 23886 4 vdd
rlabel metal1 s 1167 9995 1556 10026 4 vdd
rlabel metal1 s 18283 19234 18672 19265 4 vdd
rlabel metal1 s 4279 23854 4668 23885 4 vdd
rlabel metal1 s 2334 14615 2723 14646 4 vdd
rlabel metal1 s 3112 9994 3501 10025 4 vdd
rlabel metal1 s 22562 2295 22951 2326 4 vdd
rlabel metal1 s 5835 3835 6224 3866 4 vdd
rlabel metal1 s 17116 17695 17505 17726 4 vdd
rlabel metal1 s 16727 17695 17116 17726 4 vdd
rlabel metal1 s 15560 22315 15949 22346 4 vdd
rlabel metal1 s 11670 8455 12059 8486 4 vdd
rlabel metal1 s 11281 8455 11670 8486 4 vdd
rlabel metal1 s 17894 3834 18283 3865 4 vdd
rlabel metal1 s 1556 9995 1945 10026 4 vdd
rlabel metal1 s 10114 13074 10503 13105 4 vdd
rlabel metal1 s 13615 13075 14004 13106 4 vdd
rlabel metal1 s 9336 19235 9725 19266 4 vdd
rlabel metal1 s 1945 20774 2334 20805 4 vdd
rlabel metal1 s 1945 20775 2334 20806 4 vdd
rlabel metal1 s 1556 13074 1945 13105 4 vdd
rlabel metal1 s 22951 755 23340 786 4 vdd
rlabel metal1 s 8169 9994 8558 10025 4 vdd
rlabel metal1 s 22173 13075 22562 13106 4 vdd
rlabel metal1 s 8169 19234 8558 19265 4 vdd
rlabel metal1 s 13615 9994 14004 10025 4 vdd
rlabel metal1 s 21006 2295 21395 2326 4 vdd
rlabel metal1 s 20228 13074 20617 13105 4 vdd
rlabel metal1 s 24507 5375 24896 5406 4 vdd
rlabel metal1 s 11670 3834 12059 3865 4 vdd
rlabel metal1 s 18283 13074 18672 13105 4 vdd
rlabel metal1 s 7391 11534 7780 11565 4 vdd
rlabel metal1 s 4279 8454 4668 8485 4 vdd
rlabel metal1 s 12059 13074 12448 13105 4 vdd
rlabel metal1 s 23340 17695 23729 17726 4 vdd
rlabel metal1 s 7002 19235 7391 19266 4 vdd
rlabel metal1 s 10892 17694 11281 17725 4 vdd
rlabel metal1 s 14004 5374 14393 5405 4 vdd
rlabel metal1 s 778 13074 1167 13105 4 vdd
rlabel metal1 s 23340 23855 23729 23886 4 vdd
rlabel metal1 s 15949 8455 16338 8486 4 vdd
rlabel metal1 s 22562 755 22951 786 4 vdd
rlabel metal1 s 24507 11534 24896 11565 4 vdd
rlabel metal1 s 3112 11535 3501 11566 4 vdd
rlabel metal1 s 12059 16155 12448 16186 4 vdd
rlabel metal1 s 0 6914 389 6945 4 vdd
rlabel metal1 s 2334 16155 2723 16186 4 vdd
rlabel metal1 s 9336 22315 9725 22346 4 vdd
rlabel metal1 s 13615 8455 14004 8486 4 vdd
rlabel metal1 s 18283 13075 18672 13106 4 vdd
rlabel metal1 s 22562 5375 22951 5406 4 vdd
rlabel metal1 s 22951 9995 23340 10026 4 vdd
rlabel metal1 s 9725 23854 10114 23885 4 vdd
rlabel metal1 s 7391 2295 7780 2326 4 vdd
rlabel metal1 s 19061 3835 19450 3866 4 vdd
rlabel metal1 s 12059 2295 12448 2326 4 vdd
rlabel metal1 s 7780 16154 8169 16185 4 vdd
rlabel metal1 s 15560 19234 15949 19265 4 vdd
rlabel metal1 s 16338 19235 16727 19266 4 vdd
rlabel metal1 s 8558 3835 8947 3866 4 vdd
rlabel metal1 s 3112 9995 3501 10026 4 vdd
rlabel metal1 s 3890 23854 4279 23885 4 vdd
rlabel metal1 s 15560 13074 15949 13105 4 vdd
rlabel metal1 s 15949 2295 16338 2326 4 vdd
rlabel metal1 s 11670 6915 12059 6946 4 vdd
rlabel metal1 s 21784 14614 22173 14645 4 vdd
rlabel metal1 s 15560 3835 15949 3866 4 vdd
rlabel metal1 s 7002 11535 7391 11566 4 vdd
rlabel metal1 s 0 13075 389 13106 4 vdd
rlabel metal1 s 13226 8454 13615 8485 4 vdd
rlabel metal1 s 16727 9994 17116 10025 4 vdd
rlabel metal1 s 3890 16154 4279 16185 4 vdd
rlabel metal1 s 20617 9994 21006 10025 4 vdd
rlabel metal1 s 7002 17694 7391 17725 4 vdd
rlabel metal1 s 4279 2295 4668 2326 4 vdd
rlabel metal1 s 21395 755 21784 786 4 vdd
rlabel metal1 s 6613 14614 7002 14645 4 vdd
rlabel metal1 s 22173 17694 22562 17725 4 vdd
rlabel metal1 s 9336 23854 9725 23885 4 vdd
rlabel metal1 s 10503 16154 10892 16185 4 vdd
rlabel metal1 s 21784 8454 22173 8485 4 vdd
rlabel metal1 s 5835 20775 6224 20806 4 vdd
rlabel metal1 s 7780 2294 8169 2325 4 vdd
rlabel metal1 s 4279 22315 4668 22346 4 vdd
rlabel metal1 s 14004 17694 14393 17725 4 vdd
rlabel metal1 s 13615 16154 14004 16185 4 vdd
rlabel metal1 s 22562 6914 22951 6945 4 vdd
rlabel metal1 s 12448 13075 12837 13106 4 vdd
rlabel metal1 s 10892 6914 11281 6945 4 vdd
rlabel metal1 s 17505 754 17894 785 4 vdd
rlabel metal1 s 7002 8454 7391 8485 4 vdd
rlabel metal1 s 2334 11535 2723 11566 4 vdd
rlabel metal1 s 9336 3834 9725 3865 4 vdd
rlabel metal1 s 10114 3835 10503 3866 4 vdd
rlabel metal1 s 18283 16155 18672 16186 4 vdd
rlabel metal1 s 15171 20774 15560 20805 4 vdd
rlabel metal1 s 8558 23854 8947 23885 4 vdd
rlabel metal1 s 2723 11535 3112 11566 4 vdd
rlabel metal1 s 13226 3834 13615 3865 4 vdd
rlabel metal1 s 20228 5374 20617 5405 4 vdd
rlabel metal1 s 0 17694 389 17725 4 vdd
rlabel metal1 s 18283 2294 18672 2325 4 vdd
rlabel metal1 s 21784 3834 22173 3865 4 vdd
rlabel metal1 s 18672 19234 19061 19265 4 vdd
rlabel metal1 s 778 19235 1167 19266 4 vdd
rlabel metal1 s 16338 13075 16727 13106 4 vdd
rlabel metal1 s 21784 5375 22173 5406 4 vdd
rlabel metal1 s 22173 8455 22562 8486 4 vdd
rlabel metal1 s 12448 8454 12837 8485 4 vdd
rlabel metal1 s 24507 22315 24896 22346 4 vdd
rlabel metal1 s 19061 22315 19450 22346 4 vdd
rlabel metal1 s 11281 11535 11670 11566 4 vdd
rlabel metal1 s 15560 6915 15949 6946 4 vdd
rlabel metal1 s 15171 755 15560 786 4 vdd
rlabel metal1 s 10503 754 10892 785 4 vdd
rlabel metal1 s 9725 16155 10114 16186 4 vdd
rlabel metal1 s 17505 755 17894 786 4 vdd
rlabel metal1 s 7391 13075 7780 13106 4 vdd
rlabel metal1 s 4279 11534 4668 11565 4 vdd
rlabel metal1 s 13226 11535 13615 11566 4 vdd
rlabel metal1 s 8558 5374 8947 5405 4 vdd
rlabel metal1 s 13615 20775 14004 20806 4 vdd
rlabel metal1 s 8558 8455 8947 8486 4 vdd
rlabel metal1 s 20617 13075 21006 13106 4 vdd
rlabel metal1 s 19450 8455 19839 8486 4 vdd
rlabel metal1 s 22562 13075 22951 13106 4 vdd
rlabel metal1 s 15171 17695 15560 17726 4 vdd
rlabel metal1 s 17116 23854 17505 23885 4 vdd
rlabel metal1 s 21784 22314 22173 22345 4 vdd
rlabel metal1 s 19061 8455 19450 8486 4 vdd
rlabel metal1 s 15949 22315 16338 22346 4 vdd
rlabel metal1 s 22562 3834 22951 3865 4 vdd
rlabel metal1 s 11281 19235 11670 19266 4 vdd
rlabel metal1 s 22173 11535 22562 11566 4 vdd
rlabel metal1 s 1556 19235 1945 19266 4 vdd
rlabel metal1 s 778 3835 1167 3866 4 vdd
rlabel metal1 s 8558 22314 8947 22345 4 vdd
rlabel metal1 s 8947 3834 9336 3865 4 vdd
rlabel metal1 s 19450 19235 19839 19266 4 vdd
rlabel metal1 s 23340 2294 23729 2325 4 vdd
rlabel metal1 s 15560 23855 15949 23886 4 vdd
rlabel metal1 s 1945 2295 2334 2326 4 vdd
rlabel metal1 s 5446 5374 5835 5405 4 vdd
rlabel metal1 s 21395 16155 21784 16186 4 vdd
rlabel metal1 s 5446 20775 5835 20806 4 vdd
rlabel metal1 s 19839 22315 20228 22346 4 vdd
rlabel metal1 s 778 22315 1167 22346 4 vdd
rlabel metal1 s 23729 3834 24118 3865 4 vdd
rlabel metal1 s 2334 8455 2723 8486 4 vdd
rlabel metal1 s 24507 8454 24896 8485 4 vdd
rlabel metal1 s 1556 5375 1945 5406 4 vdd
rlabel metal1 s 1945 8454 2334 8485 4 vdd
rlabel metal1 s 2334 13075 2723 13106 4 vdd
rlabel metal1 s 12448 17694 12837 17725 4 vdd
rlabel metal1 s 19061 2294 19450 2325 4 vdd
rlabel metal1 s 7391 9994 7780 10025 4 vdd
rlabel metal1 s 22951 14615 23340 14646 4 vdd
rlabel metal1 s 389 19234 778 19265 4 vdd
rlabel metal1 s 5446 22315 5835 22346 4 vdd
rlabel metal1 s 5057 23854 5446 23885 4 vdd
rlabel metal1 s 3501 6914 3890 6945 4 vdd
rlabel metal1 s 3890 6915 4279 6946 4 vdd
rlabel metal1 s 21395 22315 21784 22346 4 vdd
rlabel metal1 s 10503 13075 10892 13106 4 vdd
rlabel metal1 s 14004 19234 14393 19265 4 vdd
rlabel metal1 s 1945 19234 2334 19265 4 vdd
rlabel metal1 s 7780 3835 8169 3866 4 vdd
rlabel metal1 s 389 23855 778 23886 4 vdd
rlabel metal1 s 1167 20775 1556 20806 4 vdd
rlabel metal1 s 6613 6915 7002 6946 4 vdd
rlabel metal1 s 5835 8454 6224 8485 4 vdd
rlabel metal1 s 22173 8454 22562 8485 4 vdd
rlabel metal1 s 14782 6915 15171 6946 4 vdd
rlabel metal1 s 22173 13074 22562 13105 4 vdd
rlabel metal1 s 17894 2295 18283 2326 4 vdd
rlabel metal1 s 16338 3834 16727 3865 4 vdd
rlabel metal1 s 7002 3835 7391 3866 4 vdd
rlabel metal1 s 12448 22314 12837 22345 4 vdd
rlabel metal1 s 23340 8455 23729 8486 4 vdd
rlabel metal1 s 15560 5375 15949 5406 4 vdd
rlabel metal1 s 6613 17695 7002 17726 4 vdd
rlabel metal1 s 3890 11534 4279 11565 4 vdd
rlabel metal1 s 15949 19235 16338 19266 4 vdd
rlabel metal1 s 778 9995 1167 10026 4 vdd
rlabel metal1 s 6224 2294 6613 2325 4 vdd
rlabel metal1 s 24507 14615 24896 14646 4 vdd
rlabel metal1 s 17894 20774 18283 20805 4 vdd
rlabel metal1 s 22173 20775 22562 20806 4 vdd
rlabel metal1 s 5835 9995 6224 10026 4 vdd
rlabel metal1 s 11670 17694 12059 17725 4 vdd
rlabel metal1 s 16727 2294 17116 2325 4 vdd
rlabel metal1 s 1945 3835 2334 3866 4 vdd
rlabel metal1 s 14393 19235 14782 19266 4 vdd
rlabel metal1 s 14782 20775 15171 20806 4 vdd
rlabel metal1 s 20617 23854 21006 23885 4 vdd
rlabel metal1 s 22562 20774 22951 20805 4 vdd
rlabel metal1 s 19061 16155 19450 16186 4 vdd
rlabel metal1 s 19061 17695 19450 17726 4 vdd
rlabel metal1 s 24507 9994 24896 10025 4 vdd
rlabel metal1 s 14004 16155 14393 16186 4 vdd
rlabel metal1 s 5446 3834 5835 3865 4 vdd
rlabel metal1 s 3112 8454 3501 8485 4 vdd
rlabel metal1 s 12837 23854 13226 23885 4 vdd
rlabel metal1 s 21784 14615 22173 14646 4 vdd
rlabel metal1 s 2334 16154 2723 16185 4 vdd
rlabel metal1 s 8169 8454 8558 8485 4 vdd
rlabel metal1 s 19450 9995 19839 10026 4 vdd
rlabel metal1 s 15171 20775 15560 20806 4 vdd
rlabel metal1 s 12059 9995 12448 10026 4 vdd
rlabel metal1 s 7391 14615 7780 14646 4 vdd
rlabel metal1 s 778 2294 1167 2325 4 vdd
rlabel metal1 s 20617 2294 21006 2325 4 vdd
rlabel metal1 s 19450 14614 19839 14645 4 vdd
rlabel metal1 s 12059 20775 12448 20806 4 vdd
rlabel metal1 s 12059 9994 12448 10025 4 vdd
rlabel metal1 s 21006 11534 21395 11565 4 vdd
rlabel metal1 s 12059 5375 12448 5406 4 vdd
rlabel metal1 s 9725 6915 10114 6946 4 vdd
rlabel metal1 s 12448 11534 12837 11565 4 vdd
rlabel metal1 s 16727 13074 17116 13105 4 vdd
rlabel metal1 s 23729 6914 24118 6945 4 vdd
rlabel metal1 s 7002 11534 7391 11565 4 vdd
rlabel metal1 s 3501 11535 3890 11566 4 vdd
rlabel metal1 s 21784 23855 22173 23886 4 vdd
rlabel metal1 s 14393 22314 14782 22345 4 vdd
rlabel metal1 s 21006 754 21395 785 4 vdd
rlabel metal1 s 19450 22314 19839 22345 4 vdd
rlabel metal1 s 3890 755 4279 786 4 vdd
rlabel metal1 s 389 3834 778 3865 4 vdd
rlabel metal1 s 11670 14615 12059 14646 4 vdd
rlabel metal1 s 12448 6914 12837 6945 4 vdd
rlabel metal1 s 4279 13075 4668 13106 4 vdd
rlabel metal1 s 8558 9994 8947 10025 4 vdd
rlabel metal1 s 9336 2294 9725 2325 4 vdd
rlabel metal1 s 4279 3834 4668 3865 4 vdd
rlabel metal1 s 17505 11535 17894 11566 4 vdd
rlabel metal1 s 10503 5374 10892 5405 4 vdd
rlabel metal1 s 2723 3834 3112 3865 4 vdd
rlabel metal1 s 14004 11535 14393 11566 4 vdd
rlabel metal1 s 22951 754 23340 785 4 vdd
rlabel metal1 s 3112 13074 3501 13105 4 vdd
rlabel metal1 s 11281 11534 11670 11565 4 vdd
rlabel metal1 s 12837 17694 13226 17725 4 vdd
rlabel metal1 s 22173 755 22562 786 4 vdd
rlabel metal1 s 8169 754 8558 785 4 vdd
rlabel metal1 s 10114 13075 10503 13106 4 vdd
rlabel metal1 s 17505 14615 17894 14646 4 vdd
rlabel metal1 s 3501 20774 3890 20805 4 vdd
rlabel metal1 s 3890 14614 4279 14645 4 vdd
rlabel metal1 s 17505 22314 17894 22345 4 vdd
rlabel metal1 s 21395 20775 21784 20806 4 vdd
rlabel metal1 s 24507 6915 24896 6946 4 vdd
rlabel metal1 s 7391 2294 7780 2325 4 vdd
rlabel metal1 s 24118 23855 24507 23886 4 vdd
rlabel metal1 s 7780 13074 8169 13105 4 vdd
rlabel metal1 s 0 14614 389 14645 4 vdd
rlabel metal1 s 18283 11535 18672 11566 4 vdd
rlabel metal1 s 5057 13075 5446 13106 4 vdd
rlabel metal1 s 20228 14615 20617 14646 4 vdd
rlabel metal1 s 5446 5375 5835 5406 4 vdd
rlabel metal1 s 16338 9995 16727 10026 4 vdd
rlabel metal1 s 11670 23855 12059 23886 4 vdd
rlabel metal1 s 0 3834 389 3865 4 vdd
rlabel metal1 s 15171 3834 15560 3865 4 vdd
rlabel metal1 s 5057 754 5446 785 4 vdd
rlabel metal1 s 19839 6915 20228 6946 4 vdd
rlabel metal1 s 4279 2294 4668 2325 4 vdd
rlabel metal1 s 23729 9995 24118 10026 4 vdd
rlabel metal1 s 3890 6914 4279 6945 4 vdd
rlabel metal1 s 19450 16155 19839 16186 4 vdd
rlabel metal1 s 14393 9995 14782 10026 4 vdd
rlabel metal1 s 21006 13074 21395 13105 4 vdd
rlabel metal1 s 11281 16155 11670 16186 4 vdd
rlabel metal1 s 23340 6915 23729 6946 4 vdd
rlabel metal1 s 7391 5375 7780 5406 4 vdd
rlabel metal1 s 14393 20775 14782 20806 4 vdd
rlabel metal1 s 11281 22315 11670 22346 4 vdd
rlabel metal1 s 15949 2294 16338 2325 4 vdd
rlabel metal1 s 7780 13075 8169 13106 4 vdd
rlabel metal1 s 9725 2295 10114 2326 4 vdd
rlabel metal1 s 24507 16154 24896 16185 4 vdd
rlabel metal1 s 7780 22314 8169 22345 4 vdd
rlabel metal1 s 12837 19234 13226 19265 4 vdd
rlabel metal1 s 17505 19234 17894 19265 4 vdd
rlabel metal1 s 21395 754 21784 785 4 vdd
rlabel metal1 s 23729 16155 24118 16186 4 vdd
rlabel metal1 s 5835 17694 6224 17725 4 vdd
rlabel metal1 s 7391 6914 7780 6945 4 vdd
rlabel metal1 s 11670 8454 12059 8485 4 vdd
rlabel metal1 s 19450 5374 19839 5405 4 vdd
rlabel metal1 s 15560 9994 15949 10025 4 vdd
rlabel metal1 s 7780 8454 8169 8485 4 vdd
rlabel metal1 s 16727 3834 17116 3865 4 vdd
rlabel metal1 s 10503 9995 10892 10026 4 vdd
rlabel metal1 s 16338 5374 16727 5405 4 vdd
rlabel metal1 s 14004 13075 14393 13106 4 vdd
rlabel metal1 s 21006 9994 21395 10025 4 vdd
rlabel metal1 s 7780 20775 8169 20806 4 vdd
rlabel metal1 s 7391 23855 7780 23886 4 vdd
rlabel metal1 s 3501 16154 3890 16185 4 vdd
rlabel metal1 s 19450 3834 19839 3865 4 vdd
rlabel metal1 s 21395 23854 21784 23885 4 vdd
rlabel metal1 s 16727 8455 17116 8486 4 vdd
rlabel metal1 s 10503 20774 10892 20805 4 vdd
rlabel metal1 s 3890 9995 4279 10026 4 vdd
rlabel metal1 s 16338 3835 16727 3866 4 vdd
rlabel metal1 s 20617 11535 21006 11566 4 vdd
rlabel metal1 s 6224 754 6613 785 4 vdd
rlabel metal1 s 3890 11535 4279 11566 4 vdd
rlabel metal1 s 15171 16154 15560 16185 4 vdd
rlabel metal1 s 17894 23855 18283 23886 4 vdd
rlabel metal1 s 16727 16154 17116 16185 4 vdd
rlabel metal1 s 6224 14615 6613 14646 4 vdd
rlabel metal1 s 21395 13074 21784 13105 4 vdd
rlabel metal1 s 15171 19234 15560 19265 4 vdd
rlabel metal1 s 3890 20774 4279 20805 4 vdd
rlabel metal1 s 16727 14614 17116 14645 4 vdd
rlabel metal1 s 21006 6914 21395 6945 4 vdd
rlabel metal1 s 13615 22315 14004 22346 4 vdd
rlabel metal1 s 7002 6915 7391 6946 4 vdd
rlabel metal1 s 5057 8455 5446 8486 4 vdd
rlabel metal1 s 4668 20774 5057 20805 4 vdd
rlabel metal1 s 1167 755 1556 786 4 vdd
rlabel metal1 s 19061 9994 19450 10025 4 vdd
rlabel metal1 s 1167 6915 1556 6946 4 vdd
rlabel metal1 s 22951 9994 23340 10025 4 vdd
rlabel metal1 s 3112 13075 3501 13106 4 vdd
rlabel metal1 s 12059 13075 12448 13106 4 vdd
rlabel metal1 s 2723 5374 3112 5405 4 vdd
rlabel metal1 s 22173 5374 22562 5405 4 vdd
rlabel metal1 s 19061 20774 19450 20805 4 vdd
rlabel metal1 s 6613 23854 7002 23885 4 vdd
rlabel metal1 s 19061 3834 19450 3865 4 vdd
rlabel metal1 s 11281 23855 11670 23886 4 vdd
rlabel metal1 s 15560 8455 15949 8486 4 vdd
rlabel metal1 s 20228 22315 20617 22346 4 vdd
rlabel metal1 s 1945 13075 2334 13106 4 vdd
rlabel metal1 s 0 9995 389 10026 4 vdd
rlabel metal1 s 22562 5374 22951 5405 4 vdd
rlabel metal1 s 15171 22314 15560 22345 4 vdd
rlabel metal1 s 16338 23854 16727 23885 4 vdd
rlabel metal1 s 4279 8455 4668 8486 4 vdd
rlabel metal1 s 10892 5374 11281 5405 4 vdd
rlabel metal1 s 10503 22314 10892 22345 4 vdd
rlabel metal1 s 6613 3835 7002 3866 4 vdd
rlabel metal1 s 21006 19235 21395 19266 4 vdd
rlabel metal1 s 24507 2294 24896 2325 4 vdd
rlabel metal1 s 1945 23855 2334 23886 4 vdd
rlabel metal1 s 20228 9995 20617 10026 4 vdd
rlabel metal1 s 9725 755 10114 786 4 vdd
rlabel metal1 s 7780 754 8169 785 4 vdd
rlabel metal1 s 1556 14615 1945 14646 4 vdd
rlabel metal1 s 22173 9995 22562 10026 4 vdd
rlabel metal1 s 21784 19234 22173 19265 4 vdd
rlabel metal1 s 6613 23855 7002 23886 4 vdd
rlabel metal1 s 11281 3834 11670 3865 4 vdd
rlabel metal1 s 11670 5375 12059 5406 4 vdd
rlabel metal1 s 1556 9994 1945 10025 4 vdd
rlabel metal1 s 8558 5375 8947 5406 4 vdd
rlabel metal1 s 23340 3835 23729 3866 4 vdd
rlabel metal1 s 20228 20775 20617 20806 4 vdd
rlabel metal1 s 11670 5374 12059 5405 4 vdd
rlabel metal1 s 12837 13075 13226 13106 4 vdd
rlabel metal1 s 19450 20775 19839 20806 4 vdd
rlabel metal1 s 6613 19234 7002 19265 4 vdd
rlabel metal1 s 24118 19235 24507 19266 4 vdd
rlabel metal1 s 1556 20775 1945 20806 4 vdd
rlabel metal1 s 3890 20775 4279 20806 4 vdd
rlabel metal1 s 18672 755 19061 786 4 vdd
rlabel metal1 s 10503 14614 10892 14645 4 vdd
rlabel metal1 s 11281 14614 11670 14645 4 vdd
rlabel metal1 s 22562 13074 22951 13105 4 vdd
rlabel metal1 s 11281 2294 11670 2325 4 vdd
rlabel metal1 s 5446 9994 5835 10025 4 vdd
rlabel metal1 s 20617 19234 21006 19265 4 vdd
rlabel metal1 s 12837 8455 13226 8486 4 vdd
rlabel metal1 s 6224 14614 6613 14645 4 vdd
rlabel metal1 s 20228 11535 20617 11566 4 vdd
rlabel metal1 s 2723 13075 3112 13106 4 vdd
rlabel metal1 s 19839 22314 20228 22345 4 vdd
rlabel metal1 s 0 755 389 786 4 vdd
rlabel metal1 s 23340 754 23729 785 4 vdd
rlabel metal1 s 24507 20775 24896 20806 4 vdd
rlabel metal1 s 19839 20775 20228 20806 4 vdd
rlabel metal1 s 14782 5374 15171 5405 4 vdd
rlabel metal1 s 14004 755 14393 786 4 vdd
rlabel metal1 s 13226 20774 13615 20805 4 vdd
rlabel metal1 s 8947 8454 9336 8485 4 vdd
rlabel metal1 s 22951 2294 23340 2325 4 vdd
rlabel metal1 s 23340 9994 23729 10025 4 vdd
rlabel metal1 s 20617 11534 21006 11565 4 vdd
rlabel metal1 s 14782 3835 15171 3866 4 vdd
rlabel metal1 s 22951 6914 23340 6945 4 vdd
rlabel metal1 s 6224 13074 6613 13105 4 vdd
rlabel metal1 s 14004 9994 14393 10025 4 vdd
rlabel metal1 s 2723 5375 3112 5406 4 vdd
rlabel metal1 s 2723 14615 3112 14646 4 vdd
rlabel metal1 s 12448 16155 12837 16186 4 vdd
rlabel metal1 s 10503 19234 10892 19265 4 vdd
rlabel metal1 s 9725 754 10114 785 4 vdd
rlabel metal1 s 16338 2294 16727 2325 4 vdd
rlabel metal1 s 5446 3835 5835 3866 4 vdd
rlabel metal1 s 8947 9994 9336 10025 4 vdd
rlabel metal1 s 21395 16154 21784 16185 4 vdd
rlabel metal1 s 10503 3835 10892 3866 4 vdd
rlabel metal1 s 8558 16154 8947 16185 4 vdd
rlabel metal1 s 9725 23855 10114 23886 4 vdd
rlabel metal1 s 4668 755 5057 786 4 vdd
rlabel metal1 s 14004 17695 14393 17726 4 vdd
rlabel metal1 s 12448 20775 12837 20806 4 vdd
rlabel metal1 s 14393 11535 14782 11566 4 vdd
rlabel metal1 s 4668 13074 5057 13105 4 vdd
rlabel metal1 s 5057 755 5446 786 4 vdd
rlabel metal1 s 21395 9995 21784 10026 4 vdd
rlabel metal1 s 9725 6914 10114 6945 4 vdd
rlabel metal1 s 6224 20775 6613 20806 4 vdd
rlabel metal1 s 4279 6915 4668 6946 4 vdd
rlabel metal1 s 10114 16155 10503 16186 4 vdd
rlabel metal1 s 8169 16155 8558 16186 4 vdd
rlabel metal1 s 5446 755 5835 786 4 vdd
rlabel metal1 s 11281 20774 11670 20805 4 vdd
rlabel metal1 s 9336 754 9725 785 4 vdd
rlabel metal1 s 19839 13074 20228 13105 4 vdd
rlabel metal1 s 8947 754 9336 785 4 vdd
rlabel metal1 s 9336 5375 9725 5406 4 vdd
rlabel metal1 s 19061 754 19450 785 4 vdd
rlabel metal1 s 1167 17694 1556 17725 4 vdd
rlabel metal1 s 18672 19235 19061 19266 4 vdd
rlabel metal1 s 14782 9994 15171 10025 4 vdd
rlabel metal1 s 778 23855 1167 23886 4 vdd
rlabel metal1 s 23340 11534 23729 11565 4 vdd
rlabel metal1 s 7002 16155 7391 16186 4 vdd
rlabel metal1 s 24118 8454 24507 8485 4 vdd
rlabel metal1 s 7391 22314 7780 22345 4 vdd
rlabel metal1 s 778 2295 1167 2326 4 vdd
rlabel metal1 s 20228 13075 20617 13106 4 vdd
rlabel metal1 s 14782 3834 15171 3865 4 vdd
rlabel metal1 s 6613 20774 7002 20805 4 vdd
rlabel metal1 s 17116 19234 17505 19265 4 vdd
rlabel metal1 s 18283 2295 18672 2326 4 vdd
rlabel metal1 s 1167 5374 1556 5405 4 vdd
rlabel metal1 s 15171 8455 15560 8486 4 vdd
rlabel metal1 s 20228 8455 20617 8486 4 vdd
rlabel metal1 s 21006 19234 21395 19265 4 vdd
rlabel metal1 s 7780 14615 8169 14646 4 vdd
rlabel metal1 s 9336 13075 9725 13106 4 vdd
rlabel metal1 s 1556 16154 1945 16185 4 vdd
rlabel metal1 s 22562 2294 22951 2325 4 vdd
rlabel metal1 s 6613 16155 7002 16186 4 vdd
rlabel metal1 s 21395 17695 21784 17726 4 vdd
rlabel metal1 s 11281 14615 11670 14646 4 vdd
rlabel metal1 s 22173 11534 22562 11565 4 vdd
rlabel metal1 s 1167 13074 1556 13105 4 vdd
rlabel metal1 s 5446 19234 5835 19265 4 vdd
rlabel metal1 s 17505 23855 17894 23886 4 vdd
rlabel metal1 s 778 20775 1167 20806 4 vdd
rlabel metal1 s 9725 20774 10114 20805 4 vdd
rlabel metal1 s 389 6915 778 6946 4 vdd
rlabel metal1 s 1167 8455 1556 8486 4 vdd
rlabel metal1 s 19450 13074 19839 13105 4 vdd
rlabel metal1 s 5446 8455 5835 8486 4 vdd
rlabel metal1 s 10114 20775 10503 20806 4 vdd
rlabel metal1 s 15171 14614 15560 14645 4 vdd
rlabel metal1 s 6613 6914 7002 6945 4 vdd
rlabel metal1 s 19061 22314 19450 22345 4 vdd
rlabel metal1 s 3501 3835 3890 3866 4 vdd
rlabel metal1 s 24118 5374 24507 5405 4 vdd
rlabel metal1 s 19839 9995 20228 10026 4 vdd
rlabel metal1 s 13615 8454 14004 8485 4 vdd
rlabel metal1 s 10892 8454 11281 8485 4 vdd
rlabel metal1 s 17116 14614 17505 14645 4 vdd
rlabel metal1 s 14004 20774 14393 20805 4 vdd
rlabel metal1 s 22173 3834 22562 3865 4 vdd
rlabel metal1 s 6613 3834 7002 3865 4 vdd
rlabel metal1 s 4668 14614 5057 14645 4 vdd
rlabel metal1 s 4279 17695 4668 17726 4 vdd
rlabel metal1 s 1945 6915 2334 6946 4 vdd
rlabel metal1 s 24507 14614 24896 14645 4 vdd
rlabel metal1 s 22173 22315 22562 22346 4 vdd
rlabel metal1 s 9336 17694 9725 17725 4 vdd
rlabel metal1 s 8169 5375 8558 5406 4 vdd
rlabel metal1 s 15560 23854 15949 23885 4 vdd
rlabel metal1 s 18283 17694 18672 17725 4 vdd
rlabel metal1 s 11670 13075 12059 13106 4 vdd
rlabel metal1 s 15171 9994 15560 10025 4 vdd
rlabel metal1 s 21006 20775 21395 20806 4 vdd
rlabel metal1 s 3890 2294 4279 2325 4 vdd
rlabel metal1 s 22173 22314 22562 22345 4 vdd
rlabel metal1 s 19450 17694 19839 17725 4 vdd
rlabel metal1 s 2334 22314 2723 22345 4 vdd
rlabel metal1 s 6613 13074 7002 13105 4 vdd
rlabel metal1 s 22562 17695 22951 17726 4 vdd
rlabel metal1 s 3501 5375 3890 5406 4 vdd
rlabel metal1 s 6613 2294 7002 2325 4 vdd
rlabel metal1 s 11281 8454 11670 8485 4 vdd
rlabel metal1 s 10503 6914 10892 6945 4 vdd
rlabel metal1 s 13226 754 13615 785 4 vdd
rlabel metal1 s 16727 19235 17116 19266 4 vdd
rlabel metal1 s 10503 20775 10892 20806 4 vdd
rlabel metal1 s 10503 9994 10892 10025 4 vdd
rlabel metal1 s 4279 16155 4668 16186 4 vdd
rlabel metal1 s 19839 16155 20228 16186 4 vdd
rlabel metal1 s 7002 17695 7391 17726 4 vdd
rlabel metal1 s 22562 3835 22951 3866 4 vdd
rlabel metal1 s 19450 6915 19839 6946 4 vdd
rlabel metal1 s 14004 8455 14393 8486 4 vdd
rlabel metal1 s 11670 9994 12059 10025 4 vdd
rlabel metal1 s 15560 16155 15949 16186 4 vdd
rlabel metal1 s 9336 20775 9725 20806 4 vdd
rlabel metal1 s 14004 22314 14393 22345 4 vdd
rlabel metal1 s 14004 2295 14393 2326 4 vdd
rlabel metal1 s 389 9995 778 10026 4 vdd
rlabel metal1 s 22173 5375 22562 5406 4 vdd
rlabel metal1 s 21395 19235 21784 19266 4 vdd
rlabel metal1 s 19061 16154 19450 16185 4 vdd
rlabel metal1 s 20617 16154 21006 16185 4 vdd
rlabel metal1 s 17505 16155 17894 16186 4 vdd
rlabel metal1 s 11281 13074 11670 13105 4 vdd
rlabel metal1 s 18283 19235 18672 19266 4 vdd
rlabel metal1 s 17116 3835 17505 3866 4 vdd
rlabel metal1 s 22562 754 22951 785 4 vdd
rlabel metal1 s 8947 16155 9336 16186 4 vdd
rlabel metal1 s 16727 755 17116 786 4 vdd
rlabel metal1 s 19839 17694 20228 17725 4 vdd
rlabel metal1 s 5057 6914 5446 6945 4 vdd
rlabel metal1 s 19450 755 19839 786 4 vdd
rlabel metal1 s 19450 19234 19839 19265 4 vdd
rlabel metal1 s 18283 23855 18672 23886 4 vdd
rlabel metal1 s 13226 16154 13615 16185 4 vdd
rlabel metal1 s 1945 19235 2334 19266 4 vdd
rlabel metal1 s 1945 13074 2334 13105 4 vdd
rlabel metal1 s 15171 6914 15560 6945 4 vdd
rlabel metal1 s 21784 17694 22173 17725 4 vdd
rlabel metal1 s 5057 17694 5446 17725 4 vdd
rlabel metal1 s 389 9994 778 10025 4 vdd
rlabel metal1 s 3890 9994 4279 10025 4 vdd
rlabel metal1 s 778 3834 1167 3865 4 vdd
rlabel metal1 s 12837 3835 13226 3866 4 vdd
rlabel metal1 s 20228 755 20617 786 4 vdd
rlabel metal1 s 18672 6915 19061 6946 4 vdd
rlabel metal1 s 16727 6915 17116 6946 4 vdd
rlabel metal1 s 10892 14614 11281 14645 4 vdd
rlabel metal1 s 10114 8455 10503 8486 4 vdd
rlabel metal1 s 22951 6915 23340 6946 4 vdd
rlabel metal1 s 7002 755 7391 786 4 vdd
rlabel metal1 s 7391 5374 7780 5405 4 vdd
rlabel metal1 s 4668 14615 5057 14646 4 vdd
rlabel metal1 s 16338 754 16727 785 4 vdd
rlabel metal1 s 24507 17695 24896 17726 4 vdd
rlabel metal1 s 5835 5375 6224 5406 4 vdd
rlabel metal1 s 15949 3835 16338 3866 4 vdd
rlabel metal1 s 21784 17695 22173 17726 4 vdd
rlabel metal1 s 8558 13074 8947 13105 4 vdd
rlabel metal1 s 0 16155 389 16186 4 vdd
rlabel metal1 s 12059 8454 12448 8485 4 vdd
rlabel metal1 s 19839 8455 20228 8486 4 vdd
rlabel metal1 s 21006 23855 21395 23886 4 vdd
rlabel metal1 s 7780 755 8169 786 4 vdd
rlabel metal1 s 12059 19235 12448 19266 4 vdd
rlabel metal1 s 7391 3835 7780 3866 4 vdd
rlabel metal1 s 5057 22314 5446 22345 4 vdd
rlabel metal1 s 22562 11534 22951 11565 4 vdd
rlabel metal1 s 14393 2295 14782 2326 4 vdd
rlabel metal1 s 20617 8455 21006 8486 4 vdd
rlabel metal1 s 23729 13074 24118 13105 4 vdd
rlabel metal1 s 4668 23855 5057 23886 4 vdd
rlabel metal1 s 24118 11535 24507 11566 4 vdd
rlabel metal1 s 1556 5374 1945 5405 4 vdd
rlabel metal1 s 3890 8455 4279 8486 4 vdd
rlabel metal1 s 778 6915 1167 6946 4 vdd
rlabel metal1 s 14393 23854 14782 23885 4 vdd
rlabel metal1 s 19061 6914 19450 6945 4 vdd
rlabel metal1 s 5835 6914 6224 6945 4 vdd
rlabel metal1 s 19450 16154 19839 16185 4 vdd
rlabel metal1 s 10892 23855 11281 23886 4 vdd
rlabel metal1 s 10892 3835 11281 3866 4 vdd
rlabel metal1 s 1167 2295 1556 2326 4 vdd
rlabel metal1 s 20228 2294 20617 2325 4 vdd
rlabel metal1 s 18672 9995 19061 10026 4 vdd
rlabel metal1 s 10503 14615 10892 14646 4 vdd
rlabel metal1 s 7391 13074 7780 13105 4 vdd
rlabel metal1 s 11670 16154 12059 16185 4 vdd
rlabel metal1 s 12448 17695 12837 17726 4 vdd
rlabel metal1 s 7780 17694 8169 17725 4 vdd
rlabel metal1 s 2723 2295 3112 2326 4 vdd
rlabel metal1 s 24118 9994 24507 10025 4 vdd
rlabel metal1 s 21006 755 21395 786 4 vdd
rlabel metal1 s 7002 9994 7391 10025 4 vdd
rlabel metal1 s 7002 2295 7391 2326 4 vdd
rlabel metal1 s 13615 23854 14004 23885 4 vdd
rlabel metal1 s 22951 3834 23340 3865 4 vdd
rlabel metal1 s 23729 8454 24118 8485 4 vdd
rlabel metal1 s 13615 19235 14004 19266 4 vdd
rlabel metal1 s 9336 11534 9725 11565 4 vdd
rlabel metal1 s 24507 11535 24896 11566 4 vdd
rlabel metal1 s 5446 14614 5835 14645 4 vdd
rlabel metal1 s 11281 6914 11670 6945 4 vdd
rlabel metal1 s 19061 5374 19450 5405 4 vdd
rlabel metal1 s 13615 755 14004 786 4 vdd
rlabel metal1 s 16727 14615 17116 14646 4 vdd
rlabel metal1 s 24118 20774 24507 20805 4 vdd
rlabel metal1 s 16727 23855 17116 23886 4 vdd
rlabel metal1 s 19061 13075 19450 13106 4 vdd
rlabel metal1 s 4668 17694 5057 17725 4 vdd
rlabel metal1 s 24118 3834 24507 3865 4 vdd
rlabel metal1 s 778 8454 1167 8485 4 vdd
rlabel metal1 s 1945 14614 2334 14645 4 vdd
rlabel metal1 s 17116 9995 17505 10026 4 vdd
rlabel metal1 s 21006 3834 21395 3865 4 vdd
rlabel metal1 s 21006 5375 21395 5406 4 vdd
rlabel metal1 s 15949 11534 16338 11565 4 vdd
rlabel metal1 s 21784 9994 22173 10025 4 vdd
rlabel metal1 s 23729 16154 24118 16185 4 vdd
rlabel metal1 s 18672 13075 19061 13106 4 vdd
rlabel metal1 s 10892 14615 11281 14646 4 vdd
rlabel metal1 s 7780 8455 8169 8486 4 vdd
rlabel metal1 s 13615 6915 14004 6946 4 vdd
rlabel metal1 s 8558 14615 8947 14646 4 vdd
rlabel metal1 s 3501 9994 3890 10025 4 vdd
rlabel metal1 s 4279 9994 4668 10025 4 vdd
rlabel metal1 s 12059 2294 12448 2325 4 vdd
rlabel metal1 s 5835 19234 6224 19265 4 vdd
rlabel metal1 s 7391 19234 7780 19265 4 vdd
rlabel metal1 s 2723 9994 3112 10025 4 vdd
rlabel metal1 s 3112 6914 3501 6945 4 vdd
rlabel metal1 s 8947 16154 9336 16185 4 vdd
rlabel metal1 s 1167 6914 1556 6945 4 vdd
rlabel metal1 s 19839 17695 20228 17726 4 vdd
rlabel metal1 s 21006 23854 21395 23885 4 vdd
rlabel metal1 s 10892 23854 11281 23885 4 vdd
rlabel metal1 s 22951 22315 23340 22346 4 vdd
rlabel metal1 s 0 23854 389 23885 4 vdd
rlabel metal1 s 17505 8454 17894 8485 4 vdd
rlabel metal1 s 5057 6915 5446 6946 4 vdd
rlabel metal1 s 3501 14615 3890 14646 4 vdd
rlabel metal1 s 16338 17694 16727 17725 4 vdd
rlabel metal1 s 5835 17695 6224 17726 4 vdd
rlabel metal1 s 778 22314 1167 22345 4 vdd
rlabel metal1 s 23340 11535 23729 11566 4 vdd
rlabel metal1 s 1945 9994 2334 10025 4 vdd
rlabel metal1 s 19839 3835 20228 3866 4 vdd
rlabel metal1 s 11281 13075 11670 13106 4 vdd
rlabel metal1 s 13226 9994 13615 10025 4 vdd
rlabel metal1 s 10114 11535 10503 11566 4 vdd
rlabel metal1 s 12059 19234 12448 19265 4 vdd
rlabel metal1 s 15949 8454 16338 8485 4 vdd
rlabel metal1 s 7780 6915 8169 6946 4 vdd
rlabel metal1 s 21006 5374 21395 5405 4 vdd
rlabel metal1 s 16338 11534 16727 11565 4 vdd
rlabel metal1 s 23729 5375 24118 5406 4 vdd
rlabel metal1 s 23340 5374 23729 5405 4 vdd
rlabel metal1 s 15949 6914 16338 6945 4 vdd
rlabel metal1 s 10892 19235 11281 19266 4 vdd
rlabel metal1 s 15171 3835 15560 3866 4 vdd
rlabel metal1 s 4279 23855 4668 23886 4 vdd
rlabel metal1 s 12448 22315 12837 22346 4 vdd
rlabel metal1 s 24507 19234 24896 19265 4 vdd
rlabel metal1 s 22562 9994 22951 10025 4 vdd
rlabel metal1 s 10892 8455 11281 8486 4 vdd
rlabel metal1 s 3501 22314 3890 22345 4 vdd
rlabel metal1 s 22951 8454 23340 8485 4 vdd
rlabel metal1 s 1556 6914 1945 6945 4 vdd
rlabel metal1 s 17116 754 17505 785 4 vdd
rlabel metal1 s 18672 2294 19061 2325 4 vdd
rlabel metal1 s 7780 11535 8169 11566 4 vdd
rlabel metal1 s 389 13074 778 13105 4 vdd
rlabel metal1 s 9336 9994 9725 10025 4 vdd
rlabel metal1 s 7002 13074 7391 13105 4 vdd
rlabel metal1 s 23729 14614 24118 14645 4 vdd
rlabel metal1 s 18672 17694 19061 17725 4 vdd
rlabel metal1 s 14004 6914 14393 6945 4 vdd
rlabel metal1 s 10114 20774 10503 20805 4 vdd
rlabel metal1 s 11281 23854 11670 23885 4 vdd
rlabel metal1 s 14004 11534 14393 11565 4 vdd
rlabel metal1 s 15560 19235 15949 19266 4 vdd
rlabel metal1 s 18672 6914 19061 6945 4 vdd
rlabel metal1 s 4668 19235 5057 19266 4 vdd
rlabel metal1 s 1556 22314 1945 22345 4 vdd
rlabel metal1 s 7002 23855 7391 23886 4 vdd
rlabel metal1 s 13615 11534 14004 11565 4 vdd
rlabel metal1 s 19450 11535 19839 11566 4 vdd
rlabel metal1 s 22173 9994 22562 10025 4 vdd
rlabel metal1 s 10892 9994 11281 10025 4 vdd
rlabel metal1 s 17116 11535 17505 11566 4 vdd
rlabel metal1 s 17894 9994 18283 10025 4 vdd
rlabel metal1 s 2334 9994 2723 10025 4 vdd
rlabel metal1 s 2334 14614 2723 14645 4 vdd
rlabel metal1 s 17116 22315 17505 22346 4 vdd
rlabel metal1 s 2723 6915 3112 6946 4 vdd
rlabel metal1 s 15171 9995 15560 10026 4 vdd
rlabel metal1 s 8169 16154 8558 16185 4 vdd
rlabel metal1 s 22173 23855 22562 23886 4 vdd
rlabel metal1 s 8169 2294 8558 2325 4 vdd
rlabel metal1 s 19839 6914 20228 6945 4 vdd
rlabel metal1 s 21395 3835 21784 3866 4 vdd
rlabel metal1 s 778 17695 1167 17726 4 vdd
rlabel metal1 s 18672 23854 19061 23885 4 vdd
rlabel metal1 s 10114 22314 10503 22345 4 vdd
rlabel metal1 s 14782 11535 15171 11566 4 vdd
rlabel metal1 s 7391 17695 7780 17726 4 vdd
rlabel metal1 s 15949 3834 16338 3865 4 vdd
rlabel metal1 s 16727 20774 17116 20805 4 vdd
rlabel metal1 s 13615 3834 14004 3865 4 vdd
rlabel metal1 s 22562 14614 22951 14645 4 vdd
rlabel metal1 s 12837 2294 13226 2325 4 vdd
rlabel metal1 s 18672 2295 19061 2326 4 vdd
rlabel metal1 s 389 23854 778 23885 4 vdd
rlabel metal1 s 5446 6915 5835 6946 4 vdd
rlabel metal1 s 20617 9995 21006 10026 4 vdd
rlabel metal1 s 19450 22315 19839 22346 4 vdd
rlabel metal1 s 6224 3835 6613 3866 4 vdd
rlabel metal1 s 22562 22315 22951 22346 4 vdd
rlabel metal1 s 7780 20774 8169 20805 4 vdd
rlabel metal1 s 8169 13075 8558 13106 4 vdd
rlabel metal1 s 14782 2294 15171 2325 4 vdd
rlabel metal1 s 3890 754 4279 785 4 vdd
rlabel metal1 s 3501 11534 3890 11565 4 vdd
rlabel metal1 s 8169 19235 8558 19266 4 vdd
rlabel metal1 s 2723 11534 3112 11565 4 vdd
rlabel metal1 s 19061 19234 19450 19265 4 vdd
rlabel metal1 s 19450 14615 19839 14646 4 vdd
rlabel metal1 s 7780 11534 8169 11565 4 vdd
rlabel metal1 s 11670 6914 12059 6945 4 vdd
rlabel metal1 s 1945 754 2334 785 4 vdd
rlabel metal1 s 8947 20774 9336 20805 4 vdd
rlabel metal1 s 7002 23854 7391 23885 4 vdd
rlabel metal1 s 16338 20774 16727 20805 4 vdd
rlabel metal1 s 8558 17694 8947 17725 4 vdd
rlabel metal1 s 13226 17695 13615 17726 4 vdd
rlabel metal1 s 21784 754 22173 785 4 vdd
rlabel metal1 s 8947 2295 9336 2326 4 vdd
rlabel metal1 s 6224 2295 6613 2326 4 vdd
rlabel metal1 s 15171 11534 15560 11565 4 vdd
rlabel metal1 s 12837 16154 13226 16185 4 vdd
rlabel metal1 s 19839 2294 20228 2325 4 vdd
rlabel metal1 s 6613 8454 7002 8485 4 vdd
rlabel metal1 s 14393 5375 14782 5406 4 vdd
rlabel metal1 s 3890 5374 4279 5405 4 vdd
rlabel metal1 s 6613 19235 7002 19266 4 vdd
rlabel metal1 s 10503 16155 10892 16186 4 vdd
rlabel metal1 s 2334 9995 2723 10026 4 vdd
rlabel metal1 s 17894 14615 18283 14646 4 vdd
rlabel metal1 s 14393 11534 14782 11565 4 vdd
rlabel metal1 s 21784 16155 22173 16186 4 vdd
rlabel metal1 s 24118 16155 24507 16186 4 vdd
rlabel metal1 s 778 13075 1167 13106 4 vdd
rlabel metal1 s 13615 6914 14004 6945 4 vdd
rlabel metal1 s 2334 23854 2723 23885 4 vdd
rlabel metal1 s 3501 5374 3890 5405 4 vdd
rlabel metal1 s 21006 9995 21395 10026 4 vdd
rlabel metal1 s 11670 14614 12059 14645 4 vdd
rlabel metal1 s 8169 5374 8558 5405 4 vdd
rlabel metal1 s 18283 5374 18672 5405 4 vdd
rlabel metal1 s 8947 22314 9336 22345 4 vdd
rlabel metal1 s 8169 8455 8558 8486 4 vdd
rlabel metal1 s 22562 6915 22951 6946 4 vdd
rlabel metal1 s 12448 13074 12837 13105 4 vdd
rlabel metal1 s 22951 2295 23340 2326 4 vdd
rlabel metal1 s 15560 20775 15949 20806 4 vdd
rlabel metal1 s 15949 17694 16338 17725 4 vdd
rlabel metal1 s 11670 19234 12059 19265 4 vdd
rlabel metal1 s 16338 13074 16727 13105 4 vdd
rlabel metal1 s 8169 17695 8558 17726 4 vdd
rlabel metal1 s 1167 19235 1556 19266 4 vdd
rlabel metal1 s 12059 6914 12448 6945 4 vdd
rlabel metal1 s 6224 13075 6613 13106 4 vdd
rlabel metal1 s 2334 11534 2723 11565 4 vdd
rlabel metal1 s 1167 17695 1556 17726 4 vdd
rlabel metal1 s 23729 755 24118 786 4 vdd
rlabel metal1 s 1945 755 2334 786 4 vdd
rlabel metal1 s 21784 2294 22173 2325 4 vdd
rlabel metal1 s 8947 11535 9336 11566 4 vdd
rlabel metal1 s 12837 5374 13226 5405 4 vdd
rlabel metal1 s 5057 2295 5446 2326 4 vdd
rlabel metal1 s 12059 22314 12448 22345 4 vdd
rlabel metal1 s 21395 19234 21784 19265 4 vdd
rlabel metal1 s 6224 20774 6613 20805 4 vdd
rlabel metal1 s 18283 22314 18672 22345 4 vdd
rlabel metal1 s 10114 9995 10503 10026 4 vdd
rlabel metal1 s 9336 11535 9725 11566 4 vdd
rlabel metal1 s 17894 5375 18283 5406 4 vdd
rlabel metal1 s 6613 22315 7002 22346 4 vdd
rlabel metal1 s 8558 22315 8947 22346 4 vdd
rlabel metal1 s 17116 6915 17505 6946 4 vdd
rlabel metal1 s 21784 16154 22173 16185 4 vdd
rlabel metal1 s 1945 17695 2334 17726 4 vdd
rlabel metal1 s 17894 22315 18283 22346 4 vdd
rlabel metal1 s 23729 2295 24118 2326 4 vdd
rlabel metal1 s 18672 9994 19061 10025 4 vdd
rlabel metal1 s 23729 11535 24118 11566 4 vdd
rlabel metal1 s 21784 9995 22173 10026 4 vdd
rlabel metal1 s 5057 16155 5446 16186 4 vdd
rlabel metal1 s 5835 20774 6224 20805 4 vdd
rlabel metal1 s 18283 755 18672 786 4 vdd
rlabel metal1 s 2334 8454 2723 8485 4 vdd
rlabel metal1 s 12448 19234 12837 19265 4 vdd
rlabel metal1 s 22951 19234 23340 19265 4 vdd
rlabel metal1 s 14393 17694 14782 17725 4 vdd
rlabel metal1 s 3890 2295 4279 2326 4 vdd
rlabel metal1 s 20617 23855 21006 23886 4 vdd
rlabel metal1 s 23340 22314 23729 22345 4 vdd
rlabel metal1 s 17894 2294 18283 2325 4 vdd
rlabel metal1 s 1167 11534 1556 11565 4 vdd
rlabel metal1 s 5835 11534 6224 11565 4 vdd
rlabel metal1 s 10114 5375 10503 5406 4 vdd
rlabel metal1 s 14004 13074 14393 13105 4 vdd
rlabel metal1 s 1167 11535 1556 11566 4 vdd
rlabel metal1 s 10114 23854 10503 23885 4 vdd
rlabel metal1 s 19061 9995 19450 10026 4 vdd
rlabel metal1 s 16338 19234 16727 19265 4 vdd
rlabel metal1 s 6613 20775 7002 20806 4 vdd
rlabel metal1 s 4279 754 4668 785 4 vdd
rlabel metal1 s 14782 5375 15171 5406 4 vdd
rlabel metal1 s 2723 8455 3112 8486 4 vdd
rlabel metal1 s 15949 22314 16338 22345 4 vdd
rlabel metal1 s 21395 22314 21784 22345 4 vdd
rlabel metal1 s 5835 9994 6224 10025 4 vdd
rlabel metal1 s 2723 17695 3112 17726 4 vdd
rlabel metal1 s 21006 17694 21395 17725 4 vdd
rlabel metal1 s 7391 14614 7780 14645 4 vdd
rlabel metal1 s 13226 11534 13615 11565 4 vdd
rlabel metal1 s 8947 13075 9336 13106 4 vdd
rlabel metal1 s 22951 3835 23340 3866 4 vdd
rlabel metal1 s 3112 19234 3501 19265 4 vdd
rlabel metal1 s 12837 20775 13226 20806 4 vdd
rlabel metal1 s 6613 17694 7002 17725 4 vdd
rlabel metal1 s 11670 22315 12059 22346 4 vdd
rlabel metal1 s 18672 11534 19061 11565 4 vdd
rlabel metal1 s 5835 6915 6224 6946 4 vdd
rlabel metal1 s 21395 8455 21784 8486 4 vdd
rlabel metal1 s 18283 23854 18672 23885 4 vdd
rlabel metal1 s 24118 13074 24507 13105 4 vdd
rlabel metal1 s 15560 2294 15949 2325 4 vdd
rlabel metal1 s 20228 9994 20617 10025 4 vdd
rlabel metal1 s 10892 20774 11281 20805 4 vdd
rlabel metal1 s 5446 9995 5835 10026 4 vdd
rlabel metal1 s 11281 17694 11670 17725 4 vdd
rlabel metal1 s 17894 755 18283 786 4 vdd
rlabel metal1 s 24507 9995 24896 10026 4 vdd
rlabel metal1 s 389 20774 778 20805 4 vdd
rlabel metal1 s 1167 23855 1556 23886 4 vdd
rlabel metal1 s 20617 754 21006 785 4 vdd
rlabel metal1 s 11670 13074 12059 13105 4 vdd
rlabel metal1 s 0 16154 389 16185 4 vdd
rlabel metal1 s 1945 9995 2334 10026 4 vdd
rlabel metal1 s 1167 8454 1556 8485 4 vdd
rlabel metal1 s 4668 6914 5057 6945 4 vdd
rlabel metal1 s 17894 8454 18283 8485 4 vdd
rlabel metal1 s 18672 23855 19061 23886 4 vdd
rlabel metal1 s 5057 22315 5446 22346 4 vdd
rlabel metal1 s 19061 14615 19450 14646 4 vdd
rlabel metal1 s 16338 17695 16727 17726 4 vdd
rlabel metal1 s 389 5374 778 5405 4 vdd
rlabel metal1 s 13615 2294 14004 2325 4 vdd
rlabel metal1 s 11281 3835 11670 3866 4 vdd
rlabel metal1 s 3112 6915 3501 6946 4 vdd
rlabel metal1 s 5835 13075 6224 13106 4 vdd
rlabel metal1 s 5446 13074 5835 13105 4 vdd
rlabel metal1 s 15560 14614 15949 14645 4 vdd
rlabel metal1 s 18672 8454 19061 8485 4 vdd
rlabel metal1 s 17894 13075 18283 13106 4 vdd
rlabel metal1 s 1556 754 1945 785 4 vdd
rlabel metal1 s 12448 19235 12837 19266 4 vdd
rlabel metal1 s 12059 14615 12448 14646 4 vdd
rlabel metal1 s 23340 22315 23729 22346 4 vdd
rlabel metal1 s 17116 9994 17505 10025 4 vdd
rlabel metal1 s 5446 754 5835 785 4 vdd
rlabel metal1 s 9336 14614 9725 14645 4 vdd
rlabel metal1 s 12837 16155 13226 16186 4 vdd
rlabel metal1 s 10892 11535 11281 11566 4 vdd
rlabel metal1 s 7002 22314 7391 22345 4 vdd
rlabel metal1 s 0 11534 389 11565 4 vdd
rlabel metal1 s 15560 16154 15949 16185 4 vdd
rlabel metal1 s 15949 20774 16338 20805 4 vdd
rlabel metal1 s 13615 17695 14004 17726 4 vdd
rlabel metal1 s 7002 19234 7391 19265 4 vdd
rlabel metal1 s 19450 13075 19839 13106 4 vdd
rlabel metal1 s 10114 22315 10503 22346 4 vdd
rlabel metal1 s 20617 14615 21006 14646 4 vdd
rlabel metal1 s 13615 20774 14004 20805 4 vdd
rlabel metal1 s 20617 6914 21006 6945 4 vdd
rlabel metal1 s 12837 3834 13226 3865 4 vdd
rlabel metal1 s 10892 17695 11281 17726 4 vdd
rlabel metal1 s 12448 23854 12837 23885 4 vdd
rlabel metal1 s 18672 11535 19061 11566 4 vdd
rlabel metal1 s 20228 2295 20617 2326 4 vdd
rlabel metal1 s 8947 22315 9336 22346 4 vdd
rlabel metal1 s 12837 22315 13226 22346 4 vdd
rlabel metal1 s 17116 2294 17505 2325 4 vdd
rlabel metal1 s 21784 11535 22173 11566 4 vdd
rlabel metal1 s 16727 20775 17116 20806 4 vdd
rlabel metal1 s 24507 13075 24896 13106 4 vdd
rlabel metal1 s 778 754 1167 785 4 vdd
rlabel metal1 s 12448 8455 12837 8486 4 vdd
rlabel metal1 s 5446 11535 5835 11566 4 vdd
rlabel metal1 s 3112 22315 3501 22346 4 vdd
rlabel metal1 s 21006 13075 21395 13106 4 vdd
rlabel metal1 s 22951 11534 23340 11565 4 vdd
rlabel metal1 s 14393 9994 14782 10025 4 vdd
rlabel metal1 s 3112 2294 3501 2325 4 vdd
rlabel metal1 s 23340 16154 23729 16185 4 vdd
rlabel metal1 s 19450 5375 19839 5406 4 vdd
rlabel metal1 s 20228 19234 20617 19265 4 vdd
rlabel metal1 s 12059 5374 12448 5405 4 vdd
rlabel metal1 s 6224 755 6613 786 4 vdd
rlabel metal1 s 778 11534 1167 11565 4 vdd
rlabel metal1 s 2723 6914 3112 6945 4 vdd
rlabel metal1 s 21006 16154 21395 16185 4 vdd
rlabel metal1 s 11670 755 12059 786 4 vdd
rlabel metal1 s 8558 9995 8947 10026 4 vdd
rlabel metal1 s 2334 2294 2723 2325 4 vdd
rlabel metal1 s 2334 23855 2723 23886 4 vdd
rlabel metal1 s 12059 8455 12448 8486 4 vdd
rlabel metal1 s 23340 19235 23729 19266 4 vdd
rlabel metal1 s 22173 6914 22562 6945 4 vdd
rlabel metal1 s 14782 14615 15171 14646 4 vdd
rlabel metal1 s 1167 2294 1556 2325 4 vdd
rlabel metal1 s 6224 8454 6613 8485 4 vdd
rlabel metal1 s 17894 8455 18283 8486 4 vdd
rlabel metal1 s 14393 754 14782 785 4 vdd
rlabel metal1 s 4668 754 5057 785 4 vdd
rlabel metal1 s 8947 755 9336 786 4 vdd
rlabel metal1 s 8947 23855 9336 23886 4 vdd
rlabel metal1 s 7780 3834 8169 3865 4 vdd
rlabel metal1 s 3112 5374 3501 5405 4 vdd
rlabel metal1 s 18672 22314 19061 22345 4 vdd
rlabel metal1 s 12059 16154 12448 16185 4 vdd
rlabel metal1 s 12448 9994 12837 10025 4 vdd
rlabel metal1 s 19450 2295 19839 2326 4 vdd
rlabel metal1 s 3112 11534 3501 11565 4 vdd
rlabel metal1 s 4668 16154 5057 16185 4 vdd
rlabel metal1 s 4668 8455 5057 8486 4 vdd
rlabel metal1 s 21395 14615 21784 14646 4 vdd
rlabel metal1 s 16727 17694 17116 17725 4 vdd
rlabel metal1 s 15949 17695 16338 17726 4 vdd
rlabel metal1 s 7780 6914 8169 6945 4 vdd
rlabel metal1 s 1556 16155 1945 16186 4 vdd
rlabel metal1 s 1167 16155 1556 16186 4 vdd
rlabel metal1 s 13226 3835 13615 3866 4 vdd
rlabel metal1 s 5057 9995 5446 10026 4 vdd
rlabel metal1 s 21784 5374 22173 5405 4 vdd
rlabel metal1 s 11670 16155 12059 16186 4 vdd
rlabel metal1 s 12059 22315 12448 22346 4 vdd
rlabel metal1 s 16338 16155 16727 16186 4 vdd
rlabel metal1 s 3890 16155 4279 16186 4 vdd
rlabel metal1 s 22173 2294 22562 2325 4 vdd
rlabel metal1 s 778 5374 1167 5405 4 vdd
rlabel metal1 s 20617 2295 21006 2326 4 vdd
rlabel metal1 s 14782 14614 15171 14645 4 vdd
rlabel metal1 s 778 755 1167 786 4 vdd
rlabel metal1 s 23340 13075 23729 13106 4 vdd
rlabel metal1 s 24118 754 24507 785 4 vdd
rlabel metal1 s 20617 6915 21006 6946 4 vdd
rlabel metal1 s 8947 17695 9336 17726 4 vdd
rlabel metal1 s 18672 13074 19061 13105 4 vdd
rlabel metal1 s 17505 6914 17894 6945 4 vdd
rlabel metal1 s 1556 6915 1945 6946 4 vdd
rlabel metal1 s 21006 6915 21395 6946 4 vdd
rlabel metal1 s 13226 16155 13615 16186 4 vdd
rlabel metal1 s 4279 14615 4668 14646 4 vdd
rlabel metal1 s 20228 11534 20617 11565 4 vdd
rlabel metal1 s 8558 11535 8947 11566 4 vdd
rlabel metal1 s 14004 16154 14393 16185 4 vdd
rlabel metal1 s 9725 17695 10114 17726 4 vdd
rlabel metal1 s 5446 16154 5835 16185 4 vdd
rlabel metal1 s 21395 6915 21784 6946 4 vdd
rlabel metal1 s 12837 13074 13226 13105 4 vdd
rlabel metal1 s 21006 8454 21395 8485 4 vdd
rlabel metal1 s 20617 3835 21006 3866 4 vdd
rlabel metal1 s 11281 17695 11670 17726 4 vdd
rlabel metal1 s 12837 11535 13226 11566 4 vdd
rlabel metal1 s 2723 13074 3112 13105 4 vdd
rlabel metal1 s 3501 754 3890 785 4 vdd
rlabel metal1 s 10114 17694 10503 17725 4 vdd
rlabel metal1 s 3501 17695 3890 17726 4 vdd
rlabel metal1 s 17116 755 17505 786 4 vdd
rlabel metal1 s 18283 8454 18672 8485 4 vdd
rlabel metal1 s 16727 22315 17116 22346 4 vdd
rlabel metal1 s 15949 11535 16338 11566 4 vdd
rlabel metal1 s 24118 19234 24507 19265 4 vdd
rlabel metal1 s 14393 16154 14782 16185 4 vdd
rlabel metal1 s 13615 3835 14004 3866 4 vdd
rlabel metal1 s 24118 9995 24507 10026 4 vdd
rlabel metal1 s 12059 14614 12448 14645 4 vdd
rlabel metal1 s 17894 17695 18283 17726 4 vdd
rlabel metal1 s 12837 9995 13226 10026 4 vdd
rlabel metal1 s 4279 20774 4668 20805 4 vdd
rlabel metal1 s 22951 17695 23340 17726 4 vdd
rlabel metal1 s 19839 8454 20228 8485 4 vdd
rlabel metal1 s 24507 5374 24896 5405 4 vdd
rlabel metal1 s 1167 9994 1556 10025 4 vdd
rlabel metal1 s 3112 2295 3501 2326 4 vdd
rlabel metal1 s 0 9994 389 10025 4 vdd
rlabel metal1 s 9725 9995 10114 10026 4 vdd
rlabel metal1 s 17894 19235 18283 19266 4 vdd
rlabel metal1 s 1167 22315 1556 22346 4 vdd
rlabel metal1 s 13226 22315 13615 22346 4 vdd
rlabel metal1 s 9725 8454 10114 8485 4 vdd
rlabel metal1 s 15949 9995 16338 10026 4 vdd
rlabel metal1 s 10892 16155 11281 16186 4 vdd
rlabel metal1 s 15560 13075 15949 13106 4 vdd
rlabel metal1 s 19061 5375 19450 5406 4 vdd
rlabel metal1 s 9725 13074 10114 13105 4 vdd
rlabel metal1 s 2334 755 2723 786 4 vdd
rlabel metal1 s 17505 6915 17894 6946 4 vdd
rlabel metal1 s 21395 2294 21784 2325 4 vdd
rlabel metal1 s 12059 755 12448 786 4 vdd
rlabel metal1 s 17116 13075 17505 13106 4 vdd
rlabel metal1 s 2334 19235 2723 19266 4 vdd
rlabel metal1 s 15171 8454 15560 8485 4 vdd
rlabel metal1 s 17894 22314 18283 22345 4 vdd
rlabel metal1 s 389 22314 778 22345 4 vdd
rlabel metal1 s 9725 17694 10114 17725 4 vdd
rlabel metal1 s 13615 16155 14004 16186 4 vdd
rlabel metal1 s 23340 6914 23729 6945 4 vdd
rlabel metal1 s 5446 22314 5835 22345 4 vdd
rlabel metal1 s 20617 5374 21006 5405 4 vdd
rlabel metal1 s 18672 16154 19061 16185 4 vdd
rlabel metal1 s 4279 17694 4668 17725 4 vdd
rlabel metal1 s 15949 16154 16338 16185 4 vdd
rlabel metal1 s 2723 8454 3112 8485 4 vdd
rlabel metal1 s 12837 6915 13226 6946 4 vdd
rlabel metal1 s 16338 8454 16727 8485 4 vdd
rlabel metal1 s 7002 8455 7391 8486 4 vdd
rlabel metal1 s 15560 11534 15949 11565 4 vdd
rlabel metal1 s 1945 5375 2334 5406 4 vdd
rlabel metal1 s 13226 13075 13615 13106 4 vdd
rlabel metal1 s 12059 754 12448 785 4 vdd
rlabel metal1 s 5446 11534 5835 11565 4 vdd
rlabel metal1 s 10503 23854 10892 23885 4 vdd
rlabel metal1 s 19061 755 19450 786 4 vdd
rlabel metal1 s 12448 6915 12837 6946 4 vdd
rlabel metal1 s 1167 23854 1556 23885 4 vdd
rlabel metal1 s 3890 3835 4279 3866 4 vdd
rlabel metal1 s 21784 2295 22173 2326 4 vdd
rlabel metal1 s 18283 17695 18672 17726 4 vdd
rlabel metal1 s 11670 17695 12059 17726 4 vdd
rlabel metal1 s 15171 22315 15560 22346 4 vdd
rlabel metal1 s 14393 23855 14782 23886 4 vdd
rlabel metal1 s 24118 5375 24507 5406 4 vdd
rlabel metal1 s 14004 3834 14393 3865 4 vdd
rlabel metal1 s 2334 19234 2723 19265 4 vdd
rlabel metal1 s 16338 22314 16727 22345 4 vdd
rlabel metal1 s 20617 20774 21006 20805 4 vdd
rlabel metal1 s 15171 14615 15560 14646 4 vdd
rlabel metal1 s 389 16154 778 16185 4 vdd
rlabel metal1 s 3890 3834 4279 3865 4 vdd
rlabel metal1 s 15949 20775 16338 20806 4 vdd
rlabel metal1 s 8169 11534 8558 11565 4 vdd
rlabel metal1 s 1945 11535 2334 11566 4 vdd
rlabel metal1 s 389 11534 778 11565 4 vdd
rlabel metal1 s 5835 19235 6224 19266 4 vdd
rlabel metal1 s 5057 19234 5446 19265 4 vdd
rlabel metal1 s 5835 23854 6224 23885 4 vdd
rlabel metal1 s 22562 16154 22951 16185 4 vdd
rlabel metal1 s 10114 9994 10503 10025 4 vdd
rlabel metal1 s 10892 13075 11281 13106 4 vdd
rlabel metal1 s 17505 14614 17894 14645 4 vdd
rlabel metal1 s 7780 17695 8169 17726 4 vdd
rlabel metal1 s 14004 754 14393 785 4 vdd
rlabel metal1 s 4279 6914 4668 6945 4 vdd
rlabel metal1 s 4668 19234 5057 19265 4 vdd
rlabel metal1 s 3501 6915 3890 6946 4 vdd
rlabel metal1 s 0 2294 389 2325 4 vdd
rlabel metal1 s 6613 755 7002 786 4 vdd
rlabel metal1 s 9725 3834 10114 3865 4 vdd
rlabel metal1 s 3112 22314 3501 22345 4 vdd
rlabel metal1 s 24507 3835 24896 3866 4 vdd
rlabel metal1 s 12059 17694 12448 17725 4 vdd
rlabel metal1 s 13226 19234 13615 19265 4 vdd
rlabel metal1 s 14393 20774 14782 20805 4 vdd
rlabel metal1 s 4668 11534 5057 11565 4 vdd
rlabel metal1 s 11670 2294 12059 2325 4 vdd
rlabel metal1 s 1945 3834 2334 3865 4 vdd
rlabel metal1 s 1167 14614 1556 14645 4 vdd
rlabel metal1 s 0 23855 389 23886 4 vdd
rlabel metal1 s 0 19234 389 19265 4 vdd
rlabel metal1 s 22951 16154 23340 16185 4 vdd
rlabel metal1 s 15949 14614 16338 14645 4 vdd
rlabel metal1 s 5057 19235 5446 19266 4 vdd
rlabel metal1 s 23340 17694 23729 17725 4 vdd
rlabel metal1 s 10114 11534 10503 11565 4 vdd
rlabel metal1 s 20617 22315 21006 22346 4 vdd
rlabel metal1 s 13615 754 14004 785 4 vdd
rlabel metal1 s 3890 14615 4279 14646 4 vdd
rlabel metal1 s 16727 11535 17116 11566 4 vdd
rlabel metal1 s 12837 14615 13226 14646 4 vdd
rlabel metal1 s 18672 14615 19061 14646 4 vdd
rlabel metal1 s 14393 16155 14782 16186 4 vdd
rlabel metal1 s 19839 3834 20228 3865 4 vdd
rlabel metal1 s 14004 23854 14393 23885 4 vdd
rlabel metal1 s 15949 19234 16338 19265 4 vdd
rlabel metal1 s 18283 3834 18672 3865 4 vdd
rlabel metal1 s 23729 11534 24118 11565 4 vdd
rlabel metal1 s 3501 23854 3890 23885 4 vdd
rlabel metal1 s 15560 11535 15949 11566 4 vdd
rlabel metal1 s 4279 22314 4668 22345 4 vdd
rlabel metal1 s 23340 755 23729 786 4 vdd
rlabel metal1 s 14782 17694 15171 17725 4 vdd
rlabel metal1 s 3501 17694 3890 17725 4 vdd
rlabel metal1 s 13226 13074 13615 13105 4 vdd
rlabel metal1 s 2723 9995 3112 10026 4 vdd
rlabel metal1 s 5835 2295 6224 2326 4 vdd
rlabel metal1 s 8558 19234 8947 19265 4 vdd
rlabel metal1 s 20228 22314 20617 22345 4 vdd
rlabel metal1 s 23340 16155 23729 16186 4 vdd
rlabel metal1 s 6224 9994 6613 10025 4 vdd
rlabel metal1 s 10114 2295 10503 2326 4 vdd
rlabel metal1 s 14393 14614 14782 14645 4 vdd
rlabel metal1 s 15949 14615 16338 14646 4 vdd
rlabel metal1 s 3501 9995 3890 10026 4 vdd
rlabel metal1 s 23729 5374 24118 5405 4 vdd
rlabel metal1 s 17894 3835 18283 3866 4 vdd
rlabel metal1 s 19839 14615 20228 14646 4 vdd
rlabel metal1 s 1945 16155 2334 16186 4 vdd
rlabel metal1 s 21784 22315 22173 22346 4 vdd
rlabel metal1 s 8558 2294 8947 2325 4 vdd
rlabel metal1 s 12837 9994 13226 10025 4 vdd
rlabel metal1 s 20228 754 20617 785 4 vdd
rlabel metal1 s 14004 22315 14393 22346 4 vdd
rlabel metal1 s 13615 19234 14004 19265 4 vdd
rlabel metal1 s 2723 755 3112 786 4 vdd
rlabel metal1 s 16338 5375 16727 5406 4 vdd
rlabel metal1 s 10892 22314 11281 22345 4 vdd
rlabel metal1 s 22951 22314 23340 22345 4 vdd
rlabel metal1 s 778 6914 1167 6945 4 vdd
rlabel metal1 s 24507 755 24896 786 4 vdd
rlabel metal1 s 9336 23855 9725 23886 4 vdd
rlabel metal1 s 19839 5375 20228 5406 4 vdd
rlabel metal1 s 24118 23854 24507 23885 4 vdd
rlabel metal1 s 5446 17694 5835 17725 4 vdd
rlabel metal1 s 9725 11534 10114 11565 4 vdd
rlabel metal1 s 5057 14615 5446 14646 4 vdd
rlabel metal1 s 17894 20775 18283 20806 4 vdd
rlabel metal1 s 5057 5374 5446 5405 4 vdd
rlabel metal1 s 23729 17694 24118 17725 4 vdd
rlabel metal1 s 1945 22314 2334 22345 4 vdd
rlabel metal1 s 9336 19234 9725 19265 4 vdd
rlabel metal1 s 22951 20774 23340 20805 4 vdd
rlabel metal1 s 6224 23854 6613 23885 4 vdd
rlabel metal1 s 21395 20774 21784 20805 4 vdd
rlabel metal1 s 14782 13074 15171 13105 4 vdd
rlabel metal1 s 20617 8454 21006 8485 4 vdd
rlabel metal1 s 19839 11535 20228 11566 4 vdd
rlabel metal1 s 4279 3835 4668 3866 4 vdd
rlabel metal1 s 12448 3834 12837 3865 4 vdd
rlabel metal1 s 19839 11534 20228 11565 4 vdd
rlabel metal1 s 8558 2295 8947 2326 4 vdd
rlabel metal1 s 12059 6915 12448 6946 4 vdd
rlabel metal1 s 9725 5374 10114 5405 4 vdd
rlabel metal1 s 1945 14615 2334 14646 4 vdd
rlabel metal1 s 10892 20775 11281 20806 4 vdd
rlabel metal1 s 14782 9995 15171 10026 4 vdd
rlabel metal1 s 13615 11535 14004 11566 4 vdd
rlabel metal1 s 778 16155 1167 16186 4 vdd
rlabel metal1 s 24118 13075 24507 13106 4 vdd
rlabel metal1 s 12059 23854 12448 23885 4 vdd
rlabel metal1 s 21395 23855 21784 23886 4 vdd
rlabel metal1 s 12448 754 12837 785 4 vdd
rlabel metal1 s 18672 17695 19061 17726 4 vdd
rlabel metal1 s 19061 11535 19450 11566 4 vdd
rlabel metal1 s 8558 17695 8947 17726 4 vdd
rlabel metal1 s 24507 19235 24896 19266 4 vdd
rlabel metal1 s 22562 19234 22951 19265 4 vdd
rlabel metal1 s 7391 19235 7780 19266 4 vdd
rlabel metal1 s 10892 755 11281 786 4 vdd
rlabel metal1 s 8169 20774 8558 20805 4 vdd
rlabel metal1 s 3501 19235 3890 19266 4 vdd
rlabel metal1 s 4668 23854 5057 23885 4 vdd
rlabel metal1 s 23729 8455 24118 8486 4 vdd
rlabel metal1 s 24118 20775 24507 20806 4 vdd
rlabel metal1 s 14393 6914 14782 6945 4 vdd
rlabel metal1 s 12448 5374 12837 5405 4 vdd
rlabel metal1 s 24507 22314 24896 22345 4 vdd
rlabel metal1 s 21395 8454 21784 8485 4 vdd
rlabel metal1 s 389 11535 778 11566 4 vdd
rlabel metal1 s 17116 13074 17505 13105 4 vdd
rlabel metal1 s 389 14615 778 14646 4 vdd
rlabel metal1 s 5446 23855 5835 23886 4 vdd
rlabel metal1 s 22173 19234 22562 19265 4 vdd
rlabel metal1 s 19061 14614 19450 14645 4 vdd
rlabel metal1 s 19839 5374 20228 5405 4 vdd
rlabel metal1 s 7780 9995 8169 10026 4 vdd
rlabel metal1 s 14393 8454 14782 8485 4 vdd
rlabel metal1 s 13226 6915 13615 6946 4 vdd
rlabel metal1 s 12448 20774 12837 20805 4 vdd
rlabel metal1 s 13226 19235 13615 19266 4 vdd
rlabel metal1 s 22951 8455 23340 8486 4 vdd
rlabel metal1 s 4668 13075 5057 13106 4 vdd
rlabel metal1 s 21784 19235 22173 19266 4 vdd
rlabel metal1 s 1556 13075 1945 13106 4 vdd
rlabel metal1 s 11281 754 11670 785 4 vdd
rlabel metal1 s 15171 23855 15560 23886 4 vdd
rlabel metal1 s 11670 11534 12059 11565 4 vdd
rlabel metal1 s 0 5374 389 5405 4 vdd
rlabel metal1 s 10503 2295 10892 2326 4 vdd
rlabel metal1 s 18672 5375 19061 5406 4 vdd
rlabel metal1 s 17505 20774 17894 20805 4 vdd
rlabel metal1 s 13226 14614 13615 14645 4 vdd
rlabel metal1 s 21395 2295 21784 2326 4 vdd
rlabel metal1 s 22562 16155 22951 16186 4 vdd
rlabel metal1 s 778 8455 1167 8486 4 vdd
rlabel metal1 s 8558 754 8947 785 4 vdd
rlabel metal1 s 0 754 389 785 4 vdd
rlabel metal1 s 22951 5374 23340 5405 4 vdd
rlabel metal1 s 22951 17694 23340 17725 4 vdd
rlabel metal1 s 778 17694 1167 17725 4 vdd
rlabel metal1 s 9336 2295 9725 2326 4 vdd
rlabel metal1 s 12837 23855 13226 23886 4 vdd
rlabel metal1 s 11281 16154 11670 16185 4 vdd
rlabel metal1 s 9725 2294 10114 2325 4 vdd
rlabel metal1 s 3112 17695 3501 17726 4 vdd
rlabel metal1 s 7391 16155 7780 16186 4 vdd
rlabel metal1 s 14782 6914 15171 6945 4 vdd
rlabel metal1 s 17505 13074 17894 13105 4 vdd
rlabel metal1 s 2723 23854 3112 23885 4 vdd
rlabel metal1 s 19450 6914 19839 6945 4 vdd
rlabel metal1 s 6224 5374 6613 5405 4 vdd
rlabel metal1 s 9725 3835 10114 3866 4 vdd
rlabel metal1 s 14004 23855 14393 23886 4 vdd
rlabel metal1 s 2334 3834 2723 3865 4 vdd
rlabel metal1 s 12448 2294 12837 2325 4 vdd
rlabel metal1 s 23340 19234 23729 19265 4 vdd
rlabel metal1 s 1167 14615 1556 14646 4 vdd
rlabel metal1 s 19839 23855 20228 23886 4 vdd
rlabel metal1 s 17505 22315 17894 22346 4 vdd
rlabel metal1 s 19839 754 20228 785 4 vdd
rlabel metal1 s 7780 2295 8169 2326 4 vdd
rlabel metal1 s 14004 14615 14393 14646 4 vdd
rlabel metal1 s 15171 6915 15560 6946 4 vdd
rlabel metal1 s 17505 2295 17894 2326 4 vdd
rlabel metal1 s 15560 17694 15949 17725 4 vdd
rlabel metal1 s 23729 17695 24118 17726 4 vdd
rlabel metal1 s 24118 755 24507 786 4 vdd
rlabel metal1 s 18283 16154 18672 16185 4 vdd
rlabel metal1 s 19450 2294 19839 2325 4 vdd
rlabel metal1 s 5057 17695 5446 17726 4 vdd
rlabel metal1 s 22562 14615 22951 14646 4 vdd
rlabel metal1 s 0 8454 389 8485 4 vdd
rlabel metal1 s 4279 11535 4668 11566 4 vdd
rlabel metal1 s 19839 19235 20228 19266 4 vdd
rlabel metal1 s 389 8454 778 8485 4 vdd
rlabel metal1 s 389 20775 778 20806 4 vdd
rlabel metal1 s 11281 9995 11670 10026 4 vdd
rlabel metal1 s 11281 5374 11670 5405 4 vdd
rlabel metal1 s 12837 8454 13226 8485 4 vdd
rlabel metal1 s 3112 14614 3501 14645 4 vdd
rlabel metal1 s 1167 22314 1556 22345 4 vdd
rlabel metal1 s 10503 5375 10892 5406 4 vdd
rlabel metal1 s 17894 6915 18283 6946 4 vdd
rlabel metal1 s 22562 8454 22951 8485 4 vdd
rlabel metal1 s 5835 3834 6224 3865 4 vdd
rlabel metal1 s 11281 19234 11670 19265 4 vdd
rlabel metal1 s 12448 3835 12837 3866 4 vdd
rlabel metal1 s 5057 16154 5446 16185 4 vdd
rlabel metal1 s 11670 754 12059 785 4 vdd
rlabel metal1 s 5835 11535 6224 11566 4 vdd
rlabel metal1 s 15949 6915 16338 6946 4 vdd
rlabel metal1 s 6224 11534 6613 11565 4 vdd
rlabel metal1 s 0 5375 389 5406 4 vdd
rlabel metal1 s 21395 9994 21784 10025 4 vdd
rlabel metal1 s 5835 14615 6224 14646 4 vdd
rlabel metal1 s 10114 2294 10503 2325 4 vdd
rlabel metal1 s 5446 8454 5835 8485 4 vdd
rlabel metal1 s 3112 5375 3501 5406 4 vdd
rlabel metal1 s 20228 6915 20617 6946 4 vdd
rlabel metal1 s 16727 16155 17116 16186 4 vdd
rlabel metal1 s 15560 20774 15949 20805 4 vdd
rlabel metal1 s 17505 2294 17894 2325 4 vdd
rlabel metal1 s 19450 3835 19839 3866 4 vdd
rlabel metal1 s 5835 13074 6224 13105 4 vdd
rlabel metal1 s 15560 14615 15949 14646 4 vdd
rlabel metal1 s 11670 22314 12059 22345 4 vdd
rlabel metal1 s 778 5375 1167 5406 4 vdd
rlabel metal1 s 18672 8455 19061 8486 4 vdd
rlabel metal1 s 3501 13075 3890 13106 4 vdd
rlabel metal1 s 8558 3834 8947 3865 4 vdd
rlabel metal1 s 19061 23855 19450 23886 4 vdd
rlabel metal1 s 5835 16155 6224 16186 4 vdd
rlabel metal1 s 8169 13074 8558 13105 4 vdd
rlabel metal1 s 11670 3835 12059 3866 4 vdd
rlabel metal1 s 22173 14615 22562 14646 4 vdd
rlabel metal1 s 18672 3834 19061 3865 4 vdd
rlabel metal1 s 16338 14615 16727 14646 4 vdd
rlabel metal1 s 10114 8454 10503 8485 4 vdd
rlabel metal1 s 1167 16154 1556 16185 4 vdd
rlabel metal1 s 22173 17695 22562 17726 4 vdd
rlabel metal1 s 3501 22315 3890 22346 4 vdd
rlabel metal1 s 13615 5374 14004 5405 4 vdd
rlabel metal1 s 12448 2295 12837 2326 4 vdd
rlabel metal1 s 3112 3834 3501 3865 4 vdd
rlabel metal1 s 20228 23855 20617 23886 4 vdd
rlabel metal1 s 2723 19235 3112 19266 4 vdd
rlabel metal1 s 21006 14615 21395 14646 4 vdd
rlabel metal1 s 15949 23855 16338 23886 4 vdd
rlabel metal1 s 13226 5374 13615 5405 4 vdd
rlabel metal1 s 9336 17695 9725 17726 4 vdd
rlabel metal1 s 8558 14614 8947 14645 4 vdd
rlabel metal1 s 21784 20774 22173 20805 4 vdd
rlabel metal1 s 4279 16154 4668 16185 4 vdd
rlabel metal1 s 389 13075 778 13106 4 vdd
rlabel metal1 s 4668 5374 5057 5405 4 vdd
rlabel metal1 s 3501 2295 3890 2326 4 vdd
rlabel metal1 s 22562 11535 22951 11566 4 vdd
rlabel metal1 s 389 754 778 785 4 vdd
rlabel metal1 s 24507 17694 24896 17725 4 vdd
rlabel metal1 s 14004 6915 14393 6946 4 vdd
rlabel metal1 s 16727 9995 17116 10026 4 vdd
rlabel metal1 s 1945 16154 2334 16185 4 vdd
rlabel metal1 s 7391 22315 7780 22346 4 vdd
rlabel metal1 s 19061 23854 19450 23885 4 vdd
rlabel metal1 s 2723 17694 3112 17725 4 vdd
rlabel metal1 s 14782 17695 15171 17726 4 vdd
rlabel metal1 s 9725 16154 10114 16185 4 vdd
rlabel metal1 s 14393 13075 14782 13106 4 vdd
rlabel metal1 s 18283 9995 18672 10026 4 vdd
rlabel metal1 s 4279 9995 4668 10026 4 vdd
rlabel metal1 s 5057 5375 5446 5406 4 vdd
rlabel metal1 s 8947 20775 9336 20806 4 vdd
rlabel metal1 s 11670 2295 12059 2326 4 vdd
rlabel metal1 s 6224 5375 6613 5406 4 vdd
rlabel metal1 s 13226 5375 13615 5406 4 vdd
rlabel metal1 s 11670 19235 12059 19266 4 vdd
rlabel metal1 s 19839 23854 20228 23885 4 vdd
rlabel metal1 s 13615 22314 14004 22345 4 vdd
rlabel metal1 s 13226 23855 13615 23886 4 vdd
rlabel metal1 s 17505 19235 17894 19266 4 vdd
rlabel metal1 s 16338 9994 16727 10025 4 vdd
rlabel metal1 s 19839 13075 20228 13106 4 vdd
rlabel metal1 s 389 3835 778 3866 4 vdd
rlabel metal1 s 8558 20774 8947 20805 4 vdd
rlabel metal1 s 14004 5375 14393 5406 4 vdd
rlabel metal1 s 12059 3834 12448 3865 4 vdd
rlabel metal1 s 12837 22314 13226 22345 4 vdd
rlabel metal1 s 17116 3834 17505 3865 4 vdd
rlabel metal1 s 16727 8454 17116 8485 4 vdd
rlabel metal1 s 24507 13074 24896 13105 4 vdd
rlabel metal1 s 15171 13074 15560 13105 4 vdd
rlabel metal1 s 13615 14615 14004 14646 4 vdd
rlabel metal1 s 14782 23854 15171 23885 4 vdd
rlabel metal1 s 1167 5375 1556 5406 4 vdd
rlabel metal1 s 7780 14614 8169 14645 4 vdd
rlabel metal1 s 5057 8454 5446 8485 4 vdd
rlabel metal1 s 10114 19234 10503 19265 4 vdd
rlabel metal1 s 5446 2295 5835 2326 4 vdd
rlabel metal1 s 2334 5374 2723 5405 4 vdd
rlabel metal1 s 14782 22315 15171 22346 4 vdd
rlabel metal1 s 7391 9995 7780 10026 4 vdd
rlabel metal1 s 778 9994 1167 10025 4 vdd
rlabel metal1 s 1945 11534 2334 11565 4 vdd
rlabel metal1 s 3890 22314 4279 22345 4 vdd
rlabel metal1 s 13226 755 13615 786 4 vdd
rlabel metal1 s 13226 9995 13615 10026 4 vdd
rlabel metal1 s 6224 16155 6613 16186 4 vdd
rlabel metal1 s 17894 754 18283 785 4 vdd
rlabel metal1 s 8947 23854 9336 23885 4 vdd
rlabel metal1 s 4668 11535 5057 11566 4 vdd
rlabel metal1 s 5835 23855 6224 23886 4 vdd
rlabel metal1 s 3890 23855 4279 23886 4 vdd
rlabel metal1 s 12837 6914 13226 6945 4 vdd
rlabel metal1 s 7002 5375 7391 5406 4 vdd
rlabel metal1 s 11281 22314 11670 22345 4 vdd
rlabel metal1 s 11281 755 11670 786 4 vdd
rlabel metal1 s 3112 14615 3501 14646 4 vdd
rlabel metal1 s 7391 6915 7780 6946 4 vdd
rlabel metal1 s 0 22315 389 22346 4 vdd
rlabel metal1 s 21784 23854 22173 23885 4 vdd
rlabel metal1 s 21784 8455 22173 8486 4 vdd
rlabel metal1 s 17116 8455 17505 8486 4 vdd
rlabel metal1 s 9725 22314 10114 22345 4 vdd
rlabel metal1 s 18283 9994 18672 10025 4 vdd
rlabel metal1 s 17894 9995 18283 10026 4 vdd
rlabel metal1 s 3501 19234 3890 19265 4 vdd
rlabel metal1 s 1167 13075 1556 13106 4 vdd
rlabel metal1 s 7002 16154 7391 16185 4 vdd
rlabel metal1 s 1556 17694 1945 17725 4 vdd
rlabel metal1 s 1167 19234 1556 19265 4 vdd
rlabel metal1 s 24507 2295 24896 2326 4 vdd
rlabel metal1 s 23729 19234 24118 19265 4 vdd
rlabel metal1 s 20228 3835 20617 3866 4 vdd
rlabel metal1 s 22562 20775 22951 20806 4 vdd
rlabel metal1 s 7780 9994 8169 10025 4 vdd
rlabel metal1 s 21006 17695 21395 17726 4 vdd
rlabel metal1 s 6613 754 7002 785 4 vdd
rlabel metal1 s 2723 22314 3112 22345 4 vdd
rlabel metal1 s 3112 23854 3501 23885 4 vdd
rlabel metal1 s 10892 2295 11281 2326 4 vdd
rlabel metal1 s 10503 23855 10892 23886 4 vdd
rlabel metal1 s 21006 22314 21395 22345 4 vdd
rlabel metal1 s 22562 17694 22951 17725 4 vdd
rlabel metal1 s 24118 11534 24507 11565 4 vdd
rlabel metal1 s 3112 8455 3501 8486 4 vdd
rlabel metal1 s 19450 754 19839 785 4 vdd
rlabel metal1 s 14004 14614 14393 14645 4 vdd
rlabel metal1 s 2334 17695 2723 17726 4 vdd
rlabel metal1 s 22173 23854 22562 23885 4 vdd
rlabel metal1 s 8169 3834 8558 3865 4 vdd
rlabel metal1 s 11281 5375 11670 5406 4 vdd
rlabel metal1 s 2723 2294 3112 2325 4 vdd
rlabel metal1 s 12837 754 13226 785 4 vdd
rlabel metal1 s 5835 755 6224 786 4 vdd
rlabel metal1 s 0 6915 389 6946 4 vdd
rlabel metal1 s 20228 14614 20617 14645 4 vdd
rlabel metal1 s 7002 754 7391 785 4 vdd
rlabel metal1 s 19450 11534 19839 11565 4 vdd
rlabel metal1 s 15171 754 15560 785 4 vdd
rlabel metal1 s 9336 20774 9725 20805 4 vdd
rlabel metal1 s 22951 16155 23340 16186 4 vdd
rlabel metal1 s 6224 8455 6613 8486 4 vdd
rlabel metal1 s 17116 14615 17505 14646 4 vdd
rlabel metal1 s 24507 6914 24896 6945 4 vdd
rlabel metal1 s 7391 16154 7780 16185 4 vdd
rlabel metal1 s 15949 13075 16338 13106 4 vdd
rlabel metal1 s 10503 19235 10892 19266 4 vdd
rlabel metal1 s 17505 20775 17894 20806 4 vdd
rlabel metal1 s 9336 14615 9725 14646 4 vdd
rlabel metal1 s 19450 20774 19839 20805 4 vdd
rlabel metal1 s 22562 9995 22951 10026 4 vdd
rlabel metal1 s 21395 17694 21784 17725 4 vdd
rlabel metal1 s 4668 2295 5057 2326 4 vdd
rlabel metal1 s 23340 2295 23729 2326 4 vdd
rlabel metal1 s 10503 13074 10892 13105 4 vdd
rlabel metal1 s 3112 19235 3501 19266 4 vdd
rlabel metal1 s 8558 19235 8947 19266 4 vdd
rlabel metal1 s 22173 14614 22562 14645 4 vdd
rlabel metal1 s 4668 2294 5057 2325 4 vdd
rlabel metal1 s 5446 13075 5835 13106 4 vdd
rlabel metal1 s 13226 14615 13615 14646 4 vdd
rlabel metal1 s 8169 22315 8558 22346 4 vdd
rlabel metal1 s 12837 11534 13226 11565 4 vdd
rlabel metal1 s 3890 19234 4279 19265 4 vdd
rlabel metal1 s 4668 22314 5057 22345 4 vdd
rlabel metal1 s 14393 19234 14782 19265 4 vdd
rlabel metal1 s 10114 5374 10503 5405 4 vdd
rlabel metal1 s 13615 13074 14004 13105 4 vdd
rlabel metal1 s 3890 8454 4279 8485 4 vdd
rlabel metal1 s 22562 8455 22951 8486 4 vdd
rlabel metal1 s 0 14615 389 14646 4 vdd
rlabel metal1 s 0 13074 389 13105 4 vdd
rlabel metal1 s 13226 22314 13615 22345 4 vdd
rlabel metal1 s 23340 8454 23729 8485 4 vdd
rlabel metal1 s 6613 13075 7002 13106 4 vdd
rlabel metal1 s 7780 5375 8169 5406 4 vdd
rlabel metal1 s 10892 6915 11281 6946 4 vdd
rlabel metal1 s 13226 2294 13615 2325 4 vdd
rlabel metal1 s 17505 8455 17894 8486 4 vdd
rlabel metal1 s 24118 14615 24507 14646 4 vdd
rlabel metal1 s 17116 17694 17505 17725 4 vdd
rlabel metal1 s 17894 13074 18283 13105 4 vdd
rlabel metal1 s 7780 16155 8169 16186 4 vdd
rlabel metal1 s 20617 17694 21006 17725 4 vdd
rlabel metal1 s 10114 755 10503 786 4 vdd
rlabel metal1 s 14004 20775 14393 20806 4 vdd
rlabel metal1 s 4279 19234 4668 19265 4 vdd
rlabel metal1 s 20228 17694 20617 17725 4 vdd
rlabel metal1 s 4668 8454 5057 8485 4 vdd
rlabel metal1 s 9725 14615 10114 14646 4 vdd
rlabel metal1 s 2723 19234 3112 19265 4 vdd
rlabel metal1 s 1556 23855 1945 23886 4 vdd
rlabel metal1 s 7002 20774 7391 20805 4 vdd
rlabel metal1 s 16727 3835 17116 3866 4 vdd
rlabel metal1 s 3112 23855 3501 23886 4 vdd
rlabel metal1 s 17116 2295 17505 2326 4 vdd
rlabel metal1 s 2334 20775 2723 20806 4 vdd
rlabel metal1 s 19839 2295 20228 2326 4 vdd
rlabel metal1 s 15560 9995 15949 10026 4 vdd
rlabel metal1 s 23729 14615 24118 14646 4 vdd
rlabel metal1 s 3112 754 3501 785 4 vdd
rlabel metal1 s 8947 19235 9336 19266 4 vdd
rlabel metal1 s 17505 16154 17894 16185 4 vdd
rlabel metal1 s 21395 14614 21784 14645 4 vdd
rlabel metal1 s 22562 23854 22951 23885 4 vdd
rlabel metal1 s 17116 16155 17505 16186 4 vdd
rlabel metal1 s 12837 19235 13226 19266 4 vdd
rlabel metal1 s 9336 9995 9725 10026 4 vdd
rlabel metal1 s 10892 11534 11281 11565 4 vdd
rlabel metal1 s 14004 2294 14393 2325 4 vdd
rlabel metal1 s 11670 20775 12059 20806 4 vdd
rlabel metal1 s 5446 2294 5835 2325 4 vdd
rlabel metal1 s 9725 22315 10114 22346 4 vdd
rlabel metal1 s 14782 13075 15171 13106 4 vdd
rlabel metal1 s 3890 17695 4279 17726 4 vdd
rlabel metal1 s 21784 13075 22173 13106 4 vdd
rlabel metal1 s 18672 754 19061 785 4 vdd
rlabel metal1 s 15171 19235 15560 19266 4 vdd
rlabel metal1 s 778 11535 1167 11566 4 vdd
rlabel metal1 s 5057 20775 5446 20806 4 vdd
rlabel metal1 s 19061 8454 19450 8485 4 vdd
rlabel metal1 s 8558 11534 8947 11565 4 vdd
rlabel metal1 s 389 16155 778 16186 4 vdd
rlabel metal1 s 20617 19235 21006 19266 4 vdd
rlabel metal1 s 14393 3835 14782 3866 4 vdd
rlabel metal1 s 17505 9994 17894 10025 4 vdd
rlabel metal1 s 22173 6915 22562 6946 4 vdd
rlabel metal1 s 14393 17695 14782 17726 4 vdd
rlabel metal1 s 7002 9995 7391 10026 4 vdd
rlabel metal1 s 14782 19235 15171 19266 4 vdd
rlabel metal1 s 5446 23854 5835 23885 4 vdd
rlabel metal1 s 14393 13074 14782 13105 4 vdd
rlabel metal1 s 20228 16155 20617 16186 4 vdd
rlabel metal1 s 17894 17694 18283 17725 4 vdd
rlabel metal1 s 9336 6914 9725 6945 4 vdd
rlabel metal1 s 19839 9994 20228 10025 4 vdd
rlabel metal1 s 12448 755 12837 786 4 vdd
rlabel metal1 s 22951 11535 23340 11566 4 vdd
rlabel metal1 s 6613 5375 7002 5406 4 vdd
rlabel metal1 s 17116 5374 17505 5405 4 vdd
rlabel metal1 s 19839 20774 20228 20805 4 vdd
rlabel metal1 s 10892 19234 11281 19265 4 vdd
rlabel metal1 s 21395 5375 21784 5406 4 vdd
rlabel metal1 s 12837 17695 13226 17726 4 vdd
rlabel metal1 s 3501 755 3890 786 4 vdd
rlabel metal1 s 8558 13075 8947 13106 4 vdd
rlabel metal1 s 8558 755 8947 786 4 vdd
rlabel metal1 s 22951 14614 23340 14645 4 vdd
rlabel metal1 s 10503 17695 10892 17726 4 vdd
rlabel metal1 s 22173 16155 22562 16186 4 vdd
rlabel metal1 s 21006 14614 21395 14645 4 vdd
rlabel metal1 s 389 2295 778 2326 4 vdd
rlabel metal1 s 778 14615 1167 14646 4 vdd
rlabel metal1 s 17894 16155 18283 16186 4 vdd
rlabel metal1 s 8947 13074 9336 13105 4 vdd
rlabel metal1 s 10892 13074 11281 13105 4 vdd
rlabel metal1 s 18283 5375 18672 5406 4 vdd
rlabel metal1 s 11670 9995 12059 10026 4 vdd
rlabel metal1 s 19839 14614 20228 14645 4 vdd
rlabel metal1 s 17505 13075 17894 13106 4 vdd
rlabel metal1 s 20617 16155 21006 16186 4 vdd
rlabel metal1 s 18672 5374 19061 5405 4 vdd
rlabel metal1 s 19839 16154 20228 16185 4 vdd
rlabel metal1 s 9336 13074 9725 13105 4 vdd
rlabel metal1 s 17894 6914 18283 6945 4 vdd
rlabel metal1 s 15171 5375 15560 5406 4 vdd
rlabel metal1 s 1556 19234 1945 19265 4 vdd
rlabel metal1 s 19061 11534 19450 11565 4 vdd
rlabel metal1 s 10892 5375 11281 5406 4 vdd
rlabel metal1 s 5057 3835 5446 3866 4 vdd
rlabel metal1 s 2723 20774 3112 20805 4 vdd
rlabel metal1 s 7391 11535 7780 11566 4 vdd
rlabel metal1 s 18283 3835 18672 3866 4 vdd
rlabel metal1 s 8169 20775 8558 20806 4 vdd
rlabel metal1 s 21006 2294 21395 2325 4 vdd
rlabel metal1 s 1556 3834 1945 3865 4 vdd
rlabel metal1 s 23729 9994 24118 10025 4 vdd
rlabel metal1 s 20617 5375 21006 5406 4 vdd
rlabel metal1 s 389 22315 778 22346 4 vdd
rlabel metal1 s 14393 3834 14782 3865 4 vdd
rlabel metal1 s 8947 6915 9336 6946 4 vdd
rlabel metal1 s 778 23854 1167 23885 4 vdd
rlabel metal1 s 2334 6915 2723 6946 4 vdd
rlabel metal1 s 14393 2294 14782 2325 4 vdd
rlabel metal1 s 21784 6915 22173 6946 4 vdd
rlabel metal1 s 14004 19235 14393 19266 4 vdd
rlabel metal1 s 17505 5375 17894 5406 4 vdd
rlabel metal1 s 6613 16154 7002 16185 4 vdd
rlabel metal1 s 16727 5375 17116 5406 4 vdd
rlabel metal1 s 15949 16155 16338 16186 4 vdd
rlabel metal1 s 17894 19234 18283 19265 4 vdd
rlabel metal1 s 16338 16154 16727 16185 4 vdd
rlabel metal1 s 7780 5374 8169 5405 4 vdd
rlabel metal1 s 10892 2294 11281 2325 4 vdd
rlabel metal1 s 22562 22314 22951 22345 4 vdd
rlabel metal1 s 20617 3834 21006 3865 4 vdd
rlabel metal1 s 3112 755 3501 786 4 vdd
rlabel metal1 s 6224 11535 6613 11566 4 vdd
rlabel metal1 s 24507 3834 24896 3865 4 vdd
rlabel metal1 s 6613 22314 7002 22345 4 vdd
rlabel metal1 s 8947 5375 9336 5406 4 vdd
rlabel metal1 s 1556 11535 1945 11566 4 vdd
rlabel metal1 s 4279 19235 4668 19266 4 vdd
rlabel metal1 s 15560 17695 15949 17726 4 vdd
rlabel metal1 s 7002 13075 7391 13106 4 vdd
rlabel metal1 s 21395 11535 21784 11566 4 vdd
rlabel metal1 s 14782 23855 15171 23886 4 vdd
rlabel metal1 s 15949 9994 16338 10025 4 vdd
rlabel metal1 s 19450 8454 19839 8485 4 vdd
rlabel metal1 s 389 8455 778 8486 4 vdd
rlabel metal1 s 24118 14614 24507 14645 4 vdd
rlabel metal1 s 14393 755 14782 786 4 vdd
rlabel metal1 s 6224 16154 6613 16185 4 vdd
rlabel metal1 s 3112 20775 3501 20806 4 vdd
rlabel metal1 s 12837 20774 13226 20805 4 vdd
rlabel metal1 s 5835 5374 6224 5405 4 vdd
rlabel metal1 s 11670 11535 12059 11566 4 vdd
rlabel metal1 s 20617 13074 21006 13105 4 vdd
rlabel metal1 s 0 3835 389 3866 4 vdd
rlabel metal1 s 23729 3835 24118 3866 4 vdd
rlabel metal1 s 22951 13074 23340 13105 4 vdd
rlabel metal1 s 14393 8455 14782 8486 4 vdd
rlabel metal1 s 6224 17694 6613 17725 4 vdd
rlabel metal1 s 5057 2294 5446 2325 4 vdd
rlabel metal1 s 24507 754 24896 785 4 vdd
rlabel metal1 s 778 14614 1167 14645 4 vdd
rlabel metal1 s 4279 5374 4668 5405 4 vdd
rlabel metal1 s 16727 5374 17116 5405 4 vdd
rlabel metal1 s 389 14614 778 14645 4 vdd
rlabel metal1 s 3501 2294 3890 2325 4 vdd
rlabel metal1 s 19061 17694 19450 17725 4 vdd
rlabel metal1 s 22951 5375 23340 5406 4 vdd
rlabel metal1 s 8947 11534 9336 11565 4 vdd
rlabel metal1 s 23729 2294 24118 2325 4 vdd
rlabel metal1 s 23340 5375 23729 5406 4 vdd
rlabel metal1 s 12059 11534 12448 11565 4 vdd
rlabel metal1 s 9336 16155 9725 16186 4 vdd
rlabel metal1 s 14782 16154 15171 16185 4 vdd
rlabel metal1 s 15560 6914 15949 6945 4 vdd
rlabel metal1 s 3112 16154 3501 16185 4 vdd
rlabel metal1 s 389 19235 778 19266 4 vdd
rlabel metal1 s 21395 13075 21784 13106 4 vdd
rlabel metal1 s 18672 14614 19061 14645 4 vdd
rlabel metal1 s 6224 17695 6613 17726 4 vdd
rlabel metal1 s 21784 20775 22173 20806 4 vdd
rlabel metal1 s 13615 17694 14004 17725 4 vdd
rlabel metal1 s 778 19234 1167 19265 4 vdd
rlabel metal1 s 16338 6915 16727 6946 4 vdd
rlabel metal1 s 9336 22314 9725 22345 4 vdd
rlabel metal1 s 389 6914 778 6945 4 vdd
rlabel metal1 s 14782 11534 15171 11565 4 vdd
rlabel metal1 s 14782 19234 15171 19265 4 vdd
rlabel metal1 s 6224 19235 6613 19266 4 vdd
rlabel metal1 s 14782 2295 15171 2326 4 vdd
rlabel metal1 s 4279 755 4668 786 4 vdd
rlabel metal1 s 21006 20774 21395 20805 4 vdd
rlabel metal1 s 23340 14615 23729 14646 4 vdd
rlabel metal1 s 5835 16154 6224 16185 4 vdd
rlabel metal1 s 13615 5375 14004 5406 4 vdd
rlabel metal1 s 8558 6914 8947 6945 4 vdd
rlabel metal1 s 15171 13075 15560 13106 4 vdd
rlabel metal1 s 21006 22315 21395 22346 4 vdd
rlabel metal1 s 2723 14614 3112 14645 4 vdd
rlabel metal1 s 18672 3835 19061 3866 4 vdd
rlabel metal1 s 8169 14614 8558 14645 4 vdd
rlabel metal1 s 15560 755 15949 786 4 vdd
rlabel metal1 s 17116 8454 17505 8485 4 vdd
rlabel metal1 s 13615 14614 14004 14645 4 vdd
rlabel metal1 s 10503 2294 10892 2325 4 vdd
rlabel metal1 s 15949 755 16338 786 4 vdd
rlabel metal1 s 3501 3834 3890 3865 4 vdd
rlabel metal1 s 6224 22314 6613 22345 4 vdd
rlabel metal1 s 17116 16154 17505 16185 4 vdd
rlabel metal1 s 16727 11534 17116 11565 4 vdd
rlabel metal1 s 1167 3834 1556 3865 4 vdd
rlabel metal1 s 2334 3835 2723 3866 4 vdd
rlabel metal1 s 9725 19234 10114 19265 4 vdd
rlabel metal1 s 16338 23855 16727 23886 4 vdd
rlabel metal1 s 18672 20774 19061 20805 4 vdd
rlabel metal1 s 13226 17694 13615 17725 4 vdd
rlabel metal1 s 3501 16155 3890 16186 4 vdd
rlabel metal1 s 21006 3835 21395 3866 4 vdd
rlabel metal1 s 15560 22314 15949 22345 4 vdd
rlabel metal1 s 17505 11534 17894 11565 4 vdd
rlabel metal1 s 4279 5375 4668 5406 4 vdd
rlabel metal1 s 2334 5375 2723 5406 4 vdd
rlabel metal1 s 23340 14614 23729 14645 4 vdd
rlabel metal1 s 6224 3834 6613 3865 4 vdd
rlabel metal1 s 2334 20774 2723 20805 4 vdd
rlabel metal1 s 4668 9994 5057 10025 4 vdd
rlabel metal1 s 10892 16154 11281 16185 4 vdd
rlabel metal1 s 14782 755 15171 786 4 vdd
rlabel metal1 s 10892 3834 11281 3865 4 vdd
rlabel metal1 s 23729 6915 24118 6946 4 vdd
rlabel metal1 s 15171 5374 15560 5405 4 vdd
rlabel metal1 s 13615 23855 14004 23886 4 vdd
rlabel metal1 s 21395 6914 21784 6945 4 vdd
rlabel metal1 s 3501 14614 3890 14645 4 vdd
rlabel metal1 s 7391 23854 7780 23885 4 vdd
rlabel metal1 s 6224 19234 6613 19265 4 vdd
rlabel metal1 s 22173 19235 22562 19266 4 vdd
rlabel metal1 s 9725 5375 10114 5406 4 vdd
rlabel metal1 s 8169 22314 8558 22345 4 vdd
rlabel metal1 s 15171 2294 15560 2325 4 vdd
rlabel metal1 s 4668 3834 5057 3865 4 vdd
rlabel metal1 s 21006 11535 21395 11566 4 vdd
rlabel metal1 s 7391 20774 7780 20805 4 vdd
rlabel metal1 s 6613 9995 7002 10026 4 vdd
rlabel metal1 s 13615 9995 14004 10026 4 vdd
rlabel metal1 s 10114 3834 10503 3865 4 vdd
rlabel metal1 s 3112 16155 3501 16186 4 vdd
rlabel metal1 s 6224 22315 6613 22346 4 vdd
rlabel metal1 s 10114 754 10503 785 4 vdd
rlabel metal1 s 5057 13074 5446 13105 4 vdd
rlabel metal1 s 6224 6914 6613 6945 4 vdd
rlabel metal1 s 22173 20774 22562 20805 4 vdd
rlabel metal1 s 3501 8455 3890 8486 4 vdd
rlabel metal1 s 2723 754 3112 785 4 vdd
rlabel metal1 s 4668 5375 5057 5406 4 vdd
rlabel metal1 s 10503 8454 10892 8485 4 vdd
rlabel metal1 s 24118 17694 24507 17725 4 vdd
rlabel metal1 s 8169 6914 8558 6945 4 vdd
rlabel metal1 s 5057 14614 5446 14645 4 vdd
rlabel metal1 s 20228 17695 20617 17726 4 vdd
rlabel metal1 s 18283 20774 18672 20805 4 vdd
rlabel metal1 s 22173 2295 22562 2326 4 vdd
rlabel metal1 s 10503 6915 10892 6946 4 vdd
rlabel metal1 s 12059 23855 12448 23886 4 vdd
rlabel metal1 s 5446 6914 5835 6945 4 vdd
rlabel metal1 s 10114 19235 10503 19266 4 vdd
rlabel metal1 s 15560 5374 15949 5405 4 vdd
rlabel metal1 s 17116 19235 17505 19266 4 vdd
rlabel metal1 s 3890 22315 4279 22346 4 vdd
rlabel metal1 s 20617 17695 21006 17726 4 vdd
rlabel metal1 s 7002 14615 7391 14646 4 vdd
rlabel metal1 s 3890 5375 4279 5406 4 vdd
rlabel metal1 s 7391 8455 7780 8486 4 vdd
rlabel metal1 s 6613 5374 7002 5405 4 vdd
rlabel metal1 s 9725 20775 10114 20806 4 vdd
rlabel metal1 s 12059 20774 12448 20805 4 vdd
rlabel metal1 s 2723 16154 3112 16185 4 vdd
rlabel metal1 s 389 17694 778 17725 4 vdd
rlabel metal1 s 17505 3834 17894 3865 4 vdd
rlabel metal1 s 7780 23854 8169 23885 4 vdd
rlabel metal1 s 389 17695 778 17726 4 vdd
rlabel metal1 s 0 20775 389 20806 4 vdd
rlabel metal1 s 23729 23854 24118 23885 4 vdd
rlabel metal1 s 17505 9995 17894 10026 4 vdd
rlabel metal1 s 15949 754 16338 785 4 vdd
rlabel metal1 s 23340 20775 23729 20806 4 vdd
rlabel metal1 s 12448 14614 12837 14645 4 vdd
rlabel metal1 s 19839 755 20228 786 4 vdd
rlabel metal1 s 4279 14614 4668 14645 4 vdd
rlabel metal1 s 17505 5374 17894 5405 4 vdd
rlabel metal1 s 10892 22315 11281 22346 4 vdd
rlabel metal1 s 24507 16155 24896 16186 4 vdd
rlabel metal1 s 14004 8454 14393 8485 4 vdd
rlabel metal1 s 15171 17694 15560 17725 4 vdd
rlabel metal1 s 6224 6915 6613 6946 4 vdd
rlabel metal1 s 1556 23854 1945 23885 4 vdd
rlabel metal1 s 24507 8455 24896 8486 4 vdd
rlabel metal1 s 21784 11534 22173 11565 4 vdd
rlabel metal1 s 17116 5375 17505 5406 4 vdd
rlabel metal1 s 5835 2294 6224 2325 4 vdd
rlabel metal1 s 7391 8454 7780 8485 4 vdd
rlabel metal1 s 7002 20775 7391 20806 4 vdd
rlabel metal1 s 5057 23855 5446 23886 4 vdd
rlabel metal1 s 17116 20774 17505 20805 4 vdd
rlabel metal1 s 8169 17694 8558 17725 4 vdd
rlabel metal1 s 1556 8455 1945 8486 4 vdd
rlabel metal1 s 10503 11535 10892 11566 4 vdd
rlabel metal1 s 8558 8454 8947 8485 4 vdd
rlabel metal1 s 23729 22314 24118 22345 4 vdd
rlabel metal1 s 10503 755 10892 786 4 vdd
rlabel metal1 s 1556 8454 1945 8485 4 vdd
rlabel metal1 s 9725 11535 10114 11566 4 vdd
rlabel metal1 s 19061 2295 19450 2326 4 vdd
rlabel metal1 s 6613 2295 7002 2326 4 vdd
rlabel metal1 s 14782 22314 15171 22345 4 vdd
rlabel metal1 s 18283 6914 18672 6945 4 vdd
rlabel metal1 s 15560 754 15949 785 4 vdd
rlabel metal1 s 9336 16154 9725 16185 4 vdd
rlabel metal1 s 1556 17695 1945 17726 4 vdd
rlabel metal1 s 0 17695 389 17726 4 vdd
rlabel metal1 s 12448 11535 12837 11566 4 vdd
rlabel metal1 s 1556 2294 1945 2325 4 vdd
rlabel metal1 s 1167 754 1556 785 4 vdd
rlabel metal1 s 18283 6915 18672 6946 4 vdd
rlabel metal1 s 11670 20774 12059 20805 4 vdd
rlabel metal1 s 10114 14614 10503 14645 4 vdd
rlabel metal1 s 22951 19235 23340 19266 4 vdd
rlabel metal1 s 16338 22315 16727 22346 4 vdd
rlabel metal1 s 7002 5374 7391 5405 4 vdd
rlabel metal1 s 24118 17695 24507 17726 4 vdd
rlabel metal1 s 3890 13075 4279 13106 4 vdd
rlabel metal1 s 18283 8455 18672 8486 4 vdd
rlabel metal1 s 6224 23855 6613 23886 4 vdd
rlabel metal1 s 15949 10764 16338 10795 4 gnd
rlabel metal1 s 8169 3064 8558 3095 4 gnd
rlabel metal1 s 21395 24625 21784 24656 4 gnd
rlabel metal1 s 9336 21545 9725 21576 4 gnd
rlabel metal1 s 24507 9224 24896 9255 4 gnd
rlabel metal1 s 7002 12304 7391 12335 4 gnd
rlabel metal1 s 13615 21544 14004 21575 4 gnd
rlabel metal1 s 23729 21545 24118 21576 4 gnd
rlabel metal1 s 22562 3065 22951 3096 4 gnd
rlabel metal1 s 16338 10765 16727 10796 4 gnd
rlabel metal1 s 14004 6144 14393 6175 4 gnd
rlabel metal1 s 7780 18464 8169 18495 4 gnd
rlabel metal1 s 15171 4604 15560 4635 4 gnd
rlabel metal1 s 17505 9225 17894 9256 4 gnd
rlabel metal1 s 20617 10764 21006 10795 4 gnd
rlabel metal1 s 18672 6145 19061 6176 4 gnd
rlabel metal1 s 11670 13844 12059 13875 4 gnd
rlabel metal1 s 22173 23085 22562 23116 4 gnd
rlabel metal1 s 16338 16925 16727 16956 4 gnd
rlabel metal1 s 5446 21545 5835 21576 4 gnd
rlabel metal1 s 22951 23084 23340 23115 4 gnd
rlabel metal1 s 15949 13844 16338 13875 4 gnd
rlabel metal1 s 21395 12304 21784 12335 4 gnd
rlabel metal1 s 2723 7685 3112 7716 4 gnd
rlabel metal1 s 5835 9225 6224 9256 4 gnd
rlabel metal1 s 0 12304 389 12335 4 gnd
rlabel metal1 s 3501 7684 3890 7715 4 gnd
rlabel metal1 s 11670 20005 12059 20036 4 gnd
rlabel metal1 s 1167 -16 1556 15 4 gnd
rlabel metal1 s 3501 20005 3890 20036 4 gnd
rlabel metal1 s 22173 10765 22562 10796 4 gnd
rlabel metal1 s 6613 23084 7002 23115 4 gnd
rlabel metal1 s 10114 15385 10503 15416 4 gnd
rlabel metal1 s 12059 4604 12448 4635 4 gnd
rlabel metal1 s 13226 6145 13615 6176 4 gnd
rlabel metal1 s 0 6144 389 6175 4 gnd
rlabel metal1 s 8558 6145 8947 6176 4 gnd
rlabel metal1 s 3501 4604 3890 4635 4 gnd
rlabel metal1 s 18283 12304 18672 12335 4 gnd
rlabel metal1 s 23729 6144 24118 6175 4 gnd
rlabel metal1 s 20228 6144 20617 6175 4 gnd
rlabel metal1 s 10503 10764 10892 10795 4 gnd
rlabel metal1 s 12837 24625 13226 24656 4 gnd
rlabel metal1 s 1556 13844 1945 13875 4 gnd
rlabel metal1 s 17505 20005 17894 20036 4 gnd
rlabel metal1 s 3890 15384 4279 15415 4 gnd
rlabel metal1 s 7002 9225 7391 9256 4 gnd
rlabel metal1 s 18672 18464 19061 18495 4 gnd
rlabel metal1 s 20617 4605 21006 4636 4 gnd
rlabel metal1 s 16727 24625 17116 24656 4 gnd
rlabel metal1 s 22562 7685 22951 7716 4 gnd
rlabel metal1 s 19061 4605 19450 4636 4 gnd
rlabel metal1 s 18283 1524 18672 1555 4 gnd
rlabel metal1 s 10892 12304 11281 12335 4 gnd
rlabel metal1 s 8558 16924 8947 16955 4 gnd
rlabel metal1 s 13226 20005 13615 20036 4 gnd
rlabel metal1 s 3890 15385 4279 15416 4 gnd
rlabel metal1 s 11670 21545 12059 21576 4 gnd
rlabel metal1 s 12059 10764 12448 10795 4 gnd
rlabel metal1 s 5446 9225 5835 9256 4 gnd
rlabel metal1 s 1556 21544 1945 21575 4 gnd
rlabel metal1 s 7002 7685 7391 7716 4 gnd
rlabel metal1 s 13615 20005 14004 20036 4 gnd
rlabel metal1 s 11281 9225 11670 9256 4 gnd
rlabel metal1 s 21395 3065 21784 3096 4 gnd
rlabel metal1 s 13226 4605 13615 4636 4 gnd
rlabel metal1 s 13226 12305 13615 12336 4 gnd
rlabel metal1 s 9336 15384 9725 15415 4 gnd
rlabel metal1 s 24118 20005 24507 20036 4 gnd
rlabel metal1 s 13615 10765 14004 10796 4 gnd
rlabel metal1 s 5057 21545 5446 21576 4 gnd
rlabel metal1 s 23729 -16 24118 15 4 gnd
rlabel metal1 s 18672 13845 19061 13876 4 gnd
rlabel metal1 s 5835 4604 6224 4635 4 gnd
rlabel metal1 s 6613 9224 7002 9255 4 gnd
rlabel metal1 s 4668 20004 5057 20035 4 gnd
rlabel metal1 s 14782 21545 15171 21576 4 gnd
rlabel metal1 s 17894 4604 18283 4635 4 gnd
rlabel metal1 s 4279 10765 4668 10796 4 gnd
rlabel metal1 s 6224 -16 6613 15 4 gnd
rlabel metal1 s 11670 7685 12059 7716 4 gnd
rlabel metal1 s 8558 20005 8947 20036 4 gnd
rlabel metal1 s 16727 23085 17116 23116 4 gnd
rlabel metal1 s 24507 12305 24896 12336 4 gnd
rlabel metal1 s 20617 13845 21006 13876 4 gnd
rlabel metal1 s 5057 16925 5446 16956 4 gnd
rlabel metal1 s 15560 6144 15949 6175 4 gnd
rlabel metal1 s 24118 1524 24507 1555 4 gnd
rlabel metal1 s 21006 20005 21395 20036 4 gnd
rlabel metal1 s 1167 13844 1556 13875 4 gnd
rlabel metal1 s 18672 21544 19061 21575 4 gnd
rlabel metal1 s 4279 20004 4668 20035 4 gnd
rlabel metal1 s 19450 10764 19839 10795 4 gnd
rlabel metal1 s 4668 4605 5057 4636 4 gnd
rlabel metal1 s 16727 16924 17116 16955 4 gnd
rlabel metal1 s 14004 6145 14393 6176 4 gnd
rlabel metal1 s 20617 20005 21006 20036 4 gnd
rlabel metal1 s 4279 15384 4668 15415 4 gnd
rlabel metal1 s 6224 24625 6613 24656 4 gnd
rlabel metal1 s 8558 10764 8947 10795 4 gnd
rlabel metal1 s 18283 4605 18672 4636 4 gnd
rlabel metal1 s 10503 3065 10892 3096 4 gnd
rlabel metal1 s 13615 18464 14004 18495 4 gnd
rlabel metal1 s 18672 10764 19061 10795 4 gnd
rlabel metal1 s 13226 16925 13615 16956 4 gnd
rlabel metal1 s 9336 18464 9725 18495 4 gnd
rlabel metal1 s 5835 24625 6224 24656 4 gnd
rlabel metal1 s 21006 4605 21395 4636 4 gnd
rlabel metal1 s 9336 4605 9725 4636 4 gnd
rlabel metal1 s 16338 20005 16727 20036 4 gnd
rlabel metal1 s 19061 21545 19450 21576 4 gnd
rlabel metal1 s 21395 7685 21784 7716 4 gnd
rlabel metal1 s 8947 21544 9336 21575 4 gnd
rlabel metal1 s 16338 18464 16727 18495 4 gnd
rlabel metal1 s 24118 4604 24507 4635 4 gnd
rlabel metal1 s 18283 20004 18672 20035 4 gnd
rlabel metal1 s 15949 23084 16338 23115 4 gnd
rlabel metal1 s 19450 16924 19839 16955 4 gnd
rlabel metal1 s 24118 13845 24507 13876 4 gnd
rlabel metal1 s 21395 21544 21784 21575 4 gnd
rlabel metal1 s 10503 23085 10892 23116 4 gnd
rlabel metal1 s 24507 24625 24896 24656 4 gnd
rlabel metal1 s 22173 7685 22562 7716 4 gnd
rlabel metal1 s 13226 7685 13615 7716 4 gnd
rlabel metal1 s 17505 3065 17894 3096 4 gnd
rlabel metal1 s 11670 23085 12059 23116 4 gnd
rlabel metal1 s 778 -16 1167 15 4 gnd
rlabel metal1 s 12448 21545 12837 21576 4 gnd
rlabel metal1 s 778 3064 1167 3095 4 gnd
rlabel metal1 s 14782 7684 15171 7715 4 gnd
rlabel metal1 s 1167 1525 1556 1556 4 gnd
rlabel metal1 s 13226 13845 13615 13876 4 gnd
rlabel metal1 s 6224 16924 6613 16955 4 gnd
rlabel metal1 s 15949 1524 16338 1555 4 gnd
rlabel metal1 s 14004 12304 14393 12335 4 gnd
rlabel metal1 s 19450 13844 19839 13875 4 gnd
rlabel metal1 s 17116 21544 17505 21575 4 gnd
rlabel metal1 s 3112 3064 3501 3095 4 gnd
rlabel metal1 s 1945 3064 2334 3095 4 gnd
rlabel metal1 s 8558 7684 8947 7715 4 gnd
rlabel metal1 s 6224 1524 6613 1555 4 gnd
rlabel metal1 s 8169 13845 8558 13876 4 gnd
rlabel metal1 s 8558 13845 8947 13876 4 gnd
rlabel metal1 s 6224 12304 6613 12335 4 gnd
rlabel metal1 s 4668 23084 5057 23115 4 gnd
rlabel metal1 s 15560 1524 15949 1555 4 gnd
rlabel metal1 s 7780 1525 8169 1556 4 gnd
rlabel metal1 s 4668 3065 5057 3096 4 gnd
rlabel metal1 s 21006 21545 21395 21576 4 gnd
rlabel metal1 s 14393 9224 14782 9255 4 gnd
rlabel metal1 s 10892 18465 11281 18496 4 gnd
rlabel metal1 s 4279 9225 4668 9256 4 gnd
rlabel metal1 s 21784 12305 22173 12336 4 gnd
rlabel metal1 s 22173 12305 22562 12336 4 gnd
rlabel metal1 s 10892 10765 11281 10796 4 gnd
rlabel metal1 s 23729 6145 24118 6176 4 gnd
rlabel metal1 s 17505 21545 17894 21576 4 gnd
rlabel metal1 s 15949 -16 16338 15 4 gnd
rlabel metal1 s 2723 12305 3112 12336 4 gnd
rlabel metal1 s 7780 3065 8169 3096 4 gnd
rlabel metal1 s 4279 9224 4668 9255 4 gnd
rlabel metal1 s 14004 9224 14393 9255 4 gnd
rlabel metal1 s 22951 12305 23340 12336 4 gnd
rlabel metal1 s 16727 12305 17116 12336 4 gnd
rlabel metal1 s 0 20004 389 20035 4 gnd
rlabel metal1 s 6613 18464 7002 18495 4 gnd
rlabel metal1 s 20617 18465 21006 18496 4 gnd
rlabel metal1 s 17505 12304 17894 12335 4 gnd
rlabel metal1 s 5057 15385 5446 15416 4 gnd
rlabel metal1 s 7391 6145 7780 6176 4 gnd
rlabel metal1 s 9336 20005 9725 20036 4 gnd
rlabel metal1 s 389 6144 778 6175 4 gnd
rlabel metal1 s 14782 4605 15171 4636 4 gnd
rlabel metal1 s 8947 1524 9336 1555 4 gnd
rlabel metal1 s 6224 16925 6613 16956 4 gnd
rlabel metal1 s 7780 18465 8169 18496 4 gnd
rlabel metal1 s 15560 13845 15949 13876 4 gnd
rlabel metal1 s 9725 7685 10114 7716 4 gnd
rlabel metal1 s 8947 16925 9336 16956 4 gnd
rlabel metal1 s 19839 24625 20228 24656 4 gnd
rlabel metal1 s 11670 10764 12059 10795 4 gnd
rlabel metal1 s 4279 3064 4668 3095 4 gnd
rlabel metal1 s 19450 12305 19839 12336 4 gnd
rlabel metal1 s 24118 24625 24507 24656 4 gnd
rlabel metal1 s 15171 9224 15560 9255 4 gnd
rlabel metal1 s 9725 3064 10114 3095 4 gnd
rlabel metal1 s 1945 9224 2334 9255 4 gnd
rlabel metal1 s 12059 23084 12448 23115 4 gnd
rlabel metal1 s 16727 3064 17116 3095 4 gnd
rlabel metal1 s 9725 6145 10114 6176 4 gnd
rlabel metal1 s 5057 13844 5446 13875 4 gnd
rlabel metal1 s 23340 15385 23729 15416 4 gnd
rlabel metal1 s 23340 13844 23729 13875 4 gnd
rlabel metal1 s 21395 13844 21784 13875 4 gnd
rlabel metal1 s 23729 15384 24118 15415 4 gnd
rlabel metal1 s 2723 12304 3112 12335 4 gnd
rlabel metal1 s 778 10764 1167 10795 4 gnd
rlabel metal1 s 4279 1524 4668 1555 4 gnd
rlabel metal1 s 7391 20004 7780 20035 4 gnd
rlabel metal1 s 7780 20004 8169 20035 4 gnd
rlabel metal1 s 6613 20005 7002 20036 4 gnd
rlabel metal1 s 23729 23084 24118 23115 4 gnd
rlabel metal1 s 20617 15385 21006 15416 4 gnd
rlabel metal1 s 1167 15385 1556 15416 4 gnd
rlabel metal1 s 6224 15385 6613 15416 4 gnd
rlabel metal1 s 11281 4605 11670 4636 4 gnd
rlabel metal1 s 389 4604 778 4635 4 gnd
rlabel metal1 s 0 3065 389 3096 4 gnd
rlabel metal1 s 21784 9224 22173 9255 4 gnd
rlabel metal1 s 17505 4604 17894 4635 4 gnd
rlabel metal1 s 7780 13845 8169 13876 4 gnd
rlabel metal1 s 9725 4604 10114 4635 4 gnd
rlabel metal1 s 10892 1524 11281 1555 4 gnd
rlabel metal1 s 23340 7684 23729 7715 4 gnd
rlabel metal1 s 21006 10764 21395 10795 4 gnd
rlabel metal1 s 10892 7685 11281 7716 4 gnd
rlabel metal1 s 10114 -16 10503 15 4 gnd
rlabel metal1 s 7780 7684 8169 7715 4 gnd
rlabel metal1 s 16338 6144 16727 6175 4 gnd
rlabel metal1 s 7780 20005 8169 20036 4 gnd
rlabel metal1 s 14004 -16 14393 15 4 gnd
rlabel metal1 s 389 23084 778 23115 4 gnd
rlabel metal1 s 3501 1525 3890 1556 4 gnd
rlabel metal1 s 23729 10765 24118 10796 4 gnd
rlabel metal1 s 11281 20004 11670 20035 4 gnd
rlabel metal1 s 10503 13844 10892 13875 4 gnd
rlabel metal1 s 4668 24625 5057 24656 4 gnd
rlabel metal1 s 11281 12304 11670 12335 4 gnd
rlabel metal1 s 6613 1525 7002 1556 4 gnd
rlabel metal1 s 15171 4605 15560 4636 4 gnd
rlabel metal1 s 7780 24625 8169 24656 4 gnd
rlabel metal1 s 7780 10764 8169 10795 4 gnd
rlabel metal1 s 21006 7684 21395 7715 4 gnd
rlabel metal1 s 15560 13844 15949 13875 4 gnd
rlabel metal1 s 14004 3064 14393 3095 4 gnd
rlabel metal1 s 16338 20004 16727 20035 4 gnd
rlabel metal1 s 20617 13844 21006 13875 4 gnd
rlabel metal1 s 778 4604 1167 4635 4 gnd
rlabel metal1 s 23340 12305 23729 12336 4 gnd
rlabel metal1 s 8169 12304 8558 12335 4 gnd
rlabel metal1 s 2723 9225 3112 9256 4 gnd
rlabel metal1 s 3501 16925 3890 16956 4 gnd
rlabel metal1 s 4668 1524 5057 1555 4 gnd
rlabel metal1 s 389 1525 778 1556 4 gnd
rlabel metal1 s 2723 23084 3112 23115 4 gnd
rlabel metal1 s 778 6145 1167 6176 4 gnd
rlabel metal1 s 24118 6145 24507 6176 4 gnd
rlabel metal1 s 16338 7684 16727 7715 4 gnd
rlabel metal1 s 5835 15384 6224 15415 4 gnd
rlabel metal1 s 18283 13844 18672 13875 4 gnd
rlabel metal1 s 18672 23085 19061 23116 4 gnd
rlabel metal1 s 4279 -16 4668 15 4 gnd
rlabel metal1 s 8947 18464 9336 18495 4 gnd
rlabel metal1 s 15171 23084 15560 23115 4 gnd
rlabel metal1 s 21784 10764 22173 10795 4 gnd
rlabel metal1 s 1556 18464 1945 18495 4 gnd
rlabel metal1 s 5446 20004 5835 20035 4 gnd
rlabel metal1 s 15949 21544 16338 21575 4 gnd
rlabel metal1 s 22173 7684 22562 7715 4 gnd
rlabel metal1 s 8558 9224 8947 9255 4 gnd
rlabel metal1 s 24507 18465 24896 18496 4 gnd
rlabel metal1 s 11670 15384 12059 15415 4 gnd
rlabel metal1 s 3890 10765 4279 10796 4 gnd
rlabel metal1 s 21395 9225 21784 9256 4 gnd
rlabel metal1 s 14393 16925 14782 16956 4 gnd
rlabel metal1 s 7002 1524 7391 1555 4 gnd
rlabel metal1 s 13615 13845 14004 13876 4 gnd
rlabel metal1 s 1167 23085 1556 23116 4 gnd
rlabel metal1 s 19450 3064 19839 3095 4 gnd
rlabel metal1 s 2723 16924 3112 16955 4 gnd
rlabel metal1 s 3112 16925 3501 16956 4 gnd
rlabel metal1 s 21395 6145 21784 6176 4 gnd
rlabel metal1 s 7391 7685 7780 7716 4 gnd
rlabel metal1 s 10114 13844 10503 13875 4 gnd
rlabel metal1 s 778 23085 1167 23116 4 gnd
rlabel metal1 s 9336 16925 9725 16956 4 gnd
rlabel metal1 s 20228 20004 20617 20035 4 gnd
rlabel metal1 s 20228 21545 20617 21576 4 gnd
rlabel metal1 s 10503 18464 10892 18495 4 gnd
rlabel metal1 s 5057 6145 5446 6176 4 gnd
rlabel metal1 s 3501 21544 3890 21575 4 gnd
rlabel metal1 s 18672 4604 19061 4635 4 gnd
rlabel metal1 s 19450 1525 19839 1556 4 gnd
rlabel metal1 s 22951 3065 23340 3096 4 gnd
rlabel metal1 s 1556 3064 1945 3095 4 gnd
rlabel metal1 s 21395 23085 21784 23116 4 gnd
rlabel metal1 s 11670 15385 12059 15416 4 gnd
rlabel metal1 s 17116 7685 17505 7716 4 gnd
rlabel metal1 s 20228 23084 20617 23115 4 gnd
rlabel metal1 s 15560 4605 15949 4636 4 gnd
rlabel metal1 s 9336 12305 9725 12336 4 gnd
rlabel metal1 s 8558 16925 8947 16956 4 gnd
rlabel metal1 s 14393 24625 14782 24656 4 gnd
rlabel metal1 s 20617 16924 21006 16955 4 gnd
rlabel metal1 s 7780 12304 8169 12335 4 gnd
rlabel metal1 s 20228 6145 20617 6176 4 gnd
rlabel metal1 s 11281 20005 11670 20036 4 gnd
rlabel metal1 s 12448 4604 12837 4635 4 gnd
rlabel metal1 s 3501 10765 3890 10796 4 gnd
rlabel metal1 s 15560 20005 15949 20036 4 gnd
rlabel metal1 s 10892 9224 11281 9255 4 gnd
rlabel metal1 s 13615 16924 14004 16955 4 gnd
rlabel metal1 s 12059 9224 12448 9255 4 gnd
rlabel metal1 s 1556 9225 1945 9256 4 gnd
rlabel metal1 s 14393 20005 14782 20036 4 gnd
rlabel metal1 s 11670 21544 12059 21575 4 gnd
rlabel metal1 s 17894 23085 18283 23116 4 gnd
rlabel metal1 s 12837 12304 13226 12335 4 gnd
rlabel metal1 s 1167 7684 1556 7715 4 gnd
rlabel metal1 s 5446 13845 5835 13876 4 gnd
rlabel metal1 s 10503 24625 10892 24656 4 gnd
rlabel metal1 s 2334 12304 2723 12335 4 gnd
rlabel metal1 s 14782 7685 15171 7716 4 gnd
rlabel metal1 s 3112 4605 3501 4636 4 gnd
rlabel metal1 s 11670 6144 12059 6175 4 gnd
rlabel metal1 s 15560 18464 15949 18495 4 gnd
rlabel metal1 s 1167 10765 1556 10796 4 gnd
rlabel metal1 s 8947 15385 9336 15416 4 gnd
rlabel metal1 s 1945 10765 2334 10796 4 gnd
rlabel metal1 s 10503 16924 10892 16955 4 gnd
rlabel metal1 s 6613 1524 7002 1555 4 gnd
rlabel metal1 s 9725 1524 10114 1555 4 gnd
rlabel metal1 s 16338 21545 16727 21576 4 gnd
rlabel metal1 s 10114 18464 10503 18495 4 gnd
rlabel metal1 s 3112 20005 3501 20036 4 gnd
rlabel metal1 s 19061 3065 19450 3096 4 gnd
rlabel metal1 s 21006 20004 21395 20035 4 gnd
rlabel metal1 s 8169 24625 8558 24656 4 gnd
rlabel metal1 s 22562 9224 22951 9255 4 gnd
rlabel metal1 s 23729 1524 24118 1555 4 gnd
rlabel metal1 s 12059 3065 12448 3096 4 gnd
rlabel metal1 s 4279 3065 4668 3096 4 gnd
rlabel metal1 s 8169 6144 8558 6175 4 gnd
rlabel metal1 s 17505 10765 17894 10796 4 gnd
rlabel metal1 s 10503 6144 10892 6175 4 gnd
rlabel metal1 s 5835 -16 6224 15 4 gnd
rlabel metal1 s 9336 21544 9725 21575 4 gnd
rlabel metal1 s 4668 18465 5057 18496 4 gnd
rlabel metal1 s 13226 15384 13615 15415 4 gnd
rlabel metal1 s 12059 -16 12448 15 4 gnd
rlabel metal1 s 17894 20005 18283 20036 4 gnd
rlabel metal1 s 12448 21544 12837 21575 4 gnd
rlabel metal1 s 6224 20005 6613 20036 4 gnd
rlabel metal1 s 23340 16925 23729 16956 4 gnd
rlabel metal1 s 12448 6145 12837 6176 4 gnd
rlabel metal1 s 3112 9225 3501 9256 4 gnd
rlabel metal1 s 23340 1524 23729 1555 4 gnd
rlabel metal1 s 15949 23085 16338 23116 4 gnd
rlabel metal1 s 17894 9224 18283 9255 4 gnd
rlabel metal1 s 21784 13844 22173 13875 4 gnd
rlabel metal1 s 4668 20005 5057 20036 4 gnd
rlabel metal1 s 778 7685 1167 7716 4 gnd
rlabel metal1 s 14393 13844 14782 13875 4 gnd
rlabel metal1 s 19450 1524 19839 1555 4 gnd
rlabel metal1 s 389 20004 778 20035 4 gnd
rlabel metal1 s 6224 3065 6613 3096 4 gnd
rlabel metal1 s 2723 18465 3112 18496 4 gnd
rlabel metal1 s 17505 1525 17894 1556 4 gnd
rlabel metal1 s 2334 3065 2723 3096 4 gnd
rlabel metal1 s 12448 12305 12837 12336 4 gnd
rlabel metal1 s 19061 3064 19450 3095 4 gnd
rlabel metal1 s 9336 9225 9725 9256 4 gnd
rlabel metal1 s 24507 23085 24896 23116 4 gnd
rlabel metal1 s 4668 15385 5057 15416 4 gnd
rlabel metal1 s 1167 18464 1556 18495 4 gnd
rlabel metal1 s 7780 9224 8169 9255 4 gnd
rlabel metal1 s 21784 15384 22173 15415 4 gnd
rlabel metal1 s 2334 15384 2723 15415 4 gnd
rlabel metal1 s 23340 18465 23729 18496 4 gnd
rlabel metal1 s 21784 16924 22173 16955 4 gnd
rlabel metal1 s 2723 4605 3112 4636 4 gnd
rlabel metal1 s 13615 3064 14004 3095 4 gnd
rlabel metal1 s 21395 1525 21784 1556 4 gnd
rlabel metal1 s 2334 9224 2723 9255 4 gnd
rlabel metal1 s 5835 21545 6224 21576 4 gnd
rlabel metal1 s 17505 18464 17894 18495 4 gnd
rlabel metal1 s 14004 13845 14393 13876 4 gnd
rlabel metal1 s 13226 -16 13615 15 4 gnd
rlabel metal1 s 16338 23085 16727 23116 4 gnd
rlabel metal1 s 14004 24625 14393 24656 4 gnd
rlabel metal1 s 10503 20005 10892 20036 4 gnd
rlabel metal1 s 13615 9224 14004 9255 4 gnd
rlabel metal1 s 5446 18465 5835 18496 4 gnd
rlabel metal1 s 7391 20005 7780 20036 4 gnd
rlabel metal1 s 3112 1524 3501 1555 4 gnd
rlabel metal1 s 3890 23085 4279 23116 4 gnd
rlabel metal1 s 21784 6145 22173 6176 4 gnd
rlabel metal1 s 24118 21544 24507 21575 4 gnd
rlabel metal1 s 19061 23085 19450 23116 4 gnd
rlabel metal1 s 3112 16924 3501 16955 4 gnd
rlabel metal1 s 12837 21545 13226 21576 4 gnd
rlabel metal1 s 389 15385 778 15416 4 gnd
rlabel metal1 s 12059 15384 12448 15415 4 gnd
rlabel metal1 s 7780 12305 8169 12336 4 gnd
rlabel metal1 s 24507 4604 24896 4635 4 gnd
rlabel metal1 s 1556 3065 1945 3096 4 gnd
rlabel metal1 s 21006 1525 21395 1556 4 gnd
rlabel metal1 s 3112 6144 3501 6175 4 gnd
rlabel metal1 s 17116 20004 17505 20035 4 gnd
rlabel metal1 s 15949 3065 16338 3096 4 gnd
rlabel metal1 s 9725 -16 10114 15 4 gnd
rlabel metal1 s 13226 10765 13615 10796 4 gnd
rlabel metal1 s 14782 23085 15171 23116 4 gnd
rlabel metal1 s 19839 21545 20228 21576 4 gnd
rlabel metal1 s 10503 20004 10892 20035 4 gnd
rlabel metal1 s 20617 3064 21006 3095 4 gnd
rlabel metal1 s 7002 4604 7391 4635 4 gnd
rlabel metal1 s 389 9225 778 9256 4 gnd
rlabel metal1 s 16727 6144 17116 6175 4 gnd
rlabel metal1 s 21395 9224 21784 9255 4 gnd
rlabel metal1 s 17116 -16 17505 15 4 gnd
rlabel metal1 s 8169 21545 8558 21576 4 gnd
rlabel metal1 s 14393 9225 14782 9256 4 gnd
rlabel metal1 s 18283 7685 18672 7716 4 gnd
rlabel metal1 s 8558 6144 8947 6175 4 gnd
rlabel metal1 s 21784 4604 22173 4635 4 gnd
rlabel metal1 s 3890 20005 4279 20036 4 gnd
rlabel metal1 s 19450 10765 19839 10796 4 gnd
rlabel metal1 s 1945 1525 2334 1556 4 gnd
rlabel metal1 s 22951 6144 23340 6175 4 gnd
rlabel metal1 s 3112 7685 3501 7716 4 gnd
rlabel metal1 s 4668 12304 5057 12335 4 gnd
rlabel metal1 s 12059 23085 12448 23116 4 gnd
rlabel metal1 s 23729 23085 24118 23116 4 gnd
rlabel metal1 s 22951 23085 23340 23116 4 gnd
rlabel metal1 s 9336 1524 9725 1555 4 gnd
rlabel metal1 s 22173 23084 22562 23115 4 gnd
rlabel metal1 s 20617 15384 21006 15415 4 gnd
rlabel metal1 s 0 21544 389 21575 4 gnd
rlabel metal1 s 778 16924 1167 16955 4 gnd
rlabel metal1 s 17116 3065 17505 3096 4 gnd
rlabel metal1 s 1945 12305 2334 12336 4 gnd
rlabel metal1 s 18672 6144 19061 6175 4 gnd
rlabel metal1 s 6613 12305 7002 12336 4 gnd
rlabel metal1 s 24507 13845 24896 13876 4 gnd
rlabel metal1 s 13615 4604 14004 4635 4 gnd
rlabel metal1 s 20228 16925 20617 16956 4 gnd
rlabel metal1 s 3890 16924 4279 16955 4 gnd
rlabel metal1 s 24118 -16 24507 15 4 gnd
rlabel metal1 s 14393 23085 14782 23116 4 gnd
rlabel metal1 s 18283 18465 18672 18496 4 gnd
rlabel metal1 s 15560 10764 15949 10795 4 gnd
rlabel metal1 s 5835 18465 6224 18496 4 gnd
rlabel metal1 s 15949 16924 16338 16955 4 gnd
rlabel metal1 s 10892 6145 11281 6176 4 gnd
rlabel metal1 s 17116 20005 17505 20036 4 gnd
rlabel metal1 s 22173 9225 22562 9256 4 gnd
rlabel metal1 s 24507 9225 24896 9256 4 gnd
rlabel metal1 s 8169 9224 8558 9255 4 gnd
rlabel metal1 s 18672 12305 19061 12336 4 gnd
rlabel metal1 s 20617 10765 21006 10796 4 gnd
rlabel metal1 s 5057 24625 5446 24656 4 gnd
rlabel metal1 s 12837 20005 13226 20036 4 gnd
rlabel metal1 s 24507 15385 24896 15416 4 gnd
rlabel metal1 s 11670 9225 12059 9256 4 gnd
rlabel metal1 s 15949 21545 16338 21576 4 gnd
rlabel metal1 s 1556 4604 1945 4635 4 gnd
rlabel metal1 s 24507 3064 24896 3095 4 gnd
rlabel metal1 s 778 7684 1167 7715 4 gnd
rlabel metal1 s 19839 23085 20228 23116 4 gnd
rlabel metal1 s 13226 3065 13615 3096 4 gnd
rlabel metal1 s 14393 18464 14782 18495 4 gnd
rlabel metal1 s 10503 7685 10892 7716 4 gnd
rlabel metal1 s 16338 1524 16727 1555 4 gnd
rlabel metal1 s 10114 15384 10503 15415 4 gnd
rlabel metal1 s 13226 13844 13615 13875 4 gnd
rlabel metal1 s 389 24625 778 24656 4 gnd
rlabel metal1 s 5835 10765 6224 10796 4 gnd
rlabel metal1 s 22951 7685 23340 7716 4 gnd
rlabel metal1 s 21006 15384 21395 15415 4 gnd
rlabel metal1 s 14004 21545 14393 21576 4 gnd
rlabel metal1 s 18283 15385 18672 15416 4 gnd
rlabel metal1 s 21006 21544 21395 21575 4 gnd
rlabel metal1 s 18283 12305 18672 12336 4 gnd
rlabel metal1 s 21784 12304 22173 12335 4 gnd
rlabel metal1 s 18672 15384 19061 15415 4 gnd
rlabel metal1 s 14782 12305 15171 12336 4 gnd
rlabel metal1 s 18283 20005 18672 20036 4 gnd
rlabel metal1 s 6613 12304 7002 12335 4 gnd
rlabel metal1 s 17894 6145 18283 6176 4 gnd
rlabel metal1 s 10892 16925 11281 16956 4 gnd
rlabel metal1 s 4279 24625 4668 24656 4 gnd
rlabel metal1 s 20617 12305 21006 12336 4 gnd
rlabel metal1 s 12059 20004 12448 20035 4 gnd
rlabel metal1 s 22951 7684 23340 7715 4 gnd
rlabel metal1 s 5057 9225 5446 9256 4 gnd
rlabel metal1 s 2334 1524 2723 1555 4 gnd
rlabel metal1 s 23729 3065 24118 3096 4 gnd
rlabel metal1 s 22562 16924 22951 16955 4 gnd
rlabel metal1 s 17894 7685 18283 7716 4 gnd
rlabel metal1 s 1556 20005 1945 20036 4 gnd
rlabel metal1 s 19061 -16 19450 15 4 gnd
rlabel metal1 s 5835 3065 6224 3096 4 gnd
rlabel metal1 s 21395 20004 21784 20035 4 gnd
rlabel metal1 s 24118 3065 24507 3096 4 gnd
rlabel metal1 s 18283 23084 18672 23115 4 gnd
rlabel metal1 s 4668 1525 5057 1556 4 gnd
rlabel metal1 s 15171 24625 15560 24656 4 gnd
rlabel metal1 s 10114 16925 10503 16956 4 gnd
rlabel metal1 s 1945 13844 2334 13875 4 gnd
rlabel metal1 s 3501 9225 3890 9256 4 gnd
rlabel metal1 s 11670 -16 12059 15 4 gnd
rlabel metal1 s 4668 12305 5057 12336 4 gnd
rlabel metal1 s 23340 10764 23729 10795 4 gnd
rlabel metal1 s 1167 7685 1556 7716 4 gnd
rlabel metal1 s 10503 1524 10892 1555 4 gnd
rlabel metal1 s 11670 4605 12059 4636 4 gnd
rlabel metal1 s 16727 23084 17116 23115 4 gnd
rlabel metal1 s 14782 18464 15171 18495 4 gnd
rlabel metal1 s 389 7684 778 7715 4 gnd
rlabel metal1 s 15560 15384 15949 15415 4 gnd
rlabel metal1 s 3501 15385 3890 15416 4 gnd
rlabel metal1 s 6613 7684 7002 7715 4 gnd
rlabel metal1 s 8558 3065 8947 3096 4 gnd
rlabel metal1 s 10503 7684 10892 7715 4 gnd
rlabel metal1 s 19061 1525 19450 1556 4 gnd
rlabel metal1 s 13226 10764 13615 10795 4 gnd
rlabel metal1 s 1556 16924 1945 16955 4 gnd
rlabel metal1 s 8947 23084 9336 23115 4 gnd
rlabel metal1 s 5835 6145 6224 6176 4 gnd
rlabel metal1 s 3501 4605 3890 4636 4 gnd
rlabel metal1 s 9336 15385 9725 15416 4 gnd
rlabel metal1 s 2723 1525 3112 1556 4 gnd
rlabel metal1 s 21784 9225 22173 9256 4 gnd
rlabel metal1 s 4668 6144 5057 6175 4 gnd
rlabel metal1 s 18672 1524 19061 1555 4 gnd
rlabel metal1 s 11670 16925 12059 16956 4 gnd
rlabel metal1 s 1556 10765 1945 10796 4 gnd
rlabel metal1 s 7391 24625 7780 24656 4 gnd
rlabel metal1 s 19839 3065 20228 3096 4 gnd
rlabel metal1 s 4279 7684 4668 7715 4 gnd
rlabel metal1 s 20228 -16 20617 15 4 gnd
rlabel metal1 s 21784 24625 22173 24656 4 gnd
rlabel metal1 s 23340 6144 23729 6175 4 gnd
rlabel metal1 s 16727 1525 17116 1556 4 gnd
rlabel metal1 s 21006 10765 21395 10796 4 gnd
rlabel metal1 s 0 9224 389 9255 4 gnd
rlabel metal1 s 22562 20005 22951 20036 4 gnd
rlabel metal1 s 9725 18464 10114 18495 4 gnd
rlabel metal1 s 0 1525 389 1556 4 gnd
rlabel metal1 s 4668 18464 5057 18495 4 gnd
rlabel metal1 s 24118 10765 24507 10796 4 gnd
rlabel metal1 s 23340 7685 23729 7716 4 gnd
rlabel metal1 s 21784 3064 22173 3095 4 gnd
rlabel metal1 s 17894 21544 18283 21575 4 gnd
rlabel metal1 s 7002 4605 7391 4636 4 gnd
rlabel metal1 s 13615 15384 14004 15415 4 gnd
rlabel metal1 s 21395 7684 21784 7715 4 gnd
rlabel metal1 s 17894 13845 18283 13876 4 gnd
rlabel metal1 s 19061 10764 19450 10795 4 gnd
rlabel metal1 s 15949 12304 16338 12335 4 gnd
rlabel metal1 s 11670 9224 12059 9255 4 gnd
rlabel metal1 s 3112 21545 3501 21576 4 gnd
rlabel metal1 s 4668 3064 5057 3095 4 gnd
rlabel metal1 s 15171 3064 15560 3095 4 gnd
rlabel metal1 s 18672 23084 19061 23115 4 gnd
rlabel metal1 s 21395 4604 21784 4635 4 gnd
rlabel metal1 s 7391 18465 7780 18496 4 gnd
rlabel metal1 s 20617 4604 21006 4635 4 gnd
rlabel metal1 s 11281 18465 11670 18496 4 gnd
rlabel metal1 s 19450 4605 19839 4636 4 gnd
rlabel metal1 s 3501 7685 3890 7716 4 gnd
rlabel metal1 s 8169 18464 8558 18495 4 gnd
rlabel metal1 s 7780 9225 8169 9256 4 gnd
rlabel metal1 s 20228 4605 20617 4636 4 gnd
rlabel metal1 s 11281 16924 11670 16955 4 gnd
rlabel metal1 s 5446 23085 5835 23116 4 gnd
rlabel metal1 s 10503 -16 10892 15 4 gnd
rlabel metal1 s 7002 10764 7391 10795 4 gnd
rlabel metal1 s 14393 12305 14782 12336 4 gnd
rlabel metal1 s 18283 9225 18672 9256 4 gnd
rlabel metal1 s 5057 15384 5446 15415 4 gnd
rlabel metal1 s 14393 15384 14782 15415 4 gnd
rlabel metal1 s 21006 7685 21395 7716 4 gnd
rlabel metal1 s 14782 1524 15171 1555 4 gnd
rlabel metal1 s 12837 23084 13226 23115 4 gnd
rlabel metal1 s 14004 1525 14393 1556 4 gnd
rlabel metal1 s 22173 9224 22562 9255 4 gnd
rlabel metal1 s 3112 6145 3501 6176 4 gnd
rlabel metal1 s 2723 23085 3112 23116 4 gnd
rlabel metal1 s 11281 10764 11670 10795 4 gnd
rlabel metal1 s 15949 3064 16338 3095 4 gnd
rlabel metal1 s 17116 4604 17505 4635 4 gnd
rlabel metal1 s 21006 15385 21395 15416 4 gnd
rlabel metal1 s 7391 23085 7780 23116 4 gnd
rlabel metal1 s 2334 4604 2723 4635 4 gnd
rlabel metal1 s 17894 20004 18283 20035 4 gnd
rlabel metal1 s 18283 23085 18672 23116 4 gnd
rlabel metal1 s 5057 13845 5446 13876 4 gnd
rlabel metal1 s 18283 18464 18672 18495 4 gnd
rlabel metal1 s 24118 13844 24507 13875 4 gnd
rlabel metal1 s 14782 24625 15171 24656 4 gnd
rlabel metal1 s 9336 23084 9725 23115 4 gnd
rlabel metal1 s 21784 18465 22173 18496 4 gnd
rlabel metal1 s 14782 13845 15171 13876 4 gnd
rlabel metal1 s 3890 21544 4279 21575 4 gnd
rlabel metal1 s 2334 21545 2723 21576 4 gnd
rlabel metal1 s 14393 10764 14782 10795 4 gnd
rlabel metal1 s 17505 9224 17894 9255 4 gnd
rlabel metal1 s 14782 10764 15171 10795 4 gnd
rlabel metal1 s 21395 10764 21784 10795 4 gnd
rlabel metal1 s 16338 23084 16727 23115 4 gnd
rlabel metal1 s 1556 4605 1945 4636 4 gnd
rlabel metal1 s 21006 13845 21395 13876 4 gnd
rlabel metal1 s 3501 15384 3890 15415 4 gnd
rlabel metal1 s 17116 13844 17505 13875 4 gnd
rlabel metal1 s 12837 1524 13226 1555 4 gnd
rlabel metal1 s 16338 12304 16727 12335 4 gnd
rlabel metal1 s 19839 18464 20228 18495 4 gnd
rlabel metal1 s 23340 21545 23729 21576 4 gnd
rlabel metal1 s 6224 18464 6613 18495 4 gnd
rlabel metal1 s 8169 6145 8558 6176 4 gnd
rlabel metal1 s 4668 4604 5057 4635 4 gnd
rlabel metal1 s 20228 1525 20617 1556 4 gnd
rlabel metal1 s 1167 18465 1556 18496 4 gnd
rlabel metal1 s 11281 9224 11670 9255 4 gnd
rlabel metal1 s 6613 13844 7002 13875 4 gnd
rlabel metal1 s 8169 23085 8558 23116 4 gnd
rlabel metal1 s 13615 -16 14004 15 4 gnd
rlabel metal1 s 7780 23084 8169 23115 4 gnd
rlabel metal1 s 14782 1525 15171 1556 4 gnd
rlabel metal1 s 15171 15385 15560 15416 4 gnd
rlabel metal1 s 15949 18464 16338 18495 4 gnd
rlabel metal1 s 21784 3065 22173 3096 4 gnd
rlabel metal1 s 23340 3064 23729 3095 4 gnd
rlabel metal1 s 20228 12304 20617 12335 4 gnd
rlabel metal1 s 6224 9225 6613 9256 4 gnd
rlabel metal1 s 22173 1524 22562 1555 4 gnd
rlabel metal1 s 14782 4604 15171 4635 4 gnd
rlabel metal1 s 2334 -16 2723 15 4 gnd
rlabel metal1 s 19061 7684 19450 7715 4 gnd
rlabel metal1 s 13615 20004 14004 20035 4 gnd
rlabel metal1 s 14004 23084 14393 23115 4 gnd
rlabel metal1 s 18283 3065 18672 3096 4 gnd
rlabel metal1 s 14782 6145 15171 6176 4 gnd
rlabel metal1 s 3112 13844 3501 13875 4 gnd
rlabel metal1 s 5446 13844 5835 13875 4 gnd
rlabel metal1 s 22562 21544 22951 21575 4 gnd
rlabel metal1 s 23340 4605 23729 4636 4 gnd
rlabel metal1 s 2334 16924 2723 16955 4 gnd
rlabel metal1 s 12059 21544 12448 21575 4 gnd
rlabel metal1 s 17505 23084 17894 23115 4 gnd
rlabel metal1 s 23729 16925 24118 16956 4 gnd
rlabel metal1 s 22173 24625 22562 24656 4 gnd
rlabel metal1 s 1167 16925 1556 16956 4 gnd
rlabel metal1 s 21784 10765 22173 10796 4 gnd
rlabel metal1 s 13226 18465 13615 18496 4 gnd
rlabel metal1 s 2334 18465 2723 18496 4 gnd
rlabel metal1 s 19450 18465 19839 18496 4 gnd
rlabel metal1 s 22951 18464 23340 18495 4 gnd
rlabel metal1 s 15171 6145 15560 6176 4 gnd
rlabel metal1 s 7391 1524 7780 1555 4 gnd
rlabel metal1 s 4668 7685 5057 7716 4 gnd
rlabel metal1 s 7002 20004 7391 20035 4 gnd
rlabel metal1 s 12837 21544 13226 21575 4 gnd
rlabel metal1 s 17505 16924 17894 16955 4 gnd
rlabel metal1 s 389 16925 778 16956 4 gnd
rlabel metal1 s 10892 18464 11281 18495 4 gnd
rlabel metal1 s 21006 3064 21395 3095 4 gnd
rlabel metal1 s 389 18465 778 18496 4 gnd
rlabel metal1 s 3112 18464 3501 18495 4 gnd
rlabel metal1 s 10114 1524 10503 1555 4 gnd
rlabel metal1 s 6224 20004 6613 20035 4 gnd
rlabel metal1 s 20228 20005 20617 20036 4 gnd
rlabel metal1 s 24507 1525 24896 1556 4 gnd
rlabel metal1 s 20228 7684 20617 7715 4 gnd
rlabel metal1 s 6613 15384 7002 15415 4 gnd
rlabel metal1 s 5057 16924 5446 16955 4 gnd
rlabel metal1 s 2723 20005 3112 20036 4 gnd
rlabel metal1 s 15949 4604 16338 4635 4 gnd
rlabel metal1 s 7391 12305 7780 12336 4 gnd
rlabel metal1 s 8169 4605 8558 4636 4 gnd
rlabel metal1 s 6224 21545 6613 21576 4 gnd
rlabel metal1 s 7780 6145 8169 6176 4 gnd
rlabel metal1 s 23729 21544 24118 21575 4 gnd
rlabel metal1 s 19061 18465 19450 18496 4 gnd
rlabel metal1 s 11670 3064 12059 3095 4 gnd
rlabel metal1 s 12837 6145 13226 6176 4 gnd
rlabel metal1 s 1556 9224 1945 9255 4 gnd
rlabel metal1 s 4668 16925 5057 16956 4 gnd
rlabel metal1 s 8947 9225 9336 9256 4 gnd
rlabel metal1 s 15949 12305 16338 12336 4 gnd
rlabel metal1 s 13226 21545 13615 21576 4 gnd
rlabel metal1 s 19061 15385 19450 15416 4 gnd
rlabel metal1 s 12448 -16 12837 15 4 gnd
rlabel metal1 s 17505 3064 17894 3095 4 gnd
rlabel metal1 s 23340 21544 23729 21575 4 gnd
rlabel metal1 s 20228 7685 20617 7716 4 gnd
rlabel metal1 s 12448 15385 12837 15416 4 gnd
rlabel metal1 s 7391 16925 7780 16956 4 gnd
rlabel metal1 s 24507 20004 24896 20035 4 gnd
rlabel metal1 s 22562 12305 22951 12336 4 gnd
rlabel metal1 s 17894 13844 18283 13875 4 gnd
rlabel metal1 s 7391 3065 7780 3096 4 gnd
rlabel metal1 s 3890 24625 4279 24656 4 gnd
rlabel metal1 s 17894 12305 18283 12336 4 gnd
rlabel metal1 s 21784 7684 22173 7715 4 gnd
rlabel metal1 s 3112 15385 3501 15416 4 gnd
rlabel metal1 s 6224 4605 6613 4636 4 gnd
rlabel metal1 s 17116 6144 17505 6175 4 gnd
rlabel metal1 s 2334 15385 2723 15416 4 gnd
rlabel metal1 s 22562 4604 22951 4635 4 gnd
rlabel metal1 s 13226 9224 13615 9255 4 gnd
rlabel metal1 s 18672 16925 19061 16956 4 gnd
rlabel metal1 s 5835 7685 6224 7716 4 gnd
rlabel metal1 s 8947 10765 9336 10796 4 gnd
rlabel metal1 s 22951 15384 23340 15415 4 gnd
rlabel metal1 s 18283 16925 18672 16956 4 gnd
rlabel metal1 s 11670 23084 12059 23115 4 gnd
rlabel metal1 s 12837 13845 13226 13876 4 gnd
rlabel metal1 s 0 4604 389 4635 4 gnd
rlabel metal1 s 22562 10764 22951 10795 4 gnd
rlabel metal1 s 12059 7684 12448 7715 4 gnd
rlabel metal1 s 9725 16924 10114 16955 4 gnd
rlabel metal1 s 14393 21545 14782 21576 4 gnd
rlabel metal1 s 20617 9224 21006 9255 4 gnd
rlabel metal1 s 17894 6144 18283 6175 4 gnd
rlabel metal1 s 24118 7685 24507 7716 4 gnd
rlabel metal1 s 1945 21545 2334 21576 4 gnd
rlabel metal1 s 778 9224 1167 9255 4 gnd
rlabel metal1 s 1945 7684 2334 7715 4 gnd
rlabel metal1 s 10114 21545 10503 21576 4 gnd
rlabel metal1 s 23729 1525 24118 1556 4 gnd
rlabel metal1 s 17116 6145 17505 6176 4 gnd
rlabel metal1 s 3890 1524 4279 1555 4 gnd
rlabel metal1 s 4279 21544 4668 21575 4 gnd
rlabel metal1 s 24507 21544 24896 21575 4 gnd
rlabel metal1 s 15949 13845 16338 13876 4 gnd
rlabel metal1 s 12059 9225 12448 9256 4 gnd
rlabel metal1 s 14393 15385 14782 15416 4 gnd
rlabel metal1 s 12837 10765 13226 10796 4 gnd
rlabel metal1 s 8558 23085 8947 23116 4 gnd
rlabel metal1 s 13615 16925 14004 16956 4 gnd
rlabel metal1 s 14004 7685 14393 7716 4 gnd
rlabel metal1 s 389 21544 778 21575 4 gnd
rlabel metal1 s 8947 -16 9336 15 4 gnd
rlabel metal1 s 17894 10764 18283 10795 4 gnd
rlabel metal1 s 17894 18465 18283 18496 4 gnd
rlabel metal1 s 21395 18464 21784 18495 4 gnd
rlabel metal1 s 19450 -16 19839 15 4 gnd
rlabel metal1 s 8169 15385 8558 15416 4 gnd
rlabel metal1 s 15171 15384 15560 15415 4 gnd
rlabel metal1 s 7391 12304 7780 12335 4 gnd
rlabel metal1 s 15171 9225 15560 9256 4 gnd
rlabel metal1 s 778 12305 1167 12336 4 gnd
rlabel metal1 s 3112 15384 3501 15415 4 gnd
rlabel metal1 s 7002 6145 7391 6176 4 gnd
rlabel metal1 s 20617 20004 21006 20035 4 gnd
rlabel metal1 s 20228 10765 20617 10796 4 gnd
rlabel metal1 s 11670 18465 12059 18496 4 gnd
rlabel metal1 s 23340 18464 23729 18495 4 gnd
rlabel metal1 s 18283 21545 18672 21576 4 gnd
rlabel metal1 s 7780 3064 8169 3095 4 gnd
rlabel metal1 s 4279 6145 4668 6176 4 gnd
rlabel metal1 s 15560 9224 15949 9255 4 gnd
rlabel metal1 s 10503 10765 10892 10796 4 gnd
rlabel metal1 s 8169 21544 8558 21575 4 gnd
rlabel metal1 s 15171 12304 15560 12335 4 gnd
rlabel metal1 s 18672 -16 19061 15 4 gnd
rlabel metal1 s 19061 20005 19450 20036 4 gnd
rlabel metal1 s 21784 20005 22173 20036 4 gnd
rlabel metal1 s 4668 13844 5057 13875 4 gnd
rlabel metal1 s 3112 12304 3501 12335 4 gnd
rlabel metal1 s 9336 3064 9725 3095 4 gnd
rlabel metal1 s 4279 4604 4668 4635 4 gnd
rlabel metal1 s 778 16925 1167 16956 4 gnd
rlabel metal1 s 24507 13844 24896 13875 4 gnd
rlabel metal1 s 21784 15385 22173 15416 4 gnd
rlabel metal1 s 12448 18465 12837 18496 4 gnd
rlabel metal1 s 4668 15384 5057 15415 4 gnd
rlabel metal1 s 18672 21545 19061 21576 4 gnd
rlabel metal1 s 14782 3065 15171 3096 4 gnd
rlabel metal1 s 8558 7685 8947 7716 4 gnd
rlabel metal1 s 16727 4604 17116 4635 4 gnd
rlabel metal1 s 16727 4605 17116 4636 4 gnd
rlabel metal1 s 22173 3065 22562 3096 4 gnd
rlabel metal1 s 11281 -16 11670 15 4 gnd
rlabel metal1 s 17116 1524 17505 1555 4 gnd
rlabel metal1 s 7002 24625 7391 24656 4 gnd
rlabel metal1 s 22173 13845 22562 13876 4 gnd
rlabel metal1 s 3890 20004 4279 20035 4 gnd
rlabel metal1 s 4668 9225 5057 9256 4 gnd
rlabel metal1 s 24118 12305 24507 12336 4 gnd
rlabel metal1 s 1945 20005 2334 20036 4 gnd
rlabel metal1 s 12837 15384 13226 15415 4 gnd
rlabel metal1 s 15560 3064 15949 3095 4 gnd
rlabel metal1 s 3890 4605 4279 4636 4 gnd
rlabel metal1 s 10892 7684 11281 7715 4 gnd
rlabel metal1 s 22951 21545 23340 21576 4 gnd
rlabel metal1 s 19450 9224 19839 9255 4 gnd
rlabel metal1 s 3501 23085 3890 23116 4 gnd
rlabel metal1 s 7391 6144 7780 6175 4 gnd
rlabel metal1 s 14393 7685 14782 7716 4 gnd
rlabel metal1 s 16338 16924 16727 16955 4 gnd
rlabel metal1 s 21784 21544 22173 21575 4 gnd
rlabel metal1 s 389 15384 778 15415 4 gnd
rlabel metal1 s 5057 1524 5446 1555 4 gnd
rlabel metal1 s 19839 6144 20228 6175 4 gnd
rlabel metal1 s 16338 4604 16727 4635 4 gnd
rlabel metal1 s 0 9225 389 9256 4 gnd
rlabel metal1 s 10892 13845 11281 13876 4 gnd
rlabel metal1 s 22951 20004 23340 20035 4 gnd
rlabel metal1 s 14004 4604 14393 4635 4 gnd
rlabel metal1 s 3112 21544 3501 21575 4 gnd
rlabel metal1 s 8558 20004 8947 20035 4 gnd
rlabel metal1 s 2334 9225 2723 9256 4 gnd
rlabel metal1 s 10503 15384 10892 15415 4 gnd
rlabel metal1 s 19839 10765 20228 10796 4 gnd
rlabel metal1 s 778 1525 1167 1556 4 gnd
rlabel metal1 s 22562 10765 22951 10796 4 gnd
rlabel metal1 s 14004 15384 14393 15415 4 gnd
rlabel metal1 s 17505 6145 17894 6176 4 gnd
rlabel metal1 s 19839 15385 20228 15416 4 gnd
rlabel metal1 s 14004 20004 14393 20035 4 gnd
rlabel metal1 s 24507 10765 24896 10796 4 gnd
rlabel metal1 s 10114 21544 10503 21575 4 gnd
rlabel metal1 s 17116 10765 17505 10796 4 gnd
rlabel metal1 s 9336 10765 9725 10796 4 gnd
rlabel metal1 s 3501 24625 3890 24656 4 gnd
rlabel metal1 s 7391 23084 7780 23115 4 gnd
rlabel metal1 s 21784 1524 22173 1555 4 gnd
rlabel metal1 s 13615 7685 14004 7716 4 gnd
rlabel metal1 s 10892 3065 11281 3096 4 gnd
rlabel metal1 s 10503 16925 10892 16956 4 gnd
rlabel metal1 s 23340 9225 23729 9256 4 gnd
rlabel metal1 s 24507 4605 24896 4636 4 gnd
rlabel metal1 s 18672 18465 19061 18496 4 gnd
rlabel metal1 s 19839 13845 20228 13876 4 gnd
rlabel metal1 s 11281 3064 11670 3095 4 gnd
rlabel metal1 s 8558 4605 8947 4636 4 gnd
rlabel metal1 s 24118 4605 24507 4636 4 gnd
rlabel metal1 s 8169 16925 8558 16956 4 gnd
rlabel metal1 s 22951 10765 23340 10796 4 gnd
rlabel metal1 s 13615 15385 14004 15416 4 gnd
rlabel metal1 s 13226 18464 13615 18495 4 gnd
rlabel metal1 s 3501 6145 3890 6176 4 gnd
rlabel metal1 s 14782 15384 15171 15415 4 gnd
rlabel metal1 s 13226 24625 13615 24656 4 gnd
rlabel metal1 s 3890 9225 4279 9256 4 gnd
rlabel metal1 s 14004 1524 14393 1555 4 gnd
rlabel metal1 s 17505 1524 17894 1555 4 gnd
rlabel metal1 s 17894 3064 18283 3095 4 gnd
rlabel metal1 s 19839 4605 20228 4636 4 gnd
rlabel metal1 s 3501 12305 3890 12336 4 gnd
rlabel metal1 s 6224 18465 6613 18496 4 gnd
rlabel metal1 s 13615 23084 14004 23115 4 gnd
rlabel metal1 s 15949 20005 16338 20036 4 gnd
rlabel metal1 s 19061 20004 19450 20035 4 gnd
rlabel metal1 s 3890 16925 4279 16956 4 gnd
rlabel metal1 s 1556 1525 1945 1556 4 gnd
rlabel metal1 s 22951 18465 23340 18496 4 gnd
rlabel metal1 s 6224 10764 6613 10795 4 gnd
rlabel metal1 s 8169 15384 8558 15415 4 gnd
rlabel metal1 s 16727 -16 17116 15 4 gnd
rlabel metal1 s 22951 12304 23340 12335 4 gnd
rlabel metal1 s 18283 10764 18672 10795 4 gnd
rlabel metal1 s 4279 21545 4668 21576 4 gnd
rlabel metal1 s 5057 21544 5446 21575 4 gnd
rlabel metal1 s 1945 13845 2334 13876 4 gnd
rlabel metal1 s 18672 16924 19061 16955 4 gnd
rlabel metal1 s 1167 10764 1556 10795 4 gnd
rlabel metal1 s 1167 15384 1556 15415 4 gnd
rlabel metal1 s 778 18465 1167 18496 4 gnd
rlabel metal1 s 23340 20005 23729 20036 4 gnd
rlabel metal1 s 23340 12304 23729 12335 4 gnd
rlabel metal1 s 14782 9224 15171 9255 4 gnd
rlabel metal1 s 20617 21545 21006 21576 4 gnd
rlabel metal1 s 17116 7684 17505 7715 4 gnd
rlabel metal1 s 14004 4605 14393 4636 4 gnd
rlabel metal1 s 3890 21545 4279 21576 4 gnd
rlabel metal1 s 778 4605 1167 4636 4 gnd
rlabel metal1 s 5835 15385 6224 15416 4 gnd
rlabel metal1 s 17116 18464 17505 18495 4 gnd
rlabel metal1 s 8947 1525 9336 1556 4 gnd
rlabel metal1 s 10503 15385 10892 15416 4 gnd
rlabel metal1 s 3501 12304 3890 12335 4 gnd
rlabel metal1 s 12448 10765 12837 10796 4 gnd
rlabel metal1 s 12059 7685 12448 7716 4 gnd
rlabel metal1 s 24118 18465 24507 18496 4 gnd
rlabel metal1 s 19839 20005 20228 20036 4 gnd
rlabel metal1 s 8947 20005 9336 20036 4 gnd
rlabel metal1 s 8169 10765 8558 10796 4 gnd
rlabel metal1 s 13226 23085 13615 23116 4 gnd
rlabel metal1 s 23729 4605 24118 4636 4 gnd
rlabel metal1 s 3501 3065 3890 3096 4 gnd
rlabel metal1 s 21784 1525 22173 1556 4 gnd
rlabel metal1 s 0 -16 389 15 4 gnd
rlabel metal1 s 10114 23085 10503 23116 4 gnd
rlabel metal1 s 19450 24625 19839 24656 4 gnd
rlabel metal1 s 9725 20005 10114 20036 4 gnd
rlabel metal1 s 12837 10764 13226 10795 4 gnd
rlabel metal1 s 2723 13844 3112 13875 4 gnd
rlabel metal1 s 10892 23085 11281 23116 4 gnd
rlabel metal1 s 13615 12304 14004 12335 4 gnd
rlabel metal1 s 22173 20005 22562 20036 4 gnd
rlabel metal1 s 8169 16924 8558 16955 4 gnd
rlabel metal1 s 13226 12304 13615 12335 4 gnd
rlabel metal1 s 19061 15384 19450 15415 4 gnd
rlabel metal1 s 11281 21544 11670 21575 4 gnd
rlabel metal1 s 9725 23084 10114 23115 4 gnd
rlabel metal1 s 23729 18464 24118 18495 4 gnd
rlabel metal1 s 1945 16924 2334 16955 4 gnd
rlabel metal1 s 2723 1524 3112 1555 4 gnd
rlabel metal1 s 23340 10765 23729 10796 4 gnd
rlabel metal1 s 12837 20004 13226 20035 4 gnd
rlabel metal1 s 7780 6144 8169 6175 4 gnd
rlabel metal1 s 21784 23084 22173 23115 4 gnd
rlabel metal1 s 8169 4604 8558 4635 4 gnd
rlabel metal1 s 22173 12304 22562 12335 4 gnd
rlabel metal1 s 9725 16925 10114 16956 4 gnd
rlabel metal1 s 21395 15385 21784 15416 4 gnd
rlabel metal1 s 12059 12305 12448 12336 4 gnd
rlabel metal1 s 3501 13844 3890 13875 4 gnd
rlabel metal1 s 10503 23084 10892 23115 4 gnd
rlabel metal1 s 5446 18464 5835 18495 4 gnd
rlabel metal1 s 1167 9225 1556 9256 4 gnd
rlabel metal1 s 16727 10764 17116 10795 4 gnd
rlabel metal1 s 20228 1524 20617 1555 4 gnd
rlabel metal1 s 1556 10764 1945 10795 4 gnd
rlabel metal1 s 4668 13845 5057 13876 4 gnd
rlabel metal1 s 21395 6144 21784 6175 4 gnd
rlabel metal1 s 14004 7684 14393 7715 4 gnd
rlabel metal1 s 2723 21545 3112 21576 4 gnd
rlabel metal1 s 22562 15384 22951 15415 4 gnd
rlabel metal1 s 19450 12304 19839 12335 4 gnd
rlabel metal1 s 7780 15384 8169 15415 4 gnd
rlabel metal1 s 8169 1525 8558 1556 4 gnd
rlabel metal1 s 2723 20004 3112 20035 4 gnd
rlabel metal1 s 1167 24625 1556 24656 4 gnd
rlabel metal1 s 22951 9225 23340 9256 4 gnd
rlabel metal1 s 389 4605 778 4636 4 gnd
rlabel metal1 s 4668 10764 5057 10795 4 gnd
rlabel metal1 s 6224 12305 6613 12336 4 gnd
rlabel metal1 s 22562 24625 22951 24656 4 gnd
rlabel metal1 s 10503 4605 10892 4636 4 gnd
rlabel metal1 s 15949 15385 16338 15416 4 gnd
rlabel metal1 s 8947 9224 9336 9255 4 gnd
rlabel metal1 s 11281 10765 11670 10796 4 gnd
rlabel metal1 s 8169 1524 8558 1555 4 gnd
rlabel metal1 s 18672 1525 19061 1556 4 gnd
rlabel metal1 s 6224 7684 6613 7715 4 gnd
rlabel metal1 s 15560 16925 15949 16956 4 gnd
rlabel metal1 s 21006 3065 21395 3096 4 gnd
rlabel metal1 s 9336 13845 9725 13876 4 gnd
rlabel metal1 s 9725 18465 10114 18496 4 gnd
rlabel metal1 s 15949 18465 16338 18496 4 gnd
rlabel metal1 s 8169 3065 8558 3096 4 gnd
rlabel metal1 s 20617 6144 21006 6175 4 gnd
rlabel metal1 s 18283 10765 18672 10796 4 gnd
rlabel metal1 s 4279 10764 4668 10795 4 gnd
rlabel metal1 s 19061 4604 19450 4635 4 gnd
rlabel metal1 s 22562 3064 22951 3095 4 gnd
rlabel metal1 s 24507 -16 24896 15 4 gnd
rlabel metal1 s 3501 23084 3890 23115 4 gnd
rlabel metal1 s 12059 1525 12448 1556 4 gnd
rlabel metal1 s 23729 20005 24118 20036 4 gnd
rlabel metal1 s 15171 16924 15560 16955 4 gnd
rlabel metal1 s 20228 24625 20617 24656 4 gnd
rlabel metal1 s 0 13844 389 13875 4 gnd
rlabel metal1 s 20228 21544 20617 21575 4 gnd
rlabel metal1 s 7002 1525 7391 1556 4 gnd
rlabel metal1 s 6613 16924 7002 16955 4 gnd
rlabel metal1 s 15560 1525 15949 1556 4 gnd
rlabel metal1 s 8558 -16 8947 15 4 gnd
rlabel metal1 s 1945 18465 2334 18496 4 gnd
rlabel metal1 s 22562 1525 22951 1556 4 gnd
rlabel metal1 s 20228 3065 20617 3096 4 gnd
rlabel metal1 s 24118 3064 24507 3095 4 gnd
rlabel metal1 s 17116 24625 17505 24656 4 gnd
rlabel metal1 s 17116 23085 17505 23116 4 gnd
rlabel metal1 s 9725 12304 10114 12335 4 gnd
rlabel metal1 s 0 3064 389 3095 4 gnd
rlabel metal1 s 6224 3064 6613 3095 4 gnd
rlabel metal1 s 18672 7685 19061 7716 4 gnd
rlabel metal1 s 1945 9225 2334 9256 4 gnd
rlabel metal1 s 1945 20004 2334 20035 4 gnd
rlabel metal1 s 13615 23085 14004 23116 4 gnd
rlabel metal1 s 18283 -16 18672 15 4 gnd
rlabel metal1 s 8558 13844 8947 13875 4 gnd
rlabel metal1 s 7780 4604 8169 4635 4 gnd
rlabel metal1 s 8169 7684 8558 7715 4 gnd
rlabel metal1 s 7391 4605 7780 4636 4 gnd
rlabel metal1 s 19839 12304 20228 12335 4 gnd
rlabel metal1 s 6613 10764 7002 10795 4 gnd
rlabel metal1 s 3501 18465 3890 18496 4 gnd
rlabel metal1 s 3890 12304 4279 12335 4 gnd
rlabel metal1 s 24118 23084 24507 23115 4 gnd
rlabel metal1 s 5835 23084 6224 23115 4 gnd
rlabel metal1 s 4279 16925 4668 16956 4 gnd
rlabel metal1 s 9725 15384 10114 15415 4 gnd
rlabel metal1 s 2334 23085 2723 23116 4 gnd
rlabel metal1 s 17505 16925 17894 16956 4 gnd
rlabel metal1 s 15949 1525 16338 1556 4 gnd
rlabel metal1 s 19061 12304 19450 12335 4 gnd
rlabel metal1 s 22562 23085 22951 23116 4 gnd
rlabel metal1 s 5446 12305 5835 12336 4 gnd
rlabel metal1 s 12448 6144 12837 6175 4 gnd
rlabel metal1 s 22173 21544 22562 21575 4 gnd
rlabel metal1 s 18672 9225 19061 9256 4 gnd
rlabel metal1 s 14782 20005 15171 20036 4 gnd
rlabel metal1 s 7002 23084 7391 23115 4 gnd
rlabel metal1 s 22951 6145 23340 6176 4 gnd
rlabel metal1 s 12837 16924 13226 16955 4 gnd
rlabel metal1 s 7002 -16 7391 15 4 gnd
rlabel metal1 s 24118 10764 24507 10795 4 gnd
rlabel metal1 s 16727 15385 17116 15416 4 gnd
rlabel metal1 s 3501 21545 3890 21576 4 gnd
rlabel metal1 s 21395 12305 21784 12336 4 gnd
rlabel metal1 s 15171 6144 15560 6175 4 gnd
rlabel metal1 s 20228 4604 20617 4635 4 gnd
rlabel metal1 s 7002 21544 7391 21575 4 gnd
rlabel metal1 s 9725 23085 10114 23116 4 gnd
rlabel metal1 s 24118 9225 24507 9256 4 gnd
rlabel metal1 s 19839 4604 20228 4635 4 gnd
rlabel metal1 s 19061 21544 19450 21575 4 gnd
rlabel metal1 s 11670 10765 12059 10796 4 gnd
rlabel metal1 s 9725 13845 10114 13876 4 gnd
rlabel metal1 s 18283 21544 18672 21575 4 gnd
rlabel metal1 s 6613 6145 7002 6176 4 gnd
rlabel metal1 s 5057 12304 5446 12335 4 gnd
rlabel metal1 s 8947 10764 9336 10795 4 gnd
rlabel metal1 s 9336 7685 9725 7716 4 gnd
rlabel metal1 s 13226 7684 13615 7715 4 gnd
rlabel metal1 s 22951 16924 23340 16955 4 gnd
rlabel metal1 s 22562 13845 22951 13876 4 gnd
rlabel metal1 s 5835 16924 6224 16955 4 gnd
rlabel metal1 s 16727 21545 17116 21576 4 gnd
rlabel metal1 s 17116 15385 17505 15416 4 gnd
rlabel metal1 s 12448 3065 12837 3096 4 gnd
rlabel metal1 s 3890 -16 4279 15 4 gnd
rlabel metal1 s 15171 1524 15560 1555 4 gnd
rlabel metal1 s 14393 7684 14782 7715 4 gnd
rlabel metal1 s 16338 15384 16727 15415 4 gnd
rlabel metal1 s 22562 9225 22951 9256 4 gnd
rlabel metal1 s 5446 10765 5835 10796 4 gnd
rlabel metal1 s 6613 23085 7002 23116 4 gnd
rlabel metal1 s 18283 1525 18672 1556 4 gnd
rlabel metal1 s 21006 1524 21395 1555 4 gnd
rlabel metal1 s 7391 -16 7780 15 4 gnd
rlabel metal1 s 12448 1525 12837 1556 4 gnd
rlabel metal1 s 21784 -16 22173 15 4 gnd
rlabel metal1 s 2723 3064 3112 3095 4 gnd
rlabel metal1 s 6613 9225 7002 9256 4 gnd
rlabel metal1 s 389 23085 778 23116 4 gnd
rlabel metal1 s 4668 6145 5057 6176 4 gnd
rlabel metal1 s 13615 9225 14004 9256 4 gnd
rlabel metal1 s 4279 23084 4668 23115 4 gnd
rlabel metal1 s 17116 9225 17505 9256 4 gnd
rlabel metal1 s 17505 13845 17894 13876 4 gnd
rlabel metal1 s 10503 4604 10892 4635 4 gnd
rlabel metal1 s 22173 6145 22562 6176 4 gnd
rlabel metal1 s 15949 24625 16338 24656 4 gnd
rlabel metal1 s 1945 4604 2334 4635 4 gnd
rlabel metal1 s 14782 21544 15171 21575 4 gnd
rlabel metal1 s 3112 12305 3501 12336 4 gnd
rlabel metal1 s 10892 6144 11281 6175 4 gnd
rlabel metal1 s 14004 3065 14393 3096 4 gnd
rlabel metal1 s 7002 23085 7391 23116 4 gnd
rlabel metal1 s 15949 16925 16338 16956 4 gnd
rlabel metal1 s 12059 6144 12448 6175 4 gnd
rlabel metal1 s 15949 7685 16338 7716 4 gnd
rlabel metal1 s 22951 4604 23340 4635 4 gnd
rlabel metal1 s 19061 7685 19450 7716 4 gnd
rlabel metal1 s 9725 12305 10114 12336 4 gnd
rlabel metal1 s 7391 13844 7780 13875 4 gnd
rlabel metal1 s 14393 12304 14782 12335 4 gnd
rlabel metal1 s 9725 7684 10114 7715 4 gnd
rlabel metal1 s 12059 12304 12448 12335 4 gnd
rlabel metal1 s 14393 16924 14782 16955 4 gnd
rlabel metal1 s 15560 24625 15949 24656 4 gnd
rlabel metal1 s 7391 16924 7780 16955 4 gnd
rlabel metal1 s 21395 23084 21784 23115 4 gnd
rlabel metal1 s 4668 10765 5057 10796 4 gnd
rlabel metal1 s 10503 12304 10892 12335 4 gnd
rlabel metal1 s 23729 7684 24118 7715 4 gnd
rlabel metal1 s 7002 16924 7391 16955 4 gnd
rlabel metal1 s 2723 24625 3112 24656 4 gnd
rlabel metal1 s 3890 18464 4279 18495 4 gnd
rlabel metal1 s 6613 6144 7002 6175 4 gnd
rlabel metal1 s 1945 15384 2334 15415 4 gnd
rlabel metal1 s 5057 3065 5446 3096 4 gnd
rlabel metal1 s 11281 16925 11670 16956 4 gnd
rlabel metal1 s 6224 21544 6613 21575 4 gnd
rlabel metal1 s 13615 18465 14004 18496 4 gnd
rlabel metal1 s 16727 9224 17116 9255 4 gnd
rlabel metal1 s 13615 10764 14004 10795 4 gnd
rlabel metal1 s 6613 4605 7002 4636 4 gnd
rlabel metal1 s 19839 16924 20228 16955 4 gnd
rlabel metal1 s 5835 21544 6224 21575 4 gnd
rlabel metal1 s 21395 1524 21784 1555 4 gnd
rlabel metal1 s 9725 1525 10114 1556 4 gnd
rlabel metal1 s 12448 16925 12837 16956 4 gnd
rlabel metal1 s 15949 4605 16338 4636 4 gnd
rlabel metal1 s 19839 12305 20228 12336 4 gnd
rlabel metal1 s 6613 7685 7002 7716 4 gnd
rlabel metal1 s 13226 16924 13615 16955 4 gnd
rlabel metal1 s 10114 7685 10503 7716 4 gnd
rlabel metal1 s 11670 6145 12059 6176 4 gnd
rlabel metal1 s 12837 18465 13226 18496 4 gnd
rlabel metal1 s 20228 18465 20617 18496 4 gnd
rlabel metal1 s 3112 7684 3501 7715 4 gnd
rlabel metal1 s 17505 15384 17894 15415 4 gnd
rlabel metal1 s 10892 24625 11281 24656 4 gnd
rlabel metal1 s 5057 10764 5446 10795 4 gnd
rlabel metal1 s 1167 20004 1556 20035 4 gnd
rlabel metal1 s 389 7685 778 7716 4 gnd
rlabel metal1 s 5057 23085 5446 23116 4 gnd
rlabel metal1 s 1945 23084 2334 23115 4 gnd
rlabel metal1 s 23340 16924 23729 16955 4 gnd
rlabel metal1 s 8558 1525 8947 1556 4 gnd
rlabel metal1 s 9725 3065 10114 3096 4 gnd
rlabel metal1 s 9336 18465 9725 18496 4 gnd
rlabel metal1 s 10503 9224 10892 9255 4 gnd
rlabel metal1 s 5835 18464 6224 18495 4 gnd
rlabel metal1 s 11670 1524 12059 1555 4 gnd
rlabel metal1 s 22562 1524 22951 1555 4 gnd
rlabel metal1 s 3501 9224 3890 9255 4 gnd
rlabel metal1 s 6613 20004 7002 20035 4 gnd
rlabel metal1 s 4668 21544 5057 21575 4 gnd
rlabel metal1 s 8558 24625 8947 24656 4 gnd
rlabel metal1 s 3501 13845 3890 13876 4 gnd
rlabel metal1 s 10114 10764 10503 10795 4 gnd
rlabel metal1 s 20228 3064 20617 3095 4 gnd
rlabel metal1 s 18672 3064 19061 3095 4 gnd
rlabel metal1 s 10114 3065 10503 3096 4 gnd
rlabel metal1 s 23340 23085 23729 23116 4 gnd
rlabel metal1 s 5835 9224 6224 9255 4 gnd
rlabel metal1 s 9336 20004 9725 20035 4 gnd
rlabel metal1 s 10892 4604 11281 4635 4 gnd
rlabel metal1 s 5057 12305 5446 12336 4 gnd
rlabel metal1 s 21006 12305 21395 12336 4 gnd
rlabel metal1 s 11281 6144 11670 6175 4 gnd
rlabel metal1 s 1556 12305 1945 12336 4 gnd
rlabel metal1 s 8947 12304 9336 12335 4 gnd
rlabel metal1 s 1167 21544 1556 21575 4 gnd
rlabel metal1 s 1945 16925 2334 16956 4 gnd
rlabel metal1 s 389 1524 778 1555 4 gnd
rlabel metal1 s 18672 10765 19061 10796 4 gnd
rlabel metal1 s 778 20004 1167 20035 4 gnd
rlabel metal1 s 1945 6145 2334 6176 4 gnd
rlabel metal1 s 6224 1525 6613 1556 4 gnd
rlabel metal1 s 3112 9224 3501 9255 4 gnd
rlabel metal1 s 5835 1524 6224 1555 4 gnd
rlabel metal1 s 19061 13844 19450 13875 4 gnd
rlabel metal1 s 6613 -16 7002 15 4 gnd
rlabel metal1 s 13615 12305 14004 12336 4 gnd
rlabel metal1 s 5835 4605 6224 4636 4 gnd
rlabel metal1 s 11670 13845 12059 13876 4 gnd
rlabel metal1 s 5446 10764 5835 10795 4 gnd
rlabel metal1 s 23729 16924 24118 16955 4 gnd
rlabel metal1 s 389 18464 778 18495 4 gnd
rlabel metal1 s 16727 3065 17116 3096 4 gnd
rlabel metal1 s 2334 20005 2723 20036 4 gnd
rlabel metal1 s 12837 7685 13226 7716 4 gnd
rlabel metal1 s 4279 20005 4668 20036 4 gnd
rlabel metal1 s 17505 20004 17894 20035 4 gnd
rlabel metal1 s 389 12304 778 12335 4 gnd
rlabel metal1 s 8947 23085 9336 23116 4 gnd
rlabel metal1 s 7780 15385 8169 15416 4 gnd
rlabel metal1 s 7002 6144 7391 6175 4 gnd
rlabel metal1 s 21395 15384 21784 15415 4 gnd
rlabel metal1 s 11281 12305 11670 12336 4 gnd
rlabel metal1 s 0 18464 389 18495 4 gnd
rlabel metal1 s 5057 4604 5446 4635 4 gnd
rlabel metal1 s 7391 15385 7780 15416 4 gnd
rlabel metal1 s 10892 21544 11281 21575 4 gnd
rlabel metal1 s 6613 13845 7002 13876 4 gnd
rlabel metal1 s 23340 -16 23729 15 4 gnd
rlabel metal1 s 10892 3064 11281 3095 4 gnd
rlabel metal1 s 8169 20004 8558 20035 4 gnd
rlabel metal1 s 6224 6145 6613 6176 4 gnd
rlabel metal1 s 19839 9225 20228 9256 4 gnd
rlabel metal1 s 8947 3064 9336 3095 4 gnd
rlabel metal1 s 2723 6144 3112 6175 4 gnd
rlabel metal1 s 389 12305 778 12336 4 gnd
rlabel metal1 s 7002 15385 7391 15416 4 gnd
rlabel metal1 s 8558 12305 8947 12336 4 gnd
rlabel metal1 s 15560 6145 15949 6176 4 gnd
rlabel metal1 s 19061 12305 19450 12336 4 gnd
rlabel metal1 s 15171 7684 15560 7715 4 gnd
rlabel metal1 s 2334 13844 2723 13875 4 gnd
rlabel metal1 s 12837 1525 13226 1556 4 gnd
rlabel metal1 s 24507 18464 24896 18495 4 gnd
rlabel metal1 s 19839 15384 20228 15415 4 gnd
rlabel metal1 s 15171 21545 15560 21576 4 gnd
rlabel metal1 s 22951 1525 23340 1556 4 gnd
rlabel metal1 s 778 15384 1167 15415 4 gnd
rlabel metal1 s 19450 9225 19839 9256 4 gnd
rlabel metal1 s 5446 24625 5835 24656 4 gnd
rlabel metal1 s 10114 12304 10503 12335 4 gnd
rlabel metal1 s 12837 4604 13226 4635 4 gnd
rlabel metal1 s 19450 20005 19839 20036 4 gnd
rlabel metal1 s 16338 4605 16727 4636 4 gnd
rlabel metal1 s 20617 7684 21006 7715 4 gnd
rlabel metal1 s 3890 13844 4279 13875 4 gnd
rlabel metal1 s 17116 21545 17505 21576 4 gnd
rlabel metal1 s 0 4605 389 4636 4 gnd
rlabel metal1 s 24507 20005 24896 20036 4 gnd
rlabel metal1 s 24507 7685 24896 7716 4 gnd
rlabel metal1 s 1945 1524 2334 1555 4 gnd
rlabel metal1 s 389 6145 778 6176 4 gnd
rlabel metal1 s 16727 7685 17116 7716 4 gnd
rlabel metal1 s 23729 3064 24118 3095 4 gnd
rlabel metal1 s 18283 13845 18672 13876 4 gnd
rlabel metal1 s 15560 18465 15949 18496 4 gnd
rlabel metal1 s 13226 20004 13615 20035 4 gnd
rlabel metal1 s 11281 24625 11670 24656 4 gnd
rlabel metal1 s 3501 10764 3890 10795 4 gnd
rlabel metal1 s 14393 10765 14782 10796 4 gnd
rlabel metal1 s 13226 3064 13615 3095 4 gnd
rlabel metal1 s 2334 16925 2723 16956 4 gnd
rlabel metal1 s 12448 13845 12837 13876 4 gnd
rlabel metal1 s 1945 7685 2334 7716 4 gnd
rlabel metal1 s 2723 15385 3112 15416 4 gnd
rlabel metal1 s 2334 6144 2723 6175 4 gnd
rlabel metal1 s 5835 20004 6224 20035 4 gnd
rlabel metal1 s 1945 4605 2334 4636 4 gnd
rlabel metal1 s 17894 10765 18283 10796 4 gnd
rlabel metal1 s 15560 23084 15949 23115 4 gnd
rlabel metal1 s 0 13845 389 13876 4 gnd
rlabel metal1 s 23340 15384 23729 15415 4 gnd
rlabel metal1 s 2723 -16 3112 15 4 gnd
rlabel metal1 s 24118 23085 24507 23116 4 gnd
rlabel metal1 s 4279 16924 4668 16955 4 gnd
rlabel metal1 s 14782 15385 15171 15416 4 gnd
rlabel metal1 s 13615 4605 14004 4636 4 gnd
rlabel metal1 s 22173 13844 22562 13875 4 gnd
rlabel metal1 s 8947 12305 9336 12336 4 gnd
rlabel metal1 s 12448 9225 12837 9256 4 gnd
rlabel metal1 s 7002 10765 7391 10796 4 gnd
rlabel metal1 s 10892 -16 11281 15 4 gnd
rlabel metal1 s 2723 10765 3112 10796 4 gnd
rlabel metal1 s 7002 16925 7391 16956 4 gnd
rlabel metal1 s 13226 1524 13615 1555 4 gnd
rlabel metal1 s 18283 15384 18672 15415 4 gnd
rlabel metal1 s 12837 13844 13226 13875 4 gnd
rlabel metal1 s 14004 15385 14393 15416 4 gnd
rlabel metal1 s 24118 16924 24507 16955 4 gnd
rlabel metal1 s 9725 10765 10114 10796 4 gnd
rlabel metal1 s 7780 23085 8169 23116 4 gnd
rlabel metal1 s 21006 16924 21395 16955 4 gnd
rlabel metal1 s 21006 23084 21395 23115 4 gnd
rlabel metal1 s 19839 9224 20228 9255 4 gnd
rlabel metal1 s 5057 4605 5446 4636 4 gnd
rlabel metal1 s 10892 9225 11281 9256 4 gnd
rlabel metal1 s 17116 16925 17505 16956 4 gnd
rlabel metal1 s 10503 21545 10892 21576 4 gnd
rlabel metal1 s 9725 15385 10114 15416 4 gnd
rlabel metal1 s 17894 1524 18283 1555 4 gnd
rlabel metal1 s 22173 15385 22562 15416 4 gnd
rlabel metal1 s 22173 1525 22562 1556 4 gnd
rlabel metal1 s 23340 4604 23729 4635 4 gnd
rlabel metal1 s 13226 4604 13615 4635 4 gnd
rlabel metal1 s 24507 21545 24896 21576 4 gnd
rlabel metal1 s 389 16924 778 16955 4 gnd
rlabel metal1 s 22562 4605 22951 4636 4 gnd
rlabel metal1 s 2334 3064 2723 3095 4 gnd
rlabel metal1 s 20617 -16 21006 15 4 gnd
rlabel metal1 s 11670 16924 12059 16955 4 gnd
rlabel metal1 s 6224 13844 6613 13875 4 gnd
rlabel metal1 s 17505 10764 17894 10795 4 gnd
rlabel metal1 s 21395 10765 21784 10796 4 gnd
rlabel metal1 s 19450 15384 19839 15415 4 gnd
rlabel metal1 s 6224 4604 6613 4635 4 gnd
rlabel metal1 s 4279 13844 4668 13875 4 gnd
rlabel metal1 s 15171 12305 15560 12336 4 gnd
rlabel metal1 s 778 20005 1167 20036 4 gnd
rlabel metal1 s 12059 16924 12448 16955 4 gnd
rlabel metal1 s 22951 21544 23340 21575 4 gnd
rlabel metal1 s 21006 9225 21395 9256 4 gnd
rlabel metal1 s 6224 9224 6613 9255 4 gnd
rlabel metal1 s 10114 18465 10503 18496 4 gnd
rlabel metal1 s 4668 16924 5057 16955 4 gnd
rlabel metal1 s 0 12305 389 12336 4 gnd
rlabel metal1 s 5446 16924 5835 16955 4 gnd
rlabel metal1 s 14782 6144 15171 6175 4 gnd
rlabel metal1 s 12837 18464 13226 18495 4 gnd
rlabel metal1 s 5446 9224 5835 9255 4 gnd
rlabel metal1 s 778 21545 1167 21576 4 gnd
rlabel metal1 s 1556 6145 1945 6176 4 gnd
rlabel metal1 s 389 13845 778 13876 4 gnd
rlabel metal1 s 15560 7684 15949 7715 4 gnd
rlabel metal1 s 21784 4605 22173 4636 4 gnd
rlabel metal1 s 19839 7684 20228 7715 4 gnd
rlabel metal1 s 22562 16925 22951 16956 4 gnd
rlabel metal1 s 11281 7684 11670 7715 4 gnd
rlabel metal1 s 23729 13845 24118 13876 4 gnd
rlabel metal1 s 10114 20005 10503 20036 4 gnd
rlabel metal1 s 16727 20005 17116 20036 4 gnd
rlabel metal1 s 3890 7685 4279 7716 4 gnd
rlabel metal1 s 10892 12305 11281 12336 4 gnd
rlabel metal1 s 18672 7684 19061 7715 4 gnd
rlabel metal1 s 5446 16925 5835 16956 4 gnd
rlabel metal1 s 20617 18464 21006 18495 4 gnd
rlabel metal1 s 389 10765 778 10796 4 gnd
rlabel metal1 s 8558 12304 8947 12335 4 gnd
rlabel metal1 s 15949 10765 16338 10796 4 gnd
rlabel metal1 s 24507 16925 24896 16956 4 gnd
rlabel metal1 s 14393 1525 14782 1556 4 gnd
rlabel metal1 s 0 1524 389 1555 4 gnd
rlabel metal1 s 21784 20004 22173 20035 4 gnd
rlabel metal1 s 4279 18464 4668 18495 4 gnd
rlabel metal1 s 18283 7684 18672 7715 4 gnd
rlabel metal1 s 23340 13845 23729 13876 4 gnd
rlabel metal1 s 15560 20004 15949 20035 4 gnd
rlabel metal1 s 5446 21544 5835 21575 4 gnd
rlabel metal1 s 16727 6145 17116 6176 4 gnd
rlabel metal1 s 21784 23085 22173 23116 4 gnd
rlabel metal1 s 8558 3064 8947 3095 4 gnd
rlabel metal1 s 3501 3064 3890 3095 4 gnd
rlabel metal1 s 22173 18465 22562 18496 4 gnd
rlabel metal1 s 19839 7685 20228 7716 4 gnd
rlabel metal1 s 6613 3065 7002 3096 4 gnd
rlabel metal1 s 16338 24625 16727 24656 4 gnd
rlabel metal1 s 14393 13845 14782 13876 4 gnd
rlabel metal1 s 389 13844 778 13875 4 gnd
rlabel metal1 s 19061 1524 19450 1555 4 gnd
rlabel metal1 s 22562 18465 22951 18496 4 gnd
rlabel metal1 s 14004 12305 14393 12336 4 gnd
rlabel metal1 s 4668 9224 5057 9255 4 gnd
rlabel metal1 s 3890 10764 4279 10795 4 gnd
rlabel metal1 s 2334 1525 2723 1556 4 gnd
rlabel metal1 s 22173 16924 22562 16955 4 gnd
rlabel metal1 s 16727 15384 17116 15415 4 gnd
rlabel metal1 s 12059 16925 12448 16956 4 gnd
rlabel metal1 s 4279 1525 4668 1556 4 gnd
rlabel metal1 s 2334 10765 2723 10796 4 gnd
rlabel metal1 s 22951 9224 23340 9255 4 gnd
rlabel metal1 s 8558 21545 8947 21576 4 gnd
rlabel metal1 s 18672 20004 19061 20035 4 gnd
rlabel metal1 s 24507 10764 24896 10795 4 gnd
rlabel metal1 s 10503 13845 10892 13876 4 gnd
rlabel metal1 s 8947 15384 9336 15415 4 gnd
rlabel metal1 s 5057 -16 5446 15 4 gnd
rlabel metal1 s 4279 6144 4668 6175 4 gnd
rlabel metal1 s 3890 18465 4279 18496 4 gnd
rlabel metal1 s 9336 3065 9725 3096 4 gnd
rlabel metal1 s 24507 1524 24896 1555 4 gnd
rlabel metal1 s 14393 18465 14782 18496 4 gnd
rlabel metal1 s 8947 6144 9336 6175 4 gnd
rlabel metal1 s 3890 1525 4279 1556 4 gnd
rlabel metal1 s 17505 7684 17894 7715 4 gnd
rlabel metal1 s 22562 6145 22951 6176 4 gnd
rlabel metal1 s 5835 16925 6224 16956 4 gnd
rlabel metal1 s 15560 15385 15949 15416 4 gnd
rlabel metal1 s 17116 4605 17505 4636 4 gnd
rlabel metal1 s 15560 7685 15949 7716 4 gnd
rlabel metal1 s 11670 3065 12059 3096 4 gnd
rlabel metal1 s 14393 4604 14782 4635 4 gnd
rlabel metal1 s 21784 6144 22173 6175 4 gnd
rlabel metal1 s 778 23084 1167 23115 4 gnd
rlabel metal1 s 8169 20005 8558 20036 4 gnd
rlabel metal1 s 12448 24625 12837 24656 4 gnd
rlabel metal1 s 9336 10764 9725 10795 4 gnd
rlabel metal1 s 9336 12304 9725 12335 4 gnd
rlabel metal1 s 3501 6144 3890 6175 4 gnd
rlabel metal1 s 23340 20004 23729 20035 4 gnd
rlabel metal1 s 22951 3064 23340 3095 4 gnd
rlabel metal1 s 3112 4604 3501 4635 4 gnd
rlabel metal1 s 12059 18465 12448 18496 4 gnd
rlabel metal1 s 7391 4604 7780 4635 4 gnd
rlabel metal1 s 19450 20004 19839 20035 4 gnd
rlabel metal1 s 1167 3065 1556 3096 4 gnd
rlabel metal1 s 13615 1524 14004 1555 4 gnd
rlabel metal1 s 12059 13844 12448 13875 4 gnd
rlabel metal1 s 14004 13844 14393 13875 4 gnd
rlabel metal1 s 24507 7684 24896 7715 4 gnd
rlabel metal1 s 12059 20005 12448 20036 4 gnd
rlabel metal1 s 4668 23085 5057 23116 4 gnd
rlabel metal1 s 17505 23085 17894 23116 4 gnd
rlabel metal1 s 19450 13845 19839 13876 4 gnd
rlabel metal1 s 3112 10764 3501 10795 4 gnd
rlabel metal1 s 5835 13844 6224 13875 4 gnd
rlabel metal1 s 18283 6145 18672 6176 4 gnd
rlabel metal1 s 6224 15384 6613 15415 4 gnd
rlabel metal1 s 10892 21545 11281 21576 4 gnd
rlabel metal1 s 12448 12304 12837 12335 4 gnd
rlabel metal1 s 10114 20004 10503 20035 4 gnd
rlabel metal1 s 5446 20005 5835 20036 4 gnd
rlabel metal1 s 778 13845 1167 13876 4 gnd
rlabel metal1 s 14004 10764 14393 10795 4 gnd
rlabel metal1 s 7780 16924 8169 16955 4 gnd
rlabel metal1 s 3890 4604 4279 4635 4 gnd
rlabel metal1 s 8169 13844 8558 13875 4 gnd
rlabel metal1 s 0 16925 389 16956 4 gnd
rlabel metal1 s 0 7685 389 7716 4 gnd
rlabel metal1 s 21006 -16 21395 15 4 gnd
rlabel metal1 s 17894 -16 18283 15 4 gnd
rlabel metal1 s 22951 10764 23340 10795 4 gnd
rlabel metal1 s 12059 21545 12448 21576 4 gnd
rlabel metal1 s 1556 -16 1945 15 4 gnd
rlabel metal1 s 11281 13845 11670 13876 4 gnd
rlabel metal1 s 778 1524 1167 1555 4 gnd
rlabel metal1 s 16727 1524 17116 1555 4 gnd
rlabel metal1 s 24507 16924 24896 16955 4 gnd
rlabel metal1 s 18283 16924 18672 16955 4 gnd
rlabel metal1 s 20617 21544 21006 21575 4 gnd
rlabel metal1 s 1945 -16 2334 15 4 gnd
rlabel metal1 s 2723 7684 3112 7715 4 gnd
rlabel metal1 s 17894 16925 18283 16956 4 gnd
rlabel metal1 s 8947 16924 9336 16955 4 gnd
rlabel metal1 s 24118 6144 24507 6175 4 gnd
rlabel metal1 s 21395 16924 21784 16955 4 gnd
rlabel metal1 s 14393 6145 14782 6176 4 gnd
rlabel metal1 s 778 3065 1167 3096 4 gnd
rlabel metal1 s 21006 6145 21395 6176 4 gnd
rlabel metal1 s 2334 7684 2723 7715 4 gnd
rlabel metal1 s 24507 6145 24896 6176 4 gnd
rlabel metal1 s 7002 21545 7391 21576 4 gnd
rlabel metal1 s 10503 18465 10892 18496 4 gnd
rlabel metal1 s 7002 20005 7391 20036 4 gnd
rlabel metal1 s 21784 13845 22173 13876 4 gnd
rlabel metal1 s 10503 12305 10892 12336 4 gnd
rlabel metal1 s 1945 10764 2334 10795 4 gnd
rlabel metal1 s 12059 3064 12448 3095 4 gnd
rlabel metal1 s 12448 23085 12837 23116 4 gnd
rlabel metal1 s 22951 4605 23340 4636 4 gnd
rlabel metal1 s 1167 9224 1556 9255 4 gnd
rlabel metal1 s 7002 7684 7391 7715 4 gnd
rlabel metal1 s 18672 9224 19061 9255 4 gnd
rlabel metal1 s 10114 24625 10503 24656 4 gnd
rlabel metal1 s 1556 6144 1945 6175 4 gnd
rlabel metal1 s 21006 9224 21395 9255 4 gnd
rlabel metal1 s 16338 13845 16727 13876 4 gnd
rlabel metal1 s 22173 4605 22562 4636 4 gnd
rlabel metal1 s 21395 18465 21784 18496 4 gnd
rlabel metal1 s 4279 12304 4668 12335 4 gnd
rlabel metal1 s 8947 21545 9336 21576 4 gnd
rlabel metal1 s 19839 21544 20228 21575 4 gnd
rlabel metal1 s 17894 16924 18283 16955 4 gnd
rlabel metal1 s 12448 7684 12837 7715 4 gnd
rlabel metal1 s 5446 -16 5835 15 4 gnd
rlabel metal1 s 11281 23085 11670 23116 4 gnd
rlabel metal1 s 8558 15385 8947 15416 4 gnd
rlabel metal1 s 16727 10765 17116 10796 4 gnd
rlabel metal1 s 22173 15384 22562 15415 4 gnd
rlabel metal1 s 16727 20004 17116 20035 4 gnd
rlabel metal1 s 7780 10765 8169 10796 4 gnd
rlabel metal1 s 11281 3065 11670 3096 4 gnd
rlabel metal1 s 2334 6145 2723 6176 4 gnd
rlabel metal1 s 0 15384 389 15415 4 gnd
rlabel metal1 s 18672 15385 19061 15416 4 gnd
rlabel metal1 s 15949 9224 16338 9255 4 gnd
rlabel metal1 s 17505 12305 17894 12336 4 gnd
rlabel metal1 s 1556 13845 1945 13876 4 gnd
rlabel metal1 s 6224 23084 6613 23115 4 gnd
rlabel metal1 s 20228 13845 20617 13876 4 gnd
rlabel metal1 s 21006 16925 21395 16956 4 gnd
rlabel metal1 s 10892 16924 11281 16955 4 gnd
rlabel metal1 s 20228 9224 20617 9255 4 gnd
rlabel metal1 s 1556 7684 1945 7715 4 gnd
rlabel metal1 s 5057 9224 5446 9255 4 gnd
rlabel metal1 s 12837 16925 13226 16956 4 gnd
rlabel metal1 s 22562 23084 22951 23115 4 gnd
rlabel metal1 s 8947 7685 9336 7716 4 gnd
rlabel metal1 s 15560 12304 15949 12335 4 gnd
rlabel metal1 s 15171 10764 15560 10795 4 gnd
rlabel metal1 s 22562 -16 22951 15 4 gnd
rlabel metal1 s 16727 9225 17116 9256 4 gnd
rlabel metal1 s 6613 18465 7002 18496 4 gnd
rlabel metal1 s 5446 15384 5835 15415 4 gnd
rlabel metal1 s 9725 21544 10114 21575 4 gnd
rlabel metal1 s 7002 3065 7391 3096 4 gnd
rlabel metal1 s 3890 6144 4279 6175 4 gnd
rlabel metal1 s 9725 9225 10114 9256 4 gnd
rlabel metal1 s 3890 3064 4279 3095 4 gnd
rlabel metal1 s 778 6144 1167 6175 4 gnd
rlabel metal1 s 8169 9225 8558 9256 4 gnd
rlabel metal1 s 5446 6144 5835 6175 4 gnd
rlabel metal1 s 1945 24625 2334 24656 4 gnd
rlabel metal1 s 1167 20005 1556 20036 4 gnd
rlabel metal1 s 22562 7684 22951 7715 4 gnd
rlabel metal1 s 10114 23084 10503 23115 4 gnd
rlabel metal1 s 1167 3064 1556 3095 4 gnd
rlabel metal1 s 10892 10764 11281 10795 4 gnd
rlabel metal1 s 7002 13845 7391 13876 4 gnd
rlabel metal1 s 2723 15384 3112 15415 4 gnd
rlabel metal1 s 15171 23085 15560 23116 4 gnd
rlabel metal1 s 0 10764 389 10795 4 gnd
rlabel metal1 s 20617 24625 21006 24656 4 gnd
rlabel metal1 s 19061 13845 19450 13876 4 gnd
rlabel metal1 s 14004 16925 14393 16956 4 gnd
rlabel metal1 s 16338 9225 16727 9256 4 gnd
rlabel metal1 s 11670 24625 12059 24656 4 gnd
rlabel metal1 s 9336 9224 9725 9255 4 gnd
rlabel metal1 s 19450 4604 19839 4635 4 gnd
rlabel metal1 s 22562 18464 22951 18495 4 gnd
rlabel metal1 s 0 24625 389 24656 4 gnd
rlabel metal1 s 20617 9225 21006 9256 4 gnd
rlabel metal1 s 22951 16925 23340 16956 4 gnd
rlabel metal1 s 8947 18465 9336 18496 4 gnd
rlabel metal1 s 7391 7684 7780 7715 4 gnd
rlabel metal1 s 5835 12304 6224 12335 4 gnd
rlabel metal1 s 13226 15385 13615 15416 4 gnd
rlabel metal1 s 24507 3065 24896 3096 4 gnd
rlabel metal1 s 17505 15385 17894 15416 4 gnd
rlabel metal1 s 9336 16924 9725 16955 4 gnd
rlabel metal1 s 24118 20004 24507 20035 4 gnd
rlabel metal1 s 17894 4605 18283 4636 4 gnd
rlabel metal1 s 9725 9224 10114 9255 4 gnd
rlabel metal1 s 23729 15385 24118 15416 4 gnd
rlabel metal1 s 24507 23084 24896 23115 4 gnd
rlabel metal1 s 10503 6145 10892 6176 4 gnd
rlabel metal1 s 6224 7685 6613 7716 4 gnd
rlabel metal1 s 17505 13844 17894 13875 4 gnd
rlabel metal1 s 1167 6144 1556 6175 4 gnd
rlabel metal1 s 18283 24625 18672 24656 4 gnd
rlabel metal1 s 14782 9225 15171 9256 4 gnd
rlabel metal1 s 1167 12305 1556 12336 4 gnd
rlabel metal1 s 389 10764 778 10795 4 gnd
rlabel metal1 s 4668 -16 5057 15 4 gnd
rlabel metal1 s 1167 4605 1556 4636 4 gnd
rlabel metal1 s 15560 4604 15949 4635 4 gnd
rlabel metal1 s 12837 -16 13226 15 4 gnd
rlabel metal1 s 6224 13845 6613 13876 4 gnd
rlabel metal1 s 21784 18464 22173 18495 4 gnd
rlabel metal1 s 12448 20004 12837 20035 4 gnd
rlabel metal1 s 20617 1525 21006 1556 4 gnd
rlabel metal1 s 24507 12304 24896 12335 4 gnd
rlabel metal1 s 15560 21545 15949 21576 4 gnd
rlabel metal1 s 17116 3064 17505 3095 4 gnd
rlabel metal1 s 3112 13845 3501 13876 4 gnd
rlabel metal1 s 1556 12304 1945 12335 4 gnd
rlabel metal1 s 21006 12304 21395 12335 4 gnd
rlabel metal1 s 24118 15384 24507 15415 4 gnd
rlabel metal1 s 9725 13844 10114 13875 4 gnd
rlabel metal1 s 6224 23085 6613 23116 4 gnd
rlabel metal1 s 22562 12304 22951 12335 4 gnd
rlabel metal1 s 5446 23084 5835 23115 4 gnd
rlabel metal1 s 1167 1524 1556 1555 4 gnd
rlabel metal1 s 12448 23084 12837 23115 4 gnd
rlabel metal1 s 12059 18464 12448 18495 4 gnd
rlabel metal1 s 2334 18464 2723 18495 4 gnd
rlabel metal1 s 12448 9224 12837 9255 4 gnd
rlabel metal1 s 8947 20004 9336 20035 4 gnd
rlabel metal1 s 15560 9225 15949 9256 4 gnd
rlabel metal1 s 4279 15385 4668 15416 4 gnd
rlabel metal1 s 7002 18465 7391 18496 4 gnd
rlabel metal1 s 15171 20004 15560 20035 4 gnd
rlabel metal1 s 7002 12305 7391 12336 4 gnd
rlabel metal1 s 7002 9224 7391 9255 4 gnd
rlabel metal1 s 7780 1524 8169 1555 4 gnd
rlabel metal1 s 3112 1525 3501 1556 4 gnd
rlabel metal1 s 13615 1525 14004 1556 4 gnd
rlabel metal1 s 10114 9224 10503 9255 4 gnd
rlabel metal1 s 11281 7685 11670 7716 4 gnd
rlabel metal1 s 11281 13844 11670 13875 4 gnd
rlabel metal1 s 14393 -16 14782 15 4 gnd
rlabel metal1 s 389 9224 778 9255 4 gnd
rlabel metal1 s 7391 10764 7780 10795 4 gnd
rlabel metal1 s 19450 7685 19839 7716 4 gnd
rlabel metal1 s 2723 16925 3112 16956 4 gnd
rlabel metal1 s 21006 18464 21395 18495 4 gnd
rlabel metal1 s 6613 21545 7002 21576 4 gnd
rlabel metal1 s 12059 10765 12448 10796 4 gnd
rlabel metal1 s 2334 24625 2723 24656 4 gnd
rlabel metal1 s 20228 16924 20617 16955 4 gnd
rlabel metal1 s 9725 24625 10114 24656 4 gnd
rlabel metal1 s 11670 18464 12059 18495 4 gnd
rlabel metal1 s 3112 18465 3501 18496 4 gnd
rlabel metal1 s 8169 23084 8558 23115 4 gnd
rlabel metal1 s 6613 4604 7002 4635 4 gnd
rlabel metal1 s 17116 16924 17505 16955 4 gnd
rlabel metal1 s 10114 1525 10503 1556 4 gnd
rlabel metal1 s 778 12304 1167 12335 4 gnd
rlabel metal1 s 12448 1524 12837 1555 4 gnd
rlabel metal1 s 2334 7685 2723 7716 4 gnd
rlabel metal1 s 10503 3064 10892 3095 4 gnd
rlabel metal1 s 5446 7685 5835 7716 4 gnd
rlabel metal1 s 12837 7684 13226 7715 4 gnd
rlabel metal1 s 15171 21544 15560 21575 4 gnd
rlabel metal1 s 15171 7685 15560 7716 4 gnd
rlabel metal1 s 24118 1525 24507 1556 4 gnd
rlabel metal1 s 4279 12305 4668 12336 4 gnd
rlabel metal1 s 16338 6145 16727 6176 4 gnd
rlabel metal1 s 6224 6144 6613 6175 4 gnd
rlabel metal1 s 16338 18465 16727 18496 4 gnd
rlabel metal1 s 3501 16924 3890 16955 4 gnd
rlabel metal1 s 23729 10764 24118 10795 4 gnd
rlabel metal1 s 15171 20005 15560 20036 4 gnd
rlabel metal1 s 16727 21544 17116 21575 4 gnd
rlabel metal1 s 6613 10765 7002 10796 4 gnd
rlabel metal1 s 16338 9224 16727 9255 4 gnd
rlabel metal1 s 24118 7684 24507 7715 4 gnd
rlabel metal1 s 12837 12305 13226 12336 4 gnd
rlabel metal1 s 5057 7685 5446 7716 4 gnd
rlabel metal1 s 15949 6144 16338 6175 4 gnd
rlabel metal1 s 8558 9225 8947 9256 4 gnd
rlabel metal1 s 6613 24625 7002 24656 4 gnd
rlabel metal1 s 8558 1524 8947 1555 4 gnd
rlabel metal1 s 19450 3065 19839 3096 4 gnd
rlabel metal1 s 1556 15385 1945 15416 4 gnd
rlabel metal1 s 14782 20004 15171 20035 4 gnd
rlabel metal1 s 21006 13844 21395 13875 4 gnd
rlabel metal1 s 10892 23084 11281 23115 4 gnd
rlabel metal1 s 9336 13844 9725 13875 4 gnd
rlabel metal1 s 12837 9224 13226 9255 4 gnd
rlabel metal1 s 24118 15385 24507 15416 4 gnd
rlabel metal1 s 3890 6145 4279 6176 4 gnd
rlabel metal1 s 5057 20004 5446 20035 4 gnd
rlabel metal1 s 19839 13844 20228 13875 4 gnd
rlabel metal1 s 23729 4604 24118 4635 4 gnd
rlabel metal1 s 8558 21544 8947 21575 4 gnd
rlabel metal1 s 3501 20004 3890 20035 4 gnd
rlabel metal1 s 7002 3064 7391 3095 4 gnd
rlabel metal1 s 1556 15384 1945 15415 4 gnd
rlabel metal1 s 11670 7684 12059 7715 4 gnd
rlabel metal1 s 19839 18465 20228 18496 4 gnd
rlabel metal1 s 23729 9225 24118 9256 4 gnd
rlabel metal1 s 17505 18465 17894 18496 4 gnd
rlabel metal1 s 21784 16925 22173 16956 4 gnd
rlabel metal1 s 11281 15384 11670 15415 4 gnd
rlabel metal1 s 7391 9225 7780 9256 4 gnd
rlabel metal1 s 5446 12304 5835 12335 4 gnd
rlabel metal1 s 21006 18465 21395 18496 4 gnd
rlabel metal1 s 22951 1524 23340 1555 4 gnd
rlabel metal1 s 16338 3064 16727 3095 4 gnd
rlabel metal1 s 22951 20005 23340 20036 4 gnd
rlabel metal1 s 1556 23085 1945 23116 4 gnd
rlabel metal1 s 20228 23085 20617 23116 4 gnd
rlabel metal1 s 14782 10765 15171 10796 4 gnd
rlabel metal1 s 3890 7684 4279 7715 4 gnd
rlabel metal1 s 14004 21544 14393 21575 4 gnd
rlabel metal1 s 7780 7685 8169 7716 4 gnd
rlabel metal1 s 22562 21545 22951 21576 4 gnd
rlabel metal1 s 8558 10765 8947 10796 4 gnd
rlabel metal1 s 5446 15385 5835 15416 4 gnd
rlabel metal1 s 23340 1525 23729 1556 4 gnd
rlabel metal1 s 389 21545 778 21576 4 gnd
rlabel metal1 s 3890 23084 4279 23115 4 gnd
rlabel metal1 s 5446 3064 5835 3095 4 gnd
rlabel metal1 s 2723 13845 3112 13876 4 gnd
rlabel metal1 s 17505 24625 17894 24656 4 gnd
rlabel metal1 s 16338 1525 16727 1556 4 gnd
rlabel metal1 s 5835 20005 6224 20036 4 gnd
rlabel metal1 s 22173 -16 22562 15 4 gnd
rlabel metal1 s 5057 20005 5446 20036 4 gnd
rlabel metal1 s 5057 18465 5446 18496 4 gnd
rlabel metal1 s 19839 10764 20228 10795 4 gnd
rlabel metal1 s 19061 23084 19450 23115 4 gnd
rlabel metal1 s 9336 7684 9725 7715 4 gnd
rlabel metal1 s 22562 13844 22951 13875 4 gnd
rlabel metal1 s 20617 12304 21006 12335 4 gnd
rlabel metal1 s 14393 21544 14782 21575 4 gnd
rlabel metal1 s 5057 6144 5446 6175 4 gnd
rlabel metal1 s 5446 6145 5835 6176 4 gnd
rlabel metal1 s 21006 23085 21395 23116 4 gnd
rlabel metal1 s 15560 12305 15949 12336 4 gnd
rlabel metal1 s 10892 15385 11281 15416 4 gnd
rlabel metal1 s 11670 12304 12059 12335 4 gnd
rlabel metal1 s 15171 10765 15560 10796 4 gnd
rlabel metal1 s 9336 24625 9725 24656 4 gnd
rlabel metal1 s 8947 7684 9336 7715 4 gnd
rlabel metal1 s 23729 24625 24118 24656 4 gnd
rlabel metal1 s 1945 6144 2334 6175 4 gnd
rlabel metal1 s 24118 21545 24507 21576 4 gnd
rlabel metal1 s 3112 23085 3501 23116 4 gnd
rlabel metal1 s 1556 23084 1945 23115 4 gnd
rlabel metal1 s 16727 16925 17116 16956 4 gnd
rlabel metal1 s 0 20005 389 20036 4 gnd
rlabel metal1 s 22562 6144 22951 6175 4 gnd
rlabel metal1 s 7391 13845 7780 13876 4 gnd
rlabel metal1 s 15560 23085 15949 23116 4 gnd
rlabel metal1 s 11281 1524 11670 1555 4 gnd
rlabel metal1 s 5057 1525 5446 1556 4 gnd
rlabel metal1 s 3112 24625 3501 24656 4 gnd
rlabel metal1 s 1945 3065 2334 3096 4 gnd
rlabel metal1 s 19061 24625 19450 24656 4 gnd
rlabel metal1 s 778 9225 1167 9256 4 gnd
rlabel metal1 s 3890 13845 4279 13876 4 gnd
rlabel metal1 s 9725 21545 10114 21576 4 gnd
rlabel metal1 s 11281 15385 11670 15416 4 gnd
rlabel metal1 s 12837 23085 13226 23116 4 gnd
rlabel metal1 s 1556 1524 1945 1555 4 gnd
rlabel metal1 s 21395 13845 21784 13876 4 gnd
rlabel metal1 s 19061 6145 19450 6176 4 gnd
rlabel metal1 s 22173 21545 22562 21576 4 gnd
rlabel metal1 s 4668 7684 5057 7715 4 gnd
rlabel metal1 s 11281 4604 11670 4635 4 gnd
rlabel metal1 s 16727 18464 17116 18495 4 gnd
rlabel metal1 s 3501 -16 3890 15 4 gnd
rlabel metal1 s 9336 1525 9725 1556 4 gnd
rlabel metal1 s 24507 6144 24896 6175 4 gnd
rlabel metal1 s 3112 23084 3501 23115 4 gnd
rlabel metal1 s 13226 1525 13615 1556 4 gnd
rlabel metal1 s 20617 16925 21006 16956 4 gnd
rlabel metal1 s 2334 20004 2723 20035 4 gnd
rlabel metal1 s 15171 13845 15560 13876 4 gnd
rlabel metal1 s 17116 10764 17505 10795 4 gnd
rlabel metal1 s 10503 21544 10892 21575 4 gnd
rlabel metal1 s 12837 6144 13226 6175 4 gnd
rlabel metal1 s 23340 3065 23729 3096 4 gnd
rlabel metal1 s 5057 3064 5446 3095 4 gnd
rlabel metal1 s 11281 1525 11670 1556 4 gnd
rlabel metal1 s 10892 20005 11281 20036 4 gnd
rlabel metal1 s 15949 6145 16338 6176 4 gnd
rlabel metal1 s 14782 12304 15171 12335 4 gnd
rlabel metal1 s 5446 1525 5835 1556 4 gnd
rlabel metal1 s 20228 12305 20617 12336 4 gnd
rlabel metal1 s 21395 -16 21784 15 4 gnd
rlabel metal1 s 10114 9225 10503 9256 4 gnd
rlabel metal1 s 2334 10764 2723 10795 4 gnd
rlabel metal1 s 2723 18464 3112 18495 4 gnd
rlabel metal1 s 18672 3065 19061 3096 4 gnd
rlabel metal1 s 2334 23084 2723 23115 4 gnd
rlabel metal1 s 13615 24625 14004 24656 4 gnd
rlabel metal1 s 16727 18465 17116 18496 4 gnd
rlabel metal1 s 13226 23084 13615 23115 4 gnd
rlabel metal1 s 9725 6144 10114 6175 4 gnd
rlabel metal1 s 5057 7684 5446 7715 4 gnd
rlabel metal1 s 12448 10764 12837 10795 4 gnd
rlabel metal1 s 11670 12305 12059 12336 4 gnd
rlabel metal1 s 24118 12304 24507 12335 4 gnd
rlabel metal1 s 5446 1524 5835 1555 4 gnd
rlabel metal1 s 5835 23085 6224 23116 4 gnd
rlabel metal1 s 15560 3065 15949 3096 4 gnd
rlabel metal1 s 8169 -16 8558 15 4 gnd
rlabel metal1 s 2334 21544 2723 21575 4 gnd
rlabel metal1 s 14393 1524 14782 1555 4 gnd
rlabel metal1 s 15949 9225 16338 9256 4 gnd
rlabel metal1 s 9336 4604 9725 4635 4 gnd
rlabel metal1 s 13615 6144 14004 6175 4 gnd
rlabel metal1 s 7391 9224 7780 9255 4 gnd
rlabel metal1 s 12059 15385 12448 15416 4 gnd
rlabel metal1 s 1945 23085 2334 23116 4 gnd
rlabel metal1 s 15560 21544 15949 21575 4 gnd
rlabel metal1 s 8169 12305 8558 12336 4 gnd
rlabel metal1 s 15171 18464 15560 18495 4 gnd
rlabel metal1 s 17505 7685 17894 7716 4 gnd
rlabel metal1 s 12837 4605 13226 4636 4 gnd
rlabel metal1 s 7780 21545 8169 21576 4 gnd
rlabel metal1 s 20228 15385 20617 15416 4 gnd
rlabel metal1 s 21006 6144 21395 6175 4 gnd
rlabel metal1 s 20617 1524 21006 1555 4 gnd
rlabel metal1 s 10114 4605 10503 4636 4 gnd
rlabel metal1 s 5446 4604 5835 4635 4 gnd
rlabel metal1 s 13226 21544 13615 21575 4 gnd
rlabel metal1 s 15171 13844 15560 13875 4 gnd
rlabel metal1 s 8947 13844 9336 13875 4 gnd
rlabel metal1 s 10892 20004 11281 20035 4 gnd
rlabel metal1 s 778 24625 1167 24656 4 gnd
rlabel metal1 s 10503 1525 10892 1556 4 gnd
rlabel metal1 s 17116 12304 17505 12335 4 gnd
rlabel metal1 s 22951 13844 23340 13875 4 gnd
rlabel metal1 s 15171 -16 15560 15 4 gnd
rlabel metal1 s 6613 15385 7002 15416 4 gnd
rlabel metal1 s 17894 9225 18283 9256 4 gnd
rlabel metal1 s 14782 -16 15171 15 4 gnd
rlabel metal1 s 13615 6145 14004 6176 4 gnd
rlabel metal1 s 1556 24625 1945 24656 4 gnd
rlabel metal1 s 20617 23085 21006 23116 4 gnd
rlabel metal1 s 8947 4604 9336 4635 4 gnd
rlabel metal1 s 1556 7685 1945 7716 4 gnd
rlabel metal1 s 2723 9224 3112 9255 4 gnd
rlabel metal1 s 23729 20004 24118 20035 4 gnd
rlabel metal1 s 11281 18464 11670 18495 4 gnd
rlabel metal1 s 19061 16925 19450 16956 4 gnd
rlabel metal1 s 18672 24625 19061 24656 4 gnd
rlabel metal1 s 14393 3065 14782 3096 4 gnd
rlabel metal1 s 19450 7684 19839 7715 4 gnd
rlabel metal1 s 12448 13844 12837 13875 4 gnd
rlabel metal1 s 10892 13844 11281 13875 4 gnd
rlabel metal1 s 5446 4605 5835 4636 4 gnd
rlabel metal1 s 8169 7685 8558 7716 4 gnd
rlabel metal1 s 9725 4605 10114 4636 4 gnd
rlabel metal1 s 19061 16924 19450 16955 4 gnd
rlabel metal1 s 15949 20004 16338 20035 4 gnd
rlabel metal1 s 10114 13845 10503 13876 4 gnd
rlabel metal1 s 1167 13845 1556 13876 4 gnd
rlabel metal1 s 17116 13845 17505 13876 4 gnd
rlabel metal1 s 19450 15385 19839 15416 4 gnd
rlabel metal1 s 17894 18464 18283 18495 4 gnd
rlabel metal1 s 22173 18464 22562 18495 4 gnd
rlabel metal1 s 23729 7685 24118 7716 4 gnd
rlabel metal1 s 15560 -16 15949 15 4 gnd
rlabel metal1 s 15171 16925 15560 16956 4 gnd
rlabel metal1 s 16338 21544 16727 21575 4 gnd
rlabel metal1 s 14782 13844 15171 13875 4 gnd
rlabel metal1 s 8947 4605 9336 4636 4 gnd
rlabel metal1 s 13615 7684 14004 7715 4 gnd
rlabel metal1 s 2723 21544 3112 21575 4 gnd
rlabel metal1 s 14782 18465 15171 18496 4 gnd
rlabel metal1 s 16727 13844 17116 13875 4 gnd
rlabel metal1 s 18283 6144 18672 6175 4 gnd
rlabel metal1 s 24118 9224 24507 9255 4 gnd
rlabel metal1 s 20617 3065 21006 3096 4 gnd
rlabel metal1 s 14782 16925 15171 16956 4 gnd
rlabel metal1 s 23729 12305 24118 12336 4 gnd
rlabel metal1 s 19450 6145 19839 6176 4 gnd
rlabel metal1 s 8947 6145 9336 6176 4 gnd
rlabel metal1 s 21006 24625 21395 24656 4 gnd
rlabel metal1 s 12448 16924 12837 16955 4 gnd
rlabel metal1 s 14004 16924 14393 16955 4 gnd
rlabel metal1 s 22951 13845 23340 13876 4 gnd
rlabel metal1 s 0 18465 389 18496 4 gnd
rlabel metal1 s 11670 20004 12059 20035 4 gnd
rlabel metal1 s 22173 10764 22562 10795 4 gnd
rlabel metal1 s 17894 12304 18283 12335 4 gnd
rlabel metal1 s 0 23085 389 23116 4 gnd
rlabel metal1 s 12448 3064 12837 3095 4 gnd
rlabel metal1 s 7391 21545 7780 21576 4 gnd
rlabel metal1 s 20228 9225 20617 9256 4 gnd
rlabel metal1 s 7780 21544 8169 21575 4 gnd
rlabel metal1 s 7780 13844 8169 13875 4 gnd
rlabel metal1 s 2334 12305 2723 12336 4 gnd
rlabel metal1 s 12448 18464 12837 18495 4 gnd
rlabel metal1 s 7391 1525 7780 1556 4 gnd
rlabel metal1 s 21395 21545 21784 21576 4 gnd
rlabel metal1 s 0 7684 389 7715 4 gnd
rlabel metal1 s 17116 9224 17505 9255 4 gnd
rlabel metal1 s 20228 13844 20617 13875 4 gnd
rlabel metal1 s 3112 -16 3501 15 4 gnd
rlabel metal1 s 17505 4605 17894 4636 4 gnd
rlabel metal1 s 5835 10764 6224 10795 4 gnd
rlabel metal1 s 14393 6144 14782 6175 4 gnd
rlabel metal1 s 8947 24625 9336 24656 4 gnd
rlabel metal1 s 7002 18464 7391 18495 4 gnd
rlabel metal1 s 12059 4605 12448 4636 4 gnd
rlabel metal1 s 5835 12305 6224 12336 4 gnd
rlabel metal1 s 14004 9225 14393 9256 4 gnd
rlabel metal1 s 17894 15384 18283 15415 4 gnd
rlabel metal1 s 1556 20004 1945 20035 4 gnd
rlabel metal1 s 778 21544 1167 21575 4 gnd
rlabel metal1 s 16338 -16 16727 15 4 gnd
rlabel metal1 s 4279 7685 4668 7716 4 gnd
rlabel metal1 s 10114 7684 10503 7715 4 gnd
rlabel metal1 s 19450 21544 19839 21575 4 gnd
rlabel metal1 s 10114 6144 10503 6175 4 gnd
rlabel metal1 s 4668 21545 5057 21576 4 gnd
rlabel metal1 s 3501 1524 3890 1555 4 gnd
rlabel metal1 s 22951 -16 23340 15 4 gnd
rlabel metal1 s 10114 4604 10503 4635 4 gnd
rlabel metal1 s 5057 18464 5446 18495 4 gnd
rlabel metal1 s 13615 21545 14004 21576 4 gnd
rlabel metal1 s 19450 23084 19839 23115 4 gnd
rlabel metal1 s 5057 23084 5446 23115 4 gnd
rlabel metal1 s 19061 18464 19450 18495 4 gnd
rlabel metal1 s 7780 16925 8169 16956 4 gnd
rlabel metal1 s 19839 6145 20228 6176 4 gnd
rlabel metal1 s 20228 10764 20617 10795 4 gnd
rlabel metal1 s 7391 15384 7780 15415 4 gnd
rlabel metal1 s 3501 18464 3890 18495 4 gnd
rlabel metal1 s 1556 18465 1945 18496 4 gnd
rlabel metal1 s 15171 1525 15560 1556 4 gnd
rlabel metal1 s 10892 1525 11281 1556 4 gnd
rlabel metal1 s 1945 15385 2334 15416 4 gnd
rlabel metal1 s 5446 3065 5835 3096 4 gnd
rlabel metal1 s 7002 15384 7391 15415 4 gnd
rlabel metal1 s 10114 10765 10503 10796 4 gnd
rlabel metal1 s 14004 10765 14393 10796 4 gnd
rlabel metal1 s 19839 1524 20228 1555 4 gnd
rlabel metal1 s 16338 12305 16727 12336 4 gnd
rlabel metal1 s 20228 15384 20617 15415 4 gnd
rlabel metal1 s 389 20005 778 20036 4 gnd
rlabel metal1 s 12448 7685 12837 7716 4 gnd
rlabel metal1 s 389 3065 778 3096 4 gnd
rlabel metal1 s 18672 20005 19061 20036 4 gnd
rlabel metal1 s 18283 9224 18672 9255 4 gnd
rlabel metal1 s 19839 20004 20228 20035 4 gnd
rlabel metal1 s 22173 20004 22562 20035 4 gnd
rlabel metal1 s 3890 12305 4279 12336 4 gnd
rlabel metal1 s 5835 3064 6224 3095 4 gnd
rlabel metal1 s 17894 7684 18283 7715 4 gnd
rlabel metal1 s 1556 16925 1945 16956 4 gnd
rlabel metal1 s 18672 12304 19061 12335 4 gnd
rlabel metal1 s 2334 13845 2723 13876 4 gnd
rlabel metal1 s 16338 3065 16727 3096 4 gnd
rlabel metal1 s 2334 4605 2723 4636 4 gnd
rlabel metal1 s 9725 10764 10114 10795 4 gnd
rlabel metal1 s 10114 16924 10503 16955 4 gnd
rlabel metal1 s 1167 21545 1556 21576 4 gnd
rlabel metal1 s 8169 10764 8558 10795 4 gnd
rlabel metal1 s 10892 15384 11281 15415 4 gnd
rlabel metal1 s 12448 4605 12837 4636 4 gnd
rlabel metal1 s 13226 6144 13615 6175 4 gnd
rlabel metal1 s 1167 12304 1556 12335 4 gnd
rlabel metal1 s 22562 20004 22951 20035 4 gnd
rlabel metal1 s 18283 3064 18672 3095 4 gnd
rlabel metal1 s 11281 23084 11670 23115 4 gnd
rlabel metal1 s 16338 13844 16727 13875 4 gnd
rlabel metal1 s 7391 18464 7780 18495 4 gnd
rlabel metal1 s 17894 3065 18283 3096 4 gnd
rlabel metal1 s 7002 13844 7391 13875 4 gnd
rlabel metal1 s 15949 7684 16338 7715 4 gnd
rlabel metal1 s 5057 10765 5446 10796 4 gnd
rlabel metal1 s 778 15385 1167 15416 4 gnd
rlabel metal1 s 22951 15385 23340 15416 4 gnd
rlabel metal1 s 3112 20004 3501 20035 4 gnd
rlabel metal1 s 1945 18464 2334 18495 4 gnd
rlabel metal1 s 7780 -16 8169 15 4 gnd
rlabel metal1 s 13226 9225 13615 9256 4 gnd
rlabel metal1 s 8558 15384 8947 15415 4 gnd
rlabel metal1 s 16338 10764 16727 10795 4 gnd
rlabel metal1 s 14004 20005 14393 20036 4 gnd
rlabel metal1 s 19061 10765 19450 10796 4 gnd
rlabel metal1 s 1167 4604 1556 4635 4 gnd
rlabel metal1 s 0 10765 389 10796 4 gnd
rlabel metal1 s 23340 9224 23729 9255 4 gnd
rlabel metal1 s 4279 4605 4668 4636 4 gnd
rlabel metal1 s 0 16924 389 16955 4 gnd
rlabel metal1 s 4279 13845 4668 13876 4 gnd
rlabel metal1 s 20617 6145 21006 6176 4 gnd
rlabel metal1 s 12448 15384 12837 15415 4 gnd
rlabel metal1 s 17116 18465 17505 18496 4 gnd
rlabel metal1 s 21395 20005 21784 20036 4 gnd
rlabel metal1 s 17894 15385 18283 15416 4 gnd
rlabel metal1 s 19839 23084 20228 23115 4 gnd
rlabel metal1 s 14393 3064 14782 3095 4 gnd
rlabel metal1 s 778 18464 1167 18495 4 gnd
rlabel metal1 s 10114 6145 10503 6176 4 gnd
rlabel metal1 s 12059 24625 12448 24656 4 gnd
rlabel metal1 s 14393 20004 14782 20035 4 gnd
rlabel metal1 s 4279 18465 4668 18496 4 gnd
rlabel metal1 s 19061 9224 19450 9255 4 gnd
rlabel metal1 s 19450 16925 19839 16956 4 gnd
rlabel metal1 s 12448 20005 12837 20036 4 gnd
rlabel metal1 s 8558 23084 8947 23115 4 gnd
rlabel metal1 s 14782 23084 15171 23115 4 gnd
rlabel metal1 s 16727 7684 17116 7715 4 gnd
rlabel metal1 s 778 13844 1167 13875 4 gnd
rlabel metal1 s 5446 7684 5835 7715 4 gnd
rlabel metal1 s 22173 3064 22562 3095 4 gnd
rlabel metal1 s 11281 21545 11670 21576 4 gnd
rlabel metal1 s 22562 15385 22951 15416 4 gnd
rlabel metal1 s 20617 23084 21006 23115 4 gnd
rlabel metal1 s 22173 16925 22562 16956 4 gnd
rlabel metal1 s 17505 -16 17894 15 4 gnd
rlabel metal1 s 12837 3064 13226 3095 4 gnd
rlabel metal1 s 17894 21545 18283 21576 4 gnd
rlabel metal1 s 12059 13845 12448 13876 4 gnd
rlabel metal1 s 17116 23084 17505 23115 4 gnd
rlabel metal1 s 23729 13844 24118 13875 4 gnd
rlabel metal1 s 10892 4605 11281 4636 4 gnd
rlabel metal1 s 18672 4605 19061 4636 4 gnd
rlabel metal1 s 13615 13844 14004 13875 4 gnd
rlabel metal1 s 18672 13844 19061 13875 4 gnd
rlabel metal1 s 17116 15384 17505 15415 4 gnd
rlabel metal1 s 8947 3065 9336 3096 4 gnd
rlabel metal1 s 14782 3064 15171 3095 4 gnd
rlabel metal1 s 16727 12304 17116 12335 4 gnd
rlabel metal1 s 14393 23084 14782 23115 4 gnd
rlabel metal1 s 19839 16925 20228 16956 4 gnd
rlabel metal1 s 12059 1524 12448 1555 4 gnd
rlabel metal1 s 0 21545 389 21576 4 gnd
rlabel metal1 s 19450 21545 19839 21576 4 gnd
rlabel metal1 s 11670 4604 12059 4635 4 gnd
rlabel metal1 s 24507 15384 24896 15415 4 gnd
rlabel metal1 s 19061 9225 19450 9256 4 gnd
rlabel metal1 s 23340 6145 23729 6176 4 gnd
rlabel metal1 s 21006 4604 21395 4635 4 gnd
rlabel metal1 s 10503 9225 10892 9256 4 gnd
rlabel metal1 s 6224 10765 6613 10796 4 gnd
rlabel metal1 s 16727 13845 17116 13876 4 gnd
rlabel metal1 s 21784 7685 22173 7716 4 gnd
rlabel metal1 s 23729 12304 24118 12335 4 gnd
rlabel metal1 s 14004 18465 14393 18496 4 gnd
rlabel metal1 s 19839 -16 20228 15 4 gnd
rlabel metal1 s 5835 13845 6224 13876 4 gnd
rlabel metal1 s 21784 21545 22173 21576 4 gnd
rlabel metal1 s 14004 18464 14393 18495 4 gnd
rlabel metal1 s 0 23084 389 23115 4 gnd
rlabel metal1 s 15171 3065 15560 3096 4 gnd
rlabel metal1 s 9336 6144 9725 6175 4 gnd
rlabel metal1 s 5835 1525 6224 1556 4 gnd
rlabel metal1 s 2723 3065 3112 3096 4 gnd
rlabel metal1 s 1167 16924 1556 16955 4 gnd
rlabel metal1 s 23729 9224 24118 9255 4 gnd
rlabel metal1 s 21395 3064 21784 3095 4 gnd
rlabel metal1 s 22173 4604 22562 4635 4 gnd
rlabel metal1 s 24118 16925 24507 16956 4 gnd
rlabel metal1 s 19450 18464 19839 18495 4 gnd
rlabel metal1 s 14004 23085 14393 23116 4 gnd
rlabel metal1 s 19450 6144 19839 6175 4 gnd
rlabel metal1 s 2723 6145 3112 6176 4 gnd
rlabel metal1 s 9336 6145 9725 6176 4 gnd
rlabel metal1 s 7391 10765 7780 10796 4 gnd
rlabel metal1 s 17116 1525 17505 1556 4 gnd
rlabel metal1 s 3112 10765 3501 10796 4 gnd
rlabel metal1 s 23340 23084 23729 23115 4 gnd
rlabel metal1 s 9725 20004 10114 20035 4 gnd
rlabel metal1 s 3890 3065 4279 3096 4 gnd
rlabel metal1 s 22951 24625 23340 24656 4 gnd
rlabel metal1 s 7391 3064 7780 3095 4 gnd
rlabel metal1 s 8169 18465 8558 18496 4 gnd
rlabel metal1 s 20617 7685 21006 7716 4 gnd
rlabel metal1 s 3112 3065 3501 3096 4 gnd
rlabel metal1 s 17894 1525 18283 1556 4 gnd
rlabel metal1 s 15949 15384 16338 15415 4 gnd
rlabel metal1 s 8558 4604 8947 4635 4 gnd
rlabel metal1 s 1945 21544 2334 21575 4 gnd
rlabel metal1 s 20228 18464 20617 18495 4 gnd
rlabel metal1 s 0 15385 389 15416 4 gnd
rlabel metal1 s 10114 3064 10503 3095 4 gnd
rlabel metal1 s 9336 -16 9725 15 4 gnd
rlabel metal1 s 15560 16924 15949 16955 4 gnd
rlabel metal1 s 9336 23085 9725 23116 4 gnd
rlabel metal1 s 16338 15385 16727 15416 4 gnd
rlabel metal1 s 1167 23084 1556 23115 4 gnd
rlabel metal1 s 17894 23084 18283 23115 4 gnd
rlabel metal1 s 0 6145 389 6176 4 gnd
rlabel metal1 s 22173 6144 22562 6175 4 gnd
rlabel metal1 s 17894 24625 18283 24656 4 gnd
rlabel metal1 s 8558 18465 8947 18496 4 gnd
rlabel metal1 s 1556 21545 1945 21576 4 gnd
rlabel metal1 s 12059 6145 12448 6176 4 gnd
rlabel metal1 s 1945 12304 2334 12335 4 gnd
rlabel metal1 s 18283 4604 18672 4635 4 gnd
rlabel metal1 s 5835 7684 6224 7715 4 gnd
rlabel metal1 s 7391 21544 7780 21575 4 gnd
rlabel metal1 s 8558 18464 8947 18495 4 gnd
rlabel metal1 s 17505 6144 17894 6175 4 gnd
rlabel metal1 s 2723 4604 3112 4635 4 gnd
rlabel metal1 s 14782 16924 15171 16955 4 gnd
rlabel metal1 s 389 -16 778 15 4 gnd
rlabel metal1 s 24118 18464 24507 18495 4 gnd
rlabel metal1 s 5835 6144 6224 6175 4 gnd
rlabel metal1 s 17505 21544 17894 21575 4 gnd
rlabel metal1 s 19839 3064 20228 3095 4 gnd
rlabel metal1 s 19839 1525 20228 1556 4 gnd
rlabel metal1 s 12837 9225 13226 9256 4 gnd
rlabel metal1 s 21395 16925 21784 16956 4 gnd
rlabel metal1 s 8947 13845 9336 13876 4 gnd
rlabel metal1 s 23340 24625 23729 24656 4 gnd
rlabel metal1 s 2723 10764 3112 10795 4 gnd
rlabel metal1 s 11281 6145 11670 6176 4 gnd
rlabel metal1 s 6613 3064 7002 3095 4 gnd
rlabel metal1 s 4279 23085 4668 23116 4 gnd
rlabel metal1 s 778 10765 1167 10796 4 gnd
rlabel metal1 s 21395 4605 21784 4636 4 gnd
rlabel metal1 s 7780 4605 8169 4636 4 gnd
rlabel metal1 s 1167 6145 1556 6176 4 gnd
rlabel metal1 s 15171 18465 15560 18496 4 gnd
rlabel metal1 s 12837 15385 13226 15416 4 gnd
rlabel metal1 s 6613 21544 7002 21575 4 gnd
rlabel metal1 s 13615 3065 14004 3096 4 gnd
rlabel metal1 s 14393 4605 14782 4636 4 gnd
rlabel metal1 s 17116 12305 17505 12336 4 gnd
rlabel metal1 s 11670 1525 12059 1556 4 gnd
rlabel metal1 s 389 3064 778 3095 4 gnd
rlabel metal1 s 15560 10765 15949 10796 4 gnd
rlabel metal1 s 6613 16925 7002 16956 4 gnd
rlabel metal1 s 16338 7685 16727 7716 4 gnd
rlabel metal1 s 3890 9224 4279 9255 4 gnd
rlabel metal1 s 12837 3065 13226 3096 4 gnd
rlabel metal1 s 19061 6144 19450 6175 4 gnd
rlabel metal1 s 10114 12305 10503 12336 4 gnd
rlabel metal1 s 19450 23085 19839 23116 4 gnd
rlabel metal1 s 23729 18465 24118 18496 4 gnd
<< properties >>
string FIXED_BBOX 0 0 49792 49280
string GDS_FILE sram_0rw2r1w_16_128_sky130A.gds
string GDS_END 1294704
string GDS_START 395200
<< end >>
