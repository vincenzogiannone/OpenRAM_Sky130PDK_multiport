magic
tech sky130A
magscale 1 2
timestamp 1644951705
<< checkpaint >>
rect -1296 -1277 1664 2857
<< nwell >>
rect -36 739 404 1597
<< pwell >>
rect 258 51 308 133
<< psubdiff >>
rect 258 109 308 133
rect 258 75 266 109
rect 300 75 308 109
rect 258 51 308 75
<< nsubdiff >>
rect 258 1465 308 1489
rect 258 1431 266 1465
rect 300 1431 308 1465
rect 258 1407 308 1431
<< psubdiffcont >>
rect 266 75 300 109
<< nsubdiffcont >>
rect 266 1431 300 1465
<< poly >>
rect 114 761 144 1211
rect 48 745 144 761
rect 48 711 64 745
rect 98 711 144 745
rect 48 695 144 711
rect 114 161 144 695
<< polycont >>
rect 64 711 98 745
<< locali >>
rect 0 1523 368 1557
rect 62 1330 96 1523
rect 266 1465 300 1523
rect 266 1415 300 1431
rect 48 745 114 761
rect 48 711 64 745
rect 98 711 114 745
rect 48 695 114 711
rect 162 745 196 1396
rect 162 711 213 745
rect 162 60 196 711
rect 266 109 300 125
rect 62 17 96 60
rect 266 17 300 75
rect 0 -17 368 17
use contact_12  contact_12_0
timestamp 1644951705
transform 1 0 48 0 1 695
box 0 0 1 1
use contact_11  contact_11_0
timestamp 1644951705
transform 1 0 258 0 1 51
box 0 0 1 1
use contact_10  contact_10_0
timestamp 1644951705
transform 1 0 258 0 1 1407
box 0 0 1 1
use nmos_m1_w0_420_sli_dli_da_p  nmos_m1_w0_420_sli_dli_da_p_0
timestamp 1644951705
transform 1 0 54 0 1 51
box 0 -26 150 110
use pmos_m1_w1_260_sli_dli_da_p  pmos_m1_w1_260_sli_dli_da_p_0
timestamp 1644951705
transform 1 0 54 0 1 1237
box -59 -54 209 306
<< labels >>
rlabel locali s 81 728 81 728 4 A
rlabel locali s 196 728 196 728 4 Z
rlabel locali s 184 0 184 0 4 gnd
rlabel locali s 184 1540 184 1540 4 vdd
<< properties >>
string FIXED_BBOX 0 0 368 1540
string GDS_FILE sram_0rw2r1w_16_128_sky130A.gds
string GDS_END 1784158
string GDS_START 1782666
<< end >>
