magic
tech sky130A
magscale 1 2
timestamp 1644951705
<< checkpaint >>
rect -1260 -1302 4272 2176
<< locali >>
rect 2169 564 2170 581
rect 2169 394 2203 564
rect 2008 360 2365 394
rect 2592 360 2711 394
rect 2677 190 2711 360
<< viali >>
rect 2170 564 2204 598
rect 1872 360 1906 394
rect 2677 156 2711 190
<< metal1 >>
rect 0 808 2976 868
rect 2154 555 2160 607
rect 2212 555 2219 607
rect 1857 351 1863 403
rect 1915 351 1921 403
rect 2662 147 2668 199
rect 2720 147 2726 199
rect 0 -30 2976 30
<< via1 >>
rect 2160 598 2212 607
rect 2160 564 2170 598
rect 2170 564 2204 598
rect 2204 564 2212 598
rect 2160 555 2212 564
rect 1863 394 1915 403
rect 1863 360 1872 394
rect 1872 360 1906 394
rect 1906 360 1915 394
rect 1863 351 1915 360
rect 2668 190 2720 199
rect 2668 156 2677 190
rect 2677 156 2711 190
rect 2711 156 2720 190
rect 2668 147 2720 156
<< metal2 >>
rect 2160 607 2212 613
rect 2160 549 2212 555
rect 1863 403 1915 409
rect 0 322 54 350
rect 1863 345 1915 351
rect 180 232 234 260
rect 1875 256 1903 345
rect 1287 228 1903 256
rect 2668 199 2720 205
rect 2668 141 2720 147
use contact_17  contact_17_0
timestamp 1644951705
transform 1 0 2154 0 1 549
box 0 0 1 1
use contact_13  contact_13_0
timestamp 1644951705
transform 1 0 2158 0 1 558
box 0 0 1 1
use contact_17  contact_17_1
timestamp 1644951705
transform 1 0 2662 0 1 141
box 0 0 1 1
use contact_13  contact_13_1
timestamp 1644951705
transform 1 0 2665 0 1 150
box 0 0 1 1
use contact_17  contact_17_2
timestamp 1644951705
transform 1 0 1857 0 1 345
box 0 0 1 1
use contact_13  contact_13_2
timestamp 1644951705
transform 1 0 1860 0 1 354
box 0 0 1 1
use pinv_3  pinv_3_0
timestamp 1644951705
transform 1 0 2284 0 1 0
box -36 -17 728 895
use pinv_2  pinv_2_0
timestamp 1644951705
transform 1 0 1808 0 1 0
box -36 -17 512 895
use dff  dff_0
timestamp 1644951705
transform 1 0 0 0 1 0
box 0 -42 1482 916
<< labels >>
rlabel metal1 s 0 808 2976 868 4 vdd
rlabel metal1 s 0 -30 2976 30 4 gnd
rlabel metal2 s 0 322 54 350 4 clk
rlabel metal2 s 180 232 234 260 4 D
rlabel metal2 s 2680 159 2708 187 4 Q
rlabel metal2 s 2172 567 2200 595 4 Qb
<< properties >>
string FIXED_BBOX 0 0 2976 838
string GDS_FILE sram_0rw2r1w_16_128_sky130A.gds
string GDS_END 1950486
string GDS_START 1948130
<< end >>
