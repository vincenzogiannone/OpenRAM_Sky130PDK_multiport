magic
tech sky130A
magscale 1 2
timestamp 1644969367
<< checkpaint >>
rect -1299 -1302 48684 2176
<< metal1 >>
rect 709 812 715 864
rect 767 812 773 864
rect 2191 812 2197 864
rect 2249 812 2255 864
rect 3673 812 3679 864
rect 3731 812 3737 864
rect 5155 812 5161 864
rect 5213 812 5219 864
rect 6637 812 6643 864
rect 6695 812 6701 864
rect 8119 812 8125 864
rect 8177 812 8183 864
rect 9601 812 9607 864
rect 9659 812 9665 864
rect 11083 812 11089 864
rect 11141 812 11147 864
rect 12565 812 12571 864
rect 12623 812 12629 864
rect 14047 812 14053 864
rect 14105 812 14111 864
rect 15529 812 15535 864
rect 15587 812 15593 864
rect 17011 812 17017 864
rect 17069 812 17075 864
rect 18493 812 18499 864
rect 18551 812 18557 864
rect 19975 812 19981 864
rect 20033 812 20039 864
rect 21457 812 21463 864
rect 21515 812 21521 864
rect 22939 812 22945 864
rect 22997 812 23003 864
rect 24421 812 24427 864
rect 24479 812 24485 864
rect 25903 812 25909 864
rect 25961 812 25967 864
rect 27385 812 27391 864
rect 27443 812 27449 864
rect 28867 812 28873 864
rect 28925 812 28931 864
rect 30349 812 30355 864
rect 30407 812 30413 864
rect 31831 812 31837 864
rect 31889 812 31895 864
rect 33313 812 33319 864
rect 33371 812 33377 864
rect 34795 812 34801 864
rect 34853 812 34859 864
rect 36277 812 36283 864
rect 36335 812 36341 864
rect 37759 812 37765 864
rect 37817 812 37823 864
rect 39241 812 39247 864
rect 39299 812 39305 864
rect 40723 812 40729 864
rect 40781 812 40787 864
rect 42205 812 42211 864
rect 42263 812 42269 864
rect 43687 812 43693 864
rect 43745 812 43751 864
rect 45169 812 45175 864
rect 45227 812 45233 864
rect 46651 812 46657 864
rect 46709 812 46715 864
rect 709 -26 715 26
rect 767 -26 773 26
rect 2191 -26 2197 26
rect 2249 -26 2255 26
rect 3673 -26 3679 26
rect 3731 -26 3737 26
rect 5155 -26 5161 26
rect 5213 -26 5219 26
rect 6637 -26 6643 26
rect 6695 -26 6701 26
rect 8119 -26 8125 26
rect 8177 -26 8183 26
rect 9601 -26 9607 26
rect 9659 -26 9665 26
rect 11083 -26 11089 26
rect 11141 -26 11147 26
rect 12565 -26 12571 26
rect 12623 -26 12629 26
rect 14047 -26 14053 26
rect 14105 -26 14111 26
rect 15529 -26 15535 26
rect 15587 -26 15593 26
rect 17011 -26 17017 26
rect 17069 -26 17075 26
rect 18493 -26 18499 26
rect 18551 -26 18557 26
rect 19975 -26 19981 26
rect 20033 -26 20039 26
rect 21457 -26 21463 26
rect 21515 -26 21521 26
rect 22939 -26 22945 26
rect 22997 -26 23003 26
rect 24421 -26 24427 26
rect 24479 -26 24485 26
rect 25903 -26 25909 26
rect 25961 -26 25967 26
rect 27385 -26 27391 26
rect 27443 -26 27449 26
rect 28867 -26 28873 26
rect 28925 -26 28931 26
rect 30349 -26 30355 26
rect 30407 -26 30413 26
rect 31831 -26 31837 26
rect 31889 -26 31895 26
rect 33313 -26 33319 26
rect 33371 -26 33377 26
rect 34795 -26 34801 26
rect 34853 -26 34859 26
rect 36277 -26 36283 26
rect 36335 -26 36341 26
rect 37759 -26 37765 26
rect 37817 -26 37823 26
rect 39241 -26 39247 26
rect 39299 -26 39305 26
rect 40723 -26 40729 26
rect 40781 -26 40787 26
rect 42205 -26 42211 26
rect 42263 -26 42269 26
rect 43687 -26 43693 26
rect 43745 -26 43751 26
rect 45169 -26 45175 26
rect 45227 -26 45233 26
rect 46651 -26 46657 26
rect 46709 -26 46715 26
<< via1 >>
rect 715 812 767 864
rect 2197 812 2249 864
rect 3679 812 3731 864
rect 5161 812 5213 864
rect 6643 812 6695 864
rect 8125 812 8177 864
rect 9607 812 9659 864
rect 11089 812 11141 864
rect 12571 812 12623 864
rect 14053 812 14105 864
rect 15535 812 15587 864
rect 17017 812 17069 864
rect 18499 812 18551 864
rect 19981 812 20033 864
rect 21463 812 21515 864
rect 22945 812 22997 864
rect 24427 812 24479 864
rect 25909 812 25961 864
rect 27391 812 27443 864
rect 28873 812 28925 864
rect 30355 812 30407 864
rect 31837 812 31889 864
rect 33319 812 33371 864
rect 34801 812 34853 864
rect 36283 812 36335 864
rect 37765 812 37817 864
rect 39247 812 39299 864
rect 40729 812 40781 864
rect 42211 812 42263 864
rect 43693 812 43745 864
rect 45175 812 45227 864
rect 46657 812 46709 864
rect 715 -26 767 26
rect 2197 -26 2249 26
rect 3679 -26 3731 26
rect 5161 -26 5213 26
rect 6643 -26 6695 26
rect 8125 -26 8177 26
rect 9607 -26 9659 26
rect 11089 -26 11141 26
rect 12571 -26 12623 26
rect 14053 -26 14105 26
rect 15535 -26 15587 26
rect 17017 -26 17069 26
rect 18499 -26 18551 26
rect 19981 -26 20033 26
rect 21463 -26 21515 26
rect 22945 -26 22997 26
rect 24427 -26 24479 26
rect 25909 -26 25961 26
rect 27391 -26 27443 26
rect 28873 -26 28925 26
rect 30355 -26 30407 26
rect 31837 -26 31889 26
rect 33319 -26 33371 26
rect 34801 -26 34853 26
rect 36283 -26 36335 26
rect 37765 -26 37817 26
rect 39247 -26 39299 26
rect 40729 -26 40781 26
rect 42211 -26 42263 26
rect 43693 -26 43745 26
rect 45175 -26 45227 26
rect 46657 -26 46709 26
<< metal2 >>
rect 713 866 769 875
rect 0 345 28 838
rect 2195 866 2251 875
rect 713 801 769 810
rect 1482 345 1510 838
rect 3677 866 3733 875
rect 2195 801 2251 810
rect 2964 345 2992 838
rect 5159 866 5215 875
rect 3677 801 3733 810
rect 4446 345 4474 838
rect 6641 866 6697 875
rect 5159 801 5215 810
rect 5928 345 5956 838
rect 8123 866 8179 875
rect 6641 801 6697 810
rect 7410 345 7438 838
rect 9605 866 9661 875
rect 8123 801 8179 810
rect 8892 345 8920 838
rect 11087 866 11143 875
rect 9605 801 9661 810
rect 10374 345 10402 838
rect 12569 866 12625 875
rect 11087 801 11143 810
rect 11856 345 11884 838
rect 14051 866 14107 875
rect 12569 801 12625 810
rect 13338 345 13366 838
rect 15533 866 15589 875
rect 14051 801 14107 810
rect 14820 345 14848 838
rect 17015 866 17071 875
rect 15533 801 15589 810
rect 16302 345 16330 838
rect 18497 866 18553 875
rect 17015 801 17071 810
rect 17784 345 17812 838
rect 19979 866 20035 875
rect 18497 801 18553 810
rect 19266 345 19294 838
rect 21461 866 21517 875
rect 19979 801 20035 810
rect 20748 345 20776 838
rect 22943 866 22999 875
rect 21461 801 21517 810
rect 22230 345 22258 838
rect 24425 866 24481 875
rect 22943 801 22999 810
rect 23712 345 23740 838
rect 25907 866 25963 875
rect 24425 801 24481 810
rect 25194 345 25222 838
rect 27389 866 27445 875
rect 25907 801 25963 810
rect 26676 345 26704 838
rect 28871 866 28927 875
rect 27389 801 27445 810
rect 28158 345 28186 838
rect 30353 866 30409 875
rect 28871 801 28927 810
rect 29640 345 29668 838
rect 31835 866 31891 875
rect 30353 801 30409 810
rect 31122 345 31150 838
rect 33317 866 33373 875
rect 31835 801 31891 810
rect 32604 345 32632 838
rect 34799 866 34855 875
rect 33317 801 33373 810
rect 34086 345 34114 838
rect 36281 866 36337 875
rect 34799 801 34855 810
rect 35568 345 35596 838
rect 37763 866 37819 875
rect 36281 801 36337 810
rect 37050 345 37078 838
rect 39245 866 39301 875
rect 37763 801 37819 810
rect 38532 345 38560 838
rect 40727 866 40783 875
rect 39245 801 39301 810
rect 40014 345 40042 838
rect 42209 866 42265 875
rect 40727 801 40783 810
rect 41496 345 41524 838
rect 43691 866 43747 875
rect 42209 801 42265 810
rect 42978 345 43006 838
rect 45173 866 45229 875
rect 43691 801 43747 810
rect 44460 345 44488 838
rect 46655 866 46711 875
rect 45173 801 45229 810
rect 45942 345 45970 838
rect 46655 801 46711 810
rect -1 336 55 345
rect -1 271 55 280
rect 1481 336 1537 345
rect 1481 271 1537 280
rect 2963 336 3019 345
rect 2963 271 3019 280
rect 4445 336 4501 345
rect 4445 271 4501 280
rect 5927 336 5983 345
rect 5927 271 5983 280
rect 7409 336 7465 345
rect 7409 271 7465 280
rect 8891 336 8947 345
rect 8891 271 8947 280
rect 10373 336 10429 345
rect 10373 271 10429 280
rect 11855 336 11911 345
rect 11855 271 11911 280
rect 13337 336 13393 345
rect 13337 271 13393 280
rect 14819 336 14875 345
rect 14819 271 14875 280
rect 16301 336 16357 345
rect 16301 271 16357 280
rect 17783 336 17839 345
rect 17783 271 17839 280
rect 19265 336 19321 345
rect 19265 271 19321 280
rect 20747 336 20803 345
rect 20747 271 20803 280
rect 22229 336 22285 345
rect 22229 271 22285 280
rect 23711 336 23767 345
rect 23711 271 23767 280
rect 25193 336 25249 345
rect 25193 271 25249 280
rect 26675 336 26731 345
rect 26675 271 26731 280
rect 28157 336 28213 345
rect 28157 271 28213 280
rect 29639 336 29695 345
rect 29639 271 29695 280
rect 31121 336 31177 345
rect 31121 271 31177 280
rect 32603 336 32659 345
rect 32603 271 32659 280
rect 34085 336 34141 345
rect 34085 271 34141 280
rect 35567 336 35623 345
rect 35567 271 35623 280
rect 37049 336 37105 345
rect 37049 271 37105 280
rect 38531 336 38587 345
rect 38531 271 38587 280
rect 40013 336 40069 345
rect 40013 271 40069 280
rect 41495 336 41551 345
rect 41495 271 41551 280
rect 42977 336 43033 345
rect 42977 271 43033 280
rect 44459 336 44515 345
rect 44459 271 44515 280
rect 45941 336 45997 345
rect 45941 271 45997 280
rect 0 0 28 271
rect 180 232 234 260
rect 1260 228 1314 256
rect 713 28 769 37
rect 1482 0 1510 271
rect 1662 232 1716 260
rect 2742 228 2796 256
rect 2195 28 2251 37
rect 713 -37 769 -28
rect 2964 0 2992 271
rect 3144 232 3198 260
rect 4224 228 4278 256
rect 3677 28 3733 37
rect 2195 -37 2251 -28
rect 4446 0 4474 271
rect 4626 232 4680 260
rect 5706 228 5760 256
rect 5159 28 5215 37
rect 3677 -37 3733 -28
rect 5928 0 5956 271
rect 6108 232 6162 260
rect 7188 228 7242 256
rect 6641 28 6697 37
rect 5159 -37 5215 -28
rect 7410 0 7438 271
rect 7590 232 7644 260
rect 8670 228 8724 256
rect 8123 28 8179 37
rect 6641 -37 6697 -28
rect 8892 0 8920 271
rect 9072 232 9126 260
rect 10152 228 10206 256
rect 9605 28 9661 37
rect 8123 -37 8179 -28
rect 10374 0 10402 271
rect 10554 232 10608 260
rect 11634 228 11688 256
rect 11087 28 11143 37
rect 9605 -37 9661 -28
rect 11856 0 11884 271
rect 12036 232 12090 260
rect 13116 228 13170 256
rect 12569 28 12625 37
rect 11087 -37 11143 -28
rect 13338 0 13366 271
rect 13518 232 13572 260
rect 14598 228 14652 256
rect 14051 28 14107 37
rect 12569 -37 12625 -28
rect 14820 0 14848 271
rect 15000 232 15054 260
rect 16080 228 16134 256
rect 15533 28 15589 37
rect 14051 -37 14107 -28
rect 16302 0 16330 271
rect 16482 232 16536 260
rect 17562 228 17616 256
rect 17015 28 17071 37
rect 15533 -37 15589 -28
rect 17784 0 17812 271
rect 17964 232 18018 260
rect 19044 228 19098 256
rect 18497 28 18553 37
rect 17015 -37 17071 -28
rect 19266 0 19294 271
rect 19446 232 19500 260
rect 20526 228 20580 256
rect 19979 28 20035 37
rect 18497 -37 18553 -28
rect 20748 0 20776 271
rect 20928 232 20982 260
rect 22008 228 22062 256
rect 21461 28 21517 37
rect 19979 -37 20035 -28
rect 22230 0 22258 271
rect 22410 232 22464 260
rect 23490 228 23544 256
rect 22943 28 22999 37
rect 21461 -37 21517 -28
rect 23712 0 23740 271
rect 23892 232 23946 260
rect 24972 228 25026 256
rect 24425 28 24481 37
rect 22943 -37 22999 -28
rect 25194 0 25222 271
rect 25374 232 25428 260
rect 26454 228 26508 256
rect 25907 28 25963 37
rect 24425 -37 24481 -28
rect 26676 0 26704 271
rect 26856 232 26910 260
rect 27936 228 27990 256
rect 27389 28 27445 37
rect 25907 -37 25963 -28
rect 28158 0 28186 271
rect 28338 232 28392 260
rect 29418 228 29472 256
rect 28871 28 28927 37
rect 27389 -37 27445 -28
rect 29640 0 29668 271
rect 29820 232 29874 260
rect 30900 228 30954 256
rect 30353 28 30409 37
rect 28871 -37 28927 -28
rect 31122 0 31150 271
rect 31302 232 31356 260
rect 32382 228 32436 256
rect 31835 28 31891 37
rect 30353 -37 30409 -28
rect 32604 0 32632 271
rect 32784 232 32838 260
rect 33864 228 33918 256
rect 33317 28 33373 37
rect 31835 -37 31891 -28
rect 34086 0 34114 271
rect 34266 232 34320 260
rect 35346 228 35400 256
rect 34799 28 34855 37
rect 33317 -37 33373 -28
rect 35568 0 35596 271
rect 35748 232 35802 260
rect 36828 228 36882 256
rect 36281 28 36337 37
rect 34799 -37 34855 -28
rect 37050 0 37078 271
rect 37230 232 37284 260
rect 38310 228 38364 256
rect 37763 28 37819 37
rect 36281 -37 36337 -28
rect 38532 0 38560 271
rect 38712 232 38766 260
rect 39792 228 39846 256
rect 39245 28 39301 37
rect 37763 -37 37819 -28
rect 40014 0 40042 271
rect 40194 232 40248 260
rect 41274 228 41328 256
rect 40727 28 40783 37
rect 39245 -37 39301 -28
rect 41496 0 41524 271
rect 41676 232 41730 260
rect 42756 228 42810 256
rect 42209 28 42265 37
rect 40727 -37 40783 -28
rect 42978 0 43006 271
rect 43158 232 43212 260
rect 44238 228 44292 256
rect 43691 28 43747 37
rect 42209 -37 42265 -28
rect 44460 0 44488 271
rect 44640 232 44694 260
rect 45720 228 45774 256
rect 45173 28 45229 37
rect 43691 -37 43747 -28
rect 45942 0 45970 271
rect 46122 232 46176 260
rect 47202 228 47256 256
rect 46655 28 46711 37
rect 45173 -37 45229 -28
rect 46655 -37 46711 -28
<< via2 >>
rect 713 864 769 866
rect 713 812 715 864
rect 715 812 767 864
rect 767 812 769 864
rect 2195 864 2251 866
rect 713 810 769 812
rect 2195 812 2197 864
rect 2197 812 2249 864
rect 2249 812 2251 864
rect 3677 864 3733 866
rect 2195 810 2251 812
rect 3677 812 3679 864
rect 3679 812 3731 864
rect 3731 812 3733 864
rect 5159 864 5215 866
rect 3677 810 3733 812
rect 5159 812 5161 864
rect 5161 812 5213 864
rect 5213 812 5215 864
rect 6641 864 6697 866
rect 5159 810 5215 812
rect 6641 812 6643 864
rect 6643 812 6695 864
rect 6695 812 6697 864
rect 8123 864 8179 866
rect 6641 810 6697 812
rect 8123 812 8125 864
rect 8125 812 8177 864
rect 8177 812 8179 864
rect 9605 864 9661 866
rect 8123 810 8179 812
rect 9605 812 9607 864
rect 9607 812 9659 864
rect 9659 812 9661 864
rect 11087 864 11143 866
rect 9605 810 9661 812
rect 11087 812 11089 864
rect 11089 812 11141 864
rect 11141 812 11143 864
rect 12569 864 12625 866
rect 11087 810 11143 812
rect 12569 812 12571 864
rect 12571 812 12623 864
rect 12623 812 12625 864
rect 14051 864 14107 866
rect 12569 810 12625 812
rect 14051 812 14053 864
rect 14053 812 14105 864
rect 14105 812 14107 864
rect 15533 864 15589 866
rect 14051 810 14107 812
rect 15533 812 15535 864
rect 15535 812 15587 864
rect 15587 812 15589 864
rect 17015 864 17071 866
rect 15533 810 15589 812
rect 17015 812 17017 864
rect 17017 812 17069 864
rect 17069 812 17071 864
rect 18497 864 18553 866
rect 17015 810 17071 812
rect 18497 812 18499 864
rect 18499 812 18551 864
rect 18551 812 18553 864
rect 19979 864 20035 866
rect 18497 810 18553 812
rect 19979 812 19981 864
rect 19981 812 20033 864
rect 20033 812 20035 864
rect 21461 864 21517 866
rect 19979 810 20035 812
rect 21461 812 21463 864
rect 21463 812 21515 864
rect 21515 812 21517 864
rect 22943 864 22999 866
rect 21461 810 21517 812
rect 22943 812 22945 864
rect 22945 812 22997 864
rect 22997 812 22999 864
rect 24425 864 24481 866
rect 22943 810 22999 812
rect 24425 812 24427 864
rect 24427 812 24479 864
rect 24479 812 24481 864
rect 25907 864 25963 866
rect 24425 810 24481 812
rect 25907 812 25909 864
rect 25909 812 25961 864
rect 25961 812 25963 864
rect 27389 864 27445 866
rect 25907 810 25963 812
rect 27389 812 27391 864
rect 27391 812 27443 864
rect 27443 812 27445 864
rect 28871 864 28927 866
rect 27389 810 27445 812
rect 28871 812 28873 864
rect 28873 812 28925 864
rect 28925 812 28927 864
rect 30353 864 30409 866
rect 28871 810 28927 812
rect 30353 812 30355 864
rect 30355 812 30407 864
rect 30407 812 30409 864
rect 31835 864 31891 866
rect 30353 810 30409 812
rect 31835 812 31837 864
rect 31837 812 31889 864
rect 31889 812 31891 864
rect 33317 864 33373 866
rect 31835 810 31891 812
rect 33317 812 33319 864
rect 33319 812 33371 864
rect 33371 812 33373 864
rect 34799 864 34855 866
rect 33317 810 33373 812
rect 34799 812 34801 864
rect 34801 812 34853 864
rect 34853 812 34855 864
rect 36281 864 36337 866
rect 34799 810 34855 812
rect 36281 812 36283 864
rect 36283 812 36335 864
rect 36335 812 36337 864
rect 37763 864 37819 866
rect 36281 810 36337 812
rect 37763 812 37765 864
rect 37765 812 37817 864
rect 37817 812 37819 864
rect 39245 864 39301 866
rect 37763 810 37819 812
rect 39245 812 39247 864
rect 39247 812 39299 864
rect 39299 812 39301 864
rect 40727 864 40783 866
rect 39245 810 39301 812
rect 40727 812 40729 864
rect 40729 812 40781 864
rect 40781 812 40783 864
rect 42209 864 42265 866
rect 40727 810 40783 812
rect 42209 812 42211 864
rect 42211 812 42263 864
rect 42263 812 42265 864
rect 43691 864 43747 866
rect 42209 810 42265 812
rect 43691 812 43693 864
rect 43693 812 43745 864
rect 43745 812 43747 864
rect 45173 864 45229 866
rect 43691 810 43747 812
rect 45173 812 45175 864
rect 45175 812 45227 864
rect 45227 812 45229 864
rect 46655 864 46711 866
rect 45173 810 45229 812
rect 46655 812 46657 864
rect 46657 812 46709 864
rect 46709 812 46711 864
rect 46655 810 46711 812
rect -1 280 55 336
rect 1481 280 1537 336
rect 2963 280 3019 336
rect 4445 280 4501 336
rect 5927 280 5983 336
rect 7409 280 7465 336
rect 8891 280 8947 336
rect 10373 280 10429 336
rect 11855 280 11911 336
rect 13337 280 13393 336
rect 14819 280 14875 336
rect 16301 280 16357 336
rect 17783 280 17839 336
rect 19265 280 19321 336
rect 20747 280 20803 336
rect 22229 280 22285 336
rect 23711 280 23767 336
rect 25193 280 25249 336
rect 26675 280 26731 336
rect 28157 280 28213 336
rect 29639 280 29695 336
rect 31121 280 31177 336
rect 32603 280 32659 336
rect 34085 280 34141 336
rect 35567 280 35623 336
rect 37049 280 37105 336
rect 38531 280 38587 336
rect 40013 280 40069 336
rect 41495 280 41551 336
rect 42977 280 43033 336
rect 44459 280 44515 336
rect 45941 280 45997 336
rect 713 26 769 28
rect 713 -26 715 26
rect 715 -26 767 26
rect 767 -26 769 26
rect 2195 26 2251 28
rect 713 -28 769 -26
rect 2195 -26 2197 26
rect 2197 -26 2249 26
rect 2249 -26 2251 26
rect 3677 26 3733 28
rect 2195 -28 2251 -26
rect 3677 -26 3679 26
rect 3679 -26 3731 26
rect 3731 -26 3733 26
rect 5159 26 5215 28
rect 3677 -28 3733 -26
rect 5159 -26 5161 26
rect 5161 -26 5213 26
rect 5213 -26 5215 26
rect 6641 26 6697 28
rect 5159 -28 5215 -26
rect 6641 -26 6643 26
rect 6643 -26 6695 26
rect 6695 -26 6697 26
rect 8123 26 8179 28
rect 6641 -28 6697 -26
rect 8123 -26 8125 26
rect 8125 -26 8177 26
rect 8177 -26 8179 26
rect 9605 26 9661 28
rect 8123 -28 8179 -26
rect 9605 -26 9607 26
rect 9607 -26 9659 26
rect 9659 -26 9661 26
rect 11087 26 11143 28
rect 9605 -28 9661 -26
rect 11087 -26 11089 26
rect 11089 -26 11141 26
rect 11141 -26 11143 26
rect 12569 26 12625 28
rect 11087 -28 11143 -26
rect 12569 -26 12571 26
rect 12571 -26 12623 26
rect 12623 -26 12625 26
rect 14051 26 14107 28
rect 12569 -28 12625 -26
rect 14051 -26 14053 26
rect 14053 -26 14105 26
rect 14105 -26 14107 26
rect 15533 26 15589 28
rect 14051 -28 14107 -26
rect 15533 -26 15535 26
rect 15535 -26 15587 26
rect 15587 -26 15589 26
rect 17015 26 17071 28
rect 15533 -28 15589 -26
rect 17015 -26 17017 26
rect 17017 -26 17069 26
rect 17069 -26 17071 26
rect 18497 26 18553 28
rect 17015 -28 17071 -26
rect 18497 -26 18499 26
rect 18499 -26 18551 26
rect 18551 -26 18553 26
rect 19979 26 20035 28
rect 18497 -28 18553 -26
rect 19979 -26 19981 26
rect 19981 -26 20033 26
rect 20033 -26 20035 26
rect 21461 26 21517 28
rect 19979 -28 20035 -26
rect 21461 -26 21463 26
rect 21463 -26 21515 26
rect 21515 -26 21517 26
rect 22943 26 22999 28
rect 21461 -28 21517 -26
rect 22943 -26 22945 26
rect 22945 -26 22997 26
rect 22997 -26 22999 26
rect 24425 26 24481 28
rect 22943 -28 22999 -26
rect 24425 -26 24427 26
rect 24427 -26 24479 26
rect 24479 -26 24481 26
rect 25907 26 25963 28
rect 24425 -28 24481 -26
rect 25907 -26 25909 26
rect 25909 -26 25961 26
rect 25961 -26 25963 26
rect 27389 26 27445 28
rect 25907 -28 25963 -26
rect 27389 -26 27391 26
rect 27391 -26 27443 26
rect 27443 -26 27445 26
rect 28871 26 28927 28
rect 27389 -28 27445 -26
rect 28871 -26 28873 26
rect 28873 -26 28925 26
rect 28925 -26 28927 26
rect 30353 26 30409 28
rect 28871 -28 28927 -26
rect 30353 -26 30355 26
rect 30355 -26 30407 26
rect 30407 -26 30409 26
rect 31835 26 31891 28
rect 30353 -28 30409 -26
rect 31835 -26 31837 26
rect 31837 -26 31889 26
rect 31889 -26 31891 26
rect 33317 26 33373 28
rect 31835 -28 31891 -26
rect 33317 -26 33319 26
rect 33319 -26 33371 26
rect 33371 -26 33373 26
rect 34799 26 34855 28
rect 33317 -28 33373 -26
rect 34799 -26 34801 26
rect 34801 -26 34853 26
rect 34853 -26 34855 26
rect 36281 26 36337 28
rect 34799 -28 34855 -26
rect 36281 -26 36283 26
rect 36283 -26 36335 26
rect 36335 -26 36337 26
rect 37763 26 37819 28
rect 36281 -28 36337 -26
rect 37763 -26 37765 26
rect 37765 -26 37817 26
rect 37817 -26 37819 26
rect 39245 26 39301 28
rect 37763 -28 37819 -26
rect 39245 -26 39247 26
rect 39247 -26 39299 26
rect 39299 -26 39301 26
rect 40727 26 40783 28
rect 39245 -28 39301 -26
rect 40727 -26 40729 26
rect 40729 -26 40781 26
rect 40781 -26 40783 26
rect 42209 26 42265 28
rect 40727 -28 40783 -26
rect 42209 -26 42211 26
rect 42211 -26 42263 26
rect 42263 -26 42265 26
rect 43691 26 43747 28
rect 42209 -28 42265 -26
rect 43691 -26 43693 26
rect 43693 -26 43745 26
rect 43745 -26 43747 26
rect 45173 26 45229 28
rect 43691 -28 43747 -26
rect 45173 -26 45175 26
rect 45175 -26 45227 26
rect 45227 -26 45229 26
rect 46655 26 46711 28
rect 45173 -28 45229 -26
rect 46655 -26 46657 26
rect 46657 -26 46709 26
rect 46709 -26 46711 26
rect 46655 -28 46711 -26
<< metal3 >>
rect 675 866 807 875
rect 675 810 713 866
rect 769 810 807 866
rect 675 801 807 810
rect 2157 866 2289 875
rect 2157 810 2195 866
rect 2251 810 2289 866
rect 2157 801 2289 810
rect 3639 866 3771 875
rect 3639 810 3677 866
rect 3733 810 3771 866
rect 3639 801 3771 810
rect 5121 866 5253 875
rect 5121 810 5159 866
rect 5215 810 5253 866
rect 5121 801 5253 810
rect 6603 866 6735 875
rect 6603 810 6641 866
rect 6697 810 6735 866
rect 6603 801 6735 810
rect 8085 866 8217 875
rect 8085 810 8123 866
rect 8179 810 8217 866
rect 8085 801 8217 810
rect 9567 866 9699 875
rect 9567 810 9605 866
rect 9661 810 9699 866
rect 9567 801 9699 810
rect 11049 866 11181 875
rect 11049 810 11087 866
rect 11143 810 11181 866
rect 11049 801 11181 810
rect 12531 866 12663 875
rect 12531 810 12569 866
rect 12625 810 12663 866
rect 12531 801 12663 810
rect 14013 866 14145 875
rect 14013 810 14051 866
rect 14107 810 14145 866
rect 14013 801 14145 810
rect 15495 866 15627 875
rect 15495 810 15533 866
rect 15589 810 15627 866
rect 15495 801 15627 810
rect 16977 866 17109 875
rect 16977 810 17015 866
rect 17071 810 17109 866
rect 16977 801 17109 810
rect 18459 866 18591 875
rect 18459 810 18497 866
rect 18553 810 18591 866
rect 18459 801 18591 810
rect 19941 866 20073 875
rect 19941 810 19979 866
rect 20035 810 20073 866
rect 19941 801 20073 810
rect 21423 866 21555 875
rect 21423 810 21461 866
rect 21517 810 21555 866
rect 21423 801 21555 810
rect 22905 866 23037 875
rect 22905 810 22943 866
rect 22999 810 23037 866
rect 22905 801 23037 810
rect 24387 866 24519 875
rect 24387 810 24425 866
rect 24481 810 24519 866
rect 24387 801 24519 810
rect 25869 866 26001 875
rect 25869 810 25907 866
rect 25963 810 26001 866
rect 25869 801 26001 810
rect 27351 866 27483 875
rect 27351 810 27389 866
rect 27445 810 27483 866
rect 27351 801 27483 810
rect 28833 866 28965 875
rect 28833 810 28871 866
rect 28927 810 28965 866
rect 28833 801 28965 810
rect 30315 866 30447 875
rect 30315 810 30353 866
rect 30409 810 30447 866
rect 30315 801 30447 810
rect 31797 866 31929 875
rect 31797 810 31835 866
rect 31891 810 31929 866
rect 31797 801 31929 810
rect 33279 866 33411 875
rect 33279 810 33317 866
rect 33373 810 33411 866
rect 33279 801 33411 810
rect 34761 866 34893 875
rect 34761 810 34799 866
rect 34855 810 34893 866
rect 34761 801 34893 810
rect 36243 866 36375 875
rect 36243 810 36281 866
rect 36337 810 36375 866
rect 36243 801 36375 810
rect 37725 866 37857 875
rect 37725 810 37763 866
rect 37819 810 37857 866
rect 37725 801 37857 810
rect 39207 866 39339 875
rect 39207 810 39245 866
rect 39301 810 39339 866
rect 39207 801 39339 810
rect 40689 866 40821 875
rect 40689 810 40727 866
rect 40783 810 40821 866
rect 40689 801 40821 810
rect 42171 866 42303 875
rect 42171 810 42209 866
rect 42265 810 42303 866
rect 42171 801 42303 810
rect 43653 866 43785 875
rect 43653 810 43691 866
rect 43747 810 43785 866
rect 43653 801 43785 810
rect 45135 866 45267 875
rect 45135 810 45173 866
rect 45229 810 45267 866
rect 45135 801 45267 810
rect 46617 866 46749 875
rect 46617 810 46655 866
rect 46711 810 46749 866
rect 46617 801 46749 810
rect -39 338 93 341
rect 1443 338 1575 341
rect 2925 338 3057 341
rect 4407 338 4539 341
rect 5889 338 6021 341
rect 7371 338 7503 341
rect 8853 338 8985 341
rect 10335 338 10467 341
rect 11817 338 11949 341
rect 13299 338 13431 341
rect 14781 338 14913 341
rect 16263 338 16395 341
rect 17745 338 17877 341
rect 19227 338 19359 341
rect 20709 338 20841 341
rect 22191 338 22323 341
rect 23673 338 23805 341
rect 25155 338 25287 341
rect 26637 338 26769 341
rect 28119 338 28251 341
rect 29601 338 29733 341
rect 31083 338 31215 341
rect 32565 338 32697 341
rect 34047 338 34179 341
rect 35529 338 35661 341
rect 37011 338 37143 341
rect 38493 338 38625 341
rect 39975 338 40107 341
rect 41457 338 41589 341
rect 42939 338 43071 341
rect 44421 338 44553 341
rect 45903 338 46035 341
rect -39 336 47424 338
rect -39 280 -1 336
rect 55 280 1481 336
rect 1537 280 2963 336
rect 3019 280 4445 336
rect 4501 280 5927 336
rect 5983 280 7409 336
rect 7465 280 8891 336
rect 8947 280 10373 336
rect 10429 280 11855 336
rect 11911 280 13337 336
rect 13393 280 14819 336
rect 14875 280 16301 336
rect 16357 280 17783 336
rect 17839 280 19265 336
rect 19321 280 20747 336
rect 20803 280 22229 336
rect 22285 280 23711 336
rect 23767 280 25193 336
rect 25249 280 26675 336
rect 26731 280 28157 336
rect 28213 280 29639 336
rect 29695 280 31121 336
rect 31177 280 32603 336
rect 32659 280 34085 336
rect 34141 280 35567 336
rect 35623 280 37049 336
rect 37105 280 38531 336
rect 38587 280 40013 336
rect 40069 280 41495 336
rect 41551 280 42977 336
rect 43033 280 44459 336
rect 44515 280 45941 336
rect 45997 280 47424 336
rect -39 278 47424 280
rect -39 275 93 278
rect 1443 275 1575 278
rect 2925 275 3057 278
rect 4407 275 4539 278
rect 5889 275 6021 278
rect 7371 275 7503 278
rect 8853 275 8985 278
rect 10335 275 10467 278
rect 11817 275 11949 278
rect 13299 275 13431 278
rect 14781 275 14913 278
rect 16263 275 16395 278
rect 17745 275 17877 278
rect 19227 275 19359 278
rect 20709 275 20841 278
rect 22191 275 22323 278
rect 23673 275 23805 278
rect 25155 275 25287 278
rect 26637 275 26769 278
rect 28119 275 28251 278
rect 29601 275 29733 278
rect 31083 275 31215 278
rect 32565 275 32697 278
rect 34047 275 34179 278
rect 35529 275 35661 278
rect 37011 275 37143 278
rect 38493 275 38625 278
rect 39975 275 40107 278
rect 41457 275 41589 278
rect 42939 275 43071 278
rect 44421 275 44553 278
rect 45903 275 46035 278
rect 675 28 807 37
rect 675 -28 713 28
rect 769 -28 807 28
rect 675 -37 807 -28
rect 2157 28 2289 37
rect 2157 -28 2195 28
rect 2251 -28 2289 28
rect 2157 -37 2289 -28
rect 3639 28 3771 37
rect 3639 -28 3677 28
rect 3733 -28 3771 28
rect 3639 -37 3771 -28
rect 5121 28 5253 37
rect 5121 -28 5159 28
rect 5215 -28 5253 28
rect 5121 -37 5253 -28
rect 6603 28 6735 37
rect 6603 -28 6641 28
rect 6697 -28 6735 28
rect 6603 -37 6735 -28
rect 8085 28 8217 37
rect 8085 -28 8123 28
rect 8179 -28 8217 28
rect 8085 -37 8217 -28
rect 9567 28 9699 37
rect 9567 -28 9605 28
rect 9661 -28 9699 28
rect 9567 -37 9699 -28
rect 11049 28 11181 37
rect 11049 -28 11087 28
rect 11143 -28 11181 28
rect 11049 -37 11181 -28
rect 12531 28 12663 37
rect 12531 -28 12569 28
rect 12625 -28 12663 28
rect 12531 -37 12663 -28
rect 14013 28 14145 37
rect 14013 -28 14051 28
rect 14107 -28 14145 28
rect 14013 -37 14145 -28
rect 15495 28 15627 37
rect 15495 -28 15533 28
rect 15589 -28 15627 28
rect 15495 -37 15627 -28
rect 16977 28 17109 37
rect 16977 -28 17015 28
rect 17071 -28 17109 28
rect 16977 -37 17109 -28
rect 18459 28 18591 37
rect 18459 -28 18497 28
rect 18553 -28 18591 28
rect 18459 -37 18591 -28
rect 19941 28 20073 37
rect 19941 -28 19979 28
rect 20035 -28 20073 28
rect 19941 -37 20073 -28
rect 21423 28 21555 37
rect 21423 -28 21461 28
rect 21517 -28 21555 28
rect 21423 -37 21555 -28
rect 22905 28 23037 37
rect 22905 -28 22943 28
rect 22999 -28 23037 28
rect 22905 -37 23037 -28
rect 24387 28 24519 37
rect 24387 -28 24425 28
rect 24481 -28 24519 28
rect 24387 -37 24519 -28
rect 25869 28 26001 37
rect 25869 -28 25907 28
rect 25963 -28 26001 28
rect 25869 -37 26001 -28
rect 27351 28 27483 37
rect 27351 -28 27389 28
rect 27445 -28 27483 28
rect 27351 -37 27483 -28
rect 28833 28 28965 37
rect 28833 -28 28871 28
rect 28927 -28 28965 28
rect 28833 -37 28965 -28
rect 30315 28 30447 37
rect 30315 -28 30353 28
rect 30409 -28 30447 28
rect 30315 -37 30447 -28
rect 31797 28 31929 37
rect 31797 -28 31835 28
rect 31891 -28 31929 28
rect 31797 -37 31929 -28
rect 33279 28 33411 37
rect 33279 -28 33317 28
rect 33373 -28 33411 28
rect 33279 -37 33411 -28
rect 34761 28 34893 37
rect 34761 -28 34799 28
rect 34855 -28 34893 28
rect 34761 -37 34893 -28
rect 36243 28 36375 37
rect 36243 -28 36281 28
rect 36337 -28 36375 28
rect 36243 -37 36375 -28
rect 37725 28 37857 37
rect 37725 -28 37763 28
rect 37819 -28 37857 28
rect 37725 -37 37857 -28
rect 39207 28 39339 37
rect 39207 -28 39245 28
rect 39301 -28 39339 28
rect 39207 -37 39339 -28
rect 40689 28 40821 37
rect 40689 -28 40727 28
rect 40783 -28 40821 28
rect 40689 -37 40821 -28
rect 42171 28 42303 37
rect 42171 -28 42209 28
rect 42265 -28 42303 28
rect 42171 -37 42303 -28
rect 43653 28 43785 37
rect 43653 -28 43691 28
rect 43747 -28 43785 28
rect 43653 -37 43785 -28
rect 45135 28 45267 37
rect 45135 -28 45173 28
rect 45229 -28 45267 28
rect 45135 -37 45267 -28
rect 46617 28 46749 37
rect 46617 -28 46655 28
rect 46711 -28 46749 28
rect 46617 -37 46749 -28
use contact_18  contact_18_0
timestamp 1644969367
transform 1 0 45903 0 1 271
box 0 0 1 1
use contact_18  contact_18_1
timestamp 1644969367
transform 1 0 44421 0 1 271
box 0 0 1 1
use contact_18  contact_18_2
timestamp 1644969367
transform 1 0 42939 0 1 271
box 0 0 1 1
use contact_18  contact_18_3
timestamp 1644969367
transform 1 0 41457 0 1 271
box 0 0 1 1
use contact_18  contact_18_4
timestamp 1644969367
transform 1 0 39975 0 1 271
box 0 0 1 1
use contact_18  contact_18_5
timestamp 1644969367
transform 1 0 38493 0 1 271
box 0 0 1 1
use contact_18  contact_18_6
timestamp 1644969367
transform 1 0 37011 0 1 271
box 0 0 1 1
use contact_18  contact_18_7
timestamp 1644969367
transform 1 0 35529 0 1 271
box 0 0 1 1
use contact_18  contact_18_8
timestamp 1644969367
transform 1 0 34047 0 1 271
box 0 0 1 1
use contact_18  contact_18_9
timestamp 1644969367
transform 1 0 32565 0 1 271
box 0 0 1 1
use contact_18  contact_18_10
timestamp 1644969367
transform 1 0 31083 0 1 271
box 0 0 1 1
use contact_18  contact_18_11
timestamp 1644969367
transform 1 0 29601 0 1 271
box 0 0 1 1
use contact_18  contact_18_12
timestamp 1644969367
transform 1 0 28119 0 1 271
box 0 0 1 1
use contact_18  contact_18_13
timestamp 1644969367
transform 1 0 26637 0 1 271
box 0 0 1 1
use contact_18  contact_18_14
timestamp 1644969367
transform 1 0 25155 0 1 271
box 0 0 1 1
use contact_18  contact_18_15
timestamp 1644969367
transform 1 0 23673 0 1 271
box 0 0 1 1
use contact_18  contact_18_16
timestamp 1644969367
transform 1 0 22191 0 1 271
box 0 0 1 1
use contact_18  contact_18_17
timestamp 1644969367
transform 1 0 20709 0 1 271
box 0 0 1 1
use contact_18  contact_18_18
timestamp 1644969367
transform 1 0 19227 0 1 271
box 0 0 1 1
use contact_18  contact_18_19
timestamp 1644969367
transform 1 0 17745 0 1 271
box 0 0 1 1
use contact_18  contact_18_20
timestamp 1644969367
transform 1 0 16263 0 1 271
box 0 0 1 1
use contact_18  contact_18_21
timestamp 1644969367
transform 1 0 14781 0 1 271
box 0 0 1 1
use contact_18  contact_18_22
timestamp 1644969367
transform 1 0 13299 0 1 271
box 0 0 1 1
use contact_18  contact_18_23
timestamp 1644969367
transform 1 0 11817 0 1 271
box 0 0 1 1
use contact_18  contact_18_24
timestamp 1644969367
transform 1 0 10335 0 1 271
box 0 0 1 1
use contact_18  contact_18_25
timestamp 1644969367
transform 1 0 8853 0 1 271
box 0 0 1 1
use contact_18  contact_18_26
timestamp 1644969367
transform 1 0 7371 0 1 271
box 0 0 1 1
use contact_18  contact_18_27
timestamp 1644969367
transform 1 0 5889 0 1 271
box 0 0 1 1
use contact_18  contact_18_28
timestamp 1644969367
transform 1 0 4407 0 1 271
box 0 0 1 1
use contact_18  contact_18_29
timestamp 1644969367
transform 1 0 2925 0 1 271
box 0 0 1 1
use contact_18  contact_18_30
timestamp 1644969367
transform 1 0 1443 0 1 271
box 0 0 1 1
use contact_18  contact_18_31
timestamp 1644969367
transform 1 0 -39 0 1 271
box 0 0 1 1
use contact_18  contact_18_32
timestamp 1644969367
transform 1 0 46617 0 1 -37
box 0 0 1 1
use contact_17  contact_17_0
timestamp 1644969367
transform 1 0 46651 0 1 -32
box 0 0 1 1
use contact_18  contact_18_33
timestamp 1644969367
transform 1 0 46617 0 1 801
box 0 0 1 1
use contact_17  contact_17_1
timestamp 1644969367
transform 1 0 46651 0 1 806
box 0 0 1 1
use contact_18  contact_18_34
timestamp 1644969367
transform 1 0 45135 0 1 -37
box 0 0 1 1
use contact_17  contact_17_2
timestamp 1644969367
transform 1 0 45169 0 1 -32
box 0 0 1 1
use contact_18  contact_18_35
timestamp 1644969367
transform 1 0 45135 0 1 801
box 0 0 1 1
use contact_17  contact_17_3
timestamp 1644969367
transform 1 0 45169 0 1 806
box 0 0 1 1
use contact_18  contact_18_36
timestamp 1644969367
transform 1 0 43653 0 1 -37
box 0 0 1 1
use contact_17  contact_17_4
timestamp 1644969367
transform 1 0 43687 0 1 -32
box 0 0 1 1
use contact_18  contact_18_37
timestamp 1644969367
transform 1 0 43653 0 1 801
box 0 0 1 1
use contact_17  contact_17_5
timestamp 1644969367
transform 1 0 43687 0 1 806
box 0 0 1 1
use contact_18  contact_18_38
timestamp 1644969367
transform 1 0 42171 0 1 -37
box 0 0 1 1
use contact_17  contact_17_6
timestamp 1644969367
transform 1 0 42205 0 1 -32
box 0 0 1 1
use contact_18  contact_18_39
timestamp 1644969367
transform 1 0 42171 0 1 801
box 0 0 1 1
use contact_17  contact_17_7
timestamp 1644969367
transform 1 0 42205 0 1 806
box 0 0 1 1
use contact_18  contact_18_40
timestamp 1644969367
transform 1 0 40689 0 1 -37
box 0 0 1 1
use contact_17  contact_17_8
timestamp 1644969367
transform 1 0 40723 0 1 -32
box 0 0 1 1
use contact_18  contact_18_41
timestamp 1644969367
transform 1 0 40689 0 1 801
box 0 0 1 1
use contact_17  contact_17_9
timestamp 1644969367
transform 1 0 40723 0 1 806
box 0 0 1 1
use contact_18  contact_18_42
timestamp 1644969367
transform 1 0 39207 0 1 -37
box 0 0 1 1
use contact_17  contact_17_10
timestamp 1644969367
transform 1 0 39241 0 1 -32
box 0 0 1 1
use contact_18  contact_18_43
timestamp 1644969367
transform 1 0 39207 0 1 801
box 0 0 1 1
use contact_17  contact_17_11
timestamp 1644969367
transform 1 0 39241 0 1 806
box 0 0 1 1
use contact_18  contact_18_44
timestamp 1644969367
transform 1 0 37725 0 1 -37
box 0 0 1 1
use contact_17  contact_17_12
timestamp 1644969367
transform 1 0 37759 0 1 -32
box 0 0 1 1
use contact_18  contact_18_45
timestamp 1644969367
transform 1 0 37725 0 1 801
box 0 0 1 1
use contact_17  contact_17_13
timestamp 1644969367
transform 1 0 37759 0 1 806
box 0 0 1 1
use contact_18  contact_18_46
timestamp 1644969367
transform 1 0 36243 0 1 -37
box 0 0 1 1
use contact_17  contact_17_14
timestamp 1644969367
transform 1 0 36277 0 1 -32
box 0 0 1 1
use contact_18  contact_18_47
timestamp 1644969367
transform 1 0 36243 0 1 801
box 0 0 1 1
use contact_17  contact_17_15
timestamp 1644969367
transform 1 0 36277 0 1 806
box 0 0 1 1
use contact_18  contact_18_48
timestamp 1644969367
transform 1 0 34761 0 1 -37
box 0 0 1 1
use contact_17  contact_17_16
timestamp 1644969367
transform 1 0 34795 0 1 -32
box 0 0 1 1
use contact_18  contact_18_49
timestamp 1644969367
transform 1 0 34761 0 1 801
box 0 0 1 1
use contact_17  contact_17_17
timestamp 1644969367
transform 1 0 34795 0 1 806
box 0 0 1 1
use contact_18  contact_18_50
timestamp 1644969367
transform 1 0 33279 0 1 -37
box 0 0 1 1
use contact_17  contact_17_18
timestamp 1644969367
transform 1 0 33313 0 1 -32
box 0 0 1 1
use contact_18  contact_18_51
timestamp 1644969367
transform 1 0 33279 0 1 801
box 0 0 1 1
use contact_17  contact_17_19
timestamp 1644969367
transform 1 0 33313 0 1 806
box 0 0 1 1
use contact_18  contact_18_52
timestamp 1644969367
transform 1 0 31797 0 1 -37
box 0 0 1 1
use contact_17  contact_17_20
timestamp 1644969367
transform 1 0 31831 0 1 -32
box 0 0 1 1
use contact_18  contact_18_53
timestamp 1644969367
transform 1 0 31797 0 1 801
box 0 0 1 1
use contact_17  contact_17_21
timestamp 1644969367
transform 1 0 31831 0 1 806
box 0 0 1 1
use contact_18  contact_18_54
timestamp 1644969367
transform 1 0 30315 0 1 -37
box 0 0 1 1
use contact_17  contact_17_22
timestamp 1644969367
transform 1 0 30349 0 1 -32
box 0 0 1 1
use contact_18  contact_18_55
timestamp 1644969367
transform 1 0 30315 0 1 801
box 0 0 1 1
use contact_17  contact_17_23
timestamp 1644969367
transform 1 0 30349 0 1 806
box 0 0 1 1
use contact_18  contact_18_56
timestamp 1644969367
transform 1 0 28833 0 1 -37
box 0 0 1 1
use contact_17  contact_17_24
timestamp 1644969367
transform 1 0 28867 0 1 -32
box 0 0 1 1
use contact_18  contact_18_57
timestamp 1644969367
transform 1 0 28833 0 1 801
box 0 0 1 1
use contact_17  contact_17_25
timestamp 1644969367
transform 1 0 28867 0 1 806
box 0 0 1 1
use contact_18  contact_18_58
timestamp 1644969367
transform 1 0 27351 0 1 -37
box 0 0 1 1
use contact_17  contact_17_26
timestamp 1644969367
transform 1 0 27385 0 1 -32
box 0 0 1 1
use contact_18  contact_18_59
timestamp 1644969367
transform 1 0 27351 0 1 801
box 0 0 1 1
use contact_17  contact_17_27
timestamp 1644969367
transform 1 0 27385 0 1 806
box 0 0 1 1
use contact_18  contact_18_60
timestamp 1644969367
transform 1 0 25869 0 1 -37
box 0 0 1 1
use contact_17  contact_17_28
timestamp 1644969367
transform 1 0 25903 0 1 -32
box 0 0 1 1
use contact_18  contact_18_61
timestamp 1644969367
transform 1 0 25869 0 1 801
box 0 0 1 1
use contact_17  contact_17_29
timestamp 1644969367
transform 1 0 25903 0 1 806
box 0 0 1 1
use contact_18  contact_18_62
timestamp 1644969367
transform 1 0 24387 0 1 -37
box 0 0 1 1
use contact_17  contact_17_30
timestamp 1644969367
transform 1 0 24421 0 1 -32
box 0 0 1 1
use contact_18  contact_18_63
timestamp 1644969367
transform 1 0 24387 0 1 801
box 0 0 1 1
use contact_17  contact_17_31
timestamp 1644969367
transform 1 0 24421 0 1 806
box 0 0 1 1
use contact_18  contact_18_64
timestamp 1644969367
transform 1 0 22905 0 1 -37
box 0 0 1 1
use contact_17  contact_17_32
timestamp 1644969367
transform 1 0 22939 0 1 -32
box 0 0 1 1
use contact_18  contact_18_65
timestamp 1644969367
transform 1 0 22905 0 1 801
box 0 0 1 1
use contact_17  contact_17_33
timestamp 1644969367
transform 1 0 22939 0 1 806
box 0 0 1 1
use contact_18  contact_18_66
timestamp 1644969367
transform 1 0 21423 0 1 -37
box 0 0 1 1
use contact_17  contact_17_34
timestamp 1644969367
transform 1 0 21457 0 1 -32
box 0 0 1 1
use contact_18  contact_18_67
timestamp 1644969367
transform 1 0 21423 0 1 801
box 0 0 1 1
use contact_17  contact_17_35
timestamp 1644969367
transform 1 0 21457 0 1 806
box 0 0 1 1
use contact_18  contact_18_68
timestamp 1644969367
transform 1 0 19941 0 1 -37
box 0 0 1 1
use contact_17  contact_17_36
timestamp 1644969367
transform 1 0 19975 0 1 -32
box 0 0 1 1
use contact_18  contact_18_69
timestamp 1644969367
transform 1 0 19941 0 1 801
box 0 0 1 1
use contact_17  contact_17_37
timestamp 1644969367
transform 1 0 19975 0 1 806
box 0 0 1 1
use contact_18  contact_18_70
timestamp 1644969367
transform 1 0 18459 0 1 -37
box 0 0 1 1
use contact_17  contact_17_38
timestamp 1644969367
transform 1 0 18493 0 1 -32
box 0 0 1 1
use contact_18  contact_18_71
timestamp 1644969367
transform 1 0 18459 0 1 801
box 0 0 1 1
use contact_17  contact_17_39
timestamp 1644969367
transform 1 0 18493 0 1 806
box 0 0 1 1
use contact_18  contact_18_72
timestamp 1644969367
transform 1 0 16977 0 1 -37
box 0 0 1 1
use contact_17  contact_17_40
timestamp 1644969367
transform 1 0 17011 0 1 -32
box 0 0 1 1
use contact_18  contact_18_73
timestamp 1644969367
transform 1 0 16977 0 1 801
box 0 0 1 1
use contact_17  contact_17_41
timestamp 1644969367
transform 1 0 17011 0 1 806
box 0 0 1 1
use contact_18  contact_18_74
timestamp 1644969367
transform 1 0 15495 0 1 -37
box 0 0 1 1
use contact_17  contact_17_42
timestamp 1644969367
transform 1 0 15529 0 1 -32
box 0 0 1 1
use contact_18  contact_18_75
timestamp 1644969367
transform 1 0 15495 0 1 801
box 0 0 1 1
use contact_17  contact_17_43
timestamp 1644969367
transform 1 0 15529 0 1 806
box 0 0 1 1
use contact_18  contact_18_76
timestamp 1644969367
transform 1 0 14013 0 1 -37
box 0 0 1 1
use contact_17  contact_17_44
timestamp 1644969367
transform 1 0 14047 0 1 -32
box 0 0 1 1
use contact_18  contact_18_77
timestamp 1644969367
transform 1 0 14013 0 1 801
box 0 0 1 1
use contact_17  contact_17_45
timestamp 1644969367
transform 1 0 14047 0 1 806
box 0 0 1 1
use contact_18  contact_18_78
timestamp 1644969367
transform 1 0 12531 0 1 -37
box 0 0 1 1
use contact_17  contact_17_46
timestamp 1644969367
transform 1 0 12565 0 1 -32
box 0 0 1 1
use contact_18  contact_18_79
timestamp 1644969367
transform 1 0 12531 0 1 801
box 0 0 1 1
use contact_17  contact_17_47
timestamp 1644969367
transform 1 0 12565 0 1 806
box 0 0 1 1
use contact_18  contact_18_80
timestamp 1644969367
transform 1 0 11049 0 1 -37
box 0 0 1 1
use contact_17  contact_17_48
timestamp 1644969367
transform 1 0 11083 0 1 -32
box 0 0 1 1
use contact_18  contact_18_81
timestamp 1644969367
transform 1 0 11049 0 1 801
box 0 0 1 1
use contact_17  contact_17_49
timestamp 1644969367
transform 1 0 11083 0 1 806
box 0 0 1 1
use contact_18  contact_18_82
timestamp 1644969367
transform 1 0 9567 0 1 -37
box 0 0 1 1
use contact_17  contact_17_50
timestamp 1644969367
transform 1 0 9601 0 1 -32
box 0 0 1 1
use contact_18  contact_18_83
timestamp 1644969367
transform 1 0 9567 0 1 801
box 0 0 1 1
use contact_17  contact_17_51
timestamp 1644969367
transform 1 0 9601 0 1 806
box 0 0 1 1
use contact_18  contact_18_84
timestamp 1644969367
transform 1 0 8085 0 1 -37
box 0 0 1 1
use contact_17  contact_17_52
timestamp 1644969367
transform 1 0 8119 0 1 -32
box 0 0 1 1
use contact_18  contact_18_85
timestamp 1644969367
transform 1 0 8085 0 1 801
box 0 0 1 1
use contact_17  contact_17_53
timestamp 1644969367
transform 1 0 8119 0 1 806
box 0 0 1 1
use contact_18  contact_18_86
timestamp 1644969367
transform 1 0 6603 0 1 -37
box 0 0 1 1
use contact_17  contact_17_54
timestamp 1644969367
transform 1 0 6637 0 1 -32
box 0 0 1 1
use contact_18  contact_18_87
timestamp 1644969367
transform 1 0 6603 0 1 801
box 0 0 1 1
use contact_17  contact_17_55
timestamp 1644969367
transform 1 0 6637 0 1 806
box 0 0 1 1
use contact_18  contact_18_88
timestamp 1644969367
transform 1 0 5121 0 1 -37
box 0 0 1 1
use contact_17  contact_17_56
timestamp 1644969367
transform 1 0 5155 0 1 -32
box 0 0 1 1
use contact_18  contact_18_89
timestamp 1644969367
transform 1 0 5121 0 1 801
box 0 0 1 1
use contact_17  contact_17_57
timestamp 1644969367
transform 1 0 5155 0 1 806
box 0 0 1 1
use contact_18  contact_18_90
timestamp 1644969367
transform 1 0 3639 0 1 -37
box 0 0 1 1
use contact_17  contact_17_58
timestamp 1644969367
transform 1 0 3673 0 1 -32
box 0 0 1 1
use contact_18  contact_18_91
timestamp 1644969367
transform 1 0 3639 0 1 801
box 0 0 1 1
use contact_17  contact_17_59
timestamp 1644969367
transform 1 0 3673 0 1 806
box 0 0 1 1
use contact_18  contact_18_92
timestamp 1644969367
transform 1 0 2157 0 1 -37
box 0 0 1 1
use contact_17  contact_17_60
timestamp 1644969367
transform 1 0 2191 0 1 -32
box 0 0 1 1
use contact_18  contact_18_93
timestamp 1644969367
transform 1 0 2157 0 1 801
box 0 0 1 1
use contact_17  contact_17_61
timestamp 1644969367
transform 1 0 2191 0 1 806
box 0 0 1 1
use contact_18  contact_18_94
timestamp 1644969367
transform 1 0 675 0 1 -37
box 0 0 1 1
use contact_17  contact_17_62
timestamp 1644969367
transform 1 0 709 0 1 -32
box 0 0 1 1
use contact_18  contact_18_95
timestamp 1644969367
transform 1 0 675 0 1 801
box 0 0 1 1
use contact_17  contact_17_63
timestamp 1644969367
transform 1 0 709 0 1 806
box 0 0 1 1
use dff  dff_0
timestamp 1644969367
transform 1 0 45942 0 1 0
box 0 -42 1482 916
use dff  dff_1
timestamp 1644969367
transform 1 0 44460 0 1 0
box 0 -42 1482 916
use dff  dff_2
timestamp 1644969367
transform 1 0 42978 0 1 0
box 0 -42 1482 916
use dff  dff_3
timestamp 1644969367
transform 1 0 41496 0 1 0
box 0 -42 1482 916
use dff  dff_4
timestamp 1644969367
transform 1 0 40014 0 1 0
box 0 -42 1482 916
use dff  dff_5
timestamp 1644969367
transform 1 0 38532 0 1 0
box 0 -42 1482 916
use dff  dff_6
timestamp 1644969367
transform 1 0 37050 0 1 0
box 0 -42 1482 916
use dff  dff_7
timestamp 1644969367
transform 1 0 35568 0 1 0
box 0 -42 1482 916
use dff  dff_8
timestamp 1644969367
transform 1 0 34086 0 1 0
box 0 -42 1482 916
use dff  dff_9
timestamp 1644969367
transform 1 0 32604 0 1 0
box 0 -42 1482 916
use dff  dff_10
timestamp 1644969367
transform 1 0 31122 0 1 0
box 0 -42 1482 916
use dff  dff_11
timestamp 1644969367
transform 1 0 29640 0 1 0
box 0 -42 1482 916
use dff  dff_12
timestamp 1644969367
transform 1 0 28158 0 1 0
box 0 -42 1482 916
use dff  dff_13
timestamp 1644969367
transform 1 0 26676 0 1 0
box 0 -42 1482 916
use dff  dff_14
timestamp 1644969367
transform 1 0 25194 0 1 0
box 0 -42 1482 916
use dff  dff_15
timestamp 1644969367
transform 1 0 23712 0 1 0
box 0 -42 1482 916
use dff  dff_16
timestamp 1644969367
transform 1 0 22230 0 1 0
box 0 -42 1482 916
use dff  dff_17
timestamp 1644969367
transform 1 0 20748 0 1 0
box 0 -42 1482 916
use dff  dff_18
timestamp 1644969367
transform 1 0 19266 0 1 0
box 0 -42 1482 916
use dff  dff_19
timestamp 1644969367
transform 1 0 17784 0 1 0
box 0 -42 1482 916
use dff  dff_20
timestamp 1644969367
transform 1 0 16302 0 1 0
box 0 -42 1482 916
use dff  dff_21
timestamp 1644969367
transform 1 0 14820 0 1 0
box 0 -42 1482 916
use dff  dff_22
timestamp 1644969367
transform 1 0 13338 0 1 0
box 0 -42 1482 916
use dff  dff_23
timestamp 1644969367
transform 1 0 11856 0 1 0
box 0 -42 1482 916
use dff  dff_24
timestamp 1644969367
transform 1 0 10374 0 1 0
box 0 -42 1482 916
use dff  dff_25
timestamp 1644969367
transform 1 0 8892 0 1 0
box 0 -42 1482 916
use dff  dff_26
timestamp 1644969367
transform 1 0 7410 0 1 0
box 0 -42 1482 916
use dff  dff_27
timestamp 1644969367
transform 1 0 5928 0 1 0
box 0 -42 1482 916
use dff  dff_28
timestamp 1644969367
transform 1 0 4446 0 1 0
box 0 -42 1482 916
use dff  dff_29
timestamp 1644969367
transform 1 0 2964 0 1 0
box 0 -42 1482 916
use dff  dff_30
timestamp 1644969367
transform 1 0 1482 0 1 0
box 0 -42 1482 916
use dff  dff_31
timestamp 1644969367
transform 1 0 0 0 1 0
box 0 -42 1482 916
<< labels >>
rlabel metal3 s 30315 801 30447 875 4 vdd
rlabel metal3 s 46617 801 46749 875 4 vdd
rlabel metal3 s 43653 801 43785 875 4 vdd
rlabel metal3 s 42171 801 42303 875 4 vdd
rlabel metal3 s 25869 801 26001 875 4 vdd
rlabel metal3 s 12531 801 12663 875 4 vdd
rlabel metal3 s 34761 801 34893 875 4 vdd
rlabel metal3 s 33279 801 33411 875 4 vdd
rlabel metal3 s 19941 801 20073 875 4 vdd
rlabel metal3 s 31797 801 31929 875 4 vdd
rlabel metal3 s 37725 801 37857 875 4 vdd
rlabel metal3 s 11049 801 11181 875 4 vdd
rlabel metal3 s 6603 801 6735 875 4 vdd
rlabel metal3 s 16977 801 17109 875 4 vdd
rlabel metal3 s 3639 801 3771 875 4 vdd
rlabel metal3 s 9567 801 9699 875 4 vdd
rlabel metal3 s 15495 801 15627 875 4 vdd
rlabel metal3 s 18459 801 18591 875 4 vdd
rlabel metal3 s 28833 801 28965 875 4 vdd
rlabel metal3 s 675 801 807 875 4 vdd
rlabel metal3 s 36243 801 36375 875 4 vdd
rlabel metal3 s 21423 801 21555 875 4 vdd
rlabel metal3 s 2157 801 2289 875 4 vdd
rlabel metal3 s 24387 801 24519 875 4 vdd
rlabel metal3 s 39207 801 39339 875 4 vdd
rlabel metal3 s 8085 801 8217 875 4 vdd
rlabel metal3 s 5121 801 5253 875 4 vdd
rlabel metal3 s 40689 801 40821 875 4 vdd
rlabel metal3 s 45135 801 45267 875 4 vdd
rlabel metal3 s 27351 801 27483 875 4 vdd
rlabel metal3 s 14013 801 14145 875 4 vdd
rlabel metal3 s 22905 801 23037 875 4 vdd
rlabel metal3 s 3639 -37 3771 37 4 gnd
rlabel metal3 s 30315 -37 30447 37 4 gnd
rlabel metal3 s 8085 -37 8217 37 4 gnd
rlabel metal3 s 12531 -37 12663 37 4 gnd
rlabel metal3 s 14013 -37 14145 37 4 gnd
rlabel metal3 s 5121 -37 5253 37 4 gnd
rlabel metal3 s 675 -37 807 37 4 gnd
rlabel metal3 s 24387 -37 24519 37 4 gnd
rlabel metal3 s 15495 -37 15627 37 4 gnd
rlabel metal3 s 39207 -37 39339 37 4 gnd
rlabel metal3 s 6603 -37 6735 37 4 gnd
rlabel metal3 s 34761 -37 34893 37 4 gnd
rlabel metal3 s 25869 -37 26001 37 4 gnd
rlabel metal3 s 43653 -37 43785 37 4 gnd
rlabel metal3 s 45135 -37 45267 37 4 gnd
rlabel metal3 s 28833 -37 28965 37 4 gnd
rlabel metal3 s 11049 -37 11181 37 4 gnd
rlabel metal3 s 2157 -37 2289 37 4 gnd
rlabel metal3 s 9567 -37 9699 37 4 gnd
rlabel metal3 s 37725 -37 37857 37 4 gnd
rlabel metal3 s 22905 -37 23037 37 4 gnd
rlabel metal3 s 36243 -37 36375 37 4 gnd
rlabel metal3 s 18459 -37 18591 37 4 gnd
rlabel metal3 s 31797 -37 31929 37 4 gnd
rlabel metal3 s 42171 -37 42303 37 4 gnd
rlabel metal3 s 19941 -37 20073 37 4 gnd
rlabel metal3 s 33279 -37 33411 37 4 gnd
rlabel metal3 s 46617 -37 46749 37 4 gnd
rlabel metal3 s 40689 -37 40821 37 4 gnd
rlabel metal3 s 21423 -37 21555 37 4 gnd
rlabel metal3 s 27351 -37 27483 37 4 gnd
rlabel metal3 s 16977 -37 17109 37 4 gnd
rlabel metal2 s 180 232 234 260 4 din_0
rlabel metal2 s 1260 228 1314 256 4 dout_0
rlabel metal2 s 1662 232 1716 260 4 din_1
rlabel metal2 s 2742 228 2796 256 4 dout_1
rlabel metal2 s 3144 232 3198 260 4 din_2
rlabel metal2 s 4224 228 4278 256 4 dout_2
rlabel metal2 s 4626 232 4680 260 4 din_3
rlabel metal2 s 5706 228 5760 256 4 dout_3
rlabel metal2 s 6108 232 6162 260 4 din_4
rlabel metal2 s 7188 228 7242 256 4 dout_4
rlabel metal2 s 7590 232 7644 260 4 din_5
rlabel metal2 s 8670 228 8724 256 4 dout_5
rlabel metal2 s 9072 232 9126 260 4 din_6
rlabel metal2 s 10152 228 10206 256 4 dout_6
rlabel metal2 s 10554 232 10608 260 4 din_7
rlabel metal2 s 11634 228 11688 256 4 dout_7
rlabel metal2 s 12036 232 12090 260 4 din_8
rlabel metal2 s 13116 228 13170 256 4 dout_8
rlabel metal2 s 13518 232 13572 260 4 din_9
rlabel metal2 s 14598 228 14652 256 4 dout_9
rlabel metal2 s 15000 232 15054 260 4 din_10
rlabel metal2 s 16080 228 16134 256 4 dout_10
rlabel metal2 s 16482 232 16536 260 4 din_11
rlabel metal2 s 17562 228 17616 256 4 dout_11
rlabel metal2 s 17964 232 18018 260 4 din_12
rlabel metal2 s 19044 228 19098 256 4 dout_12
rlabel metal2 s 19446 232 19500 260 4 din_13
rlabel metal2 s 20526 228 20580 256 4 dout_13
rlabel metal2 s 20928 232 20982 260 4 din_14
rlabel metal2 s 22008 228 22062 256 4 dout_14
rlabel metal2 s 22410 232 22464 260 4 din_15
rlabel metal2 s 23490 228 23544 256 4 dout_15
rlabel metal2 s 23892 232 23946 260 4 din_16
rlabel metal2 s 24972 228 25026 256 4 dout_16
rlabel metal2 s 25374 232 25428 260 4 din_17
rlabel metal2 s 26454 228 26508 256 4 dout_17
rlabel metal2 s 26856 232 26910 260 4 din_18
rlabel metal2 s 27936 228 27990 256 4 dout_18
rlabel metal2 s 28338 232 28392 260 4 din_19
rlabel metal2 s 29418 228 29472 256 4 dout_19
rlabel metal2 s 29820 232 29874 260 4 din_20
rlabel metal2 s 30900 228 30954 256 4 dout_20
rlabel metal2 s 31302 232 31356 260 4 din_21
rlabel metal2 s 32382 228 32436 256 4 dout_21
rlabel metal2 s 32784 232 32838 260 4 din_22
rlabel metal2 s 33864 228 33918 256 4 dout_22
rlabel metal2 s 34266 232 34320 260 4 din_23
rlabel metal2 s 35346 228 35400 256 4 dout_23
rlabel metal2 s 35748 232 35802 260 4 din_24
rlabel metal2 s 36828 228 36882 256 4 dout_24
rlabel metal2 s 37230 232 37284 260 4 din_25
rlabel metal2 s 38310 228 38364 256 4 dout_25
rlabel metal2 s 38712 232 38766 260 4 din_26
rlabel metal2 s 39792 228 39846 256 4 dout_26
rlabel metal2 s 40194 232 40248 260 4 din_27
rlabel metal2 s 41274 228 41328 256 4 dout_27
rlabel metal2 s 41676 232 41730 260 4 din_28
rlabel metal2 s 42756 228 42810 256 4 dout_28
rlabel metal2 s 43158 232 43212 260 4 din_29
rlabel metal2 s 44238 228 44292 256 4 dout_29
rlabel metal2 s 44640 232 44694 260 4 din_30
rlabel metal2 s 45720 228 45774 256 4 dout_30
rlabel metal2 s 46122 232 46176 260 4 din_31
rlabel metal2 s 47202 228 47256 256 4 dout_31
rlabel metal3 s 0 278 47424 338 4 clk
<< properties >>
string FIXED_BBOX 46617 -37 46749 0
string GDS_FILE sram_0rw2r1w_32_128_sky130A.gds
string GDS_END 3465540
string GDS_START 3427610
<< end >>
