magic
tech sky130A
magscale 1 2
timestamp 1644969367
<< checkpaint >>
rect -1296 -1277 5606 2155
<< locali >>
rect 0 821 4310 855
rect 196 381 262 447
rect 330 386 364 561
rect 330 352 459 386
rect 2289 352 2323 386
rect 96 257 162 323
rect 0 -17 4310 17
use pdriver_2  pdriver_2_0
timestamp 1644969367
transform 1 0 378 0 1 0
box -36 -17 3968 895
use pnand2_0  pnand2_0_0
timestamp 1644969367
transform 1 0 0 0 1 0
box -36 -17 414 895
<< labels >>
rlabel locali s 2306 369 2306 369 4 Z
rlabel locali s 129 290 129 290 4 A
rlabel locali s 229 414 229 414 4 B
rlabel locali s 2155 0 2155 0 4 gnd
rlabel locali s 2155 838 2155 838 4 vdd
<< properties >>
string FIXED_BBOX 0 0 4310 838
string GDS_FILE sram_0rw2r1w_32_128_sky130A.gds
string GDS_END 3393758
string GDS_START 3392624
<< end >>
