magic
tech sky130A
magscale 1 2
timestamp 1644969367
<< checkpaint >>
rect -1319 -1316 1685 1566
<< nwell >>
rect -54 210 420 306
rect -59 42 425 210
rect -54 -54 420 42
<< scpmos >>
rect 60 0 90 252
rect 168 0 198 252
rect 276 0 306 252
<< pdiff >>
rect 0 143 60 252
rect 0 109 8 143
rect 42 109 60 143
rect 0 0 60 109
rect 90 143 168 252
rect 90 109 112 143
rect 146 109 168 143
rect 90 0 168 109
rect 198 143 276 252
rect 198 109 220 143
rect 254 109 276 143
rect 198 0 276 109
rect 306 143 366 252
rect 306 109 324 143
rect 358 109 366 143
rect 306 0 366 109
<< pdiffc >>
rect 8 109 42 143
rect 112 109 146 143
rect 220 109 254 143
rect 324 109 358 143
<< poly >>
rect 60 252 90 278
rect 168 252 198 278
rect 276 252 306 278
rect 60 -26 90 0
rect 168 -26 198 0
rect 276 -26 306 0
rect 60 -56 306 -26
<< locali >>
rect 8 143 42 159
rect 8 93 42 109
rect 112 143 146 159
rect 112 59 146 109
rect 220 143 254 159
rect 220 93 254 109
rect 324 143 358 159
rect 324 59 358 109
rect 112 25 358 59
use contact_9  contact_9_0
timestamp 1644969367
transform 1 0 316 0 1 85
box 0 0 2 2
use contact_9  contact_9_1
timestamp 1644969367
transform 1 0 212 0 1 85
box 0 0 2 2
use contact_9  contact_9_2
timestamp 1644969367
transform 1 0 104 0 1 85
box 0 0 2 2
use contact_9  contact_9_3
timestamp 1644969367
transform 1 0 0 0 1 85
box 0 0 2 2
<< labels >>
rlabel mvvaractor s 183 -41 183 -41 4 G
rlabel locali s 25 126 25 126 4 S
rlabel locali s 237 126 237 126 4 S
rlabel locali s 235 42 235 42 4 D
<< properties >>
string FIXED_BBOX -54 -56 420 42
string GDS_FILE sram_0rw2r1w_32_128_sky130A.gds
string GDS_END 3309772
string GDS_START 3308488
<< end >>
