magic
tech sky130A
magscale 1 2
timestamp 1643671299
<< checkpaint >>
rect -1260 -1070 54316 6866
<< metal1 >>
rect 0 5222 24038 5250
rect 0 2994 24896 3022
rect 0 2936 24896 2964
rect 0 1171 25674 1199
<< metal2 >>
rect 196 5306 250 5334
rect 1752 5306 1806 5334
rect 3308 5306 3362 5334
rect 4864 5306 4918 5334
rect 6420 5306 6474 5334
rect 7976 5306 8030 5334
rect 9532 5306 9586 5334
rect 11088 5306 11142 5334
rect 12644 5306 12698 5334
rect 14200 5306 14254 5334
rect 15756 5306 15810 5334
rect 17312 5306 17366 5334
rect 18868 5306 18922 5334
rect 20424 5306 20478 5334
rect 21980 5306 22034 5334
rect 23536 5306 23590 5334
rect 630 4654 658 5284
rect 2186 4654 2214 5284
rect 4750 4210 4778 4450
rect 6306 4210 6334 4450
rect 7862 4210 7890 4450
rect 9418 4210 9446 4450
rect 10974 4210 11002 4450
rect 12530 4210 12558 4450
rect 14086 4210 14114 4450
rect 15642 4210 15670 4450
rect 17198 4210 17226 4450
rect 18754 4210 18782 4450
rect 20310 4210 20338 4450
rect 21866 4210 21894 4450
rect 23422 4210 23450 4450
rect 24978 4210 25006 4450
rect 26534 4210 26562 4450
rect 28090 4210 28118 4450
rect 68 1344 96 1398
rect 54 1316 96 1344
rect 54 204 82 1316
rect 710 1276 738 1398
rect 846 1344 874 1398
rect 532 1248 738 1276
rect 832 1316 874 1344
rect 532 204 560 1248
rect 832 204 860 1316
rect 1488 1276 1516 1398
rect 1624 1344 1652 1398
rect 1310 1248 1516 1276
rect 1610 1316 1652 1344
rect 1310 204 1338 1248
rect 1610 204 1638 1316
rect 2266 1276 2294 1398
rect 2402 1344 2430 1398
rect 2088 1248 2294 1276
rect 2388 1316 2430 1344
rect 2088 204 2116 1248
rect 2388 204 2416 1316
rect 3044 1276 3072 1398
rect 3180 1344 3208 1398
rect 2866 1248 3072 1276
rect 3166 1316 3208 1344
rect 2866 204 2894 1248
rect 3166 204 3194 1316
rect 3822 1276 3850 1398
rect 3958 1344 3986 1398
rect 3644 1248 3850 1276
rect 3944 1316 3986 1344
rect 3644 204 3672 1248
rect 3944 204 3972 1316
rect 4600 1276 4628 1398
rect 4736 1344 4764 1398
rect 4422 1248 4628 1276
rect 4722 1316 4764 1344
rect 4422 204 4450 1248
rect 4722 204 4750 1316
rect 5378 1276 5406 1398
rect 5514 1344 5542 1398
rect 5200 1248 5406 1276
rect 5500 1316 5542 1344
rect 5200 204 5228 1248
rect 5500 204 5528 1316
rect 6156 1276 6184 1398
rect 6292 1344 6320 1398
rect 5978 1248 6184 1276
rect 6278 1316 6320 1344
rect 5978 204 6006 1248
rect 6278 204 6306 1316
rect 6934 1276 6962 1398
rect 7070 1344 7098 1398
rect 6756 1248 6962 1276
rect 7056 1316 7098 1344
rect 6756 204 6784 1248
rect 7056 204 7084 1316
rect 7712 1276 7740 1398
rect 7848 1344 7876 1398
rect 7534 1248 7740 1276
rect 7834 1316 7876 1344
rect 7534 204 7562 1248
rect 7834 204 7862 1316
rect 8490 1276 8518 1398
rect 8626 1344 8654 1398
rect 8312 1248 8518 1276
rect 8612 1316 8654 1344
rect 8312 204 8340 1248
rect 8612 204 8640 1316
rect 9268 1276 9296 1398
rect 9404 1344 9432 1398
rect 9090 1248 9296 1276
rect 9390 1316 9432 1344
rect 9090 204 9118 1248
rect 9390 204 9418 1316
rect 10046 1276 10074 1398
rect 10182 1344 10210 1398
rect 9868 1248 10074 1276
rect 10168 1316 10210 1344
rect 9868 204 9896 1248
rect 10168 204 10196 1316
rect 10824 1276 10852 1398
rect 10960 1344 10988 1398
rect 10646 1248 10852 1276
rect 10946 1316 10988 1344
rect 10646 204 10674 1248
rect 10946 204 10974 1316
rect 11602 1276 11630 1398
rect 11738 1344 11766 1398
rect 11424 1248 11630 1276
rect 11724 1316 11766 1344
rect 11424 204 11452 1248
rect 11724 204 11752 1316
rect 12380 1276 12408 1398
rect 12516 1344 12544 1398
rect 12202 1248 12408 1276
rect 12502 1316 12544 1344
rect 12202 204 12230 1248
rect 12502 204 12530 1316
rect 13158 1276 13186 1398
rect 13294 1344 13322 1398
rect 12980 1248 13186 1276
rect 13280 1316 13322 1344
rect 12980 204 13008 1248
rect 13280 204 13308 1316
rect 13936 1276 13964 1398
rect 14072 1344 14100 1398
rect 13758 1248 13964 1276
rect 14058 1316 14100 1344
rect 13758 204 13786 1248
rect 14058 204 14086 1316
rect 14714 1276 14742 1398
rect 14850 1344 14878 1398
rect 14536 1248 14742 1276
rect 14836 1316 14878 1344
rect 14536 204 14564 1248
rect 14836 204 14864 1316
rect 15492 1276 15520 1398
rect 15628 1344 15656 1398
rect 15314 1248 15520 1276
rect 15614 1316 15656 1344
rect 15314 204 15342 1248
rect 15614 204 15642 1316
rect 16270 1276 16298 1398
rect 16406 1344 16434 1398
rect 16092 1248 16298 1276
rect 16392 1316 16434 1344
rect 16092 204 16120 1248
rect 16392 204 16420 1316
rect 17048 1276 17076 1398
rect 17184 1344 17212 1398
rect 16870 1248 17076 1276
rect 17170 1316 17212 1344
rect 16870 204 16898 1248
rect 17170 204 17198 1316
rect 17826 1276 17854 1398
rect 17962 1344 17990 1398
rect 17648 1248 17854 1276
rect 17948 1316 17990 1344
rect 17648 204 17676 1248
rect 17948 204 17976 1316
rect 18604 1276 18632 1398
rect 18740 1344 18768 1398
rect 18426 1248 18632 1276
rect 18726 1316 18768 1344
rect 18426 204 18454 1248
rect 18726 204 18754 1316
rect 19382 1276 19410 1398
rect 19518 1344 19546 1398
rect 19204 1248 19410 1276
rect 19504 1316 19546 1344
rect 19204 204 19232 1248
rect 19504 204 19532 1316
rect 20160 1276 20188 1398
rect 20296 1344 20324 1398
rect 19982 1248 20188 1276
rect 20282 1316 20324 1344
rect 19982 204 20010 1248
rect 20282 204 20310 1316
rect 20938 1276 20966 1398
rect 21074 1344 21102 1398
rect 20760 1248 20966 1276
rect 21060 1316 21102 1344
rect 20760 204 20788 1248
rect 21060 204 21088 1316
rect 21716 1276 21744 1398
rect 21852 1344 21880 1398
rect 21538 1248 21744 1276
rect 21838 1316 21880 1344
rect 21538 204 21566 1248
rect 21838 204 21866 1316
rect 22494 1276 22522 1398
rect 22630 1344 22658 1398
rect 22316 1248 22522 1276
rect 22616 1316 22658 1344
rect 22316 204 22344 1248
rect 22616 204 22644 1316
rect 23272 1276 23300 1398
rect 23408 1344 23436 1398
rect 23094 1248 23300 1276
rect 23394 1316 23436 1344
rect 23094 204 23122 1248
rect 23394 204 23422 1316
rect 24050 1276 24078 1398
rect 24186 1344 24214 1398
rect 23872 1248 24078 1276
rect 24172 1316 24214 1344
rect 23872 204 23900 1248
rect 24172 204 24200 1316
rect 24828 1276 24856 1398
rect 24650 1248 24856 1276
rect 24650 204 24678 1248
<< metal3 >>
rect 319 5534 379 5594
rect 1875 5534 1935 5594
rect 3431 5534 3491 5594
rect 4987 5534 5047 5594
rect 6543 5534 6603 5594
rect 8099 5534 8159 5594
rect 9655 5534 9715 5594
rect 11211 5534 11271 5594
rect 12767 5534 12827 5594
rect 14323 5534 14383 5594
rect 15879 5534 15939 5594
rect 17435 5534 17495 5594
rect 18991 5534 19051 5594
rect 20547 5534 20607 5594
rect 22103 5534 22163 5594
rect 23659 5534 23719 5594
rect 319 4702 379 4762
rect 1875 4702 1935 4762
rect 3431 4702 3491 4762
rect 4987 4702 5047 4762
rect 6543 4702 6603 4762
rect 8099 4702 8159 4762
rect 9655 4702 9715 4762
rect 11211 4702 11271 4762
rect 12767 4702 12827 4762
rect 14323 4702 14383 4762
rect 15879 4702 15939 4762
rect 17435 4702 17495 4762
rect 18991 4702 19051 4762
rect 20547 4702 20607 4762
rect 22103 4702 22163 4762
rect 23659 4702 23719 4762
rect 4654 4386 4714 4446
rect 6210 4386 6270 4446
rect 7766 4386 7826 4446
rect 9322 4386 9382 4446
rect 10878 4386 10938 4446
rect 12434 4386 12494 4446
rect 13990 4386 14050 4446
rect 15546 4386 15606 4446
rect 17102 4386 17162 4446
rect 18658 4386 18718 4446
rect 20214 4386 20274 4446
rect 21770 4386 21830 4446
rect 23326 4386 23386 4446
rect 24882 4386 24942 4446
rect 26438 4386 26498 4446
rect 27994 4386 28054 4446
rect 29550 4386 29610 4446
rect 31106 4386 31166 4446
rect 32662 4386 32722 4446
rect 34218 4386 34278 4446
rect 35774 4386 35834 4446
rect 37330 4386 37390 4446
rect 38886 4386 38946 4446
rect 40442 4386 40502 4446
rect 41998 4386 42058 4446
rect 43554 4386 43614 4446
rect 45110 4386 45170 4446
rect 46666 4386 46726 4446
rect 48222 4386 48282 4446
rect 49778 4386 49838 4446
rect 51334 4386 51394 4446
rect 52890 4386 52950 4446
rect 4654 3440 4714 3500
rect 6210 3440 6270 3500
rect 7766 3440 7826 3500
rect 9322 3440 9382 3500
rect 10878 3440 10938 3500
rect 12434 3440 12494 3500
rect 13990 3440 14050 3500
rect 15546 3440 15606 3500
rect 17102 3440 17162 3500
rect 18658 3440 18718 3500
rect 20214 3440 20274 3500
rect 21770 3440 21830 3500
rect 23326 3440 23386 3500
rect 24882 3440 24942 3500
rect 26438 3440 26498 3500
rect 27994 3440 28054 3500
rect 29550 3440 29610 3500
rect 31106 3440 31166 3500
rect 32662 3440 32722 3500
rect 34218 3440 34278 3500
rect 35774 3440 35834 3500
rect 37330 3440 37390 3500
rect 38886 3440 38946 3500
rect 40442 3440 40502 3500
rect 41998 3440 42058 3500
rect 43554 3440 43614 3500
rect 45110 3440 45170 3500
rect 46666 3440 46726 3500
rect 48222 3440 48282 3500
rect 49778 3440 49838 3500
rect 51334 3440 51394 3500
rect 52890 3440 52950 3500
rect 748 2117 808 2177
rect 1526 2117 1586 2177
rect 2304 2117 2364 2177
rect 3082 2117 3142 2177
rect 3860 2117 3920 2177
rect 4638 2117 4698 2177
rect 5416 2117 5476 2177
rect 6194 2117 6254 2177
rect 6972 2117 7032 2177
rect 7750 2117 7810 2177
rect 8528 2117 8588 2177
rect 9306 2117 9366 2177
rect 10084 2117 10144 2177
rect 10862 2117 10922 2177
rect 11640 2117 11700 2177
rect 12418 2117 12478 2177
rect 13196 2117 13256 2177
rect 13974 2117 14034 2177
rect 14752 2117 14812 2177
rect 15530 2117 15590 2177
rect 16308 2117 16368 2177
rect 17086 2117 17146 2177
rect 17864 2117 17924 2177
rect 18642 2117 18702 2177
rect 19420 2117 19480 2177
rect 20198 2117 20258 2177
rect 20976 2117 21036 2177
rect 21754 2117 21814 2177
rect 22532 2117 22592 2177
rect 23310 2117 23370 2177
rect 24088 2117 24148 2177
rect 24866 2117 24926 2177
rect 163 284 223 344
rect 941 284 1001 344
rect 1719 284 1779 344
rect 2497 284 2557 344
rect 3275 284 3335 344
rect 4053 284 4113 344
rect 4831 284 4891 344
rect 5609 284 5669 344
rect 6387 284 6447 344
rect 7165 284 7225 344
rect 7943 284 8003 344
rect 8721 284 8781 344
rect 9499 284 9559 344
rect 10277 284 10337 344
rect 11055 284 11115 344
rect 11833 284 11893 344
rect 12611 284 12671 344
rect 13389 284 13449 344
rect 14167 284 14227 344
rect 14945 284 15005 344
rect 15723 284 15783 344
rect 16501 284 16561 344
rect 17279 284 17339 344
rect 18057 284 18117 344
rect 18835 284 18895 344
rect 19613 284 19673 344
rect 20391 284 20451 344
rect 21169 284 21229 344
rect 21947 284 22007 344
rect 22725 284 22785 344
rect 23503 284 23563 344
rect 24281 284 24341 344
rect 25059 284 25119 344
use column_mux_array_multiport  column_mux_array_multiport_0
timestamp 1643671299
transform 1 0 0 0 -1 3196
box 0 32 24926 1798
use write_driver_array  write_driver_array_0
timestamp 1643671299
transform 1 0 0 0 -1 5606
box 0 0 24038 952
use sense_amp_array  sense_amp_array_0
timestamp 1643671299
transform 1 0 0 0 -1 4450
box 4548 0 53056 1050
use precharge_array_multiport  precharge_array_multiport_0
timestamp 1643671299
transform 1 0 0 0 -1 1194
box 0 -24 25674 1004
<< labels >>
rlabel metal2 s 196 5306 250 5334 4 din0_0
rlabel metal2 s 1752 5306 1806 5334 4 din0_1
rlabel metal2 s 3308 5306 3362 5334 4 din0_2
rlabel metal2 s 4864 5306 4918 5334 4 din0_3
rlabel metal2 s 6420 5306 6474 5334 4 din0_4
rlabel metal2 s 7976 5306 8030 5334 4 din0_5
rlabel metal2 s 9532 5306 9586 5334 4 din0_6
rlabel metal2 s 11088 5306 11142 5334 4 din0_7
rlabel metal2 s 12644 5306 12698 5334 4 din0_8
rlabel metal2 s 14200 5306 14254 5334 4 din0_9
rlabel metal2 s 15756 5306 15810 5334 4 din0_10
rlabel metal2 s 17312 5306 17366 5334 4 din0_11
rlabel metal2 s 18868 5306 18922 5334 4 din0_12
rlabel metal2 s 20424 5306 20478 5334 4 din0_13
rlabel metal2 s 21980 5306 22034 5334 4 din0_14
rlabel metal2 s 23536 5306 23590 5334 4 din0_15
rlabel metal2 s 4750 4210 4778 4450 4 dout0_0
rlabel metal2 s 4764 4330 4764 4330 4 dout1_0
rlabel metal2 s 6306 4210 6334 4450 4 dout0_1
rlabel metal2 s 6320 4330 6320 4330 4 dout1_1
rlabel metal2 s 7862 4210 7890 4450 4 dout0_2
rlabel metal2 s 7876 4330 7876 4330 4 dout1_2
rlabel metal2 s 9418 4210 9446 4450 4 dout0_3
rlabel metal2 s 9432 4330 9432 4330 4 dout1_3
rlabel metal2 s 10974 4210 11002 4450 4 dout0_4
rlabel metal2 s 10988 4330 10988 4330 4 dout1_4
rlabel metal2 s 12530 4210 12558 4450 4 dout0_5
rlabel metal2 s 12544 4330 12544 4330 4 dout1_5
rlabel metal2 s 14086 4210 14114 4450 4 dout0_6
rlabel metal2 s 14100 4330 14100 4330 4 dout1_6
rlabel metal2 s 15642 4210 15670 4450 4 dout0_7
rlabel metal2 s 15656 4330 15656 4330 4 dout1_7
rlabel metal2 s 17198 4210 17226 4450 4 dout0_8
rlabel metal2 s 17212 4330 17212 4330 4 dout1_8
rlabel metal2 s 18754 4210 18782 4450 4 dout0_9
rlabel metal2 s 18768 4330 18768 4330 4 dout1_9
rlabel metal2 s 20310 4210 20338 4450 4 dout0_10
rlabel metal2 s 20324 4330 20324 4330 4 dout1_10
rlabel metal2 s 21866 4210 21894 4450 4 dout0_11
rlabel metal2 s 21880 4330 21880 4330 4 dout1_11
rlabel metal2 s 23422 4210 23450 4450 4 dout0_12
rlabel metal2 s 23436 4330 23436 4330 4 dout1_12
rlabel metal2 s 24978 4210 25006 4450 4 dout0_13
rlabel metal2 s 24992 4330 24992 4330 4 dout1_13
rlabel metal2 s 26534 4210 26562 4450 4 dout0_14
rlabel metal2 s 26548 4330 26548 4330 4 dout1_14
rlabel metal2 s 28090 4210 28118 4450 4 dout0_15
rlabel metal2 s 28104 4330 28104 4330 4 dout1_15
rlabel metal2 s 54 204 82 1194 4 rbl0_0
rlabel metal2 s 532 204 560 1194 4 rbl1_0
rlabel metal2 s 832 204 860 1194 4 rbl0_1
rlabel metal2 s 1310 204 1338 1194 4 rbl1_1
rlabel metal2 s 1610 204 1638 1194 4 rbl0_2
rlabel metal2 s 2088 204 2116 1194 4 rbl1_2
rlabel metal2 s 2388 204 2416 1194 4 rbl0_3
rlabel metal2 s 2866 204 2894 1194 4 rbl1_3
rlabel metal2 s 3166 204 3194 1194 4 rbl0_4
rlabel metal2 s 3644 204 3672 1194 4 rbl1_4
rlabel metal2 s 3944 204 3972 1194 4 rbl0_5
rlabel metal2 s 4422 204 4450 1194 4 rbl1_5
rlabel metal2 s 4722 204 4750 1194 4 rbl0_6
rlabel metal2 s 5200 204 5228 1194 4 rbl1_6
rlabel metal2 s 5500 204 5528 1194 4 rbl0_7
rlabel metal2 s 5978 204 6006 1194 4 rbl1_7
rlabel metal2 s 6278 204 6306 1194 4 rbl0_8
rlabel metal2 s 6756 204 6784 1194 4 rbl1_8
rlabel metal2 s 7056 204 7084 1194 4 rbl0_9
rlabel metal2 s 7534 204 7562 1194 4 rbl1_9
rlabel metal2 s 7834 204 7862 1194 4 rbl0_10
rlabel metal2 s 8312 204 8340 1194 4 rbl1_10
rlabel metal2 s 8612 204 8640 1194 4 rbl0_11
rlabel metal2 s 9090 204 9118 1194 4 rbl1_11
rlabel metal2 s 9390 204 9418 1194 4 rbl0_12
rlabel metal2 s 9868 204 9896 1194 4 rbl1_12
rlabel metal2 s 10168 204 10196 1194 4 rbl0_13
rlabel metal2 s 10646 204 10674 1194 4 rbl1_13
rlabel metal2 s 10946 204 10974 1194 4 rbl0_14
rlabel metal2 s 11424 204 11452 1194 4 rbl1_14
rlabel metal2 s 11724 204 11752 1194 4 rbl0_15
rlabel metal2 s 12202 204 12230 1194 4 rbl1_15
rlabel metal2 s 12502 204 12530 1194 4 rbl0_16
rlabel metal2 s 12980 204 13008 1194 4 rbl1_16
rlabel metal2 s 13280 204 13308 1194 4 rbl0_17
rlabel metal2 s 13758 204 13786 1194 4 rbl1_17
rlabel metal2 s 14058 204 14086 1194 4 rbl0_18
rlabel metal2 s 14536 204 14564 1194 4 rbl1_18
rlabel metal2 s 14836 204 14864 1194 4 rbl0_19
rlabel metal2 s 15314 204 15342 1194 4 rbl1_19
rlabel metal2 s 15614 204 15642 1194 4 rbl0_20
rlabel metal2 s 16092 204 16120 1194 4 rbl1_20
rlabel metal2 s 16392 204 16420 1194 4 rbl0_21
rlabel metal2 s 16870 204 16898 1194 4 rbl1_21
rlabel metal2 s 17170 204 17198 1194 4 rbl0_22
rlabel metal2 s 17648 204 17676 1194 4 rbl1_22
rlabel metal2 s 17948 204 17976 1194 4 rbl0_23
rlabel metal2 s 18426 204 18454 1194 4 rbl1_23
rlabel metal2 s 18726 204 18754 1194 4 rbl0_24
rlabel metal2 s 19204 204 19232 1194 4 rbl1_24
rlabel metal2 s 19504 204 19532 1194 4 rbl0_25
rlabel metal2 s 19982 204 20010 1194 4 rbl1_25
rlabel metal2 s 20282 204 20310 1194 4 rbl0_26
rlabel metal2 s 20760 204 20788 1194 4 rbl1_26
rlabel metal2 s 21060 204 21088 1194 4 rbl0_27
rlabel metal2 s 21538 204 21566 1194 4 rbl1_27
rlabel metal2 s 21838 204 21866 1194 4 rbl0_28
rlabel metal2 s 22316 204 22344 1194 4 rbl1_28
rlabel metal2 s 22616 204 22644 1194 4 rbl0_29
rlabel metal2 s 23094 204 23122 1194 4 rbl1_29
rlabel metal2 s 23394 204 23422 1194 4 rbl0_30
rlabel metal2 s 23872 204 23900 1194 4 rbl1_30
rlabel metal2 s 24172 204 24200 1194 4 rbl0_31
rlabel metal2 s 24650 204 24678 1194 4 rbl1_31
rlabel metal2 s 630 4654 658 5284 4 wbl0_0
rlabel metal2 s 2186 4654 2214 5284 4 wbl0_1
rlabel metal1 s 0 1170 25674 1198 4 p_en_bar
rlabel metal1 s 0 2994 24896 3022 4 sel_0
rlabel metal1 s 0 2936 24896 2964 4 sel_1
rlabel metal1 s 0 5222 24038 5250 4 w_en
rlabel metal3 s 31106 3440 31166 3500 4 vdd
rlabel metal3 s 7942 284 8002 344 4 vdd
rlabel metal3 s 26438 3440 26498 3500 4 vdd
rlabel metal3 s 18056 284 18116 344 4 vdd
rlabel metal3 s 4830 284 4890 344 4 vdd
rlabel metal3 s 7766 3440 7826 3500 4 vdd
rlabel metal3 s 49778 3440 49838 3500 4 vdd
rlabel metal3 s 8720 284 8780 344 4 vdd
rlabel metal3 s 32662 3440 32722 3500 4 vdd
rlabel metal3 s 40442 3440 40502 3500 4 vdd
rlabel metal3 s 45110 3440 45170 3500 4 vdd
rlabel metal3 s 5608 284 5668 344 4 vdd
rlabel metal3 s 17434 4702 17494 4762 4 vdd
rlabel metal3 s 7164 284 7224 344 4 vdd
rlabel metal3 s 29550 3440 29610 3500 4 vdd
rlabel metal3 s 23502 284 23562 344 4 vdd
rlabel metal3 s 17278 284 17338 344 4 vdd
rlabel metal3 s 10878 3440 10938 3500 4 vdd
rlabel metal3 s 24280 284 24340 344 4 vdd
rlabel metal3 s 21168 284 21228 344 4 vdd
rlabel metal3 s 22102 4702 22162 4762 4 vdd
rlabel metal3 s 20390 284 20450 344 4 vdd
rlabel metal3 s 13388 284 13448 344 4 vdd
rlabel metal3 s 52890 3440 52950 3500 4 vdd
rlabel metal3 s 20546 4702 20606 4762 4 vdd
rlabel metal3 s 22724 284 22784 344 4 vdd
rlabel metal3 s 48222 3440 48282 3500 4 vdd
rlabel metal3 s 17102 3440 17162 3500 4 vdd
rlabel metal3 s 14944 284 15004 344 4 vdd
rlabel metal3 s 23326 3440 23386 3500 4 vdd
rlabel metal3 s 38886 3440 38946 3500 4 vdd
rlabel metal3 s 19612 284 19672 344 4 vdd
rlabel metal3 s 14166 284 14226 344 4 vdd
rlabel metal3 s 11210 4702 11270 4762 4 vdd
rlabel metal3 s 9498 284 9558 344 4 vdd
rlabel metal3 s 318 4702 378 4762 4 vdd
rlabel metal3 s 9654 4702 9714 4762 4 vdd
rlabel metal3 s 12434 3440 12494 3500 4 vdd
rlabel metal3 s 13990 3440 14050 3500 4 vdd
rlabel metal3 s 12766 4702 12826 4762 4 vdd
rlabel metal3 s 2496 284 2556 344 4 vdd
rlabel metal3 s 8098 4702 8158 4762 4 vdd
rlabel metal3 s 11054 284 11114 344 4 vdd
rlabel metal3 s 3274 284 3334 344 4 vdd
rlabel metal3 s 14322 4702 14382 4762 4 vdd
rlabel metal3 s 11832 284 11892 344 4 vdd
rlabel metal3 s 6210 3440 6270 3500 4 vdd
rlabel metal3 s 940 284 1000 344 4 vdd
rlabel metal3 s 3430 4702 3490 4762 4 vdd
rlabel metal3 s 43554 3440 43614 3500 4 vdd
rlabel metal3 s 18990 4702 19050 4762 4 vdd
rlabel metal3 s 9322 3440 9382 3500 4 vdd
rlabel metal3 s 15722 284 15782 344 4 vdd
rlabel metal3 s 4052 284 4112 344 4 vdd
rlabel metal3 s 6386 284 6446 344 4 vdd
rlabel metal3 s 1874 4702 1934 4762 4 vdd
rlabel metal3 s 6542 4702 6602 4762 4 vdd
rlabel metal3 s 15878 4702 15938 4762 4 vdd
rlabel metal3 s 21946 284 22006 344 4 vdd
rlabel metal3 s 41998 3440 42058 3500 4 vdd
rlabel metal3 s 23658 4702 23718 4762 4 vdd
rlabel metal3 s 51334 3440 51394 3500 4 vdd
rlabel metal3 s 21770 3440 21830 3500 4 vdd
rlabel metal3 s 37330 3440 37390 3500 4 vdd
rlabel metal3 s 46666 3440 46726 3500 4 vdd
rlabel metal3 s 15546 3440 15606 3500 4 vdd
rlabel metal3 s 20214 3440 20274 3500 4 vdd
rlabel metal3 s 24882 3440 24942 3500 4 vdd
rlabel metal3 s 18658 3440 18718 3500 4 vdd
rlabel metal3 s 162 284 222 344 4 vdd
rlabel metal3 s 27994 3440 28054 3500 4 vdd
rlabel metal3 s 12610 284 12670 344 4 vdd
rlabel metal3 s 4986 4702 5046 4762 4 vdd
rlabel metal3 s 4654 3440 4714 3500 4 vdd
rlabel metal3 s 34218 3440 34278 3500 4 vdd
rlabel metal3 s 10276 284 10336 344 4 vdd
rlabel metal3 s 35774 3440 35834 3500 4 vdd
rlabel metal3 s 25058 284 25118 344 4 vdd
rlabel metal3 s 16500 284 16560 344 4 vdd
rlabel metal3 s 18834 284 18894 344 4 vdd
rlabel metal3 s 1718 284 1778 344 4 vdd
rlabel metal3 s 46666 4386 46726 4446 4 gnd
rlabel metal3 s 18990 5534 19050 5594 4 gnd
rlabel metal3 s 8098 5534 8158 5594 4 gnd
rlabel metal3 s 7750 2116 7810 2176 4 gnd
rlabel metal3 s 6210 4386 6270 4446 4 gnd
rlabel metal3 s 20214 4386 20274 4446 4 gnd
rlabel metal3 s 32662 4386 32722 4446 4 gnd
rlabel metal3 s 37330 4386 37390 4446 4 gnd
rlabel metal3 s 13196 2116 13256 2176 4 gnd
rlabel metal3 s 21754 2116 21814 2176 4 gnd
rlabel metal3 s 21770 4386 21830 4446 4 gnd
rlabel metal3 s 49778 4386 49838 4446 4 gnd
rlabel metal3 s 748 2116 808 2176 4 gnd
rlabel metal3 s 48222 4386 48282 4446 4 gnd
rlabel metal3 s 14322 5534 14382 5594 4 gnd
rlabel metal3 s 38886 4386 38946 4446 4 gnd
rlabel metal3 s 12766 5534 12826 5594 4 gnd
rlabel metal3 s 29550 4386 29610 4446 4 gnd
rlabel metal3 s 41998 4386 42058 4446 4 gnd
rlabel metal3 s 10862 2116 10922 2176 4 gnd
rlabel metal3 s 20976 2116 21036 2176 4 gnd
rlabel metal3 s 17086 2116 17146 2176 4 gnd
rlabel metal3 s 20546 5534 20606 5594 4 gnd
rlabel metal3 s 40442 4386 40502 4446 4 gnd
rlabel metal3 s 17102 4386 17162 4446 4 gnd
rlabel metal3 s 18642 2116 18702 2176 4 gnd
rlabel metal3 s 12434 4386 12494 4446 4 gnd
rlabel metal3 s 4654 4386 4714 4446 4 gnd
rlabel metal3 s 23326 4386 23386 4446 4 gnd
rlabel metal3 s 24866 2116 24926 2176 4 gnd
rlabel metal3 s 35774 4386 35834 4446 4 gnd
rlabel metal3 s 9306 2116 9366 2176 4 gnd
rlabel metal3 s 7766 4386 7826 4446 4 gnd
rlabel metal3 s 1526 2116 1586 2176 4 gnd
rlabel metal3 s 11640 2116 11700 2176 4 gnd
rlabel metal3 s 20198 2116 20258 2176 4 gnd
rlabel metal3 s 24088 2116 24148 2176 4 gnd
rlabel metal3 s 9654 5534 9714 5594 4 gnd
rlabel metal3 s 34218 4386 34278 4446 4 gnd
rlabel metal3 s 16308 2116 16368 2176 4 gnd
rlabel metal3 s 17434 5534 17494 5594 4 gnd
rlabel metal3 s 45110 4386 45170 4446 4 gnd
rlabel metal3 s 6194 2116 6254 2176 4 gnd
rlabel metal3 s 13990 4386 14050 4446 4 gnd
rlabel metal3 s 2304 2116 2364 2176 4 gnd
rlabel metal3 s 26438 4386 26498 4446 4 gnd
rlabel metal3 s 3430 5534 3490 5594 4 gnd
rlabel metal3 s 24882 4386 24942 4446 4 gnd
rlabel metal3 s 9322 4386 9382 4446 4 gnd
rlabel metal3 s 15530 2116 15590 2176 4 gnd
rlabel metal3 s 1874 5534 1934 5594 4 gnd
rlabel metal3 s 23658 5534 23718 5594 4 gnd
rlabel metal3 s 23310 2116 23370 2176 4 gnd
rlabel metal3 s 13974 2116 14034 2176 4 gnd
rlabel metal3 s 5416 2116 5476 2176 4 gnd
rlabel metal3 s 3082 2116 3142 2176 4 gnd
rlabel metal3 s 18658 4386 18718 4446 4 gnd
rlabel metal3 s 12418 2116 12478 2176 4 gnd
rlabel metal3 s 43554 4386 43614 4446 4 gnd
rlabel metal3 s 10878 4386 10938 4446 4 gnd
rlabel metal3 s 19420 2116 19480 2176 4 gnd
rlabel metal3 s 22532 2116 22592 2176 4 gnd
rlabel metal3 s 3860 2116 3920 2176 4 gnd
rlabel metal3 s 14752 2116 14812 2176 4 gnd
rlabel metal3 s 51334 4386 51394 4446 4 gnd
rlabel metal3 s 27994 4386 28054 4446 4 gnd
rlabel metal3 s 15546 4386 15606 4446 4 gnd
rlabel metal3 s 8528 2116 8588 2176 4 gnd
rlabel metal3 s 6972 2116 7032 2176 4 gnd
rlabel metal3 s 10084 2116 10144 2176 4 gnd
rlabel metal3 s 11210 5534 11270 5594 4 gnd
rlabel metal3 s 52890 4386 52950 4446 4 gnd
rlabel metal3 s 6542 5534 6602 5594 4 gnd
rlabel metal3 s 31106 4386 31166 4446 4 gnd
rlabel metal3 s 22102 5534 22162 5594 4 gnd
rlabel metal3 s 318 5534 378 5594 4 gnd
rlabel metal3 s 15878 5534 15938 5594 4 gnd
rlabel metal3 s 4638 2116 4698 2176 4 gnd
rlabel metal3 s 17864 2116 17924 2176 4 gnd
rlabel metal3 s 4986 5534 5046 5594 4 gnd
<< properties >>
string FIXED_BBOX 0 0 53056 5606
string GDS_FILE sram_0rw2r1w_16_32_sky130A.gds
string GDS_END 749954
string GDS_START 676842
<< end >>
