magic
tech sky130A
magscale 1 2
timestamp 1643593061
<< checkpaint >>
rect -1319 -1316 2333 1594
<< nwell >>
rect -54 224 1068 334
rect -59 56 1073 224
rect -54 -54 1068 56
<< scpmos >>
rect 60 0 90 280
rect 168 0 198 280
rect 276 0 306 280
rect 384 0 414 280
rect 492 0 522 280
rect 600 0 630 280
rect 708 0 738 280
rect 816 0 846 280
rect 924 0 954 280
<< pdiff >>
rect 0 157 60 280
rect 0 123 8 157
rect 42 123 60 157
rect 0 0 60 123
rect 90 157 168 280
rect 90 123 112 157
rect 146 123 168 157
rect 90 0 168 123
rect 198 157 276 280
rect 198 123 220 157
rect 254 123 276 157
rect 198 0 276 123
rect 306 157 384 280
rect 306 123 328 157
rect 362 123 384 157
rect 306 0 384 123
rect 414 157 492 280
rect 414 123 436 157
rect 470 123 492 157
rect 414 0 492 123
rect 522 157 600 280
rect 522 123 544 157
rect 578 123 600 157
rect 522 0 600 123
rect 630 157 708 280
rect 630 123 652 157
rect 686 123 708 157
rect 630 0 708 123
rect 738 157 816 280
rect 738 123 760 157
rect 794 123 816 157
rect 738 0 816 123
rect 846 157 924 280
rect 846 123 868 157
rect 902 123 924 157
rect 846 0 924 123
rect 954 157 1014 280
rect 954 123 972 157
rect 1006 123 1014 157
rect 954 0 1014 123
<< pdiffc >>
rect 8 123 42 157
rect 112 123 146 157
rect 220 123 254 157
rect 328 123 362 157
rect 436 123 470 157
rect 544 123 578 157
rect 652 123 686 157
rect 760 123 794 157
rect 868 123 902 157
rect 972 123 1006 157
<< poly >>
rect 60 280 90 306
rect 168 280 198 306
rect 276 280 306 306
rect 384 280 414 306
rect 492 280 522 306
rect 600 280 630 306
rect 708 280 738 306
rect 816 280 846 306
rect 924 280 954 306
rect 60 -26 90 0
rect 168 -26 198 0
rect 276 -26 306 0
rect 384 -26 414 0
rect 492 -26 522 0
rect 600 -26 630 0
rect 708 -26 738 0
rect 816 -26 846 0
rect 924 -26 954 0
rect 60 -56 954 -26
<< locali >>
rect 8 157 42 173
rect 8 107 42 123
rect 112 157 146 173
rect 112 73 146 123
rect 220 157 254 173
rect 220 107 254 123
rect 328 157 362 173
rect 328 73 362 123
rect 436 157 470 173
rect 436 107 470 123
rect 544 157 578 173
rect 544 73 578 123
rect 652 157 686 173
rect 652 107 686 123
rect 760 157 794 173
rect 760 73 794 123
rect 868 157 902 173
rect 868 107 902 123
rect 972 157 1006 173
rect 972 73 1006 123
rect 112 39 1006 73
use contact_9  contact_9_0
timestamp 1643593061
transform 1 0 964 0 1 99
box 0 0 2 2
use contact_9  contact_9_1
timestamp 1643593061
transform 1 0 860 0 1 99
box 0 0 2 2
use contact_9  contact_9_2
timestamp 1643593061
transform 1 0 752 0 1 99
box 0 0 2 2
use contact_9  contact_9_3
timestamp 1643593061
transform 1 0 644 0 1 99
box 0 0 2 2
use contact_9  contact_9_4
timestamp 1643593061
transform 1 0 536 0 1 99
box 0 0 2 2
use contact_9  contact_9_5
timestamp 1643593061
transform 1 0 428 0 1 99
box 0 0 2 2
use contact_9  contact_9_6
timestamp 1643593061
transform 1 0 320 0 1 99
box 0 0 2 2
use contact_9  contact_9_7
timestamp 1643593061
transform 1 0 212 0 1 99
box 0 0 2 2
use contact_9  contact_9_8
timestamp 1643593061
transform 1 0 104 0 1 99
box 0 0 2 2
use contact_9  contact_9_9
timestamp 1643593061
transform 1 0 0 0 1 99
box 0 0 2 2
<< labels >>
rlabel mvvaractor s 507 -41 507 -41 4 G
rlabel locali s 885 140 885 140 4 S
rlabel locali s 669 140 669 140 4 S
rlabel locali s 453 140 453 140 4 S
rlabel locali s 237 140 237 140 4 S
rlabel locali s 25 140 25 140 4 S
rlabel locali s 559 56 559 56 4 D
<< properties >>
string FIXED_BBOX -54 -56 1068 56
string GDS_FILE sram_0rw2r1w_2_16_sky130A.gds
string GDS_END 564646
string GDS_START 562186
<< end >>
