magic
tech sky130A
magscale 1 2
timestamp 1644949024
<< checkpaint >>
rect -1260 -1260 25368 37452
<< metal2 >>
rect 8993 14146 9049 14155
rect 8993 14081 9049 14090
rect 10073 14150 10129 14159
rect 10073 14085 10129 14094
rect 8993 12962 9049 12971
rect 8993 12897 9049 12906
rect 10073 12958 10129 12967
rect 10073 12893 10129 12902
rect 8993 12470 9049 12479
rect 8993 12405 9049 12414
rect 10073 12474 10129 12483
rect 10073 12409 10129 12418
rect 8993 11286 9049 11295
rect 8993 11221 9049 11230
rect 10073 11282 10129 11291
rect 10073 11217 10129 11226
rect 8993 10794 9049 10803
rect 8993 10729 9049 10738
rect 10073 10798 10129 10807
rect 10073 10733 10129 10742
rect 8702 9672 8758 9681
rect 8702 9607 8758 9616
rect 8993 9610 9049 9619
rect 10482 9615 10510 21484
rect 10566 10807 10594 21484
rect 10650 11291 10678 21484
rect 10734 12483 10762 21484
rect 10818 12967 10846 21484
rect 10902 14159 10930 21484
rect 10888 14150 10944 14159
rect 10888 14085 10944 14094
rect 10804 12958 10860 12967
rect 10804 12893 10860 12902
rect 10720 12474 10776 12483
rect 10720 12409 10776 12418
rect 10636 11282 10692 11291
rect 10636 11217 10692 11226
rect 10552 10798 10608 10807
rect 10552 10733 10608 10742
rect 2919 4636 2975 4645
rect 2919 4571 2975 4580
rect 6441 4421 6497 4430
rect 8716 4401 8744 9607
rect 8993 9545 9049 9554
rect 10073 9606 10129 9615
rect 10073 9541 10129 9550
rect 10468 9606 10524 9615
rect 10468 9541 10524 9550
rect 15994 8704 16022 33776
rect 10268 8695 10324 8704
rect 10268 8630 10324 8639
rect 15980 8695 16036 8704
rect 15980 8630 16036 8639
rect 10268 7773 10324 7782
rect 10268 7708 10324 7717
rect 17116 7032 17144 8762
rect 20896 7773 20952 7782
rect 20896 7708 20952 7717
rect 17676 7620 17732 7629
rect 17676 7555 17732 7564
rect 17948 7620 18004 7629
rect 17948 7555 18004 7564
rect 18454 7620 18510 7629
rect 18454 7555 18510 7564
rect 18726 7620 18782 7629
rect 18726 7555 18782 7564
rect 10268 7023 10324 7032
rect 10268 6958 10324 6967
rect 17102 7023 17158 7032
rect 17102 6958 17158 6967
rect 20910 4938 20938 7708
rect 8716 4387 9096 4401
rect 6441 4356 6497 4365
rect 8664 4373 9096 4387
rect 2919 3452 2975 3461
rect 2919 3387 2975 3396
rect 8664 2986 8796 4373
rect 8664 2958 8702 2986
rect 8758 2958 8796 2986
rect 8702 2921 8758 2930
rect 11957 2924 12013 2933
rect 11957 2859 12013 2868
rect 13439 2924 13495 2933
rect 13439 2859 13495 2868
rect 14921 2924 14977 2933
rect 14921 2859 14977 2868
rect 16403 2924 16459 2933
rect 16403 2859 16459 2868
<< via2 >>
rect 8993 14090 9049 14146
rect 10073 14094 10129 14150
rect 8993 12906 9049 12962
rect 10073 12902 10129 12958
rect 8993 12414 9049 12470
rect 10073 12418 10129 12474
rect 8993 11230 9049 11286
rect 10073 11226 10129 11282
rect 8993 10738 9049 10794
rect 10073 10742 10129 10798
rect 8702 9616 8758 9672
rect 10888 14094 10944 14150
rect 10804 12902 10860 12958
rect 10720 12418 10776 12474
rect 10636 11226 10692 11282
rect 10552 10742 10608 10798
rect 2919 4580 2975 4636
rect 6441 4365 6497 4421
rect 8993 9554 9049 9610
rect 10073 9550 10129 9606
rect 10468 9550 10524 9606
rect 10268 8639 10324 8695
rect 15980 8639 16036 8695
rect 10268 7717 10324 7773
rect 20896 7717 20952 7773
rect 17676 7564 17732 7620
rect 17948 7564 18004 7620
rect 18454 7564 18510 7620
rect 18726 7564 18782 7620
rect 10268 6967 10324 7023
rect 17102 6967 17158 7023
rect 2919 3396 2975 3452
rect 8702 2930 8758 2986
rect 11957 2868 12013 2924
rect 13439 2868 13495 2924
rect 14921 2868 14977 2924
rect 16403 2868 16459 2924
<< metal3 >>
rect 424 36148 23684 36192
rect 424 36084 468 36148
rect 532 36084 680 36148
rect 744 36084 892 36148
rect 956 36084 23152 36148
rect 23216 36084 23364 36148
rect 23428 36084 23576 36148
rect 23640 36084 23684 36148
rect 424 35936 23684 36084
rect 424 35872 468 35936
rect 532 35872 680 35936
rect 744 35872 892 35936
rect 956 35872 23152 35936
rect 23216 35872 23364 35936
rect 23428 35872 23576 35936
rect 23640 35872 23684 35936
rect 424 35724 23684 35872
rect 424 35660 468 35724
rect 532 35660 680 35724
rect 744 35660 892 35724
rect 956 35660 12340 35724
rect 12404 35660 17004 35724
rect 17068 35660 23152 35724
rect 23216 35660 23364 35724
rect 23428 35660 23576 35724
rect 23640 35660 23684 35724
rect 424 35616 23684 35660
rect 1484 35088 22624 35132
rect 1484 35024 1528 35088
rect 1592 35024 1740 35088
rect 1804 35024 1952 35088
rect 2016 35024 22092 35088
rect 22156 35024 22304 35088
rect 22368 35024 22516 35088
rect 22580 35024 22624 35088
rect 1484 34876 22624 35024
rect 1484 34812 1528 34876
rect 1592 34812 1740 34876
rect 1804 34812 1952 34876
rect 2016 34812 22092 34876
rect 22156 34812 22304 34876
rect 22368 34812 22516 34876
rect 22580 34812 22624 34876
rect 1484 34664 22624 34812
rect 1484 34600 1528 34664
rect 1592 34600 1740 34664
rect 1804 34600 1952 34664
rect 2016 34600 11492 34664
rect 11556 34600 15520 34664
rect 15584 34600 22092 34664
rect 22156 34600 22304 34664
rect 22368 34600 22516 34664
rect 22580 34600 22624 34664
rect 1484 34556 22624 34600
rect 11236 33816 12448 33860
rect 11236 33752 12128 33816
rect 12192 33752 12340 33816
rect 12404 33752 12448 33816
rect 11236 33708 12448 33752
rect 15476 33816 17324 33860
rect 15476 33752 17004 33816
rect 17068 33752 17216 33816
rect 17280 33752 17324 33816
rect 15476 33708 17324 33752
rect 11236 32332 12448 32376
rect 11236 32268 11492 32332
rect 11556 32268 12448 32332
rect 11236 32224 12448 32268
rect 11256 32223 11600 32224
rect 11448 32012 11600 32223
rect 12084 32120 12448 32224
rect 12084 32056 12340 32120
rect 12404 32056 12448 32120
rect 12084 32012 12448 32056
rect 15476 32332 15840 32376
rect 15476 32268 15520 32332
rect 15584 32268 15840 32332
rect 15476 32164 15840 32268
rect 16960 32164 17324 32376
rect 15476 32120 17324 32164
rect 15476 32056 15732 32120
rect 15796 32056 17324 32120
rect 15476 32012 17324 32056
rect 11236 30848 12448 30892
rect 11236 30784 12128 30848
rect 12192 30784 12448 30848
rect 11236 30740 12448 30784
rect 11236 30680 11600 30740
rect 11236 30636 12024 30680
rect 11236 30572 11916 30636
rect 11980 30572 12024 30636
rect 11236 30528 12024 30572
rect 12084 30528 12448 30740
rect 15476 30848 17324 30892
rect 15476 30784 17216 30848
rect 17280 30784 17324 30848
rect 15476 30740 17324 30784
rect 15476 30636 15840 30740
rect 15476 30572 15520 30636
rect 15584 30572 15840 30636
rect 15476 30528 15840 30572
rect 16960 30528 17324 30740
rect 11448 29217 11600 29408
rect 11256 29196 11600 29217
rect 12084 29364 12448 29408
rect 12084 29300 12340 29364
rect 12404 29300 12448 29364
rect 12084 29196 12448 29300
rect 11236 29044 12448 29196
rect 15476 29364 15840 29408
rect 15476 29300 15732 29364
rect 15796 29300 15840 29364
rect 15476 29196 15840 29300
rect 16960 29196 17324 29408
rect 15476 29044 17324 29196
rect 11448 27772 12236 27924
rect 11448 27712 11600 27772
rect 12084 27712 12236 27772
rect 11236 27668 11812 27712
rect 11948 27668 12448 27712
rect 11236 27604 11704 27668
rect 11768 27604 11812 27668
rect 11872 27604 11916 27668
rect 11980 27604 12448 27668
rect 11236 27560 11812 27604
rect 11948 27560 12448 27604
rect 15476 27668 17324 27712
rect 15476 27604 15520 27668
rect 15584 27604 17004 27668
rect 17068 27604 17324 27668
rect 15476 27560 17324 27604
rect 15476 26076 17324 26228
rect 15476 25972 15840 26076
rect 15476 25908 15520 25972
rect 15584 25908 15840 25972
rect 15476 25864 15840 25908
rect 16960 25864 17324 26076
rect 11236 24532 11600 24744
rect 11736 24700 12448 24744
rect 11660 24636 11704 24700
rect 11768 24636 12448 24700
rect 11736 24592 12448 24636
rect 12084 24532 12448 24592
rect 11236 24488 12448 24532
rect 11236 24424 12128 24488
rect 12192 24424 12448 24488
rect 11236 24380 12448 24424
rect 15476 24532 15840 24744
rect 16960 24700 17324 24744
rect 16960 24636 17004 24700
rect 17068 24636 17324 24700
rect 16960 24532 17324 24636
rect 15476 24488 17324 24532
rect 15476 24424 17004 24488
rect 17068 24424 17324 24488
rect 15476 24380 17324 24424
rect 11448 23108 12448 23260
rect 11448 23061 11600 23108
rect 11256 23048 11600 23061
rect 12084 23048 12448 23108
rect 11236 22896 11600 23048
rect 11948 23004 12660 23048
rect 11872 22940 11916 23004
rect 11980 22940 12660 23004
rect 11948 22896 12660 22940
rect 12508 22836 12660 22896
rect 15476 23004 17324 23048
rect 15476 22940 15520 23004
rect 15584 22940 15732 23004
rect 15796 22940 17324 23004
rect 15476 22896 17324 22940
rect 15476 22836 15628 22896
rect 12508 22684 15628 22836
rect 11448 21732 12236 21776
rect 11448 21668 12128 21732
rect 12192 21668 12236 21732
rect 11448 21624 12236 21668
rect 11448 21564 11600 21624
rect 11236 21520 11812 21564
rect 11236 21456 11704 21520
rect 11768 21456 11812 21520
rect 11236 21412 11812 21456
rect 12084 21412 12448 21564
rect 15476 21520 17324 21564
rect 15476 21456 17004 21520
rect 17068 21456 17216 21520
rect 17280 21456 17324 21520
rect 15476 21412 17324 21456
rect 11448 21352 11600 21412
rect 12084 21352 12236 21412
rect 11448 21200 12236 21352
rect 11236 20036 12024 20080
rect 11236 19972 11916 20036
rect 11980 19972 12024 20036
rect 11236 19928 12024 19972
rect 11256 19907 11600 19928
rect 11448 19868 11600 19907
rect 12084 19868 12448 20080
rect 11448 19716 12448 19868
rect 15476 20036 15840 20080
rect 15476 19972 15732 20036
rect 15796 19972 15840 20036
rect 15476 19868 15840 19972
rect 16960 19868 17324 20080
rect 15476 19824 17324 19868
rect 15476 19760 15732 19824
rect 15796 19760 17324 19824
rect 15476 19716 17324 19760
rect 11236 18444 12448 18596
rect 11236 18340 11600 18444
rect 12084 18384 12448 18444
rect 11736 18340 12448 18384
rect 11236 18276 11280 18340
rect 11344 18276 11600 18340
rect 11660 18276 11704 18340
rect 11768 18276 12448 18340
rect 11236 18232 11600 18276
rect 11736 18232 12448 18276
rect 15476 18384 15840 18596
rect 16960 18552 17324 18596
rect 16960 18488 17216 18552
rect 17280 18488 17324 18552
rect 16960 18384 17324 18488
rect 15476 18232 17324 18384
rect 15476 16856 17324 16900
rect 15476 16792 15520 16856
rect 15584 16792 15732 16856
rect 15796 16792 17324 16856
rect 15476 16748 17324 16792
rect 9328 16220 11388 16264
rect 9328 16156 11280 16220
rect 11344 16156 11388 16220
rect 9328 16112 11388 16156
rect 9328 16008 9692 16112
rect 9328 15944 9584 16008
rect 9648 15944 9692 16008
rect 9328 15900 9692 15944
rect 9328 15160 9692 15416
rect 11236 15372 12448 15416
rect 11236 15308 11280 15372
rect 11344 15308 12448 15372
rect 11236 15264 12448 15308
rect 15476 15372 17324 15416
rect 15476 15308 17004 15372
rect 17068 15308 17324 15372
rect 15476 15264 17324 15308
rect 9328 15096 9372 15160
rect 9436 15096 9692 15160
rect 9328 15052 9692 15096
rect 9328 14524 11388 14568
rect 9328 14460 9584 14524
rect 9648 14460 11280 14524
rect 11344 14460 11388 14524
rect 9328 14416 11388 14460
rect 8904 14146 9268 14356
rect 9489 14327 9692 14416
rect 9540 14312 9692 14327
rect 9540 14248 9584 14312
rect 9648 14248 9692 14312
rect 9540 14204 9692 14248
rect 8904 14144 8993 14146
rect 0 14090 8993 14144
rect 9049 14090 9268 14146
rect 0 13992 9268 14090
rect 10035 14152 10167 14155
rect 10850 14152 10982 14155
rect 10035 14150 10982 14152
rect 10035 14094 10073 14150
rect 10129 14094 10888 14150
rect 10944 14094 10982 14150
rect 10035 14092 10982 14094
rect 10035 14089 10167 14092
rect 10850 14089 10982 14092
rect 11024 13780 12448 13932
rect 11024 13720 11176 13780
rect 11256 13751 11600 13780
rect 9328 13676 11176 13720
rect 9328 13612 9372 13676
rect 9436 13612 11176 13676
rect 9328 13568 11176 13612
rect 11448 13568 11600 13751
rect 12084 13568 12448 13780
rect 15476 13888 15840 13932
rect 15476 13824 15520 13888
rect 15584 13824 15840 13888
rect 15476 13720 15840 13824
rect 16960 13720 17324 13932
rect 15476 13676 17324 13720
rect 15476 13612 17216 13676
rect 17280 13612 17324 13676
rect 15476 13568 17324 13612
rect 9328 13464 9692 13568
rect 9328 13400 9372 13464
rect 9436 13400 9692 13464
rect 9328 13356 9692 13400
rect 8904 12962 9268 13084
rect 8904 12906 8993 12962
rect 9049 12906 9268 12962
rect 8904 12872 9268 12906
rect 10035 12960 10167 12963
rect 10766 12960 10898 12963
rect 10035 12958 10898 12960
rect 10035 12902 10073 12958
rect 10129 12902 10804 12958
rect 10860 12902 10898 12958
rect 10035 12900 10898 12902
rect 10035 12897 10167 12900
rect 10766 12897 10898 12900
rect 0 12720 9268 12872
rect 9540 12828 9692 12872
rect 9540 12764 9584 12828
rect 9648 12764 9692 12828
rect 9540 12725 9692 12764
rect 9489 12660 9692 12725
rect 8904 12470 9268 12660
rect 9489 12651 9904 12660
rect 9540 12616 9904 12651
rect 9540 12552 9584 12616
rect 9648 12552 9796 12616
rect 9860 12552 9904 12616
rect 9540 12508 9904 12552
rect 8904 12448 8993 12470
rect 0 12414 8993 12448
rect 9049 12414 9268 12470
rect 0 12296 9268 12414
rect 10035 12476 10167 12479
rect 10682 12476 10814 12479
rect 10035 12474 10814 12476
rect 10035 12418 10073 12474
rect 10129 12418 10720 12474
rect 10776 12418 10814 12474
rect 10035 12416 10814 12418
rect 10035 12413 10167 12416
rect 10682 12413 10814 12416
rect 11236 12236 11600 12448
rect 12084 12236 12448 12448
rect 9828 12192 12448 12236
rect 9752 12128 9796 12192
rect 9860 12128 12448 12192
rect 9828 12084 12448 12128
rect 15476 12404 17324 12448
rect 15476 12340 17004 12404
rect 17068 12340 17324 12404
rect 15476 12296 17324 12340
rect 15476 12192 15840 12296
rect 15476 12128 15520 12192
rect 15584 12128 15840 12192
rect 15476 12084 15840 12128
rect 16960 12084 17324 12296
rect 9328 11980 9692 12024
rect 9328 11916 9372 11980
rect 9436 11916 9692 11980
rect 9328 11768 9692 11916
rect 9328 11704 9372 11768
rect 9436 11704 9692 11768
rect 9328 11660 9692 11704
rect 8904 11286 9268 11388
rect 8904 11230 8993 11286
rect 9049 11230 9268 11286
rect 8904 11176 9268 11230
rect 10035 11284 10167 11287
rect 10598 11284 10730 11287
rect 10035 11282 10730 11284
rect 10035 11226 10073 11282
rect 10129 11226 10636 11282
rect 10692 11226 10730 11282
rect 10035 11224 10730 11226
rect 10035 11221 10167 11224
rect 10598 11221 10730 11224
rect 0 11024 9268 11176
rect 9540 11132 9692 11176
rect 9540 11068 9584 11132
rect 9648 11068 9692 11132
rect 9540 11049 9692 11068
rect 9489 10975 9692 11049
rect 8904 10794 9268 10964
rect 9540 10920 9692 10975
rect 9540 10856 9584 10920
rect 9648 10856 9692 10920
rect 9540 10812 9692 10856
rect 8904 10752 8993 10794
rect 0 10738 8993 10752
rect 9049 10738 9268 10794
rect 0 10600 9268 10738
rect 10035 10800 10167 10803
rect 10514 10800 10646 10803
rect 10035 10798 10646 10800
rect 10035 10742 10073 10798
rect 10129 10742 10552 10798
rect 10608 10742 10646 10798
rect 10035 10740 10646 10742
rect 10035 10737 10167 10740
rect 10514 10737 10646 10740
rect 11236 10708 12660 10752
rect 11236 10644 11280 10708
rect 11344 10644 12660 10708
rect 11236 10600 12660 10644
rect 12508 10540 12660 10600
rect 15476 10708 17748 10752
rect 15476 10644 17216 10708
rect 17280 10644 17640 10708
rect 17704 10644 17748 10708
rect 15476 10600 17748 10644
rect 15476 10540 15628 10600
rect 12508 10388 15628 10540
rect 9328 10284 11388 10328
rect 9328 10220 9372 10284
rect 9436 10220 11280 10284
rect 11344 10220 11388 10284
rect 9328 10176 11388 10220
rect 9328 9964 9692 10176
rect 0 9752 9056 9904
rect 8730 9677 8814 9681
rect 8664 9672 8814 9677
rect 8664 9616 8702 9672
rect 8758 9616 8814 9672
rect 8664 9611 8814 9616
rect 8730 9607 8814 9611
rect 8904 9619 9056 9752
rect 9116 9619 9268 9692
rect 8904 9610 9268 9619
rect 8904 9554 8993 9610
rect 9049 9554 9268 9610
rect 8904 9545 9268 9554
rect 10035 9608 10167 9611
rect 10430 9608 10562 9611
rect 10035 9606 10562 9608
rect 10035 9550 10073 9606
rect 10129 9550 10468 9606
rect 10524 9550 10562 9606
rect 10035 9548 10562 9550
rect 10035 9545 10167 9548
rect 10430 9545 10562 9548
rect 8904 9540 9056 9545
rect 9116 9540 9268 9545
rect 9540 9436 9692 9480
rect 9540 9373 9584 9436
rect 9489 9372 9584 9373
rect 9648 9372 9692 9436
rect 9489 9268 9692 9372
rect 9328 9116 12448 9268
rect 15476 9224 17748 9268
rect 15476 9160 15520 9224
rect 15584 9160 17748 9224
rect 15476 9116 17748 9160
rect 17596 9056 17748 9116
rect 17596 8844 17960 9056
rect 18096 9012 18808 9056
rect 18020 8948 18064 9012
rect 18128 8948 18808 9012
rect 18096 8904 18808 8948
rect 18444 8844 18808 8904
rect 19292 8904 20292 9056
rect 19292 8844 19656 8904
rect 10230 8697 10362 8700
rect 15942 8697 16074 8700
rect 10230 8695 16074 8697
rect 10230 8639 10268 8695
rect 10324 8639 15980 8695
rect 16036 8639 16074 8695
rect 17596 8692 19656 8844
rect 20140 8692 20292 8904
rect 10230 8637 16074 8639
rect 10230 8634 10362 8637
rect 15942 8634 16074 8637
rect 17596 8164 17960 8208
rect 17596 8100 17640 8164
rect 17704 8100 17960 8164
rect 17596 7996 17960 8100
rect 18444 8056 19656 8208
rect 18444 7996 18808 8056
rect 17596 7952 18808 7996
rect 17596 7888 18488 7952
rect 18552 7888 18808 7952
rect 17596 7844 18808 7888
rect 19292 7996 19656 8056
rect 20140 7996 20292 8208
rect 19292 7844 20292 7996
rect 20352 7952 23260 7996
rect 20352 7888 23152 7952
rect 23216 7888 23260 7952
rect 20352 7844 23260 7888
rect 10230 7775 10362 7778
rect 17384 7775 17536 7784
rect 17596 7775 17960 7784
rect 18020 7775 18384 7784
rect 18444 7775 18596 7784
rect 18656 7775 18808 7784
rect 19080 7775 19232 7784
rect 19292 7775 19444 7784
rect 19504 7775 19868 7784
rect 19928 7775 20292 7784
rect 20352 7775 20504 7844
rect 20858 7775 20990 7778
rect 10230 7773 20990 7775
rect 10230 7717 10268 7773
rect 10324 7740 20896 7773
rect 10324 7717 18064 7740
rect 10230 7715 18064 7717
rect 10230 7712 10362 7715
rect 17384 7676 18064 7715
rect 18128 7676 18700 7740
rect 18764 7715 19124 7740
rect 18764 7676 18808 7715
rect 17384 7641 18808 7676
rect 17384 7632 17536 7641
rect 17596 7632 17960 7641
rect 18020 7632 18384 7641
rect 18444 7632 18596 7641
rect 18656 7632 18808 7641
rect 19080 7676 19124 7715
rect 19188 7676 19336 7740
rect 19400 7676 19760 7740
rect 19824 7717 20896 7740
rect 20952 7717 20990 7773
rect 19824 7715 20990 7717
rect 19824 7676 20504 7715
rect 20858 7712 20990 7715
rect 19080 7641 20504 7676
rect 19080 7632 19232 7641
rect 19292 7632 19444 7641
rect 19504 7632 19868 7641
rect 19928 7632 20292 7641
rect 20352 7632 20504 7641
rect 17638 7620 17770 7629
rect 17638 7572 17676 7620
rect 17596 7564 17676 7572
rect 17732 7564 17770 7620
rect 17910 7620 18042 7629
rect 17910 7572 17948 7620
rect 17596 7555 17770 7564
rect 17808 7564 17948 7572
rect 18004 7572 18042 7620
rect 18416 7620 18548 7629
rect 18416 7572 18454 7620
rect 18004 7564 18172 7572
rect 17596 7528 17748 7555
rect 17596 7464 17640 7528
rect 17704 7464 17748 7528
rect 17596 7420 17748 7464
rect 17808 7528 18172 7564
rect 17808 7464 18064 7528
rect 18128 7464 18172 7528
rect 17808 7420 18172 7464
rect 18232 7564 18454 7572
rect 18510 7572 18548 7620
rect 18688 7620 18820 7629
rect 18688 7572 18726 7620
rect 18510 7564 18596 7572
rect 18232 7420 18596 7564
rect 18656 7564 18726 7572
rect 18782 7572 18820 7620
rect 18782 7564 24108 7572
rect 18656 7420 24108 7564
rect 18444 7360 18596 7420
rect 18444 7208 24108 7360
rect 18096 7104 24108 7148
rect 18020 7040 18064 7104
rect 18128 7040 24108 7104
rect 10230 7025 10362 7028
rect 17064 7025 17196 7028
rect 10230 7023 17196 7025
rect 10230 6967 10268 7023
rect 10324 6967 17102 7023
rect 17158 6967 17196 7023
rect 18096 6996 24108 7040
rect 10230 6965 17196 6967
rect 10230 6962 10362 6965
rect 17064 6962 17196 6965
rect 17384 6724 17748 6936
rect 17808 6892 18808 6936
rect 17808 6828 18064 6892
rect 18128 6828 18808 6892
rect 17808 6784 18808 6828
rect 17808 6724 18172 6784
rect 17384 6572 18172 6724
rect 18232 6724 18808 6784
rect 19080 6784 20504 6936
rect 19080 6724 19656 6784
rect 18232 6680 19656 6724
rect 18232 6616 19336 6680
rect 19400 6616 19656 6680
rect 18232 6572 19656 6616
rect 19716 6572 20080 6784
rect 20140 6572 20504 6784
rect 18020 6512 18172 6572
rect 18444 6512 18596 6572
rect 18020 6360 18596 6512
rect 19292 6512 19444 6572
rect 19716 6512 19868 6572
rect 19292 6360 19868 6512
rect 19368 5832 20080 5876
rect 19292 5768 19336 5832
rect 19400 5768 20080 5832
rect 19368 5724 20080 5768
rect 19928 5664 20080 5724
rect 17596 5452 17748 5664
rect 18232 5452 18596 5664
rect 19080 5452 19444 5664
rect 19928 5512 20928 5664
rect 19928 5452 20080 5512
rect 17596 5300 20080 5452
rect 20564 5452 20928 5512
rect 20564 5408 22200 5452
rect 20564 5344 22092 5408
rect 22156 5344 22200 5408
rect 20564 5300 22200 5344
rect 2544 4876 2908 5028
rect 2544 4817 2806 4876
rect 2544 4772 2696 4817
rect 2544 4708 2588 4772
rect 2652 4708 2696 4772
rect 2544 4664 2696 4708
rect 2881 4636 3013 4645
rect 2881 4580 2919 4636
rect 2975 4580 3013 4636
rect 2881 4571 3013 4580
rect 6360 4421 6724 4604
rect 6360 4365 6441 4421
rect 6497 4365 6724 4421
rect 6360 4348 6724 4365
rect 6360 4284 6404 4348
rect 6468 4284 6724 4348
rect 6360 4240 6724 4284
rect 2544 3968 2908 4180
rect 1908 3924 2908 3968
rect 1908 3860 1952 3924
rect 2016 3860 2908 3924
rect 1908 3816 2908 3860
rect 12296 3500 15628 3544
rect 2881 3452 3013 3461
rect 2881 3396 2919 3452
rect 2975 3396 3013 3452
rect 2881 3387 3013 3396
rect 12296 3436 15308 3500
rect 15372 3436 15628 3500
rect 12296 3392 15628 3436
rect 16748 3500 17112 3544
rect 16748 3436 16792 3500
rect 16856 3436 17112 3500
rect 16748 3392 17112 3436
rect 848 3288 2696 3332
rect 848 3224 892 3288
rect 956 3224 2588 3288
rect 2652 3224 2696 3288
rect 848 3215 2696 3224
rect 848 3180 2806 3215
rect 2544 3120 2806 3180
rect 2544 2968 2908 3120
rect 8664 2988 8796 2991
rect 8664 2986 14742 2988
rect 8664 2930 8702 2986
rect 8758 2930 14742 2986
rect 8664 2928 14742 2930
rect 8664 2925 8796 2928
rect 11919 2924 12051 2928
rect 11919 2908 11957 2924
rect 11872 2868 11957 2908
rect 12013 2868 12051 2924
rect 13401 2924 13533 2928
rect 13401 2908 13439 2924
rect 11872 2864 12051 2868
rect 11872 2800 11916 2864
rect 11980 2859 12051 2864
rect 13356 2868 13439 2908
rect 13495 2868 13533 2924
rect 14883 2924 15015 2933
rect 14883 2908 14921 2924
rect 13356 2864 13533 2868
rect 11980 2800 12024 2859
rect 11872 2756 12024 2800
rect 13356 2800 13400 2864
rect 13464 2859 13533 2864
rect 14840 2868 14921 2908
rect 14977 2868 15015 2924
rect 16365 2924 16497 2933
rect 16365 2908 16403 2924
rect 14840 2864 15015 2868
rect 13464 2800 13508 2859
rect 13356 2756 13508 2800
rect 14840 2800 14884 2864
rect 14948 2859 15015 2864
rect 16324 2868 16403 2908
rect 16459 2868 16497 2924
rect 16324 2864 16497 2868
rect 14948 2800 14992 2859
rect 14840 2756 14992 2800
rect 16324 2800 16368 2864
rect 16432 2859 16497 2864
rect 16432 2800 16476 2859
rect 16324 2756 16476 2800
rect 12296 2652 17112 2696
rect 12296 2588 14036 2652
rect 14100 2588 17112 2652
rect 12296 2544 17112 2588
rect 1484 2016 22624 2060
rect 1484 1952 1528 2016
rect 1592 1952 1740 2016
rect 1804 1952 1952 2016
rect 2016 1952 15308 2016
rect 15372 1952 16792 2016
rect 16856 1952 22092 2016
rect 22156 1952 22304 2016
rect 22368 1952 22516 2016
rect 22580 1952 22624 2016
rect 1484 1804 22624 1952
rect 1484 1740 1528 1804
rect 1592 1740 1740 1804
rect 1804 1740 1952 1804
rect 2016 1740 22092 1804
rect 22156 1740 22304 1804
rect 22368 1740 22516 1804
rect 22580 1740 22624 1804
rect 1484 1592 22624 1740
rect 1484 1528 1528 1592
rect 1592 1528 1740 1592
rect 1804 1528 1952 1592
rect 2016 1528 22092 1592
rect 22156 1528 22304 1592
rect 22368 1528 22516 1592
rect 22580 1528 22624 1592
rect 1484 1484 22624 1528
rect 424 956 23684 1000
rect 424 892 468 956
rect 532 892 680 956
rect 744 892 892 956
rect 956 892 14036 956
rect 14100 892 23152 956
rect 23216 892 23364 956
rect 23428 892 23576 956
rect 23640 892 23684 956
rect 424 744 23684 892
rect 424 680 468 744
rect 532 680 680 744
rect 744 680 892 744
rect 956 680 23152 744
rect 23216 680 23364 744
rect 23428 680 23576 744
rect 23640 680 23684 744
rect 424 532 23684 680
rect 424 468 468 532
rect 532 468 680 532
rect 744 468 892 532
rect 956 468 23152 532
rect 23216 468 23364 532
rect 23428 468 23576 532
rect 23640 468 23684 532
rect 424 424 23684 468
<< via3 >>
rect 468 36084 532 36148
rect 680 36084 744 36148
rect 892 36084 956 36148
rect 23152 36084 23216 36148
rect 23364 36084 23428 36148
rect 23576 36084 23640 36148
rect 468 35872 532 35936
rect 680 35872 744 35936
rect 892 35872 956 35936
rect 23152 35872 23216 35936
rect 23364 35872 23428 35936
rect 23576 35872 23640 35936
rect 468 35660 532 35724
rect 680 35660 744 35724
rect 892 35660 956 35724
rect 12340 35660 12404 35724
rect 17004 35660 17068 35724
rect 23152 35660 23216 35724
rect 23364 35660 23428 35724
rect 23576 35660 23640 35724
rect 1528 35024 1592 35088
rect 1740 35024 1804 35088
rect 1952 35024 2016 35088
rect 22092 35024 22156 35088
rect 22304 35024 22368 35088
rect 22516 35024 22580 35088
rect 1528 34812 1592 34876
rect 1740 34812 1804 34876
rect 1952 34812 2016 34876
rect 22092 34812 22156 34876
rect 22304 34812 22368 34876
rect 22516 34812 22580 34876
rect 1528 34600 1592 34664
rect 1740 34600 1804 34664
rect 1952 34600 2016 34664
rect 11492 34600 11556 34664
rect 15520 34600 15584 34664
rect 22092 34600 22156 34664
rect 22304 34600 22368 34664
rect 22516 34600 22580 34664
rect 12128 33752 12192 33816
rect 12340 33752 12404 33816
rect 17004 33752 17068 33816
rect 17216 33752 17280 33816
rect 11492 32268 11556 32332
rect 12340 32056 12404 32120
rect 15520 32268 15584 32332
rect 15732 32056 15796 32120
rect 12128 30784 12192 30848
rect 11916 30572 11980 30636
rect 17216 30784 17280 30848
rect 15520 30572 15584 30636
rect 12340 29300 12404 29364
rect 15732 29300 15796 29364
rect 11704 27604 11768 27668
rect 11916 27604 11980 27668
rect 15520 27604 15584 27668
rect 17004 27604 17068 27668
rect 15520 25908 15584 25972
rect 11704 24636 11768 24700
rect 12128 24424 12192 24488
rect 17004 24636 17068 24700
rect 17004 24424 17068 24488
rect 11916 22940 11980 23004
rect 15520 22940 15584 23004
rect 15732 22940 15796 23004
rect 12128 21668 12192 21732
rect 11704 21456 11768 21520
rect 17004 21456 17068 21520
rect 17216 21456 17280 21520
rect 11916 19972 11980 20036
rect 15732 19972 15796 20036
rect 15732 19760 15796 19824
rect 11280 18276 11344 18340
rect 11704 18276 11768 18340
rect 17216 18488 17280 18552
rect 15520 16792 15584 16856
rect 15732 16792 15796 16856
rect 11280 16156 11344 16220
rect 9584 15944 9648 16008
rect 11280 15308 11344 15372
rect 17004 15308 17068 15372
rect 9372 15096 9436 15160
rect 9584 14460 9648 14524
rect 11280 14460 11344 14524
rect 9584 14248 9648 14312
rect 9372 13612 9436 13676
rect 15520 13824 15584 13888
rect 17216 13612 17280 13676
rect 9372 13400 9436 13464
rect 9584 12764 9648 12828
rect 9584 12552 9648 12616
rect 9796 12552 9860 12616
rect 9796 12128 9860 12192
rect 17004 12340 17068 12404
rect 15520 12128 15584 12192
rect 9372 11916 9436 11980
rect 9372 11704 9436 11768
rect 9584 11068 9648 11132
rect 9584 10856 9648 10920
rect 11280 10644 11344 10708
rect 17216 10644 17280 10708
rect 17640 10644 17704 10708
rect 9372 10220 9436 10284
rect 11280 10220 11344 10284
rect 9584 9372 9648 9436
rect 15520 9160 15584 9224
rect 18064 8948 18128 9012
rect 17640 8100 17704 8164
rect 18488 7888 18552 7952
rect 23152 7888 23216 7952
rect 18064 7676 18128 7740
rect 18700 7676 18764 7740
rect 19124 7676 19188 7740
rect 19336 7676 19400 7740
rect 19760 7676 19824 7740
rect 17640 7464 17704 7528
rect 18064 7464 18128 7528
rect 18064 7040 18128 7104
rect 18064 6828 18128 6892
rect 19336 6616 19400 6680
rect 19336 5768 19400 5832
rect 22092 5344 22156 5408
rect 2588 4708 2652 4772
rect 6404 4284 6468 4348
rect 1952 3860 2016 3924
rect 15308 3436 15372 3500
rect 16792 3436 16856 3500
rect 892 3224 956 3288
rect 2588 3224 2652 3288
rect 11916 2800 11980 2864
rect 13400 2800 13464 2864
rect 14884 2800 14948 2864
rect 16368 2800 16432 2864
rect 14036 2588 14100 2652
rect 1528 1952 1592 2016
rect 1740 1952 1804 2016
rect 1952 1952 2016 2016
rect 15308 1952 15372 2016
rect 16792 1952 16856 2016
rect 22092 1952 22156 2016
rect 22304 1952 22368 2016
rect 22516 1952 22580 2016
rect 1528 1740 1592 1804
rect 1740 1740 1804 1804
rect 1952 1740 2016 1804
rect 22092 1740 22156 1804
rect 22304 1740 22368 1804
rect 22516 1740 22580 1804
rect 1528 1528 1592 1592
rect 1740 1528 1804 1592
rect 1952 1528 2016 1592
rect 22092 1528 22156 1592
rect 22304 1528 22368 1592
rect 22516 1528 22580 1592
rect 468 892 532 956
rect 680 892 744 956
rect 892 892 956 956
rect 14036 892 14100 956
rect 23152 892 23216 956
rect 23364 892 23428 956
rect 23576 892 23640 956
rect 468 680 532 744
rect 680 680 744 744
rect 892 680 956 744
rect 23152 680 23216 744
rect 23364 680 23428 744
rect 23576 680 23640 744
rect 468 468 532 532
rect 680 468 744 532
rect 892 468 956 532
rect 23152 468 23216 532
rect 23364 468 23428 532
rect 23576 468 23640 532
<< metal4 >>
rect 424 36148 1000 36192
rect 424 36084 468 36148
rect 532 36084 680 36148
rect 744 36084 892 36148
rect 956 36084 1000 36148
rect 424 35936 1000 36084
rect 424 35872 468 35936
rect 532 35872 680 35936
rect 744 35872 892 35936
rect 956 35872 1000 35936
rect 424 35724 1000 35872
rect 23108 36148 23684 36192
rect 23108 36084 23152 36148
rect 23216 36084 23364 36148
rect 23428 36084 23576 36148
rect 23640 36084 23684 36148
rect 23108 35936 23684 36084
rect 23108 35872 23152 35936
rect 23216 35872 23364 35936
rect 23428 35872 23576 35936
rect 23640 35872 23684 35936
rect 424 35660 468 35724
rect 532 35660 680 35724
rect 744 35660 892 35724
rect 956 35660 1000 35724
rect 424 3288 1000 35660
rect 12296 35724 12448 35768
rect 12296 35660 12340 35724
rect 12404 35660 12448 35724
rect 424 3224 892 3288
rect 956 3224 1000 3288
rect 424 956 1000 3224
rect 1484 35088 2060 35132
rect 1484 35024 1528 35088
rect 1592 35024 1740 35088
rect 1804 35024 1952 35088
rect 2016 35024 2060 35088
rect 1484 34876 2060 35024
rect 1484 34812 1528 34876
rect 1592 34812 1740 34876
rect 1804 34812 1952 34876
rect 2016 34812 2060 34876
rect 1484 34664 2060 34812
rect 1484 34600 1528 34664
rect 1592 34600 1740 34664
rect 1804 34600 1952 34664
rect 2016 34600 2060 34664
rect 1484 3924 2060 34600
rect 11448 34664 11600 34708
rect 11448 34600 11492 34664
rect 11556 34600 11600 34664
rect 11448 32332 11600 34600
rect 12114 33816 12206 33830
rect 12114 33784 12128 33816
rect 11448 32300 11492 32332
rect 11478 32268 11492 32300
rect 11556 32300 11600 32332
rect 12084 33752 12128 33784
rect 12192 33784 12206 33816
rect 12296 33816 12448 35660
rect 16960 35724 17112 35768
rect 16960 35660 17004 35724
rect 17068 35660 17112 35724
rect 12296 33784 12340 33816
rect 12192 33752 12236 33784
rect 11556 32268 11570 32300
rect 11478 32254 11570 32268
rect 12084 30848 12236 33752
rect 12326 33752 12340 33784
rect 12404 33784 12448 33816
rect 15476 34664 15628 34708
rect 15476 34600 15520 34664
rect 15584 34600 15628 34664
rect 12404 33752 12418 33784
rect 12326 33738 12418 33752
rect 15476 32332 15628 34600
rect 16960 33816 17112 35660
rect 23108 35724 23684 35872
rect 23108 35660 23152 35724
rect 23216 35660 23364 35724
rect 23428 35660 23576 35724
rect 23640 35660 23684 35724
rect 22048 35088 22624 35132
rect 22048 35024 22092 35088
rect 22156 35024 22304 35088
rect 22368 35024 22516 35088
rect 22580 35024 22624 35088
rect 22048 34876 22624 35024
rect 22048 34812 22092 34876
rect 22156 34812 22304 34876
rect 22368 34812 22516 34876
rect 22580 34812 22624 34876
rect 22048 34664 22624 34812
rect 22048 34600 22092 34664
rect 22156 34600 22304 34664
rect 22368 34600 22516 34664
rect 22580 34600 22624 34664
rect 16960 33784 17004 33816
rect 16990 33752 17004 33784
rect 17068 33784 17112 33816
rect 17172 33816 17324 33860
rect 17068 33752 17082 33784
rect 16990 33738 17082 33752
rect 17172 33752 17216 33816
rect 17280 33752 17324 33816
rect 15476 32300 15520 32332
rect 15506 32268 15520 32300
rect 15584 32300 15628 32332
rect 15584 32268 15598 32300
rect 15506 32254 15598 32268
rect 12084 30784 12128 30848
rect 12192 30784 12236 30848
rect 12084 30740 12236 30784
rect 12296 32120 12448 32164
rect 12296 32056 12340 32120
rect 12404 32056 12448 32120
rect 15718 32120 15810 32134
rect 15718 32088 15732 32120
rect 11902 30636 11994 30650
rect 11902 30604 11916 30636
rect 11872 30572 11916 30604
rect 11980 30604 11994 30636
rect 11980 30572 12024 30604
rect 11690 27668 11782 27682
rect 11690 27636 11704 27668
rect 11660 27604 11704 27636
rect 11768 27636 11782 27668
rect 11872 27668 12024 30572
rect 12296 29364 12448 32056
rect 15688 32056 15732 32088
rect 15796 32088 15810 32120
rect 15796 32056 15840 32088
rect 15506 30636 15598 30650
rect 15506 30604 15520 30636
rect 12296 29332 12340 29364
rect 12326 29300 12340 29332
rect 12404 29332 12448 29364
rect 15476 30572 15520 30604
rect 15584 30604 15598 30636
rect 15584 30572 15628 30604
rect 12404 29300 12418 29332
rect 12326 29286 12418 29300
rect 11768 27604 11812 27636
rect 11660 24700 11812 27604
rect 11872 27604 11916 27668
rect 11980 27604 12024 27668
rect 11872 27560 12024 27604
rect 15476 27668 15628 30572
rect 15688 29364 15840 32056
rect 17172 30848 17324 33752
rect 17172 30816 17216 30848
rect 17202 30784 17216 30816
rect 17280 30816 17324 30848
rect 17280 30784 17294 30816
rect 17202 30770 17294 30784
rect 15688 29300 15732 29364
rect 15796 29300 15840 29364
rect 15688 29256 15840 29300
rect 15476 27604 15520 27668
rect 15584 27604 15628 27668
rect 16990 27668 17082 27682
rect 16990 27636 17004 27668
rect 15476 27560 15628 27604
rect 16960 27604 17004 27636
rect 17068 27636 17082 27668
rect 17068 27604 17112 27636
rect 15506 25972 15598 25986
rect 15506 25940 15520 25972
rect 11660 24636 11704 24700
rect 11768 24636 11812 24700
rect 11660 24592 11812 24636
rect 15476 25908 15520 25940
rect 15584 25940 15598 25972
rect 15584 25908 15628 25940
rect 12084 24488 12236 24532
rect 12084 24424 12128 24488
rect 12192 24424 12236 24488
rect 11872 23004 12024 23048
rect 11872 22940 11916 23004
rect 11980 22940 12024 23004
rect 11690 21520 11782 21534
rect 11690 21488 11704 21520
rect 11660 21456 11704 21488
rect 11768 21488 11782 21520
rect 11768 21456 11812 21488
rect 11236 18340 11388 18384
rect 11236 18276 11280 18340
rect 11344 18276 11388 18340
rect 11236 16220 11388 18276
rect 11660 18340 11812 21456
rect 11872 20036 12024 22940
rect 12084 21732 12236 24424
rect 15476 23004 15628 25908
rect 16960 24700 17112 27604
rect 16960 24636 17004 24700
rect 17068 24636 17112 24700
rect 16960 24592 17112 24636
rect 16960 24488 17112 24532
rect 16960 24424 17004 24488
rect 17068 24424 17112 24488
rect 15476 22940 15520 23004
rect 15584 22940 15628 23004
rect 15718 23004 15810 23018
rect 15718 22972 15732 23004
rect 15476 22896 15628 22940
rect 15688 22940 15732 22972
rect 15796 22972 15810 23004
rect 15796 22940 15840 22972
rect 12084 21700 12128 21732
rect 12114 21668 12128 21700
rect 12192 21700 12236 21732
rect 12192 21668 12206 21700
rect 12114 21654 12206 21668
rect 11872 20004 11916 20036
rect 11902 19972 11916 20004
rect 11980 20004 12024 20036
rect 15688 20036 15840 22940
rect 16960 21520 17112 24424
rect 16960 21488 17004 21520
rect 16990 21456 17004 21488
rect 17068 21488 17112 21520
rect 17202 21520 17294 21534
rect 17202 21488 17216 21520
rect 17068 21456 17082 21488
rect 16990 21442 17082 21456
rect 17172 21456 17216 21488
rect 17280 21488 17294 21520
rect 17280 21456 17324 21488
rect 11980 19972 11994 20004
rect 11902 19958 11994 19972
rect 15688 19972 15732 20036
rect 15796 19972 15840 20036
rect 15688 19928 15840 19972
rect 15718 19824 15810 19838
rect 15718 19792 15732 19824
rect 11660 18276 11704 18340
rect 11768 18276 11812 18340
rect 11660 18232 11812 18276
rect 15688 19760 15732 19792
rect 15796 19792 15810 19824
rect 15796 19760 15840 19792
rect 11236 16188 11280 16220
rect 11266 16156 11280 16188
rect 11344 16188 11388 16220
rect 15476 16856 15628 16900
rect 15476 16792 15520 16856
rect 15584 16792 15628 16856
rect 11344 16156 11358 16188
rect 11266 16142 11358 16156
rect 9540 16008 9692 16052
rect 9540 15944 9584 16008
rect 9648 15944 9692 16008
rect 9358 15160 9450 15174
rect 9358 15128 9372 15160
rect 9328 15096 9372 15128
rect 9436 15128 9450 15160
rect 9436 15096 9480 15128
rect 9328 13676 9480 15096
rect 9540 14524 9692 15944
rect 9540 14492 9584 14524
rect 9570 14460 9584 14492
rect 9648 14492 9692 14524
rect 11236 15372 11388 15416
rect 11236 15308 11280 15372
rect 11344 15308 11388 15372
rect 11236 14524 11388 15308
rect 11236 14492 11280 14524
rect 9648 14460 9662 14492
rect 9570 14446 9662 14460
rect 11266 14460 11280 14492
rect 11344 14492 11388 14524
rect 11344 14460 11358 14492
rect 11266 14446 11358 14460
rect 9570 14312 9662 14326
rect 9570 14280 9584 14312
rect 9328 13612 9372 13676
rect 9436 13612 9480 13676
rect 9328 13568 9480 13612
rect 9540 14248 9584 14280
rect 9648 14280 9662 14312
rect 9648 14248 9692 14280
rect 9328 13464 9480 13508
rect 9328 13400 9372 13464
rect 9436 13400 9480 13464
rect 9328 11980 9480 13400
rect 9540 12828 9692 14248
rect 15476 13888 15628 16792
rect 15688 16856 15840 19760
rect 17172 18552 17324 21456
rect 17172 18488 17216 18552
rect 17280 18488 17324 18552
rect 17172 18444 17324 18488
rect 15688 16792 15732 16856
rect 15796 16792 15840 16856
rect 15688 16748 15840 16792
rect 16990 15372 17082 15386
rect 16990 15340 17004 15372
rect 15476 13856 15520 13888
rect 15506 13824 15520 13856
rect 15584 13856 15628 13888
rect 16960 15308 17004 15340
rect 17068 15340 17082 15372
rect 17068 15308 17112 15340
rect 15584 13824 15598 13856
rect 15506 13810 15598 13824
rect 9540 12764 9584 12828
rect 9648 12764 9692 12828
rect 9540 12720 9692 12764
rect 9328 11948 9372 11980
rect 9358 11916 9372 11948
rect 9436 11948 9480 11980
rect 9540 12616 9692 12660
rect 9540 12552 9584 12616
rect 9648 12552 9692 12616
rect 9782 12616 9874 12630
rect 9782 12584 9796 12616
rect 9436 11916 9450 11948
rect 9358 11902 9450 11916
rect 9358 11768 9450 11782
rect 9358 11736 9372 11768
rect 9328 11704 9372 11736
rect 9436 11736 9450 11768
rect 9436 11704 9480 11736
rect 9328 10284 9480 11704
rect 9540 11132 9692 12552
rect 9752 12552 9796 12584
rect 9860 12584 9874 12616
rect 9860 12552 9904 12584
rect 9752 12192 9904 12552
rect 16960 12404 17112 15308
rect 16960 12340 17004 12404
rect 17068 12340 17112 12404
rect 16960 12296 17112 12340
rect 17172 13676 17324 13720
rect 17172 13612 17216 13676
rect 17280 13612 17324 13676
rect 9752 12128 9796 12192
rect 9860 12128 9904 12192
rect 15506 12192 15598 12206
rect 15506 12160 15520 12192
rect 9752 12084 9904 12128
rect 15476 12128 15520 12160
rect 15584 12160 15598 12192
rect 15584 12128 15628 12160
rect 9540 11100 9584 11132
rect 9570 11068 9584 11100
rect 9648 11100 9692 11132
rect 9648 11068 9662 11100
rect 9570 11054 9662 11068
rect 9570 10920 9662 10934
rect 9570 10888 9584 10920
rect 9328 10220 9372 10284
rect 9436 10220 9480 10284
rect 9328 10176 9480 10220
rect 9540 10856 9584 10888
rect 9648 10888 9662 10920
rect 9648 10856 9692 10888
rect 9540 9436 9692 10856
rect 11236 10708 11388 10752
rect 11236 10644 11280 10708
rect 11344 10644 11388 10708
rect 11236 10284 11388 10644
rect 11236 10252 11280 10284
rect 11266 10220 11280 10252
rect 11344 10252 11388 10284
rect 11344 10220 11358 10252
rect 11266 10206 11358 10220
rect 9540 9372 9584 9436
rect 9648 9372 9692 9436
rect 9540 9328 9692 9372
rect 15476 9224 15628 12128
rect 17172 10708 17324 13612
rect 17172 10676 17216 10708
rect 17202 10644 17216 10676
rect 17280 10676 17324 10708
rect 17626 10708 17718 10722
rect 17626 10676 17640 10708
rect 17280 10644 17294 10676
rect 17202 10630 17294 10644
rect 17596 10644 17640 10676
rect 17704 10676 17718 10708
rect 17704 10644 17748 10676
rect 15476 9160 15520 9224
rect 15584 9160 15628 9224
rect 15476 9116 15628 9160
rect 17596 8164 17748 10644
rect 17596 8100 17640 8164
rect 17704 8100 17748 8164
rect 17596 8056 17748 8100
rect 18020 9012 18172 9056
rect 18020 8948 18064 9012
rect 18128 8948 18172 9012
rect 18020 7740 18172 8948
rect 18020 7708 18064 7740
rect 18050 7676 18064 7708
rect 18128 7708 18172 7740
rect 18232 7952 18596 7996
rect 18232 7888 18488 7952
rect 18552 7888 18596 7952
rect 18232 7844 18596 7888
rect 18128 7676 18142 7708
rect 18050 7662 18142 7676
rect 17626 7528 17718 7542
rect 17626 7496 17640 7528
rect 17596 7464 17640 7496
rect 17704 7496 17718 7528
rect 18050 7528 18142 7542
rect 18050 7496 18064 7528
rect 17704 7464 17748 7496
rect 2574 4772 2666 4786
rect 2574 4740 2588 4772
rect 1484 3860 1952 3924
rect 2016 3860 2060 3924
rect 1484 2016 2060 3860
rect 2544 4708 2588 4740
rect 2652 4740 2666 4772
rect 2652 4708 2696 4740
rect 2544 3288 2696 4708
rect 6390 4348 6482 4362
rect 6390 4316 6404 4348
rect 2544 3224 2588 3288
rect 2652 3224 2696 3288
rect 2544 3180 2696 3224
rect 6360 4284 6404 4316
rect 6468 4316 6482 4348
rect 6468 4284 6512 4316
rect 1484 1952 1528 2016
rect 1592 1952 1740 2016
rect 1804 1952 1952 2016
rect 2016 1952 2060 2016
rect 1484 1804 2060 1952
rect 1484 1740 1528 1804
rect 1592 1740 1740 1804
rect 1804 1740 1952 1804
rect 2016 1740 2060 1804
rect 1484 1592 2060 1740
rect 1484 1528 1528 1592
rect 1592 1528 1740 1592
rect 1804 1528 1952 1592
rect 2016 1528 2060 1592
rect 1484 1484 2060 1528
rect 424 892 468 956
rect 532 892 680 956
rect 744 892 892 956
rect 956 892 1000 956
rect 424 744 1000 892
rect 424 680 468 744
rect 532 680 680 744
rect 744 680 892 744
rect 956 680 1000 744
rect 424 532 1000 680
rect 424 468 468 532
rect 532 468 680 532
rect 744 468 892 532
rect 956 468 1000 532
rect 424 424 1000 468
rect 6360 0 6512 4284
rect 15294 3500 15386 3514
rect 15294 3468 15308 3500
rect 15264 3436 15308 3468
rect 15372 3468 15386 3500
rect 16778 3500 16870 3514
rect 16778 3468 16792 3500
rect 15372 3436 15416 3468
rect 11902 2864 11994 2878
rect 11902 2832 11916 2864
rect 11872 2800 11916 2832
rect 11980 2832 11994 2864
rect 13386 2864 13478 2878
rect 13386 2832 13400 2864
rect 11980 2800 12024 2832
rect 11872 0 12024 2800
rect 13356 2800 13400 2832
rect 13464 2832 13478 2864
rect 14870 2864 14962 2878
rect 14870 2832 14884 2864
rect 13464 2800 13508 2832
rect 13356 0 13508 2800
rect 14840 2800 14884 2832
rect 14948 2832 14962 2864
rect 14948 2800 14992 2832
rect 14022 2652 14114 2666
rect 14022 2620 14036 2652
rect 13992 2588 14036 2620
rect 14100 2620 14114 2652
rect 14100 2588 14144 2620
rect 13992 956 14144 2588
rect 13992 892 14036 956
rect 14100 892 14144 956
rect 13992 848 14144 892
rect 14840 0 14992 2800
rect 15264 2016 15416 3436
rect 16748 3436 16792 3468
rect 16856 3468 16870 3500
rect 16856 3436 16900 3468
rect 16354 2864 16446 2878
rect 16354 2832 16368 2864
rect 15264 1952 15308 2016
rect 15372 1952 15416 2016
rect 15264 1908 15416 1952
rect 16324 2800 16368 2832
rect 16432 2832 16446 2864
rect 16432 2800 16476 2832
rect 16324 0 16476 2800
rect 16748 2016 16900 3436
rect 16748 1952 16792 2016
rect 16856 1952 16900 2016
rect 16748 1908 16900 1952
rect 17596 0 17748 7464
rect 18020 7464 18064 7496
rect 18128 7496 18142 7528
rect 18128 7464 18172 7496
rect 18020 7104 18172 7464
rect 18020 7040 18064 7104
rect 18128 7040 18172 7104
rect 18020 6996 18172 7040
rect 18232 6936 18384 7844
rect 18732 7754 19232 7784
rect 19368 7754 19868 7784
rect 18686 7740 19232 7754
rect 18686 7676 18700 7740
rect 18764 7676 19124 7740
rect 19188 7676 19232 7740
rect 18686 7662 19232 7676
rect 19322 7740 19868 7754
rect 19322 7676 19336 7740
rect 19400 7676 19760 7740
rect 19824 7676 19868 7740
rect 19322 7662 19868 7676
rect 18732 7632 19232 7662
rect 19368 7632 19868 7662
rect 18096 6906 18384 6936
rect 18050 6892 18384 6906
rect 18050 6828 18064 6892
rect 18128 6828 18384 6892
rect 18050 6814 18384 6828
rect 18096 6784 18384 6814
rect 19322 6680 19414 6694
rect 19322 6648 19336 6680
rect 19292 6616 19336 6648
rect 19400 6648 19414 6680
rect 19400 6616 19444 6648
rect 19292 5832 19444 6616
rect 19292 5768 19336 5832
rect 19400 5768 19444 5832
rect 19292 5724 19444 5768
rect 22048 5408 22624 34600
rect 22048 5344 22092 5408
rect 22156 5344 22624 5408
rect 22048 2016 22624 5344
rect 22048 1952 22092 2016
rect 22156 1952 22304 2016
rect 22368 1952 22516 2016
rect 22580 1952 22624 2016
rect 22048 1804 22624 1952
rect 22048 1740 22092 1804
rect 22156 1740 22304 1804
rect 22368 1740 22516 1804
rect 22580 1740 22624 1804
rect 22048 1592 22624 1740
rect 22048 1528 22092 1592
rect 22156 1528 22304 1592
rect 22368 1528 22516 1592
rect 22580 1528 22624 1592
rect 22048 1484 22624 1528
rect 23108 7952 23684 35660
rect 23108 7888 23152 7952
rect 23216 7888 23684 7952
rect 23108 956 23684 7888
rect 23108 892 23152 956
rect 23216 892 23364 956
rect 23428 892 23576 956
rect 23640 892 23684 956
rect 23108 744 23684 892
rect 23108 680 23152 744
rect 23216 680 23364 744
rect 23428 680 23576 744
rect 23640 680 23684 744
rect 23108 532 23684 680
rect 23108 468 23152 532
rect 23216 468 23364 532
rect 23428 468 23576 532
rect 23640 468 23684 532
rect 23108 424 23684 468
use contact_28  contact_28_0
timestamp 1644949024
transform 1 0 23108 0 1 7874
box 0 0 1 1
use contact_28  contact_28_1
timestamp 1644949024
transform 1 0 19716 0 1 7662
box 0 0 1 1
use contact_28  contact_28_2
timestamp 1644949024
transform 1 0 19292 0 1 7662
box 0 0 1 1
use contact_28  contact_28_3
timestamp 1644949024
transform 1 0 19080 0 1 7662
box 0 0 1 1
use contact_28  contact_28_4
timestamp 1644949024
transform 1 0 18656 0 1 7662
box 0 0 1 1
use contact_28  contact_28_5
timestamp 1644949024
transform 1 0 18020 0 1 8934
box 0 0 1 1
use contact_28  contact_28_6
timestamp 1644949024
transform 1 0 18020 0 1 7662
box 0 0 1 1
use contact_28  contact_28_7
timestamp 1644949024
transform 1 0 16960 0 1 35646
box 0 0 1 1
use contact_28  contact_28_8
timestamp 1644949024
transform 1 0 16960 0 1 33738
box 0 0 1 1
use contact_28  contact_28_9
timestamp 1644949024
transform 1 0 16960 0 1 24410
box 0 0 1 1
use contact_28  contact_28_10
timestamp 1644949024
transform 1 0 16960 0 1 21442
box 0 0 1 1
use contact_28  contact_28_11
timestamp 1644949024
transform 1 0 17172 0 1 18474
box 0 0 1 1
use contact_28  contact_28_12
timestamp 1644949024
transform 1 0 17172 0 1 21442
box 0 0 1 1
use contact_28  contact_28_13
timestamp 1644949024
transform 1 0 17172 0 1 33738
box 0 0 1 1
use contact_28  contact_28_14
timestamp 1644949024
transform 1 0 17172 0 1 30770
box 0 0 1 1
use contact_28  contact_28_15
timestamp 1644949024
transform 1 0 16960 0 1 24622
box 0 0 1 1
use contact_28  contact_28_16
timestamp 1644949024
transform 1 0 16960 0 1 27590
box 0 0 1 1
use contact_28  contact_28_17
timestamp 1644949024
transform 1 0 16960 0 1 12326
box 0 0 1 1
use contact_28  contact_28_18
timestamp 1644949024
transform 1 0 16960 0 1 15294
box 0 0 1 1
use contact_28  contact_28_19
timestamp 1644949024
transform 1 0 15476 0 1 27590
box 0 0 1 1
use contact_28  contact_28_20
timestamp 1644949024
transform 1 0 15476 0 1 30558
box 0 0 1 1
use contact_28  contact_28_21
timestamp 1644949024
transform 1 0 15476 0 1 9146
box 0 0 1 1
use contact_28  contact_28_22
timestamp 1644949024
transform 1 0 15476 0 1 12114
box 0 0 1 1
use contact_28  contact_28_23
timestamp 1644949024
transform 1 0 13992 0 1 878
box 0 0 1 1
use contact_28  contact_28_24
timestamp 1644949024
transform 1 0 13992 0 1 2574
box 0 0 1 1
use contact_28  contact_28_25
timestamp 1644949024
transform 1 0 12296 0 1 35646
box 0 0 1 1
use contact_28  contact_28_26
timestamp 1644949024
transform 1 0 12296 0 1 33738
box 0 0 1 1
use contact_28  contact_28_27
timestamp 1644949024
transform 1 0 12084 0 1 30770
box 0 0 1 1
use contact_28  contact_28_28
timestamp 1644949024
transform 1 0 12084 0 1 33738
box 0 0 1 1
use contact_28  contact_28_29
timestamp 1644949024
transform 1 0 12084 0 1 24410
box 0 0 1 1
use contact_28  contact_28_30
timestamp 1644949024
transform 1 0 12084 0 1 21654
box 0 0 1 1
use contact_28  contact_28_31
timestamp 1644949024
transform 1 0 11660 0 1 18262
box 0 0 1 1
use contact_28  contact_28_32
timestamp 1644949024
transform 1 0 11660 0 1 21442
box 0 0 1 1
use contact_28  contact_28_33
timestamp 1644949024
transform 1 0 11660 0 1 24622
box 0 0 1 1
use contact_28  contact_28_34
timestamp 1644949024
transform 1 0 11660 0 1 27590
box 0 0 1 1
use contact_28  contact_28_35
timestamp 1644949024
transform 1 0 11872 0 1 27590
box 0 0 1 1
use contact_28  contact_28_36
timestamp 1644949024
transform 1 0 11872 0 1 30558
box 0 0 1 1
use contact_28  contact_28_37
timestamp 1644949024
transform 1 0 11236 0 1 18262
box 0 0 1 1
use contact_28  contact_28_38
timestamp 1644949024
transform 1 0 11236 0 1 16142
box 0 0 1 1
use contact_28  contact_28_39
timestamp 1644949024
transform 1 0 9752 0 1 12114
box 0 0 1 1
use contact_28  contact_28_40
timestamp 1644949024
transform 1 0 9752 0 1 12538
box 0 0 1 1
use contact_28  contact_28_41
timestamp 1644949024
transform 1 0 9540 0 1 9358
box 0 0 1 1
use contact_28  contact_28_42
timestamp 1644949024
transform 1 0 9540 0 1 10842
box 0 0 1 1
use contact_28  contact_28_43
timestamp 1644949024
transform 1 0 9540 0 1 12538
box 0 0 1 1
use contact_28  contact_28_44
timestamp 1644949024
transform 1 0 9540 0 1 11054
box 0 0 1 1
use contact_28  contact_28_45
timestamp 1644949024
transform 1 0 11236 0 1 15294
box 0 0 1 1
use contact_28  contact_28_46
timestamp 1644949024
transform 1 0 11236 0 1 14446
box 0 0 1 1
use contact_28  contact_28_47
timestamp 1644949024
transform 1 0 9540 0 1 15930
box 0 0 1 1
use contact_28  contact_28_48
timestamp 1644949024
transform 1 0 9540 0 1 14446
box 0 0 1 1
use contact_28  contact_28_49
timestamp 1644949024
transform 1 0 9540 0 1 12750
box 0 0 1 1
use contact_28  contact_28_50
timestamp 1644949024
transform 1 0 9540 0 1 14234
box 0 0 1 1
use contact_28  contact_28_51
timestamp 1644949024
transform 1 0 848 0 1 3210
box 0 0 1 1
use contact_28  contact_28_52
timestamp 1644949024
transform 1 0 2544 0 1 3210
box 0 0 1 1
use contact_28  contact_28_53
timestamp 1644949024
transform 1 0 2544 0 1 4694
box 0 0 1 1
use contact_28  contact_28_54
timestamp 1644949024
transform 1 0 22048 0 1 5330
box 0 0 1 1
use contact_28  contact_28_55
timestamp 1644949024
transform 1 0 19292 0 1 5754
box 0 0 1 1
use contact_28  contact_28_56
timestamp 1644949024
transform 1 0 19292 0 1 6602
box 0 0 1 1
use contact_28  contact_28_57
timestamp 1644949024
transform 1 0 18444 0 1 7874
box 0 0 1 1
use contact_28  contact_28_58
timestamp 1644949024
transform 1 0 18020 0 1 6814
box 0 0 1 1
use contact_28  contact_28_59
timestamp 1644949024
transform 1 0 17596 0 1 8086
box 0 0 1 1
use contact_28  contact_28_60
timestamp 1644949024
transform 1 0 17596 0 1 10630
box 0 0 1 1
use contact_28  contact_28_61
timestamp 1644949024
transform 1 0 17172 0 1 13598
box 0 0 1 1
use contact_28  contact_28_62
timestamp 1644949024
transform 1 0 17172 0 1 10630
box 0 0 1 1
use contact_28  contact_28_63
timestamp 1644949024
transform 1 0 16748 0 1 1938
box 0 0 1 1
use contact_28  contact_28_64
timestamp 1644949024
transform 1 0 16748 0 1 3422
box 0 0 1 1
use contact_28  contact_28_65
timestamp 1644949024
transform 1 0 15688 0 1 16778
box 0 0 1 1
use contact_28  contact_28_66
timestamp 1644949024
transform 1 0 15688 0 1 19746
box 0 0 1 1
use contact_28  contact_28_67
timestamp 1644949024
transform 1 0 15688 0 1 19958
box 0 0 1 1
use contact_28  contact_28_68
timestamp 1644949024
transform 1 0 15688 0 1 22926
box 0 0 1 1
use contact_28  contact_28_69
timestamp 1644949024
transform 1 0 15476 0 1 16778
box 0 0 1 1
use contact_28  contact_28_70
timestamp 1644949024
transform 1 0 15476 0 1 13810
box 0 0 1 1
use contact_28  contact_28_71
timestamp 1644949024
transform 1 0 15476 0 1 34586
box 0 0 1 1
use contact_28  contact_28_72
timestamp 1644949024
transform 1 0 15476 0 1 32254
box 0 0 1 1
use contact_28  contact_28_73
timestamp 1644949024
transform 1 0 15688 0 1 29286
box 0 0 1 1
use contact_28  contact_28_74
timestamp 1644949024
transform 1 0 15688 0 1 32042
box 0 0 1 1
use contact_28  contact_28_75
timestamp 1644949024
transform 1 0 15476 0 1 22926
box 0 0 1 1
use contact_28  contact_28_76
timestamp 1644949024
transform 1 0 15476 0 1 25894
box 0 0 1 1
use contact_28  contact_28_77
timestamp 1644949024
transform 1 0 15264 0 1 1938
box 0 0 1 1
use contact_28  contact_28_78
timestamp 1644949024
transform 1 0 15264 0 1 3422
box 0 0 1 1
use contact_28  contact_28_79
timestamp 1644949024
transform 1 0 12296 0 1 32042
box 0 0 1 1
use contact_28  contact_28_80
timestamp 1644949024
transform 1 0 12296 0 1 29286
box 0 0 1 1
use contact_28  contact_28_81
timestamp 1644949024
transform 1 0 11872 0 1 22926
box 0 0 1 1
use contact_28  contact_28_82
timestamp 1644949024
transform 1 0 11872 0 1 19958
box 0 0 1 1
use contact_28  contact_28_83
timestamp 1644949024
transform 1 0 11448 0 1 34586
box 0 0 1 1
use contact_28  contact_28_84
timestamp 1644949024
transform 1 0 11448 0 1 32254
box 0 0 1 1
use contact_28  contact_28_85
timestamp 1644949024
transform 1 0 11236 0 1 10630
box 0 0 1 1
use contact_28  contact_28_86
timestamp 1644949024
transform 1 0 11236 0 1 10206
box 0 0 1 1
use contact_28  contact_28_87
timestamp 1644949024
transform 1 0 9328 0 1 10206
box 0 0 1 1
use contact_28  contact_28_88
timestamp 1644949024
transform 1 0 9328 0 1 11690
box 0 0 1 1
use contact_28  contact_28_89
timestamp 1644949024
transform 1 0 9328 0 1 13386
box 0 0 1 1
use contact_28  contact_28_90
timestamp 1644949024
transform 1 0 9328 0 1 11902
box 0 0 1 1
use contact_28  contact_28_91
timestamp 1644949024
transform 1 0 9328 0 1 13598
box 0 0 1 1
use contact_28  contact_28_92
timestamp 1644949024
transform 1 0 9328 0 1 15082
box 0 0 1 1
use contact_28  contact_28_93
timestamp 1644949024
transform 1 0 1908 0 1 3846
box 0 0 1 1
use contact_30  contact_30_0
timestamp 1644949024
transform 1 0 23108 0 1 454
box 0 0 1 1
use contact_30  contact_30_1
timestamp 1644949024
transform 1 0 848 0 1 878
box 0 0 1 1
use contact_30  contact_30_2
timestamp 1644949024
transform 1 0 23532 0 1 35858
box 0 0 1 1
use contact_30  contact_30_3
timestamp 1644949024
transform 1 0 23532 0 1 878
box 0 0 1 1
use contact_30  contact_30_4
timestamp 1644949024
transform 1 0 636 0 1 878
box 0 0 1 1
use contact_30  contact_30_5
timestamp 1644949024
transform 1 0 23320 0 1 36070
box 0 0 1 1
use contact_30  contact_30_6
timestamp 1644949024
transform 1 0 848 0 1 35858
box 0 0 1 1
use contact_30  contact_30_7
timestamp 1644949024
transform 1 0 424 0 1 878
box 0 0 1 1
use contact_30  contact_30_8
timestamp 1644949024
transform 1 0 23320 0 1 666
box 0 0 1 1
use contact_30  contact_30_9
timestamp 1644949024
transform 1 0 848 0 1 454
box 0 0 1 1
use contact_30  contact_30_10
timestamp 1644949024
transform 1 0 23108 0 1 36070
box 0 0 1 1
use contact_30  contact_30_11
timestamp 1644949024
transform 1 0 636 0 1 35858
box 0 0 1 1
use contact_30  contact_30_12
timestamp 1644949024
transform 1 0 23108 0 1 666
box 0 0 1 1
use contact_30  contact_30_13
timestamp 1644949024
transform 1 0 23532 0 1 454
box 0 0 1 1
use contact_30  contact_30_14
timestamp 1644949024
transform 1 0 636 0 1 454
box 0 0 1 1
use contact_30  contact_30_15
timestamp 1644949024
transform 1 0 424 0 1 35858
box 0 0 1 1
use contact_30  contact_30_16
timestamp 1644949024
transform 1 0 23320 0 1 35646
box 0 0 1 1
use contact_30  contact_30_17
timestamp 1644949024
transform 1 0 424 0 1 454
box 0 0 1 1
use contact_30  contact_30_18
timestamp 1644949024
transform 1 0 23108 0 1 35646
box 0 0 1 1
use contact_30  contact_30_19
timestamp 1644949024
transform 1 0 848 0 1 36070
box 0 0 1 1
use contact_30  contact_30_20
timestamp 1644949024
transform 1 0 23532 0 1 36070
box 0 0 1 1
use contact_30  contact_30_21
timestamp 1644949024
transform 1 0 636 0 1 36070
box 0 0 1 1
use contact_30  contact_30_22
timestamp 1644949024
transform 1 0 23532 0 1 666
box 0 0 1 1
use contact_30  contact_30_23
timestamp 1644949024
transform 1 0 424 0 1 35646
box 0 0 1 1
use contact_30  contact_30_24
timestamp 1644949024
transform 1 0 848 0 1 666
box 0 0 1 1
use contact_30  contact_30_25
timestamp 1644949024
transform 1 0 424 0 1 36070
box 0 0 1 1
use contact_30  contact_30_26
timestamp 1644949024
transform 1 0 23320 0 1 35858
box 0 0 1 1
use contact_30  contact_30_27
timestamp 1644949024
transform 1 0 848 0 1 35646
box 0 0 1 1
use contact_30  contact_30_28
timestamp 1644949024
transform 1 0 23532 0 1 35646
box 0 0 1 1
use contact_30  contact_30_29
timestamp 1644949024
transform 1 0 23108 0 1 878
box 0 0 1 1
use contact_30  contact_30_30
timestamp 1644949024
transform 1 0 23108 0 1 35858
box 0 0 1 1
use contact_30  contact_30_31
timestamp 1644949024
transform 1 0 636 0 1 35646
box 0 0 1 1
use contact_30  contact_30_32
timestamp 1644949024
transform 1 0 636 0 1 666
box 0 0 1 1
use contact_30  contact_30_33
timestamp 1644949024
transform 1 0 23320 0 1 878
box 0 0 1 1
use contact_30  contact_30_34
timestamp 1644949024
transform 1 0 424 0 1 666
box 0 0 1 1
use contact_30  contact_30_35
timestamp 1644949024
transform 1 0 23320 0 1 454
box 0 0 1 1
use contact_30  contact_30_36
timestamp 1644949024
transform 1 0 22472 0 1 1514
box 0 0 1 1
use contact_30  contact_30_37
timestamp 1644949024
transform 1 0 1484 0 1 34586
box 0 0 1 1
use contact_30  contact_30_38
timestamp 1644949024
transform 1 0 22260 0 1 1726
box 0 0 1 1
use contact_30  contact_30_39
timestamp 1644949024
transform 1 0 1484 0 1 1938
box 0 0 1 1
use contact_30  contact_30_40
timestamp 1644949024
transform 1 0 1908 0 1 1514
box 0 0 1 1
use contact_30  contact_30_41
timestamp 1644949024
transform 1 0 1696 0 1 34798
box 0 0 1 1
use contact_30  contact_30_42
timestamp 1644949024
transform 1 0 22048 0 1 1726
box 0 0 1 1
use contact_30  contact_30_43
timestamp 1644949024
transform 1 0 1696 0 1 1726
box 0 0 1 1
use contact_30  contact_30_44
timestamp 1644949024
transform 1 0 1484 0 1 1514
box 0 0 1 1
use contact_30  contact_30_45
timestamp 1644949024
transform 1 0 22472 0 1 34798
box 0 0 1 1
use contact_30  contact_30_46
timestamp 1644949024
transform 1 0 1908 0 1 34798
box 0 0 1 1
use contact_30  contact_30_47
timestamp 1644949024
transform 1 0 22048 0 1 35010
box 0 0 1 1
use contact_30  contact_30_48
timestamp 1644949024
transform 1 0 1696 0 1 35010
box 0 0 1 1
use contact_30  contact_30_49
timestamp 1644949024
transform 1 0 22472 0 1 1726
box 0 0 1 1
use contact_30  contact_30_50
timestamp 1644949024
transform 1 0 1696 0 1 34586
box 0 0 1 1
use contact_30  contact_30_51
timestamp 1644949024
transform 1 0 1484 0 1 34798
box 0 0 1 1
use contact_30  contact_30_52
timestamp 1644949024
transform 1 0 22260 0 1 35010
box 0 0 1 1
use contact_30  contact_30_53
timestamp 1644949024
transform 1 0 22260 0 1 1938
box 0 0 1 1
use contact_30  contact_30_54
timestamp 1644949024
transform 1 0 22260 0 1 34586
box 0 0 1 1
use contact_30  contact_30_55
timestamp 1644949024
transform 1 0 1908 0 1 1726
box 0 0 1 1
use contact_30  contact_30_56
timestamp 1644949024
transform 1 0 22048 0 1 34586
box 0 0 1 1
use contact_30  contact_30_57
timestamp 1644949024
transform 1 0 22048 0 1 1938
box 0 0 1 1
use contact_30  contact_30_58
timestamp 1644949024
transform 1 0 22048 0 1 1514
box 0 0 1 1
use contact_30  contact_30_59
timestamp 1644949024
transform 1 0 1696 0 1 1938
box 0 0 1 1
use contact_30  contact_30_60
timestamp 1644949024
transform 1 0 1696 0 1 1514
box 0 0 1 1
use contact_30  contact_30_61
timestamp 1644949024
transform 1 0 1484 0 1 1726
box 0 0 1 1
use contact_30  contact_30_62
timestamp 1644949024
transform 1 0 22472 0 1 35010
box 0 0 1 1
use contact_30  contact_30_63
timestamp 1644949024
transform 1 0 22260 0 1 1514
box 0 0 1 1
use contact_30  contact_30_64
timestamp 1644949024
transform 1 0 1484 0 1 35010
box 0 0 1 1
use contact_30  contact_30_65
timestamp 1644949024
transform 1 0 1908 0 1 35010
box 0 0 1 1
use contact_30  contact_30_66
timestamp 1644949024
transform 1 0 22260 0 1 34798
box 0 0 1 1
use contact_30  contact_30_67
timestamp 1644949024
transform 1 0 1908 0 1 1938
box 0 0 1 1
use contact_30  contact_30_68
timestamp 1644949024
transform 1 0 22472 0 1 34586
box 0 0 1 1
use contact_30  contact_30_69
timestamp 1644949024
transform 1 0 1908 0 1 34586
box 0 0 1 1
use contact_30  contact_30_70
timestamp 1644949024
transform 1 0 22048 0 1 34798
box 0 0 1 1
use contact_30  contact_30_71
timestamp 1644949024
transform 1 0 22472 0 1 1938
box 0 0 1 1
use contact_28  contact_28_94
timestamp 1644949024
transform 1 0 17596 0 1 7450
box 0 0 1 1
use contact_28  contact_28_95
timestamp 1644949024
transform 1 0 18020 0 1 7026
box 0 0 1 1
use contact_28  contact_28_96
timestamp 1644949024
transform 1 0 18020 0 1 7450
box 0 0 1 1
use contact_28  contact_28_97
timestamp 1644949024
transform 1 0 6360 0 1 4270
box 0 0 1 1
use contact_28  contact_28_98
timestamp 1644949024
transform 1 0 16324 0 1 2786
box 0 0 1 1
use contact_28  contact_28_99
timestamp 1644949024
transform 1 0 14840 0 1 2786
box 0 0 1 1
use contact_28  contact_28_100
timestamp 1644949024
transform 1 0 13356 0 1 2786
box 0 0 1 1
use contact_28  contact_28_101
timestamp 1644949024
transform 1 0 11872 0 1 2786
box 0 0 1 1
use contact_18  contact_18_0
timestamp 1644949024
transform 1 0 8955 0 1 14081
box 0 0 1 1
use contact_18  contact_18_1
timestamp 1644949024
transform 1 0 8955 0 1 12897
box 0 0 1 1
use contact_18  contact_18_2
timestamp 1644949024
transform 1 0 8955 0 1 12405
box 0 0 1 1
use contact_18  contact_18_3
timestamp 1644949024
transform 1 0 8955 0 1 11221
box 0 0 1 1
use contact_18  contact_18_4
timestamp 1644949024
transform 1 0 8955 0 1 10729
box 0 0 1 1
use contact_18  contact_18_5
timestamp 1644949024
transform 1 0 8955 0 1 9545
box 0 0 1 1
use contact_18  contact_18_6
timestamp 1644949024
transform 1 0 18688 0 1 7555
box 0 0 1 1
use contact_18  contact_18_7
timestamp 1644949024
transform 1 0 18688 0 1 7555
box 0 0 1 1
use contact_18  contact_18_8
timestamp 1644949024
transform 1 0 18416 0 1 7555
box 0 0 1 1
use contact_18  contact_18_9
timestamp 1644949024
transform 1 0 18416 0 1 7555
box 0 0 1 1
use contact_18  contact_18_10
timestamp 1644949024
transform 1 0 17910 0 1 7555
box 0 0 1 1
use contact_18  contact_18_11
timestamp 1644949024
transform 1 0 17910 0 1 7555
box 0 0 1 1
use contact_18  contact_18_12
timestamp 1644949024
transform 1 0 17638 0 1 7555
box 0 0 1 1
use contact_18  contact_18_13
timestamp 1644949024
transform 1 0 17638 0 1 7555
box 0 0 1 1
use contact_18  contact_18_14
timestamp 1644949024
transform 1 0 16365 0 1 2859
box 0 0 1 1
use contact_18  contact_18_15
timestamp 1644949024
transform 1 0 14883 0 1 2859
box 0 0 1 1
use contact_18  contact_18_16
timestamp 1644949024
transform 1 0 13401 0 1 2859
box 0 0 1 1
use contact_18  contact_18_17
timestamp 1644949024
transform 1 0 11919 0 1 2859
box 0 0 1 1
use contact_18  contact_18_18
timestamp 1644949024
transform 1 0 6403 0 1 4356
box 0 0 1 1
use contact_18  contact_18_19
timestamp 1644949024
transform 1 0 2881 0 1 4571
box 0 0 1 1
use contact_18  contact_18_20
timestamp 1644949024
transform 1 0 2881 0 1 3387
box 0 0 1 1
use contact_18  contact_18_21
timestamp 1644949024
transform 1 0 10850 0 1 14085
box 0 0 1 1
use contact_18  contact_18_22
timestamp 1644949024
transform 1 0 10035 0 1 14085
box 0 0 1 1
use contact_18  contact_18_23
timestamp 1644949024
transform 1 0 10766 0 1 12893
box 0 0 1 1
use contact_18  contact_18_24
timestamp 1644949024
transform 1 0 10035 0 1 12893
box 0 0 1 1
use contact_18  contact_18_25
timestamp 1644949024
transform 1 0 10682 0 1 12409
box 0 0 1 1
use contact_18  contact_18_26
timestamp 1644949024
transform 1 0 10035 0 1 12409
box 0 0 1 1
use contact_18  contact_18_27
timestamp 1644949024
transform 1 0 10598 0 1 11217
box 0 0 1 1
use contact_18  contact_18_28
timestamp 1644949024
transform 1 0 10035 0 1 11217
box 0 0 1 1
use contact_18  contact_18_29
timestamp 1644949024
transform 1 0 10514 0 1 10733
box 0 0 1 1
use contact_18  contact_18_30
timestamp 1644949024
transform 1 0 10035 0 1 10733
box 0 0 1 1
use contact_18  contact_18_31
timestamp 1644949024
transform 1 0 10430 0 1 9541
box 0 0 1 1
use contact_18  contact_18_32
timestamp 1644949024
transform 1 0 10035 0 1 9541
box 0 0 1 1
use contact_18  contact_18_33
timestamp 1644949024
transform 1 0 15942 0 1 8630
box 0 0 1 1
use contact_18  contact_18_34
timestamp 1644949024
transform 1 0 10230 0 1 8630
box 0 0 1 1
use contact_18  contact_18_35
timestamp 1644949024
transform 1 0 20858 0 1 7708
box 0 0 1 1
use contact_18  contact_18_36
timestamp 1644949024
transform 1 0 10230 0 1 7708
box 0 0 1 1
use contact_18  contact_18_37
timestamp 1644949024
transform 1 0 17064 0 1 6958
box 0 0 1 1
use contact_18  contact_18_38
timestamp 1644949024
transform 1 0 10230 0 1 6958
box 0 0 1 1
use contact_26  contact_26_0
timestamp 1644949024
transform 1 0 8664 0 1 2921
box 0 0 1 1
use contact_26  contact_26_1
timestamp 1644949024
transform 1 0 8664 0 1 9607
box 0 0 1 1
use data_dff  data_dff_0
timestamp 1644949024
transform 1 0 11778 0 1 2650
box -39 -42 5928 916
use row_addr_dff  row_addr_dff_0
timestamp 1644949024
transform 1 0 8814 0 1 9336
box -39 -42 1482 6746
use control_logic_multiport  control_logic_multiport_0
timestamp 1644949024
transform 1 0 2740 0 1 3178
box -66 -42 7556 5906
use bank  bank_0
timestamp 1644949024
transform 1 0 10464 0 1 4952
box 0 0 10914 28960
<< labels >>
rlabel metal3 s 2880 3386 3012 3460 4 web
rlabel metal3 s 2880 4570 3012 4644 4 csb
rlabel metal4 s 6360 0 6512 364 4 clk
rlabel metal4 s 11872 0 12024 364 4 din0[0]
rlabel metal4 s 13356 0 13508 364 4 din0[1]
rlabel metal4 s 14840 0 14992 364 4 din0[2]
rlabel metal4 s 16324 0 16476 364 4 din0[3]
rlabel metal4 s 17596 0 17748 364 4 dout0[0]
rlabel metal3 s 17638 7554 17770 7628 4 dout1[0]
rlabel metal3 s 23744 6996 24108 7148 4 dout0[1]
rlabel metal3 s 17910 7554 18042 7628 4 dout1[1]
rlabel metal3 s 23744 7208 24108 7360 4 dout0[2]
rlabel metal3 s 18416 7554 18548 7628 4 dout1[2]
rlabel metal3 s 23744 7420 24108 7572 4 dout0[3]
rlabel metal3 s 18688 7554 18820 7628 4 dout1[3]
rlabel metal3 s 0 9752 364 9904 4 addr1[0]
rlabel metal3 s 0 10600 364 10752 4 addr1[1]
rlabel metal3 s 0 11024 364 11176 4 addr1[2]
rlabel metal3 s 0 12296 364 12448 4 addr1[3]
rlabel metal3 s 0 12720 364 12872 4 addr1[4]
rlabel metal3 s 0 13992 364 14144 4 addr1[5]
rlabel metal3 s 1484 1484 22624 2060 4 vdd
rlabel metal4 s 22048 1484 22624 35132 4 vdd
rlabel metal3 s 1484 34556 22624 35132 4 vdd
rlabel metal4 s 1484 1484 2060 35132 4 vdd
rlabel metal3 s 424 424 23684 1000 4 gnd
rlabel metal4 s 424 424 1000 36192 4 gnd
rlabel metal4 s 23108 424 23684 36192 4 gnd
rlabel metal3 s 424 35616 23684 36192 4 gnd
<< properties >>
string FIXED_BBOX 0 0 24108 36192
string GDS_FILE sram_0rw2r1w_4_16_sky130A.gds
string GDS_END 73180
string GDS_START 126
<< end >>
