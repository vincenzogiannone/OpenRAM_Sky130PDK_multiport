magic
tech sky130A
timestamp 1643678851
<< checkpaint >>
rect -630 -651 25526 25291
<< metal1 >>
rect 0 24304 24896 24318
rect 0 24241 24896 24255
rect 0 24128 24896 24142
rect 0 23598 24896 23612
rect 0 23485 24896 23499
rect 0 23422 24896 23436
rect 0 22764 24896 22778
rect 0 22701 24896 22715
rect 0 22588 24896 22602
rect 0 22058 24896 22072
rect 0 21945 24896 21959
rect 0 21882 24896 21896
rect 0 21224 24896 21238
rect 0 21161 24896 21175
rect 0 21048 24896 21062
rect 0 20518 24896 20532
rect 0 20405 24896 20419
rect 0 20342 24896 20356
rect 0 19684 24896 19698
rect 0 19621 24896 19635
rect 0 19508 24896 19522
rect 0 18978 24896 18992
rect 0 18865 24896 18879
rect 0 18802 24896 18816
rect 0 18144 24896 18158
rect 0 18081 24896 18095
rect 0 17968 24896 17982
rect 0 17438 24896 17452
rect 0 17325 24896 17339
rect 0 17262 24896 17276
rect 0 16604 24896 16618
rect 0 16541 24896 16555
rect 0 16428 24896 16442
rect 0 15898 24896 15912
rect 0 15785 24896 15799
rect 0 15722 24896 15736
rect 0 15064 24896 15078
rect 0 15001 24896 15015
rect 0 14888 24896 14902
rect 0 14358 24896 14372
rect 0 14245 24896 14259
rect 0 14182 24896 14196
rect 0 13524 24896 13538
rect 0 13461 24896 13475
rect 0 13348 24896 13362
rect 0 12818 24896 12832
rect 0 12705 24896 12719
rect 0 12642 24896 12656
rect 0 11984 24896 11998
rect 0 11921 24896 11935
rect 0 11808 24896 11822
rect 0 11278 24896 11292
rect 0 11165 24896 11179
rect 0 11102 24896 11116
rect 0 10444 24896 10458
rect 0 10381 24896 10395
rect 0 10268 24896 10282
rect 0 9738 24896 9752
rect 0 9625 24896 9639
rect 0 9562 24896 9576
rect 0 8904 24896 8918
rect 0 8841 24896 8855
rect 0 8728 24896 8742
rect 0 8198 24896 8212
rect 0 8085 24896 8099
rect 0 8022 24896 8036
rect 0 7364 24896 7378
rect 0 7301 24896 7315
rect 0 7188 24896 7202
rect 0 6658 24896 6672
rect 0 6545 24896 6559
rect 0 6482 24896 6496
rect 0 5824 24896 5838
rect 0 5761 24896 5775
rect 0 5648 24896 5662
rect 0 5118 24896 5132
rect 0 5005 24896 5019
rect 0 4942 24896 4956
rect 0 4284 24896 4298
rect 0 4221 24896 4235
rect 0 4108 24896 4122
rect 0 3578 24896 3592
rect 0 3465 24896 3479
rect 0 3402 24896 3416
rect 0 2744 24896 2758
rect 0 2681 24896 2695
rect 0 2568 24896 2582
rect 0 2038 24896 2052
rect 0 1925 24896 1939
rect 0 1862 24896 1876
rect 0 1204 24896 1218
rect 0 1141 24896 1155
rect 0 1028 24896 1042
rect 0 498 24896 512
rect 0 385 24896 399
rect 0 322 24896 336
<< metal2 >>
rect 96 0 110 24640
rect 222 0 236 24640
rect 313 0 327 24640
rect 485 0 499 24640
rect 611 0 625 24640
rect 702 0 716 24640
rect 874 0 888 24640
rect 1000 0 1014 24640
rect 1091 0 1105 24640
rect 1263 0 1277 24640
rect 1389 0 1403 24640
rect 1480 0 1494 24640
rect 1652 0 1666 24640
rect 1778 0 1792 24640
rect 1869 0 1883 24640
rect 2041 0 2055 24640
rect 2167 0 2181 24640
rect 2258 0 2272 24640
rect 2430 0 2444 24640
rect 2556 0 2570 24640
rect 2647 0 2661 24640
rect 2819 0 2833 24640
rect 2945 0 2959 24640
rect 3036 0 3050 24640
rect 3208 0 3222 24640
rect 3334 0 3348 24640
rect 3425 0 3439 24640
rect 3597 0 3611 24640
rect 3723 0 3737 24640
rect 3814 0 3828 24640
rect 3986 0 4000 24640
rect 4112 0 4126 24640
rect 4203 0 4217 24640
rect 4375 0 4389 24640
rect 4501 0 4515 24640
rect 4592 0 4606 24640
rect 4764 0 4778 24640
rect 4890 0 4904 24640
rect 4981 0 4995 24640
rect 5153 0 5167 24640
rect 5279 0 5293 24640
rect 5370 0 5384 24640
rect 5542 0 5556 24640
rect 5668 0 5682 24640
rect 5759 0 5773 24640
rect 5931 0 5945 24640
rect 6057 0 6071 24640
rect 6148 0 6162 24640
rect 6320 0 6334 24640
rect 6446 0 6460 24640
rect 6537 0 6551 24640
rect 6709 0 6723 24640
rect 6835 0 6849 24640
rect 6926 0 6940 24640
rect 7098 0 7112 24640
rect 7224 0 7238 24640
rect 7315 0 7329 24640
rect 7487 0 7501 24640
rect 7613 0 7627 24640
rect 7704 0 7718 24640
rect 7876 0 7890 24640
rect 8002 0 8016 24640
rect 8093 0 8107 24640
rect 8265 0 8279 24640
rect 8391 0 8405 24640
rect 8482 0 8496 24640
rect 8654 0 8668 24640
rect 8780 0 8794 24640
rect 8871 0 8885 24640
rect 9043 0 9057 24640
rect 9169 0 9183 24640
rect 9260 0 9274 24640
rect 9432 0 9446 24640
rect 9558 0 9572 24640
rect 9649 0 9663 24640
rect 9821 0 9835 24640
rect 9947 0 9961 24640
rect 10038 0 10052 24640
rect 10210 0 10224 24640
rect 10336 0 10350 24640
rect 10427 0 10441 24640
rect 10599 0 10613 24640
rect 10725 0 10739 24640
rect 10816 0 10830 24640
rect 10988 0 11002 24640
rect 11114 0 11128 24640
rect 11205 0 11219 24640
rect 11377 0 11391 24640
rect 11503 0 11517 24640
rect 11594 0 11608 24640
rect 11766 0 11780 24640
rect 11892 0 11906 24640
rect 11983 0 11997 24640
rect 12155 0 12169 24640
rect 12281 0 12295 24640
rect 12372 0 12386 24640
rect 12544 0 12558 24640
rect 12670 0 12684 24640
rect 12761 0 12775 24640
rect 12933 0 12947 24640
rect 13059 0 13073 24640
rect 13150 0 13164 24640
rect 13322 0 13336 24640
rect 13448 0 13462 24640
rect 13539 0 13553 24640
rect 13711 0 13725 24640
rect 13837 0 13851 24640
rect 13928 0 13942 24640
rect 14100 0 14114 24640
rect 14226 0 14240 24640
rect 14317 0 14331 24640
rect 14489 0 14503 24640
rect 14615 0 14629 24640
rect 14706 0 14720 24640
rect 14878 0 14892 24640
rect 15004 0 15018 24640
rect 15095 0 15109 24640
rect 15267 0 15281 24640
rect 15393 0 15407 24640
rect 15484 0 15498 24640
rect 15656 0 15670 24640
rect 15782 0 15796 24640
rect 15873 0 15887 24640
rect 16045 0 16059 24640
rect 16171 0 16185 24640
rect 16262 0 16276 24640
rect 16434 0 16448 24640
rect 16560 0 16574 24640
rect 16651 0 16665 24640
rect 16823 0 16837 24640
rect 16949 0 16963 24640
rect 17040 0 17054 24640
rect 17212 0 17226 24640
rect 17338 0 17352 24640
rect 17429 0 17443 24640
rect 17601 0 17615 24640
rect 17727 0 17741 24640
rect 17818 0 17832 24640
rect 17990 0 18004 24640
rect 18116 0 18130 24640
rect 18207 0 18221 24640
rect 18379 0 18393 24640
rect 18505 0 18519 24640
rect 18596 0 18610 24640
rect 18768 0 18782 24640
rect 18894 0 18908 24640
rect 18985 0 18999 24640
rect 19157 0 19171 24640
rect 19283 0 19297 24640
rect 19374 0 19388 24640
rect 19546 0 19560 24640
rect 19672 0 19686 24640
rect 19763 0 19777 24640
rect 19935 0 19949 24640
rect 20061 0 20075 24640
rect 20152 0 20166 24640
rect 20324 0 20338 24640
rect 20450 0 20464 24640
rect 20541 0 20555 24640
rect 20713 0 20727 24640
rect 20839 0 20853 24640
rect 20930 0 20944 24640
rect 21102 0 21116 24640
rect 21228 0 21242 24640
rect 21319 0 21333 24640
rect 21491 0 21505 24640
rect 21617 0 21631 24640
rect 21708 0 21722 24640
rect 21880 0 21894 24640
rect 22006 0 22020 24640
rect 22097 0 22111 24640
rect 22269 0 22283 24640
rect 22395 0 22409 24640
rect 22486 0 22500 24640
rect 22658 0 22672 24640
rect 22784 0 22798 24640
rect 22875 0 22889 24640
rect 23047 0 23061 24640
rect 23173 0 23187 24640
rect 23264 0 23278 24640
rect 23436 0 23450 24640
rect 23562 0 23576 24640
rect 23653 0 23667 24640
rect 23825 0 23839 24640
rect 23951 0 23965 24640
rect 24042 0 24056 24640
rect 24214 0 24228 24640
rect 24340 0 24354 24640
rect 24431 0 24445 24640
rect 24603 0 24617 24640
rect 24729 0 24743 24640
rect 24820 0 24834 24640
use bitcell_array  bitcell_array_0
timestamp 1643678851
transform 1 0 0 0 1 0
box 0 -21 24896 24661
<< labels >>
rlabel metal1 s 0 385 24896 399 4 rwl_0_0
rlabel metal1 s 0 498 24896 512 4 rwl_1_0
rlabel metal1 s 0 322 24896 336 4 wwl_0_0
rlabel metal1 s 0 1141 24896 1155 4 rwl_0_1
rlabel metal1 s 0 1028 24896 1042 4 rwl_1_1
rlabel metal1 s 0 1204 24896 1218 4 wwl_0_1
rlabel metal1 s 0 1925 24896 1939 4 rwl_0_2
rlabel metal1 s 0 2038 24896 2052 4 rwl_1_2
rlabel metal1 s 0 1862 24896 1876 4 wwl_0_2
rlabel metal1 s 0 2681 24896 2695 4 rwl_0_3
rlabel metal1 s 0 2568 24896 2582 4 rwl_1_3
rlabel metal1 s 0 2744 24896 2758 4 wwl_0_3
rlabel metal1 s 0 3465 24896 3479 4 rwl_0_4
rlabel metal1 s 0 3578 24896 3592 4 rwl_1_4
rlabel metal1 s 0 3402 24896 3416 4 wwl_0_4
rlabel metal1 s 0 4221 24896 4235 4 rwl_0_5
rlabel metal1 s 0 4108 24896 4122 4 rwl_1_5
rlabel metal1 s 0 4284 24896 4298 4 wwl_0_5
rlabel metal1 s 0 5005 24896 5019 4 rwl_0_6
rlabel metal1 s 0 5118 24896 5132 4 rwl_1_6
rlabel metal1 s 0 4942 24896 4956 4 wwl_0_6
rlabel metal1 s 0 5761 24896 5775 4 rwl_0_7
rlabel metal1 s 0 5648 24896 5662 4 rwl_1_7
rlabel metal1 s 0 5824 24896 5838 4 wwl_0_7
rlabel metal1 s 0 6545 24896 6559 4 rwl_0_8
rlabel metal1 s 0 6658 24896 6672 4 rwl_1_8
rlabel metal1 s 0 6482 24896 6496 4 wwl_0_8
rlabel metal1 s 0 7301 24896 7315 4 rwl_0_9
rlabel metal1 s 0 7188 24896 7202 4 rwl_1_9
rlabel metal1 s 0 7364 24896 7378 4 wwl_0_9
rlabel metal1 s 0 8085 24896 8099 4 rwl_0_10
rlabel metal1 s 0 8198 24896 8212 4 rwl_1_10
rlabel metal1 s 0 8022 24896 8036 4 wwl_0_10
rlabel metal1 s 0 8841 24896 8855 4 rwl_0_11
rlabel metal1 s 0 8728 24896 8742 4 rwl_1_11
rlabel metal1 s 0 8904 24896 8918 4 wwl_0_11
rlabel metal1 s 0 9625 24896 9639 4 rwl_0_12
rlabel metal1 s 0 9738 24896 9752 4 rwl_1_12
rlabel metal1 s 0 9562 24896 9576 4 wwl_0_12
rlabel metal1 s 0 10381 24896 10395 4 rwl_0_13
rlabel metal1 s 0 10268 24896 10282 4 rwl_1_13
rlabel metal1 s 0 10444 24896 10458 4 wwl_0_13
rlabel metal1 s 0 11165 24896 11179 4 rwl_0_14
rlabel metal1 s 0 11278 24896 11292 4 rwl_1_14
rlabel metal1 s 0 11102 24896 11116 4 wwl_0_14
rlabel metal1 s 0 11921 24896 11935 4 rwl_0_15
rlabel metal1 s 0 11808 24896 11822 4 rwl_1_15
rlabel metal1 s 0 11984 24896 11998 4 wwl_0_15
rlabel metal1 s 0 12705 24896 12719 4 rwl_0_16
rlabel metal1 s 0 12818 24896 12832 4 rwl_1_16
rlabel metal1 s 0 12642 24896 12656 4 wwl_0_16
rlabel metal1 s 0 13461 24896 13475 4 rwl_0_17
rlabel metal1 s 0 13348 24896 13362 4 rwl_1_17
rlabel metal1 s 0 13524 24896 13538 4 wwl_0_17
rlabel metal1 s 0 14245 24896 14259 4 rwl_0_18
rlabel metal1 s 0 14358 24896 14372 4 rwl_1_18
rlabel metal1 s 0 14182 24896 14196 4 wwl_0_18
rlabel metal1 s 0 15001 24896 15015 4 rwl_0_19
rlabel metal1 s 0 14888 24896 14902 4 rwl_1_19
rlabel metal1 s 0 15064 24896 15078 4 wwl_0_19
rlabel metal1 s 0 15785 24896 15799 4 rwl_0_20
rlabel metal1 s 0 15898 24896 15912 4 rwl_1_20
rlabel metal1 s 0 15722 24896 15736 4 wwl_0_20
rlabel metal1 s 0 16541 24896 16555 4 rwl_0_21
rlabel metal1 s 0 16428 24896 16442 4 rwl_1_21
rlabel metal1 s 0 16604 24896 16618 4 wwl_0_21
rlabel metal1 s 0 17325 24896 17339 4 rwl_0_22
rlabel metal1 s 0 17438 24896 17452 4 rwl_1_22
rlabel metal1 s 0 17262 24896 17276 4 wwl_0_22
rlabel metal1 s 0 18081 24896 18095 4 rwl_0_23
rlabel metal1 s 0 17968 24896 17982 4 rwl_1_23
rlabel metal1 s 0 18144 24896 18158 4 wwl_0_23
rlabel metal1 s 0 18865 24896 18879 4 rwl_0_24
rlabel metal1 s 0 18978 24896 18992 4 rwl_1_24
rlabel metal1 s 0 18802 24896 18816 4 wwl_0_24
rlabel metal1 s 0 19621 24896 19635 4 rwl_0_25
rlabel metal1 s 0 19508 24896 19522 4 rwl_1_25
rlabel metal1 s 0 19684 24896 19698 4 wwl_0_25
rlabel metal1 s 0 20405 24896 20419 4 rwl_0_26
rlabel metal1 s 0 20518 24896 20532 4 rwl_1_26
rlabel metal1 s 0 20342 24896 20356 4 wwl_0_26
rlabel metal1 s 0 21161 24896 21175 4 rwl_0_27
rlabel metal1 s 0 21048 24896 21062 4 rwl_1_27
rlabel metal1 s 0 21224 24896 21238 4 wwl_0_27
rlabel metal1 s 0 21945 24896 21959 4 rwl_0_28
rlabel metal1 s 0 22058 24896 22072 4 rwl_1_28
rlabel metal1 s 0 21882 24896 21896 4 wwl_0_28
rlabel metal1 s 0 22701 24896 22715 4 rwl_0_29
rlabel metal1 s 0 22588 24896 22602 4 rwl_1_29
rlabel metal1 s 0 22764 24896 22778 4 wwl_0_29
rlabel metal1 s 0 23485 24896 23499 4 rwl_0_30
rlabel metal1 s 0 23598 24896 23612 4 rwl_1_30
rlabel metal1 s 0 23422 24896 23436 4 wwl_0_30
rlabel metal1 s 0 24241 24896 24255 4 rwl_0_31
rlabel metal1 s 0 24128 24896 24142 4 rwl_1_31
rlabel metal1 s 0 24304 24896 24318 4 wwl_0_31
rlabel metal2 s 96 0 110 24640 4 read_bl_0_0
rlabel metal2 s 485 0 499 24640 4 read_bl_0_1
rlabel metal2 s 874 0 888 24640 4 read_bl_0_2
rlabel metal2 s 1263 0 1277 24640 4 read_bl_0_3
rlabel metal2 s 1652 0 1666 24640 4 read_bl_0_4
rlabel metal2 s 2041 0 2055 24640 4 read_bl_0_5
rlabel metal2 s 2430 0 2444 24640 4 read_bl_0_6
rlabel metal2 s 2819 0 2833 24640 4 read_bl_0_7
rlabel metal2 s 3208 0 3222 24640 4 read_bl_0_8
rlabel metal2 s 3597 0 3611 24640 4 read_bl_0_9
rlabel metal2 s 3986 0 4000 24640 4 read_bl_0_10
rlabel metal2 s 4375 0 4389 24640 4 read_bl_0_11
rlabel metal2 s 4764 0 4778 24640 4 read_bl_0_12
rlabel metal2 s 5153 0 5167 24640 4 read_bl_0_13
rlabel metal2 s 5542 0 5556 24640 4 read_bl_0_14
rlabel metal2 s 5931 0 5945 24640 4 read_bl_0_15
rlabel metal2 s 6320 0 6334 24640 4 read_bl_0_16
rlabel metal2 s 6709 0 6723 24640 4 read_bl_0_17
rlabel metal2 s 7098 0 7112 24640 4 read_bl_0_18
rlabel metal2 s 7487 0 7501 24640 4 read_bl_0_19
rlabel metal2 s 7876 0 7890 24640 4 read_bl_0_20
rlabel metal2 s 8265 0 8279 24640 4 read_bl_0_21
rlabel metal2 s 8654 0 8668 24640 4 read_bl_0_22
rlabel metal2 s 9043 0 9057 24640 4 read_bl_0_23
rlabel metal2 s 9432 0 9446 24640 4 read_bl_0_24
rlabel metal2 s 9821 0 9835 24640 4 read_bl_0_25
rlabel metal2 s 10210 0 10224 24640 4 read_bl_0_26
rlabel metal2 s 10599 0 10613 24640 4 read_bl_0_27
rlabel metal2 s 10988 0 11002 24640 4 read_bl_0_28
rlabel metal2 s 11377 0 11391 24640 4 read_bl_0_29
rlabel metal2 s 11766 0 11780 24640 4 read_bl_0_30
rlabel metal2 s 12155 0 12169 24640 4 read_bl_0_31
rlabel metal2 s 12544 0 12558 24640 4 read_bl_0_32
rlabel metal2 s 12933 0 12947 24640 4 read_bl_0_33
rlabel metal2 s 13322 0 13336 24640 4 read_bl_0_34
rlabel metal2 s 13711 0 13725 24640 4 read_bl_0_35
rlabel metal2 s 14100 0 14114 24640 4 read_bl_0_36
rlabel metal2 s 14489 0 14503 24640 4 read_bl_0_37
rlabel metal2 s 14878 0 14892 24640 4 read_bl_0_38
rlabel metal2 s 15267 0 15281 24640 4 read_bl_0_39
rlabel metal2 s 15656 0 15670 24640 4 read_bl_0_40
rlabel metal2 s 16045 0 16059 24640 4 read_bl_0_41
rlabel metal2 s 16434 0 16448 24640 4 read_bl_0_42
rlabel metal2 s 16823 0 16837 24640 4 read_bl_0_43
rlabel metal2 s 17212 0 17226 24640 4 read_bl_0_44
rlabel metal2 s 17601 0 17615 24640 4 read_bl_0_45
rlabel metal2 s 17990 0 18004 24640 4 read_bl_0_46
rlabel metal2 s 18379 0 18393 24640 4 read_bl_0_47
rlabel metal2 s 18768 0 18782 24640 4 read_bl_0_48
rlabel metal2 s 19157 0 19171 24640 4 read_bl_0_49
rlabel metal2 s 19546 0 19560 24640 4 read_bl_0_50
rlabel metal2 s 19935 0 19949 24640 4 read_bl_0_51
rlabel metal2 s 20324 0 20338 24640 4 read_bl_0_52
rlabel metal2 s 20713 0 20727 24640 4 read_bl_0_53
rlabel metal2 s 21102 0 21116 24640 4 read_bl_0_54
rlabel metal2 s 21491 0 21505 24640 4 read_bl_0_55
rlabel metal2 s 21880 0 21894 24640 4 read_bl_0_56
rlabel metal2 s 22269 0 22283 24640 4 read_bl_0_57
rlabel metal2 s 22658 0 22672 24640 4 read_bl_0_58
rlabel metal2 s 23047 0 23061 24640 4 read_bl_0_59
rlabel metal2 s 23436 0 23450 24640 4 read_bl_0_60
rlabel metal2 s 23825 0 23839 24640 4 read_bl_0_61
rlabel metal2 s 24214 0 24228 24640 4 read_bl_0_62
rlabel metal2 s 24603 0 24617 24640 4 read_bl_0_63
rlabel metal2 s 222 0 236 24640 4 read_bl_1_0
rlabel metal2 s 611 0 625 24640 4 read_bl_1_1
rlabel metal2 s 1000 0 1014 24640 4 read_bl_1_2
rlabel metal2 s 1389 0 1403 24640 4 read_bl_1_3
rlabel metal2 s 1778 0 1792 24640 4 read_bl_1_4
rlabel metal2 s 2167 0 2181 24640 4 read_bl_1_5
rlabel metal2 s 2556 0 2570 24640 4 read_bl_1_6
rlabel metal2 s 2945 0 2959 24640 4 read_bl_1_7
rlabel metal2 s 3334 0 3348 24640 4 read_bl_1_8
rlabel metal2 s 3723 0 3737 24640 4 read_bl_1_9
rlabel metal2 s 4112 0 4126 24640 4 read_bl_1_10
rlabel metal2 s 4501 0 4515 24640 4 read_bl_1_11
rlabel metal2 s 4890 0 4904 24640 4 read_bl_1_12
rlabel metal2 s 5279 0 5293 24640 4 read_bl_1_13
rlabel metal2 s 5668 0 5682 24640 4 read_bl_1_14
rlabel metal2 s 6057 0 6071 24640 4 read_bl_1_15
rlabel metal2 s 6446 0 6460 24640 4 read_bl_1_16
rlabel metal2 s 6835 0 6849 24640 4 read_bl_1_17
rlabel metal2 s 7224 0 7238 24640 4 read_bl_1_18
rlabel metal2 s 7613 0 7627 24640 4 read_bl_1_19
rlabel metal2 s 8002 0 8016 24640 4 read_bl_1_20
rlabel metal2 s 8391 0 8405 24640 4 read_bl_1_21
rlabel metal2 s 8780 0 8794 24640 4 read_bl_1_22
rlabel metal2 s 9169 0 9183 24640 4 read_bl_1_23
rlabel metal2 s 9558 0 9572 24640 4 read_bl_1_24
rlabel metal2 s 9947 0 9961 24640 4 read_bl_1_25
rlabel metal2 s 10336 0 10350 24640 4 read_bl_1_26
rlabel metal2 s 10725 0 10739 24640 4 read_bl_1_27
rlabel metal2 s 11114 0 11128 24640 4 read_bl_1_28
rlabel metal2 s 11503 0 11517 24640 4 read_bl_1_29
rlabel metal2 s 11892 0 11906 24640 4 read_bl_1_30
rlabel metal2 s 12281 0 12295 24640 4 read_bl_1_31
rlabel metal2 s 12670 0 12684 24640 4 read_bl_1_32
rlabel metal2 s 13059 0 13073 24640 4 read_bl_1_33
rlabel metal2 s 13448 0 13462 24640 4 read_bl_1_34
rlabel metal2 s 13837 0 13851 24640 4 read_bl_1_35
rlabel metal2 s 14226 0 14240 24640 4 read_bl_1_36
rlabel metal2 s 14615 0 14629 24640 4 read_bl_1_37
rlabel metal2 s 15004 0 15018 24640 4 read_bl_1_38
rlabel metal2 s 15393 0 15407 24640 4 read_bl_1_39
rlabel metal2 s 15782 0 15796 24640 4 read_bl_1_40
rlabel metal2 s 16171 0 16185 24640 4 read_bl_1_41
rlabel metal2 s 16560 0 16574 24640 4 read_bl_1_42
rlabel metal2 s 16949 0 16963 24640 4 read_bl_1_43
rlabel metal2 s 17338 0 17352 24640 4 read_bl_1_44
rlabel metal2 s 17727 0 17741 24640 4 read_bl_1_45
rlabel metal2 s 18116 0 18130 24640 4 read_bl_1_46
rlabel metal2 s 18505 0 18519 24640 4 read_bl_1_47
rlabel metal2 s 18894 0 18908 24640 4 read_bl_1_48
rlabel metal2 s 19283 0 19297 24640 4 read_bl_1_49
rlabel metal2 s 19672 0 19686 24640 4 read_bl_1_50
rlabel metal2 s 20061 0 20075 24640 4 read_bl_1_51
rlabel metal2 s 20450 0 20464 24640 4 read_bl_1_52
rlabel metal2 s 20839 0 20853 24640 4 read_bl_1_53
rlabel metal2 s 21228 0 21242 24640 4 read_bl_1_54
rlabel metal2 s 21617 0 21631 24640 4 read_bl_1_55
rlabel metal2 s 22006 0 22020 24640 4 read_bl_1_56
rlabel metal2 s 22395 0 22409 24640 4 read_bl_1_57
rlabel metal2 s 22784 0 22798 24640 4 read_bl_1_58
rlabel metal2 s 23173 0 23187 24640 4 read_bl_1_59
rlabel metal2 s 23562 0 23576 24640 4 read_bl_1_60
rlabel metal2 s 23951 0 23965 24640 4 read_bl_1_61
rlabel metal2 s 24340 0 24354 24640 4 read_bl_1_62
rlabel metal2 s 24729 0 24743 24640 4 read_bl_1_63
rlabel metal2 s 313 0 327 24640 4 write_bl_0_0
rlabel metal2 s 702 0 716 24640 4 write_bl_0_1
rlabel metal2 s 1091 0 1105 24640 4 write_bl_0_2
rlabel metal2 s 1480 0 1494 24640 4 write_bl_0_3
rlabel metal2 s 1869 0 1883 24640 4 write_bl_0_4
rlabel metal2 s 2258 0 2272 24640 4 write_bl_0_5
rlabel metal2 s 2647 0 2661 24640 4 write_bl_0_6
rlabel metal2 s 3036 0 3050 24640 4 write_bl_0_7
rlabel metal2 s 3425 0 3439 24640 4 write_bl_0_8
rlabel metal2 s 3814 0 3828 24640 4 write_bl_0_9
rlabel metal2 s 4203 0 4217 24640 4 write_bl_0_10
rlabel metal2 s 4592 0 4606 24640 4 write_bl_0_11
rlabel metal2 s 4981 0 4995 24640 4 write_bl_0_12
rlabel metal2 s 5370 0 5384 24640 4 write_bl_0_13
rlabel metal2 s 5759 0 5773 24640 4 write_bl_0_14
rlabel metal2 s 6148 0 6162 24640 4 write_bl_0_15
rlabel metal2 s 6537 0 6551 24640 4 write_bl_0_16
rlabel metal2 s 6926 0 6940 24640 4 write_bl_0_17
rlabel metal2 s 7315 0 7329 24640 4 write_bl_0_18
rlabel metal2 s 7704 0 7718 24640 4 write_bl_0_19
rlabel metal2 s 8093 0 8107 24640 4 write_bl_0_20
rlabel metal2 s 8482 0 8496 24640 4 write_bl_0_21
rlabel metal2 s 8871 0 8885 24640 4 write_bl_0_22
rlabel metal2 s 9260 0 9274 24640 4 write_bl_0_23
rlabel metal2 s 9649 0 9663 24640 4 write_bl_0_24
rlabel metal2 s 10038 0 10052 24640 4 write_bl_0_25
rlabel metal2 s 10427 0 10441 24640 4 write_bl_0_26
rlabel metal2 s 10816 0 10830 24640 4 write_bl_0_27
rlabel metal2 s 11205 0 11219 24640 4 write_bl_0_28
rlabel metal2 s 11594 0 11608 24640 4 write_bl_0_29
rlabel metal2 s 11983 0 11997 24640 4 write_bl_0_30
rlabel metal2 s 12372 0 12386 24640 4 write_bl_0_31
rlabel metal2 s 12761 0 12775 24640 4 write_bl_0_32
rlabel metal2 s 13150 0 13164 24640 4 write_bl_0_33
rlabel metal2 s 13539 0 13553 24640 4 write_bl_0_34
rlabel metal2 s 13928 0 13942 24640 4 write_bl_0_35
rlabel metal2 s 14317 0 14331 24640 4 write_bl_0_36
rlabel metal2 s 14706 0 14720 24640 4 write_bl_0_37
rlabel metal2 s 15095 0 15109 24640 4 write_bl_0_38
rlabel metal2 s 15484 0 15498 24640 4 write_bl_0_39
rlabel metal2 s 15873 0 15887 24640 4 write_bl_0_40
rlabel metal2 s 16262 0 16276 24640 4 write_bl_0_41
rlabel metal2 s 16651 0 16665 24640 4 write_bl_0_42
rlabel metal2 s 17040 0 17054 24640 4 write_bl_0_43
rlabel metal2 s 17429 0 17443 24640 4 write_bl_0_44
rlabel metal2 s 17818 0 17832 24640 4 write_bl_0_45
rlabel metal2 s 18207 0 18221 24640 4 write_bl_0_46
rlabel metal2 s 18596 0 18610 24640 4 write_bl_0_47
rlabel metal2 s 18985 0 18999 24640 4 write_bl_0_48
rlabel metal2 s 19374 0 19388 24640 4 write_bl_0_49
rlabel metal2 s 19763 0 19777 24640 4 write_bl_0_50
rlabel metal2 s 20152 0 20166 24640 4 write_bl_0_51
rlabel metal2 s 20541 0 20555 24640 4 write_bl_0_52
rlabel metal2 s 20930 0 20944 24640 4 write_bl_0_53
rlabel metal2 s 21319 0 21333 24640 4 write_bl_0_54
rlabel metal2 s 21708 0 21722 24640 4 write_bl_0_55
rlabel metal2 s 22097 0 22111 24640 4 write_bl_0_56
rlabel metal2 s 22486 0 22500 24640 4 write_bl_0_57
rlabel metal2 s 22875 0 22889 24640 4 write_bl_0_58
rlabel metal2 s 23264 0 23278 24640 4 write_bl_0_59
rlabel metal2 s 23653 0 23667 24640 4 write_bl_0_60
rlabel metal2 s 24042 0 24056 24640 4 write_bl_0_61
rlabel metal2 s 24431 0 24445 24640 4 write_bl_0_62
rlabel metal2 s 24820 0 24834 24640 4 write_bl_0_63
<< properties >>
string FIXED_BBOX 0 0 49792 49280
string GDS_FILE sram_0rw2r1w_16_128_sky130A.gds
string GDS_END 395154
string GDS_START 339382
<< end >>
