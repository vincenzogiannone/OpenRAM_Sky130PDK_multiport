magic
tech sky130A
timestamp 1643593061
<< checkpaint >>
rect -630 -630 631 631
<< properties >>
string GDS_FILE sram_0rw2r1w_2_16_sky130A.gds
string GDS_END 248896
string GDS_START 248444
<< end >>
