magic
tech sky130A
magscale 1 2
timestamp 1644951705
<< checkpaint >>
rect -1143 -1263 48601 2310
<< metal1 >>
rect 221 954 227 1006
rect 279 954 285 1006
rect 493 954 499 1006
rect 551 954 557 1006
rect 3333 954 3339 1006
rect 3391 954 3397 1006
rect 3605 954 3611 1006
rect 3663 954 3669 1006
rect 6445 954 6451 1006
rect 6503 954 6509 1006
rect 6717 954 6723 1006
rect 6775 954 6781 1006
rect 9557 954 9563 1006
rect 9615 954 9621 1006
rect 9829 954 9835 1006
rect 9887 954 9893 1006
rect 12669 954 12675 1006
rect 12727 954 12733 1006
rect 12941 954 12947 1006
rect 12999 954 13005 1006
rect 15781 954 15787 1006
rect 15839 954 15845 1006
rect 16053 954 16059 1006
rect 16111 954 16117 1006
rect 18893 954 18899 1006
rect 18951 954 18957 1006
rect 19165 954 19171 1006
rect 19223 954 19229 1006
rect 22005 954 22011 1006
rect 22063 954 22069 1006
rect 22277 954 22283 1006
rect 22335 954 22341 1006
rect 25117 954 25123 1006
rect 25175 954 25181 1006
rect 25389 954 25395 1006
rect 25447 954 25453 1006
rect 28229 954 28235 1006
rect 28287 954 28293 1006
rect 28501 954 28507 1006
rect 28559 954 28565 1006
rect 31341 954 31347 1006
rect 31399 954 31405 1006
rect 31613 954 31619 1006
rect 31671 954 31677 1006
rect 34453 954 34459 1006
rect 34511 954 34517 1006
rect 34725 954 34731 1006
rect 34783 954 34789 1006
rect 37565 954 37571 1006
rect 37623 954 37629 1006
rect 37837 954 37843 1006
rect 37895 954 37901 1006
rect 40677 954 40683 1006
rect 40735 954 40741 1006
rect 40949 954 40955 1006
rect 41007 954 41013 1006
rect 43789 954 43795 1006
rect 43847 954 43853 1006
rect 44061 954 44067 1006
rect 44119 954 44125 1006
rect 46901 954 46907 1006
rect 46959 954 46965 1006
rect 47173 954 47179 1006
rect 47231 954 47237 1006
rect 221 8 227 60
rect 279 8 285 60
rect 493 8 499 60
rect 551 8 557 60
rect 3333 8 3339 60
rect 3391 8 3397 60
rect 3605 8 3611 60
rect 3663 8 3669 60
rect 6445 8 6451 60
rect 6503 8 6509 60
rect 6717 8 6723 60
rect 6775 8 6781 60
rect 9557 8 9563 60
rect 9615 8 9621 60
rect 9829 8 9835 60
rect 9887 8 9893 60
rect 12669 8 12675 60
rect 12727 8 12733 60
rect 12941 8 12947 60
rect 12999 8 13005 60
rect 15781 8 15787 60
rect 15839 8 15845 60
rect 16053 8 16059 60
rect 16111 8 16117 60
rect 18893 8 18899 60
rect 18951 8 18957 60
rect 19165 8 19171 60
rect 19223 8 19229 60
rect 22005 8 22011 60
rect 22063 8 22069 60
rect 22277 8 22283 60
rect 22335 8 22341 60
rect 25117 8 25123 60
rect 25175 8 25181 60
rect 25389 8 25395 60
rect 25447 8 25453 60
rect 28229 8 28235 60
rect 28287 8 28293 60
rect 28501 8 28507 60
rect 28559 8 28565 60
rect 31341 8 31347 60
rect 31399 8 31405 60
rect 31613 8 31619 60
rect 31671 8 31677 60
rect 34453 8 34459 60
rect 34511 8 34517 60
rect 34725 8 34731 60
rect 34783 8 34789 60
rect 37565 8 37571 60
rect 37623 8 37629 60
rect 37837 8 37843 60
rect 37895 8 37901 60
rect 40677 8 40683 60
rect 40735 8 40741 60
rect 40949 8 40955 60
rect 41007 8 41013 60
rect 43789 8 43795 60
rect 43847 8 43853 60
rect 44061 8 44067 60
rect 44119 8 44125 60
rect 46901 8 46907 60
rect 46959 8 46965 60
rect 47173 8 47179 60
rect 47231 8 47237 60
<< via1 >>
rect 227 954 279 1006
rect 499 954 551 1006
rect 3339 954 3391 1006
rect 3611 954 3663 1006
rect 6451 954 6503 1006
rect 6723 954 6775 1006
rect 9563 954 9615 1006
rect 9835 954 9887 1006
rect 12675 954 12727 1006
rect 12947 954 12999 1006
rect 15787 954 15839 1006
rect 16059 954 16111 1006
rect 18899 954 18951 1006
rect 19171 954 19223 1006
rect 22011 954 22063 1006
rect 22283 954 22335 1006
rect 25123 954 25175 1006
rect 25395 954 25447 1006
rect 28235 954 28287 1006
rect 28507 954 28559 1006
rect 31347 954 31399 1006
rect 31619 954 31671 1006
rect 34459 954 34511 1006
rect 34731 954 34783 1006
rect 37571 954 37623 1006
rect 37843 954 37895 1006
rect 40683 954 40735 1006
rect 40955 954 41007 1006
rect 43795 954 43847 1006
rect 44067 954 44119 1006
rect 46907 954 46959 1006
rect 47179 954 47231 1006
rect 227 8 279 60
rect 499 8 551 60
rect 3339 8 3391 60
rect 3611 8 3663 60
rect 6451 8 6503 60
rect 6723 8 6775 60
rect 9563 8 9615 60
rect 9835 8 9887 60
rect 12675 8 12727 60
rect 12947 8 12999 60
rect 15787 8 15839 60
rect 16059 8 16111 60
rect 18899 8 18951 60
rect 19171 8 19223 60
rect 22011 8 22063 60
rect 22283 8 22335 60
rect 25123 8 25175 60
rect 25395 8 25447 60
rect 28235 8 28287 60
rect 28507 8 28559 60
rect 31347 8 31399 60
rect 31619 8 31671 60
rect 34459 8 34511 60
rect 34731 8 34783 60
rect 37571 8 37623 60
rect 37843 8 37895 60
rect 40683 8 40735 60
rect 40955 8 41007 60
rect 43795 8 43847 60
rect 44067 8 44119 60
rect 46907 8 46959 60
rect 47179 8 47231 60
<< metal2 >>
rect 225 1008 281 1017
rect 225 943 281 952
rect 497 1008 553 1017
rect 497 943 553 952
rect 3337 1008 3393 1017
rect 3337 943 3393 952
rect 3609 1008 3665 1017
rect 3609 943 3665 952
rect 6449 1008 6505 1017
rect 6449 943 6505 952
rect 6721 1008 6777 1017
rect 6721 943 6777 952
rect 9561 1008 9617 1017
rect 9561 943 9617 952
rect 9833 1008 9889 1017
rect 9833 943 9889 952
rect 12673 1008 12729 1017
rect 12673 943 12729 952
rect 12945 1008 13001 1017
rect 12945 943 13001 952
rect 15785 1008 15841 1017
rect 15785 943 15841 952
rect 16057 1008 16113 1017
rect 16057 943 16113 952
rect 18897 1008 18953 1017
rect 18897 943 18953 952
rect 19169 1008 19225 1017
rect 19169 943 19225 952
rect 22009 1008 22065 1017
rect 22009 943 22065 952
rect 22281 1008 22337 1017
rect 22281 943 22337 952
rect 25121 1008 25177 1017
rect 25121 943 25177 952
rect 25393 1008 25449 1017
rect 25393 943 25449 952
rect 28233 1008 28289 1017
rect 28233 943 28289 952
rect 28505 1008 28561 1017
rect 28505 943 28561 952
rect 31345 1008 31401 1017
rect 31345 943 31401 952
rect 31617 1008 31673 1017
rect 31617 943 31673 952
rect 34457 1008 34513 1017
rect 34457 943 34513 952
rect 34729 1008 34785 1017
rect 34729 943 34785 952
rect 37569 1008 37625 1017
rect 37569 943 37625 952
rect 37841 1008 37897 1017
rect 37841 943 37897 952
rect 40681 1008 40737 1017
rect 40681 943 40737 952
rect 40953 1008 41009 1017
rect 40953 943 41009 952
rect 43793 1008 43849 1017
rect 43793 943 43849 952
rect 44065 1008 44121 1017
rect 44065 943 44121 952
rect 46905 1008 46961 1017
rect 46905 943 46961 952
rect 47177 1008 47233 1017
rect 47177 943 47233 952
rect 131 0 159 240
rect 225 62 281 71
rect 225 -3 281 6
rect 319 0 347 240
rect 403 0 431 240
rect 497 62 553 71
rect 497 -3 553 6
rect 591 0 619 240
rect 3243 0 3271 240
rect 3337 62 3393 71
rect 3337 -3 3393 6
rect 3431 0 3459 240
rect 3515 0 3543 240
rect 3609 62 3665 71
rect 3609 -3 3665 6
rect 3703 0 3731 240
rect 6355 0 6383 240
rect 6449 62 6505 71
rect 6449 -3 6505 6
rect 6543 0 6571 240
rect 6627 0 6655 240
rect 6721 62 6777 71
rect 6721 -3 6777 6
rect 6815 0 6843 240
rect 9467 0 9495 240
rect 9561 62 9617 71
rect 9561 -3 9617 6
rect 9655 0 9683 240
rect 9739 0 9767 240
rect 9833 62 9889 71
rect 9833 -3 9889 6
rect 9927 0 9955 240
rect 12579 0 12607 240
rect 12673 62 12729 71
rect 12673 -3 12729 6
rect 12767 0 12795 240
rect 12851 0 12879 240
rect 12945 62 13001 71
rect 12945 -3 13001 6
rect 13039 0 13067 240
rect 15691 0 15719 240
rect 15785 62 15841 71
rect 15785 -3 15841 6
rect 15879 0 15907 240
rect 15963 0 15991 240
rect 16057 62 16113 71
rect 16057 -3 16113 6
rect 16151 0 16179 240
rect 18803 0 18831 240
rect 18897 62 18953 71
rect 18897 -3 18953 6
rect 18991 0 19019 240
rect 19075 0 19103 240
rect 19169 62 19225 71
rect 19169 -3 19225 6
rect 19263 0 19291 240
rect 21915 0 21943 240
rect 22009 62 22065 71
rect 22009 -3 22065 6
rect 22103 0 22131 240
rect 22187 0 22215 240
rect 22281 62 22337 71
rect 22281 -3 22337 6
rect 22375 0 22403 240
rect 25027 0 25055 240
rect 25121 62 25177 71
rect 25121 -3 25177 6
rect 25215 0 25243 240
rect 25299 0 25327 240
rect 25393 62 25449 71
rect 25393 -3 25449 6
rect 25487 0 25515 240
rect 28139 0 28167 240
rect 28233 62 28289 71
rect 28233 -3 28289 6
rect 28327 0 28355 240
rect 28411 0 28439 240
rect 28505 62 28561 71
rect 28505 -3 28561 6
rect 28599 0 28627 240
rect 31251 0 31279 240
rect 31345 62 31401 71
rect 31345 -3 31401 6
rect 31439 0 31467 240
rect 31523 0 31551 240
rect 31617 62 31673 71
rect 31617 -3 31673 6
rect 31711 0 31739 240
rect 34363 0 34391 240
rect 34457 62 34513 71
rect 34457 -3 34513 6
rect 34551 0 34579 240
rect 34635 0 34663 240
rect 34729 62 34785 71
rect 34729 -3 34785 6
rect 34823 0 34851 240
rect 37475 0 37503 240
rect 37569 62 37625 71
rect 37569 -3 37625 6
rect 37663 0 37691 240
rect 37747 0 37775 240
rect 37841 62 37897 71
rect 37841 -3 37897 6
rect 37935 0 37963 240
rect 40587 0 40615 240
rect 40681 62 40737 71
rect 40681 -3 40737 6
rect 40775 0 40803 240
rect 40859 0 40887 240
rect 40953 62 41009 71
rect 40953 -3 41009 6
rect 41047 0 41075 240
rect 43699 0 43727 240
rect 43793 62 43849 71
rect 43793 -3 43849 6
rect 43887 0 43915 240
rect 43971 0 43999 240
rect 44065 62 44121 71
rect 44065 -3 44121 6
rect 44159 0 44187 240
rect 46811 0 46839 240
rect 46905 62 46961 71
rect 46905 -3 46961 6
rect 46999 0 47027 240
rect 47083 0 47111 240
rect 47177 62 47233 71
rect 47177 -3 47233 6
rect 47271 0 47299 240
<< via2 >>
rect 225 1006 281 1008
rect 225 954 227 1006
rect 227 954 279 1006
rect 279 954 281 1006
rect 225 952 281 954
rect 497 1006 553 1008
rect 497 954 499 1006
rect 499 954 551 1006
rect 551 954 553 1006
rect 497 952 553 954
rect 3337 1006 3393 1008
rect 3337 954 3339 1006
rect 3339 954 3391 1006
rect 3391 954 3393 1006
rect 3337 952 3393 954
rect 3609 1006 3665 1008
rect 3609 954 3611 1006
rect 3611 954 3663 1006
rect 3663 954 3665 1006
rect 3609 952 3665 954
rect 6449 1006 6505 1008
rect 6449 954 6451 1006
rect 6451 954 6503 1006
rect 6503 954 6505 1006
rect 6449 952 6505 954
rect 6721 1006 6777 1008
rect 6721 954 6723 1006
rect 6723 954 6775 1006
rect 6775 954 6777 1006
rect 6721 952 6777 954
rect 9561 1006 9617 1008
rect 9561 954 9563 1006
rect 9563 954 9615 1006
rect 9615 954 9617 1006
rect 9561 952 9617 954
rect 9833 1006 9889 1008
rect 9833 954 9835 1006
rect 9835 954 9887 1006
rect 9887 954 9889 1006
rect 9833 952 9889 954
rect 12673 1006 12729 1008
rect 12673 954 12675 1006
rect 12675 954 12727 1006
rect 12727 954 12729 1006
rect 12673 952 12729 954
rect 12945 1006 13001 1008
rect 12945 954 12947 1006
rect 12947 954 12999 1006
rect 12999 954 13001 1006
rect 12945 952 13001 954
rect 15785 1006 15841 1008
rect 15785 954 15787 1006
rect 15787 954 15839 1006
rect 15839 954 15841 1006
rect 15785 952 15841 954
rect 16057 1006 16113 1008
rect 16057 954 16059 1006
rect 16059 954 16111 1006
rect 16111 954 16113 1006
rect 16057 952 16113 954
rect 18897 1006 18953 1008
rect 18897 954 18899 1006
rect 18899 954 18951 1006
rect 18951 954 18953 1006
rect 18897 952 18953 954
rect 19169 1006 19225 1008
rect 19169 954 19171 1006
rect 19171 954 19223 1006
rect 19223 954 19225 1006
rect 19169 952 19225 954
rect 22009 1006 22065 1008
rect 22009 954 22011 1006
rect 22011 954 22063 1006
rect 22063 954 22065 1006
rect 22009 952 22065 954
rect 22281 1006 22337 1008
rect 22281 954 22283 1006
rect 22283 954 22335 1006
rect 22335 954 22337 1006
rect 22281 952 22337 954
rect 25121 1006 25177 1008
rect 25121 954 25123 1006
rect 25123 954 25175 1006
rect 25175 954 25177 1006
rect 25121 952 25177 954
rect 25393 1006 25449 1008
rect 25393 954 25395 1006
rect 25395 954 25447 1006
rect 25447 954 25449 1006
rect 25393 952 25449 954
rect 28233 1006 28289 1008
rect 28233 954 28235 1006
rect 28235 954 28287 1006
rect 28287 954 28289 1006
rect 28233 952 28289 954
rect 28505 1006 28561 1008
rect 28505 954 28507 1006
rect 28507 954 28559 1006
rect 28559 954 28561 1006
rect 28505 952 28561 954
rect 31345 1006 31401 1008
rect 31345 954 31347 1006
rect 31347 954 31399 1006
rect 31399 954 31401 1006
rect 31345 952 31401 954
rect 31617 1006 31673 1008
rect 31617 954 31619 1006
rect 31619 954 31671 1006
rect 31671 954 31673 1006
rect 31617 952 31673 954
rect 34457 1006 34513 1008
rect 34457 954 34459 1006
rect 34459 954 34511 1006
rect 34511 954 34513 1006
rect 34457 952 34513 954
rect 34729 1006 34785 1008
rect 34729 954 34731 1006
rect 34731 954 34783 1006
rect 34783 954 34785 1006
rect 34729 952 34785 954
rect 37569 1006 37625 1008
rect 37569 954 37571 1006
rect 37571 954 37623 1006
rect 37623 954 37625 1006
rect 37569 952 37625 954
rect 37841 1006 37897 1008
rect 37841 954 37843 1006
rect 37843 954 37895 1006
rect 37895 954 37897 1006
rect 37841 952 37897 954
rect 40681 1006 40737 1008
rect 40681 954 40683 1006
rect 40683 954 40735 1006
rect 40735 954 40737 1006
rect 40681 952 40737 954
rect 40953 1006 41009 1008
rect 40953 954 40955 1006
rect 40955 954 41007 1006
rect 41007 954 41009 1006
rect 40953 952 41009 954
rect 43793 1006 43849 1008
rect 43793 954 43795 1006
rect 43795 954 43847 1006
rect 43847 954 43849 1006
rect 43793 952 43849 954
rect 44065 1006 44121 1008
rect 44065 954 44067 1006
rect 44067 954 44119 1006
rect 44119 954 44121 1006
rect 44065 952 44121 954
rect 46905 1006 46961 1008
rect 46905 954 46907 1006
rect 46907 954 46959 1006
rect 46959 954 46961 1006
rect 46905 952 46961 954
rect 47177 1006 47233 1008
rect 47177 954 47179 1006
rect 47179 954 47231 1006
rect 47231 954 47233 1006
rect 47177 952 47233 954
rect 225 60 281 62
rect 225 8 227 60
rect 227 8 279 60
rect 279 8 281 60
rect 225 6 281 8
rect 497 60 553 62
rect 497 8 499 60
rect 499 8 551 60
rect 551 8 553 60
rect 497 6 553 8
rect 3337 60 3393 62
rect 3337 8 3339 60
rect 3339 8 3391 60
rect 3391 8 3393 60
rect 3337 6 3393 8
rect 3609 60 3665 62
rect 3609 8 3611 60
rect 3611 8 3663 60
rect 3663 8 3665 60
rect 3609 6 3665 8
rect 6449 60 6505 62
rect 6449 8 6451 60
rect 6451 8 6503 60
rect 6503 8 6505 60
rect 6449 6 6505 8
rect 6721 60 6777 62
rect 6721 8 6723 60
rect 6723 8 6775 60
rect 6775 8 6777 60
rect 6721 6 6777 8
rect 9561 60 9617 62
rect 9561 8 9563 60
rect 9563 8 9615 60
rect 9615 8 9617 60
rect 9561 6 9617 8
rect 9833 60 9889 62
rect 9833 8 9835 60
rect 9835 8 9887 60
rect 9887 8 9889 60
rect 9833 6 9889 8
rect 12673 60 12729 62
rect 12673 8 12675 60
rect 12675 8 12727 60
rect 12727 8 12729 60
rect 12673 6 12729 8
rect 12945 60 13001 62
rect 12945 8 12947 60
rect 12947 8 12999 60
rect 12999 8 13001 60
rect 12945 6 13001 8
rect 15785 60 15841 62
rect 15785 8 15787 60
rect 15787 8 15839 60
rect 15839 8 15841 60
rect 15785 6 15841 8
rect 16057 60 16113 62
rect 16057 8 16059 60
rect 16059 8 16111 60
rect 16111 8 16113 60
rect 16057 6 16113 8
rect 18897 60 18953 62
rect 18897 8 18899 60
rect 18899 8 18951 60
rect 18951 8 18953 60
rect 18897 6 18953 8
rect 19169 60 19225 62
rect 19169 8 19171 60
rect 19171 8 19223 60
rect 19223 8 19225 60
rect 19169 6 19225 8
rect 22009 60 22065 62
rect 22009 8 22011 60
rect 22011 8 22063 60
rect 22063 8 22065 60
rect 22009 6 22065 8
rect 22281 60 22337 62
rect 22281 8 22283 60
rect 22283 8 22335 60
rect 22335 8 22337 60
rect 22281 6 22337 8
rect 25121 60 25177 62
rect 25121 8 25123 60
rect 25123 8 25175 60
rect 25175 8 25177 60
rect 25121 6 25177 8
rect 25393 60 25449 62
rect 25393 8 25395 60
rect 25395 8 25447 60
rect 25447 8 25449 60
rect 25393 6 25449 8
rect 28233 60 28289 62
rect 28233 8 28235 60
rect 28235 8 28287 60
rect 28287 8 28289 60
rect 28233 6 28289 8
rect 28505 60 28561 62
rect 28505 8 28507 60
rect 28507 8 28559 60
rect 28559 8 28561 60
rect 28505 6 28561 8
rect 31345 60 31401 62
rect 31345 8 31347 60
rect 31347 8 31399 60
rect 31399 8 31401 60
rect 31345 6 31401 8
rect 31617 60 31673 62
rect 31617 8 31619 60
rect 31619 8 31671 60
rect 31671 8 31673 60
rect 31617 6 31673 8
rect 34457 60 34513 62
rect 34457 8 34459 60
rect 34459 8 34511 60
rect 34511 8 34513 60
rect 34457 6 34513 8
rect 34729 60 34785 62
rect 34729 8 34731 60
rect 34731 8 34783 60
rect 34783 8 34785 60
rect 34729 6 34785 8
rect 37569 60 37625 62
rect 37569 8 37571 60
rect 37571 8 37623 60
rect 37623 8 37625 60
rect 37569 6 37625 8
rect 37841 60 37897 62
rect 37841 8 37843 60
rect 37843 8 37895 60
rect 37895 8 37897 60
rect 37841 6 37897 8
rect 40681 60 40737 62
rect 40681 8 40683 60
rect 40683 8 40735 60
rect 40735 8 40737 60
rect 40681 6 40737 8
rect 40953 60 41009 62
rect 40953 8 40955 60
rect 40955 8 41007 60
rect 41007 8 41009 60
rect 40953 6 41009 8
rect 43793 60 43849 62
rect 43793 8 43795 60
rect 43795 8 43847 60
rect 43847 8 43849 60
rect 43793 6 43849 8
rect 44065 60 44121 62
rect 44065 8 44067 60
rect 44067 8 44119 60
rect 44119 8 44121 60
rect 44065 6 44121 8
rect 46905 60 46961 62
rect 46905 8 46907 60
rect 46907 8 46959 60
rect 46959 8 46961 60
rect 46905 6 46961 8
rect 47177 60 47233 62
rect 47177 8 47179 60
rect 47179 8 47231 60
rect 47231 8 47233 60
rect 47177 6 47233 8
<< metal3 >>
rect 187 1008 319 1017
rect 187 952 225 1008
rect 281 952 319 1008
rect 187 943 319 952
rect 459 1008 591 1017
rect 459 952 497 1008
rect 553 952 591 1008
rect 459 943 591 952
rect 3299 1008 3431 1017
rect 3299 952 3337 1008
rect 3393 952 3431 1008
rect 3299 943 3431 952
rect 3571 1008 3703 1017
rect 3571 952 3609 1008
rect 3665 952 3703 1008
rect 3571 943 3703 952
rect 6411 1008 6543 1017
rect 6411 952 6449 1008
rect 6505 952 6543 1008
rect 6411 943 6543 952
rect 6683 1008 6815 1017
rect 6683 952 6721 1008
rect 6777 952 6815 1008
rect 6683 943 6815 952
rect 9523 1008 9655 1017
rect 9523 952 9561 1008
rect 9617 952 9655 1008
rect 9523 943 9655 952
rect 9795 1008 9927 1017
rect 9795 952 9833 1008
rect 9889 952 9927 1008
rect 9795 943 9927 952
rect 12635 1008 12767 1017
rect 12635 952 12673 1008
rect 12729 952 12767 1008
rect 12635 943 12767 952
rect 12907 1008 13039 1017
rect 12907 952 12945 1008
rect 13001 952 13039 1008
rect 12907 943 13039 952
rect 15747 1008 15879 1017
rect 15747 952 15785 1008
rect 15841 952 15879 1008
rect 15747 943 15879 952
rect 16019 1008 16151 1017
rect 16019 952 16057 1008
rect 16113 952 16151 1008
rect 16019 943 16151 952
rect 18859 1008 18991 1017
rect 18859 952 18897 1008
rect 18953 952 18991 1008
rect 18859 943 18991 952
rect 19131 1008 19263 1017
rect 19131 952 19169 1008
rect 19225 952 19263 1008
rect 19131 943 19263 952
rect 21971 1008 22103 1017
rect 21971 952 22009 1008
rect 22065 952 22103 1008
rect 21971 943 22103 952
rect 22243 1008 22375 1017
rect 22243 952 22281 1008
rect 22337 952 22375 1008
rect 22243 943 22375 952
rect 25083 1008 25215 1017
rect 25083 952 25121 1008
rect 25177 952 25215 1008
rect 25083 943 25215 952
rect 25355 1008 25487 1017
rect 25355 952 25393 1008
rect 25449 952 25487 1008
rect 25355 943 25487 952
rect 28195 1008 28327 1017
rect 28195 952 28233 1008
rect 28289 952 28327 1008
rect 28195 943 28327 952
rect 28467 1008 28599 1017
rect 28467 952 28505 1008
rect 28561 952 28599 1008
rect 28467 943 28599 952
rect 31307 1008 31439 1017
rect 31307 952 31345 1008
rect 31401 952 31439 1008
rect 31307 943 31439 952
rect 31579 1008 31711 1017
rect 31579 952 31617 1008
rect 31673 952 31711 1008
rect 31579 943 31711 952
rect 34419 1008 34551 1017
rect 34419 952 34457 1008
rect 34513 952 34551 1008
rect 34419 943 34551 952
rect 34691 1008 34823 1017
rect 34691 952 34729 1008
rect 34785 952 34823 1008
rect 34691 943 34823 952
rect 37531 1008 37663 1017
rect 37531 952 37569 1008
rect 37625 952 37663 1008
rect 37531 943 37663 952
rect 37803 1008 37935 1017
rect 37803 952 37841 1008
rect 37897 952 37935 1008
rect 37803 943 37935 952
rect 40643 1008 40775 1017
rect 40643 952 40681 1008
rect 40737 952 40775 1008
rect 40643 943 40775 952
rect 40915 1008 41047 1017
rect 40915 952 40953 1008
rect 41009 952 41047 1008
rect 40915 943 41047 952
rect 43755 1008 43887 1017
rect 43755 952 43793 1008
rect 43849 952 43887 1008
rect 43755 943 43887 952
rect 44027 1008 44159 1017
rect 44027 952 44065 1008
rect 44121 952 44159 1008
rect 44027 943 44159 952
rect 46867 1008 46999 1017
rect 46867 952 46905 1008
rect 46961 952 46999 1008
rect 46867 943 46999 952
rect 47139 1008 47271 1017
rect 47139 952 47177 1008
rect 47233 952 47271 1008
rect 47139 943 47271 952
rect 187 62 319 71
rect 187 6 225 62
rect 281 6 319 62
rect 187 -3 319 6
rect 459 62 591 71
rect 459 6 497 62
rect 553 6 591 62
rect 459 -3 591 6
rect 3299 62 3431 71
rect 3299 6 3337 62
rect 3393 6 3431 62
rect 3299 -3 3431 6
rect 3571 62 3703 71
rect 3571 6 3609 62
rect 3665 6 3703 62
rect 3571 -3 3703 6
rect 6411 62 6543 71
rect 6411 6 6449 62
rect 6505 6 6543 62
rect 6411 -3 6543 6
rect 6683 62 6815 71
rect 6683 6 6721 62
rect 6777 6 6815 62
rect 6683 -3 6815 6
rect 9523 62 9655 71
rect 9523 6 9561 62
rect 9617 6 9655 62
rect 9523 -3 9655 6
rect 9795 62 9927 71
rect 9795 6 9833 62
rect 9889 6 9927 62
rect 9795 -3 9927 6
rect 12635 62 12767 71
rect 12635 6 12673 62
rect 12729 6 12767 62
rect 12635 -3 12767 6
rect 12907 62 13039 71
rect 12907 6 12945 62
rect 13001 6 13039 62
rect 12907 -3 13039 6
rect 15747 62 15879 71
rect 15747 6 15785 62
rect 15841 6 15879 62
rect 15747 -3 15879 6
rect 16019 62 16151 71
rect 16019 6 16057 62
rect 16113 6 16151 62
rect 16019 -3 16151 6
rect 18859 62 18991 71
rect 18859 6 18897 62
rect 18953 6 18991 62
rect 18859 -3 18991 6
rect 19131 62 19263 71
rect 19131 6 19169 62
rect 19225 6 19263 62
rect 19131 -3 19263 6
rect 21971 62 22103 71
rect 21971 6 22009 62
rect 22065 6 22103 62
rect 21971 -3 22103 6
rect 22243 62 22375 71
rect 22243 6 22281 62
rect 22337 6 22375 62
rect 22243 -3 22375 6
rect 25083 62 25215 71
rect 25083 6 25121 62
rect 25177 6 25215 62
rect 25083 -3 25215 6
rect 25355 62 25487 71
rect 25355 6 25393 62
rect 25449 6 25487 62
rect 25355 -3 25487 6
rect 28195 62 28327 71
rect 28195 6 28233 62
rect 28289 6 28327 62
rect 28195 -3 28327 6
rect 28467 62 28599 71
rect 28467 6 28505 62
rect 28561 6 28599 62
rect 28467 -3 28599 6
rect 31307 62 31439 71
rect 31307 6 31345 62
rect 31401 6 31439 62
rect 31307 -3 31439 6
rect 31579 62 31711 71
rect 31579 6 31617 62
rect 31673 6 31711 62
rect 31579 -3 31711 6
rect 34419 62 34551 71
rect 34419 6 34457 62
rect 34513 6 34551 62
rect 34419 -3 34551 6
rect 34691 62 34823 71
rect 34691 6 34729 62
rect 34785 6 34823 62
rect 34691 -3 34823 6
rect 37531 62 37663 71
rect 37531 6 37569 62
rect 37625 6 37663 62
rect 37531 -3 37663 6
rect 37803 62 37935 71
rect 37803 6 37841 62
rect 37897 6 37935 62
rect 37803 -3 37935 6
rect 40643 62 40775 71
rect 40643 6 40681 62
rect 40737 6 40775 62
rect 40643 -3 40775 6
rect 40915 62 41047 71
rect 40915 6 40953 62
rect 41009 6 41047 62
rect 40915 -3 41047 6
rect 43755 62 43887 71
rect 43755 6 43793 62
rect 43849 6 43887 62
rect 43755 -3 43887 6
rect 44027 62 44159 71
rect 44027 6 44065 62
rect 44121 6 44159 62
rect 44027 -3 44159 6
rect 46867 62 46999 71
rect 46867 6 46905 62
rect 46961 6 46999 62
rect 46867 -3 46999 6
rect 47139 62 47271 71
rect 47139 6 47177 62
rect 47233 6 47271 62
rect 47139 -3 47271 6
use contact_18  contact_18_0
timestamp 1644951705
transform 1 0 47139 0 1 943
box 0 0 1 1
use contact_17  contact_17_0
timestamp 1644951705
transform 1 0 47173 0 1 948
box 0 0 1 1
use contact_18  contact_18_1
timestamp 1644951705
transform 1 0 47139 0 1 -3
box 0 0 1 1
use contact_17  contact_17_1
timestamp 1644951705
transform 1 0 47173 0 1 2
box 0 0 1 1
use contact_18  contact_18_2
timestamp 1644951705
transform 1 0 46867 0 1 943
box 0 0 1 1
use contact_17  contact_17_2
timestamp 1644951705
transform 1 0 46901 0 1 948
box 0 0 1 1
use contact_18  contact_18_3
timestamp 1644951705
transform 1 0 46867 0 1 -3
box 0 0 1 1
use contact_17  contact_17_3
timestamp 1644951705
transform 1 0 46901 0 1 2
box 0 0 1 1
use contact_18  contact_18_4
timestamp 1644951705
transform 1 0 44027 0 1 943
box 0 0 1 1
use contact_17  contact_17_4
timestamp 1644951705
transform 1 0 44061 0 1 948
box 0 0 1 1
use contact_18  contact_18_5
timestamp 1644951705
transform 1 0 44027 0 1 -3
box 0 0 1 1
use contact_17  contact_17_5
timestamp 1644951705
transform 1 0 44061 0 1 2
box 0 0 1 1
use contact_18  contact_18_6
timestamp 1644951705
transform 1 0 43755 0 1 943
box 0 0 1 1
use contact_17  contact_17_6
timestamp 1644951705
transform 1 0 43789 0 1 948
box 0 0 1 1
use contact_18  contact_18_7
timestamp 1644951705
transform 1 0 43755 0 1 -3
box 0 0 1 1
use contact_17  contact_17_7
timestamp 1644951705
transform 1 0 43789 0 1 2
box 0 0 1 1
use contact_18  contact_18_8
timestamp 1644951705
transform 1 0 40915 0 1 943
box 0 0 1 1
use contact_17  contact_17_8
timestamp 1644951705
transform 1 0 40949 0 1 948
box 0 0 1 1
use contact_18  contact_18_9
timestamp 1644951705
transform 1 0 40915 0 1 -3
box 0 0 1 1
use contact_17  contact_17_9
timestamp 1644951705
transform 1 0 40949 0 1 2
box 0 0 1 1
use contact_18  contact_18_10
timestamp 1644951705
transform 1 0 40643 0 1 943
box 0 0 1 1
use contact_17  contact_17_10
timestamp 1644951705
transform 1 0 40677 0 1 948
box 0 0 1 1
use contact_18  contact_18_11
timestamp 1644951705
transform 1 0 40643 0 1 -3
box 0 0 1 1
use contact_17  contact_17_11
timestamp 1644951705
transform 1 0 40677 0 1 2
box 0 0 1 1
use contact_18  contact_18_12
timestamp 1644951705
transform 1 0 37803 0 1 943
box 0 0 1 1
use contact_17  contact_17_12
timestamp 1644951705
transform 1 0 37837 0 1 948
box 0 0 1 1
use contact_18  contact_18_13
timestamp 1644951705
transform 1 0 37803 0 1 -3
box 0 0 1 1
use contact_17  contact_17_13
timestamp 1644951705
transform 1 0 37837 0 1 2
box 0 0 1 1
use contact_18  contact_18_14
timestamp 1644951705
transform 1 0 37531 0 1 943
box 0 0 1 1
use contact_17  contact_17_14
timestamp 1644951705
transform 1 0 37565 0 1 948
box 0 0 1 1
use contact_18  contact_18_15
timestamp 1644951705
transform 1 0 37531 0 1 -3
box 0 0 1 1
use contact_17  contact_17_15
timestamp 1644951705
transform 1 0 37565 0 1 2
box 0 0 1 1
use contact_18  contact_18_16
timestamp 1644951705
transform 1 0 34691 0 1 943
box 0 0 1 1
use contact_17  contact_17_16
timestamp 1644951705
transform 1 0 34725 0 1 948
box 0 0 1 1
use contact_18  contact_18_17
timestamp 1644951705
transform 1 0 34691 0 1 -3
box 0 0 1 1
use contact_17  contact_17_17
timestamp 1644951705
transform 1 0 34725 0 1 2
box 0 0 1 1
use contact_18  contact_18_18
timestamp 1644951705
transform 1 0 34419 0 1 943
box 0 0 1 1
use contact_17  contact_17_18
timestamp 1644951705
transform 1 0 34453 0 1 948
box 0 0 1 1
use contact_18  contact_18_19
timestamp 1644951705
transform 1 0 34419 0 1 -3
box 0 0 1 1
use contact_17  contact_17_19
timestamp 1644951705
transform 1 0 34453 0 1 2
box 0 0 1 1
use contact_18  contact_18_20
timestamp 1644951705
transform 1 0 31579 0 1 943
box 0 0 1 1
use contact_17  contact_17_20
timestamp 1644951705
transform 1 0 31613 0 1 948
box 0 0 1 1
use contact_18  contact_18_21
timestamp 1644951705
transform 1 0 31579 0 1 -3
box 0 0 1 1
use contact_17  contact_17_21
timestamp 1644951705
transform 1 0 31613 0 1 2
box 0 0 1 1
use contact_18  contact_18_22
timestamp 1644951705
transform 1 0 31307 0 1 943
box 0 0 1 1
use contact_17  contact_17_22
timestamp 1644951705
transform 1 0 31341 0 1 948
box 0 0 1 1
use contact_18  contact_18_23
timestamp 1644951705
transform 1 0 31307 0 1 -3
box 0 0 1 1
use contact_17  contact_17_23
timestamp 1644951705
transform 1 0 31341 0 1 2
box 0 0 1 1
use contact_18  contact_18_24
timestamp 1644951705
transform 1 0 28467 0 1 943
box 0 0 1 1
use contact_17  contact_17_24
timestamp 1644951705
transform 1 0 28501 0 1 948
box 0 0 1 1
use contact_18  contact_18_25
timestamp 1644951705
transform 1 0 28467 0 1 -3
box 0 0 1 1
use contact_17  contact_17_25
timestamp 1644951705
transform 1 0 28501 0 1 2
box 0 0 1 1
use contact_18  contact_18_26
timestamp 1644951705
transform 1 0 28195 0 1 943
box 0 0 1 1
use contact_17  contact_17_26
timestamp 1644951705
transform 1 0 28229 0 1 948
box 0 0 1 1
use contact_18  contact_18_27
timestamp 1644951705
transform 1 0 28195 0 1 -3
box 0 0 1 1
use contact_17  contact_17_27
timestamp 1644951705
transform 1 0 28229 0 1 2
box 0 0 1 1
use contact_18  contact_18_28
timestamp 1644951705
transform 1 0 25355 0 1 943
box 0 0 1 1
use contact_17  contact_17_28
timestamp 1644951705
transform 1 0 25389 0 1 948
box 0 0 1 1
use contact_18  contact_18_29
timestamp 1644951705
transform 1 0 25355 0 1 -3
box 0 0 1 1
use contact_17  contact_17_29
timestamp 1644951705
transform 1 0 25389 0 1 2
box 0 0 1 1
use contact_18  contact_18_30
timestamp 1644951705
transform 1 0 25083 0 1 943
box 0 0 1 1
use contact_17  contact_17_30
timestamp 1644951705
transform 1 0 25117 0 1 948
box 0 0 1 1
use contact_18  contact_18_31
timestamp 1644951705
transform 1 0 25083 0 1 -3
box 0 0 1 1
use contact_17  contact_17_31
timestamp 1644951705
transform 1 0 25117 0 1 2
box 0 0 1 1
use contact_18  contact_18_32
timestamp 1644951705
transform 1 0 22243 0 1 943
box 0 0 1 1
use contact_17  contact_17_32
timestamp 1644951705
transform 1 0 22277 0 1 948
box 0 0 1 1
use contact_18  contact_18_33
timestamp 1644951705
transform 1 0 22243 0 1 -3
box 0 0 1 1
use contact_17  contact_17_33
timestamp 1644951705
transform 1 0 22277 0 1 2
box 0 0 1 1
use contact_18  contact_18_34
timestamp 1644951705
transform 1 0 21971 0 1 943
box 0 0 1 1
use contact_17  contact_17_34
timestamp 1644951705
transform 1 0 22005 0 1 948
box 0 0 1 1
use contact_18  contact_18_35
timestamp 1644951705
transform 1 0 21971 0 1 -3
box 0 0 1 1
use contact_17  contact_17_35
timestamp 1644951705
transform 1 0 22005 0 1 2
box 0 0 1 1
use contact_18  contact_18_36
timestamp 1644951705
transform 1 0 19131 0 1 943
box 0 0 1 1
use contact_17  contact_17_36
timestamp 1644951705
transform 1 0 19165 0 1 948
box 0 0 1 1
use contact_18  contact_18_37
timestamp 1644951705
transform 1 0 19131 0 1 -3
box 0 0 1 1
use contact_17  contact_17_37
timestamp 1644951705
transform 1 0 19165 0 1 2
box 0 0 1 1
use contact_18  contact_18_38
timestamp 1644951705
transform 1 0 18859 0 1 943
box 0 0 1 1
use contact_17  contact_17_38
timestamp 1644951705
transform 1 0 18893 0 1 948
box 0 0 1 1
use contact_18  contact_18_39
timestamp 1644951705
transform 1 0 18859 0 1 -3
box 0 0 1 1
use contact_17  contact_17_39
timestamp 1644951705
transform 1 0 18893 0 1 2
box 0 0 1 1
use contact_18  contact_18_40
timestamp 1644951705
transform 1 0 16019 0 1 943
box 0 0 1 1
use contact_17  contact_17_40
timestamp 1644951705
transform 1 0 16053 0 1 948
box 0 0 1 1
use contact_18  contact_18_41
timestamp 1644951705
transform 1 0 16019 0 1 -3
box 0 0 1 1
use contact_17  contact_17_41
timestamp 1644951705
transform 1 0 16053 0 1 2
box 0 0 1 1
use contact_18  contact_18_42
timestamp 1644951705
transform 1 0 15747 0 1 943
box 0 0 1 1
use contact_17  contact_17_42
timestamp 1644951705
transform 1 0 15781 0 1 948
box 0 0 1 1
use contact_18  contact_18_43
timestamp 1644951705
transform 1 0 15747 0 1 -3
box 0 0 1 1
use contact_17  contact_17_43
timestamp 1644951705
transform 1 0 15781 0 1 2
box 0 0 1 1
use contact_18  contact_18_44
timestamp 1644951705
transform 1 0 12907 0 1 943
box 0 0 1 1
use contact_17  contact_17_44
timestamp 1644951705
transform 1 0 12941 0 1 948
box 0 0 1 1
use contact_18  contact_18_45
timestamp 1644951705
transform 1 0 12907 0 1 -3
box 0 0 1 1
use contact_17  contact_17_45
timestamp 1644951705
transform 1 0 12941 0 1 2
box 0 0 1 1
use contact_18  contact_18_46
timestamp 1644951705
transform 1 0 12635 0 1 943
box 0 0 1 1
use contact_17  contact_17_46
timestamp 1644951705
transform 1 0 12669 0 1 948
box 0 0 1 1
use contact_18  contact_18_47
timestamp 1644951705
transform 1 0 12635 0 1 -3
box 0 0 1 1
use contact_17  contact_17_47
timestamp 1644951705
transform 1 0 12669 0 1 2
box 0 0 1 1
use contact_18  contact_18_48
timestamp 1644951705
transform 1 0 9795 0 1 943
box 0 0 1 1
use contact_17  contact_17_48
timestamp 1644951705
transform 1 0 9829 0 1 948
box 0 0 1 1
use contact_18  contact_18_49
timestamp 1644951705
transform 1 0 9795 0 1 -3
box 0 0 1 1
use contact_17  contact_17_49
timestamp 1644951705
transform 1 0 9829 0 1 2
box 0 0 1 1
use contact_18  contact_18_50
timestamp 1644951705
transform 1 0 9523 0 1 943
box 0 0 1 1
use contact_17  contact_17_50
timestamp 1644951705
transform 1 0 9557 0 1 948
box 0 0 1 1
use contact_18  contact_18_51
timestamp 1644951705
transform 1 0 9523 0 1 -3
box 0 0 1 1
use contact_17  contact_17_51
timestamp 1644951705
transform 1 0 9557 0 1 2
box 0 0 1 1
use contact_18  contact_18_52
timestamp 1644951705
transform 1 0 6683 0 1 943
box 0 0 1 1
use contact_17  contact_17_52
timestamp 1644951705
transform 1 0 6717 0 1 948
box 0 0 1 1
use contact_18  contact_18_53
timestamp 1644951705
transform 1 0 6683 0 1 -3
box 0 0 1 1
use contact_17  contact_17_53
timestamp 1644951705
transform 1 0 6717 0 1 2
box 0 0 1 1
use contact_18  contact_18_54
timestamp 1644951705
transform 1 0 6411 0 1 943
box 0 0 1 1
use contact_17  contact_17_54
timestamp 1644951705
transform 1 0 6445 0 1 948
box 0 0 1 1
use contact_18  contact_18_55
timestamp 1644951705
transform 1 0 6411 0 1 -3
box 0 0 1 1
use contact_17  contact_17_55
timestamp 1644951705
transform 1 0 6445 0 1 2
box 0 0 1 1
use contact_18  contact_18_56
timestamp 1644951705
transform 1 0 3571 0 1 943
box 0 0 1 1
use contact_17  contact_17_56
timestamp 1644951705
transform 1 0 3605 0 1 948
box 0 0 1 1
use contact_18  contact_18_57
timestamp 1644951705
transform 1 0 3571 0 1 -3
box 0 0 1 1
use contact_17  contact_17_57
timestamp 1644951705
transform 1 0 3605 0 1 2
box 0 0 1 1
use contact_18  contact_18_58
timestamp 1644951705
transform 1 0 3299 0 1 943
box 0 0 1 1
use contact_17  contact_17_58
timestamp 1644951705
transform 1 0 3333 0 1 948
box 0 0 1 1
use contact_18  contact_18_59
timestamp 1644951705
transform 1 0 3299 0 1 -3
box 0 0 1 1
use contact_17  contact_17_59
timestamp 1644951705
transform 1 0 3333 0 1 2
box 0 0 1 1
use contact_18  contact_18_60
timestamp 1644951705
transform 1 0 459 0 1 943
box 0 0 1 1
use contact_17  contact_17_60
timestamp 1644951705
transform 1 0 493 0 1 948
box 0 0 1 1
use contact_18  contact_18_61
timestamp 1644951705
transform 1 0 459 0 1 -3
box 0 0 1 1
use contact_17  contact_17_61
timestamp 1644951705
transform 1 0 493 0 1 2
box 0 0 1 1
use contact_18  contact_18_62
timestamp 1644951705
transform 1 0 187 0 1 943
box 0 0 1 1
use contact_17  contact_17_62
timestamp 1644951705
transform 1 0 221 0 1 948
box 0 0 1 1
use contact_18  contact_18_63
timestamp 1644951705
transform 1 0 187 0 1 -3
box 0 0 1 1
use contact_17  contact_17_63
timestamp 1644951705
transform 1 0 221 0 1 2
box 0 0 1 1
use sense_amp_multiport  sense_amp_multiport_0
timestamp 1644951705
transform 1 0 47069 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_1
timestamp 1644951705
transform 1 0 46797 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_2
timestamp 1644951705
transform 1 0 43957 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_3
timestamp 1644951705
transform 1 0 43685 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_4
timestamp 1644951705
transform 1 0 40845 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_5
timestamp 1644951705
transform 1 0 40573 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_6
timestamp 1644951705
transform 1 0 37733 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_7
timestamp 1644951705
transform 1 0 37461 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_8
timestamp 1644951705
transform 1 0 34621 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_9
timestamp 1644951705
transform 1 0 34349 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_10
timestamp 1644951705
transform 1 0 31509 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_11
timestamp 1644951705
transform 1 0 31237 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_12
timestamp 1644951705
transform 1 0 28397 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_13
timestamp 1644951705
transform 1 0 28125 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_14
timestamp 1644951705
transform 1 0 25285 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_15
timestamp 1644951705
transform 1 0 25013 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_16
timestamp 1644951705
transform 1 0 22173 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_17
timestamp 1644951705
transform 1 0 21901 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_18
timestamp 1644951705
transform 1 0 19061 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_19
timestamp 1644951705
transform 1 0 18789 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_20
timestamp 1644951705
transform 1 0 15949 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_21
timestamp 1644951705
transform 1 0 15677 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_22
timestamp 1644951705
transform 1 0 12837 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_23
timestamp 1644951705
transform 1 0 12565 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_24
timestamp 1644951705
transform 1 0 9725 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_25
timestamp 1644951705
transform 1 0 9453 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_26
timestamp 1644951705
transform 1 0 6613 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_27
timestamp 1644951705
transform 1 0 6341 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_28
timestamp 1644951705
transform 1 0 3501 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_29
timestamp 1644951705
transform 1 0 3229 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_30
timestamp 1644951705
transform 1 0 389 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_31
timestamp 1644951705
transform 1 0 117 0 1 0
box 0 0 272 1050
<< labels >>
rlabel metal3 s 18859 -3 18991 71 4 gnd
rlabel metal3 s 44027 -3 44159 71 4 gnd
rlabel metal3 s 16019 -3 16151 71 4 gnd
rlabel metal3 s 34419 -3 34551 71 4 gnd
rlabel metal3 s 28467 -3 28599 71 4 gnd
rlabel metal3 s 31307 -3 31439 71 4 gnd
rlabel metal3 s 25083 -3 25215 71 4 gnd
rlabel metal3 s 40643 -3 40775 71 4 gnd
rlabel metal3 s 28195 -3 28327 71 4 gnd
rlabel metal3 s 6411 -3 6543 71 4 gnd
rlabel metal3 s 47139 -3 47271 71 4 gnd
rlabel metal3 s 40915 -3 41047 71 4 gnd
rlabel metal3 s 3571 -3 3703 71 4 gnd
rlabel metal3 s 6683 -3 6815 71 4 gnd
rlabel metal3 s 25355 -3 25487 71 4 gnd
rlabel metal3 s 9523 -3 9655 71 4 gnd
rlabel metal3 s 37803 -3 37935 71 4 gnd
rlabel metal3 s 187 -3 319 71 4 gnd
rlabel metal3 s 12635 -3 12767 71 4 gnd
rlabel metal3 s 15747 -3 15879 71 4 gnd
rlabel metal3 s 31579 -3 31711 71 4 gnd
rlabel metal3 s 3299 -3 3431 71 4 gnd
rlabel metal3 s 19131 -3 19263 71 4 gnd
rlabel metal3 s 22243 -3 22375 71 4 gnd
rlabel metal3 s 459 -3 591 71 4 gnd
rlabel metal3 s 34691 -3 34823 71 4 gnd
rlabel metal3 s 9795 -3 9927 71 4 gnd
rlabel metal3 s 12907 -3 13039 71 4 gnd
rlabel metal3 s 37531 -3 37663 71 4 gnd
rlabel metal3 s 43755 -3 43887 71 4 gnd
rlabel metal3 s 21971 -3 22103 71 4 gnd
rlabel metal3 s 46867 -3 46999 71 4 gnd
rlabel metal3 s 22243 943 22375 1017 4 vdd
rlabel metal3 s 16019 943 16151 1017 4 vdd
rlabel metal3 s 18859 943 18991 1017 4 vdd
rlabel metal3 s 25355 943 25487 1017 4 vdd
rlabel metal3 s 47139 943 47271 1017 4 vdd
rlabel metal3 s 31579 943 31711 1017 4 vdd
rlabel metal3 s 28467 943 28599 1017 4 vdd
rlabel metal3 s 44027 943 44159 1017 4 vdd
rlabel metal3 s 3571 943 3703 1017 4 vdd
rlabel metal3 s 6683 943 6815 1017 4 vdd
rlabel metal3 s 34691 943 34823 1017 4 vdd
rlabel metal3 s 459 943 591 1017 4 vdd
rlabel metal3 s 9523 943 9655 1017 4 vdd
rlabel metal3 s 28195 943 28327 1017 4 vdd
rlabel metal3 s 19131 943 19263 1017 4 vdd
rlabel metal3 s 37803 943 37935 1017 4 vdd
rlabel metal3 s 43755 943 43887 1017 4 vdd
rlabel metal3 s 40915 943 41047 1017 4 vdd
rlabel metal3 s 34419 943 34551 1017 4 vdd
rlabel metal3 s 187 943 319 1017 4 vdd
rlabel metal3 s 12635 943 12767 1017 4 vdd
rlabel metal3 s 6411 943 6543 1017 4 vdd
rlabel metal3 s 21971 943 22103 1017 4 vdd
rlabel metal3 s 31307 943 31439 1017 4 vdd
rlabel metal3 s 9795 943 9927 1017 4 vdd
rlabel metal3 s 46867 943 46999 1017 4 vdd
rlabel metal3 s 40643 943 40775 1017 4 vdd
rlabel metal3 s 37531 943 37663 1017 4 vdd
rlabel metal3 s 25083 943 25215 1017 4 vdd
rlabel metal3 s 15747 943 15879 1017 4 vdd
rlabel metal3 s 12907 943 13039 1017 4 vdd
rlabel metal3 s 3299 943 3431 1017 4 vdd
rlabel metal2 s 131 0 159 240 4 rbl_0
rlabel metal2 s 319 0 347 240 4 data_0
rlabel metal2 s 403 0 431 240 4 rbl_1
rlabel metal2 s 591 0 619 240 4 data_1
rlabel metal2 s 3243 0 3271 240 4 rbl_2
rlabel metal2 s 3431 0 3459 240 4 data_2
rlabel metal2 s 3515 0 3543 240 4 rbl_3
rlabel metal2 s 3703 0 3731 240 4 data_3
rlabel metal2 s 6355 0 6383 240 4 rbl_4
rlabel metal2 s 6543 0 6571 240 4 data_4
rlabel metal2 s 6627 0 6655 240 4 rbl_5
rlabel metal2 s 6815 0 6843 240 4 data_5
rlabel metal2 s 9467 0 9495 240 4 rbl_6
rlabel metal2 s 9655 0 9683 240 4 data_6
rlabel metal2 s 9739 0 9767 240 4 rbl_7
rlabel metal2 s 9927 0 9955 240 4 data_7
rlabel metal2 s 12579 0 12607 240 4 rbl_8
rlabel metal2 s 12767 0 12795 240 4 data_8
rlabel metal2 s 12851 0 12879 240 4 rbl_9
rlabel metal2 s 13039 0 13067 240 4 data_9
rlabel metal2 s 15691 0 15719 240 4 rbl_10
rlabel metal2 s 15879 0 15907 240 4 data_10
rlabel metal2 s 15963 0 15991 240 4 rbl_11
rlabel metal2 s 16151 0 16179 240 4 data_11
rlabel metal2 s 18803 0 18831 240 4 rbl_12
rlabel metal2 s 18991 0 19019 240 4 data_12
rlabel metal2 s 19075 0 19103 240 4 rbl_13
rlabel metal2 s 19263 0 19291 240 4 data_13
rlabel metal2 s 21915 0 21943 240 4 rbl_14
rlabel metal2 s 22103 0 22131 240 4 data_14
rlabel metal2 s 22187 0 22215 240 4 rbl_15
rlabel metal2 s 22375 0 22403 240 4 data_15
rlabel metal2 s 25027 0 25055 240 4 rbl_16
rlabel metal2 s 25215 0 25243 240 4 data_16
rlabel metal2 s 25299 0 25327 240 4 rbl_17
rlabel metal2 s 25487 0 25515 240 4 data_17
rlabel metal2 s 28139 0 28167 240 4 rbl_18
rlabel metal2 s 28327 0 28355 240 4 data_18
rlabel metal2 s 28411 0 28439 240 4 rbl_19
rlabel metal2 s 28599 0 28627 240 4 data_19
rlabel metal2 s 31251 0 31279 240 4 rbl_20
rlabel metal2 s 31439 0 31467 240 4 data_20
rlabel metal2 s 31523 0 31551 240 4 rbl_21
rlabel metal2 s 31711 0 31739 240 4 data_21
rlabel metal2 s 34363 0 34391 240 4 rbl_22
rlabel metal2 s 34551 0 34579 240 4 data_22
rlabel metal2 s 34635 0 34663 240 4 rbl_23
rlabel metal2 s 34823 0 34851 240 4 data_23
rlabel metal2 s 37475 0 37503 240 4 rbl_24
rlabel metal2 s 37663 0 37691 240 4 data_24
rlabel metal2 s 37747 0 37775 240 4 rbl_25
rlabel metal2 s 37935 0 37963 240 4 data_25
rlabel metal2 s 40587 0 40615 240 4 rbl_26
rlabel metal2 s 40775 0 40803 240 4 data_26
rlabel metal2 s 40859 0 40887 240 4 rbl_27
rlabel metal2 s 41047 0 41075 240 4 data_27
rlabel metal2 s 43699 0 43727 240 4 rbl_28
rlabel metal2 s 43887 0 43915 240 4 data_28
rlabel metal2 s 43971 0 43999 240 4 rbl_29
rlabel metal2 s 44159 0 44187 240 4 data_29
rlabel metal2 s 46811 0 46839 240 4 rbl_30
rlabel metal2 s 46999 0 47027 240 4 data_30
rlabel metal2 s 47083 0 47111 240 4 rbl_31
rlabel metal2 s 47271 0 47299 240 4 data_31
<< properties >>
string FIXED_BBOX 47139 -3 47271 0
string GDS_FILE sram_0rw2r1w_16_128_sky130A.gds
string GDS_END 1489918
string GDS_START 1454990
<< end >>
