magic
tech sky130A
magscale 1 2
timestamp 1644949024
<< checkpaint >>
rect -1260 -1286 1410 1370
<< scnmos >>
rect 60 0 90 84
<< ndiff >>
rect 0 59 60 84
rect 0 25 8 59
rect 42 25 60 59
rect 0 0 60 25
rect 90 59 150 84
rect 90 25 108 59
rect 142 25 150 59
rect 90 0 150 25
<< ndiffc >>
rect 8 25 42 59
rect 108 25 142 59
<< poly >>
rect 60 84 90 110
rect 60 -26 90 0
<< locali >>
rect 8 59 42 75
rect 8 9 42 25
rect 108 59 142 75
rect 108 9 142 25
use contact_8  contact_8_0
timestamp 1644949024
transform 1 0 100 0 1 1
box 0 0 1 1
use contact_8  contact_8_1
timestamp 1644949024
transform 1 0 0 0 1 1
box 0 0 1 1
<< labels >>
rlabel mvvaractor s 75 42 75 42 4 G
rlabel locali s 25 42 25 42 4 S
rlabel locali s 125 42 125 42 4 D
<< properties >>
string FIXED_BBOX -25 -26 175 110
string GDS_FILE sram_0rw2r1w_4_16_sky130A.gds
string GDS_END 339574
string GDS_START 338810
<< end >>
