magic
tech sky130A
magscale 1 2
timestamp 1644969367
<< checkpaint >>
rect -1296 -1277 1772 2155
<< nwell >>
rect -36 402 512 895
<< pwell >>
rect 366 51 416 133
<< psubdiff >>
rect 366 109 416 133
rect 366 75 374 109
rect 408 75 416 109
rect 366 51 416 75
<< nsubdiff >>
rect 366 763 416 787
rect 366 729 374 763
rect 408 729 416 763
rect 366 705 416 729
<< psubdiffcont >>
rect 374 75 408 109
<< nsubdiffcont >>
rect 374 729 408 763
<< poly >>
rect 114 410 144 479
rect 48 394 144 410
rect 48 360 64 394
rect 98 360 144 394
rect 48 344 144 360
rect 114 191 144 344
<< polycont >>
rect 64 360 98 394
<< locali >>
rect 0 821 476 855
rect 62 628 96 821
rect 48 394 114 410
rect 48 360 64 394
rect 98 360 114 394
rect 48 344 114 360
rect 166 394 200 694
rect 270 628 304 821
rect 374 763 408 821
rect 374 713 408 729
rect 166 360 217 394
rect 166 60 200 360
rect 374 109 408 125
rect 62 17 96 60
rect 270 17 304 60
rect 374 17 408 75
rect 0 -17 476 17
use contact_12  contact_12_0
timestamp 1644969367
transform 1 0 48 0 1 344
box 0 0 1 1
use contact_11  contact_11_0
timestamp 1644969367
transform 1 0 366 0 1 51
box 0 0 1 1
use contact_10  contact_10_0
timestamp 1644969367
transform 1 0 366 0 1 705
box 0 0 1 1
use nmos_m2_w0_420_sli_dli_da_p  nmos_m2_w0_420_sli_dli_da_p_0
timestamp 1644969367
transform 1 0 54 0 1 51
box 0 -26 258 140
use pmos_m2_w1_260_sli_dli_da_p  pmos_m2_w1_260_sli_dli_da_p_0
timestamp 1644969367
transform 1 0 54 0 1 535
box -59 -56 317 306
<< labels >>
rlabel locali s 81 377 81 377 4 A
rlabel locali s 200 377 200 377 4 Z
rlabel locali s 238 0 238 0 4 gnd
rlabel locali s 238 838 238 838 4 vdd
<< properties >>
string FIXED_BBOX 0 0 476 838
string GDS_FILE sram_0rw2r1w_32_128_sky130A.gds
string GDS_END 3260842
string GDS_START 3259222
<< end >>
