magic
tech sky130A
magscale 1 2
timestamp 1644969367
<< checkpaint >>
rect -1296 -1277 3500 2155
<< nwell >>
rect -36 402 2240 895
<< pwell >>
rect 2094 51 2144 133
<< psubdiff >>
rect 2094 109 2144 133
rect 2094 75 2102 109
rect 2136 75 2144 109
rect 2094 51 2144 75
<< nsubdiff >>
rect 2094 763 2144 787
rect 2094 729 2102 763
rect 2136 729 2144 763
rect 2094 705 2144 729
<< psubdiffcont >>
rect 2102 75 2136 109
<< nsubdiffcont >>
rect 2102 729 2136 763
<< poly >>
rect 114 403 144 437
rect 48 387 144 403
rect 48 353 64 387
rect 98 353 144 387
rect 48 337 144 353
rect 114 205 144 337
<< polycont >>
rect 64 353 98 387
<< locali >>
rect 0 821 2204 855
rect 62 607 96 821
rect 274 607 308 821
rect 490 607 524 821
rect 706 607 740 821
rect 922 607 956 821
rect 1138 607 1172 821
rect 1354 607 1388 821
rect 1570 607 1604 821
rect 1786 607 1820 821
rect 1998 607 2032 821
rect 2102 763 2136 821
rect 2102 713 2136 729
rect 48 387 114 403
rect 48 353 64 387
rect 98 353 114 387
rect 48 337 114 353
rect 1030 387 1064 573
rect 1030 353 1081 387
rect 1030 167 1064 353
rect 2102 109 2136 125
rect 62 17 96 67
rect 274 17 308 67
rect 490 17 524 67
rect 706 17 740 67
rect 922 17 956 67
rect 1138 17 1172 67
rect 1354 17 1388 67
rect 1570 17 1604 67
rect 1786 17 1820 67
rect 1998 17 2032 67
rect 2102 17 2136 75
rect 0 -17 2204 17
use contact_12  contact_12_0
timestamp 1644969367
transform 1 0 48 0 1 337
box 0 0 1 1
use contact_11  contact_11_0
timestamp 1644969367
transform 1 0 2094 0 1 51
box 0 0 1 1
use contact_10  contact_10_0
timestamp 1644969367
transform 1 0 2094 0 1 705
box 0 0 1 1
use nmos_m18_w0_490_sli_dli_da_p  nmos_m18_w0_490_sli_dli_da_p_0
timestamp 1644969367
transform 1 0 54 0 1 51
box 0 -26 1986 154
use pmos_m18_w1_470_sli_dli_da_p  pmos_m18_w1_470_sli_dli_da_p_0
timestamp 1644969367
transform 1 0 54 0 1 493
box -59 -56 2045 348
<< labels >>
rlabel locali s 81 370 81 370 4 A
rlabel locali s 1064 370 1064 370 4 Z
rlabel locali s 1102 0 1102 0 4 gnd
rlabel locali s 1102 838 1102 838 4 vdd
<< properties >>
string FIXED_BBOX 0 0 2204 838
string GDS_FILE sram_0rw2r1w_32_128_sky130A.gds
string GDS_END 3384024
string GDS_START 3381380
<< end >>
