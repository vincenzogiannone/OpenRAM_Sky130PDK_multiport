magic
tech sky130A
timestamp 1644915396
<< nwell >>
rect 0 559 747 808
<< nmos >>
rect 47 66 62 166
rect 95 66 110 166
rect 143 66 158 166
rect 191 66 206 166
rect 239 66 254 166
rect 287 66 302 166
rect 389 66 404 166
rect 437 66 452 166
rect 485 66 500 166
rect 537 66 552 108
rect 637 66 652 108
rect 685 66 700 108
<< pmos >>
rect 47 577 62 619
rect 95 577 110 619
rect 143 577 158 619
rect 191 577 206 619
rect 239 577 254 619
rect 287 577 302 619
rect 389 577 404 619
rect 437 577 452 619
rect 485 577 500 619
rect 537 577 552 712
rect 637 577 652 712
rect 685 577 700 712
<< ndiff >>
rect 18 149 47 166
rect 18 132 22 149
rect 39 132 47 149
rect 18 100 47 132
rect 18 83 22 100
rect 39 83 47 100
rect 18 66 47 83
rect 62 66 95 166
rect 110 66 143 166
rect 158 149 191 166
rect 158 132 166 149
rect 183 132 191 149
rect 158 100 191 132
rect 158 83 166 100
rect 183 83 191 100
rect 158 66 191 83
rect 206 66 239 166
rect 254 66 287 166
rect 302 149 331 166
rect 302 132 310 149
rect 327 132 331 149
rect 302 100 331 132
rect 302 83 310 100
rect 327 83 331 100
rect 302 66 331 83
rect 360 149 389 166
rect 360 132 364 149
rect 381 132 389 149
rect 360 100 389 132
rect 360 83 364 100
rect 381 83 389 100
rect 360 66 389 83
rect 404 66 437 166
rect 452 66 485 166
rect 500 149 529 166
rect 500 132 508 149
rect 525 132 529 149
rect 500 108 529 132
rect 500 100 537 108
rect 500 83 508 100
rect 525 83 537 100
rect 500 66 537 83
rect 552 95 581 108
rect 552 78 560 95
rect 577 78 581 95
rect 552 66 581 78
rect 608 95 637 108
rect 608 78 612 95
rect 629 78 637 95
rect 608 66 637 78
rect 652 95 685 108
rect 652 78 660 95
rect 677 78 685 95
rect 652 66 685 78
rect 700 95 729 108
rect 700 78 708 95
rect 725 78 729 95
rect 700 66 729 78
<< pdiff >>
rect 508 695 537 712
rect 508 678 512 695
rect 529 678 537 695
rect 508 653 537 678
rect 508 636 512 653
rect 529 636 537 653
rect 508 619 537 636
rect 18 606 47 619
rect 18 589 22 606
rect 39 589 47 606
rect 18 577 47 589
rect 62 606 95 619
rect 62 589 70 606
rect 87 589 95 606
rect 62 577 95 589
rect 110 606 143 619
rect 110 589 118 606
rect 135 589 143 606
rect 110 577 143 589
rect 158 606 191 619
rect 158 589 166 606
rect 183 589 191 606
rect 158 577 191 589
rect 206 606 239 619
rect 206 589 214 606
rect 231 589 239 606
rect 206 577 239 589
rect 254 606 287 619
rect 254 589 262 606
rect 279 589 287 606
rect 254 577 287 589
rect 302 606 331 619
rect 302 589 310 606
rect 327 589 331 606
rect 302 577 331 589
rect 360 606 389 619
rect 360 589 364 606
rect 381 589 389 606
rect 360 577 389 589
rect 404 606 437 619
rect 404 589 412 606
rect 429 589 437 606
rect 404 577 437 589
rect 452 606 485 619
rect 452 589 460 606
rect 477 589 485 606
rect 452 577 485 589
rect 500 611 537 619
rect 500 594 512 611
rect 529 594 537 611
rect 500 577 537 594
rect 552 695 581 712
rect 552 678 560 695
rect 577 678 581 695
rect 552 653 581 678
rect 552 636 560 653
rect 577 636 581 653
rect 552 611 581 636
rect 552 594 560 611
rect 577 594 581 611
rect 552 577 581 594
rect 608 695 637 712
rect 608 678 612 695
rect 629 678 637 695
rect 608 653 637 678
rect 608 636 612 653
rect 629 636 637 653
rect 608 611 637 636
rect 608 594 612 611
rect 629 594 637 611
rect 608 577 637 594
rect 652 695 685 712
rect 652 678 660 695
rect 677 678 685 695
rect 652 653 685 678
rect 652 636 660 653
rect 677 636 685 653
rect 652 611 685 636
rect 652 594 660 611
rect 677 594 685 611
rect 652 577 685 594
rect 700 695 729 712
rect 700 678 708 695
rect 725 678 729 695
rect 700 653 729 678
rect 700 636 708 653
rect 725 636 729 653
rect 700 611 729 636
rect 700 594 708 611
rect 725 594 729 611
rect 700 577 729 594
<< ndiffc >>
rect 22 132 39 149
rect 22 83 39 100
rect 166 132 183 149
rect 166 83 183 100
rect 310 132 327 149
rect 310 83 327 100
rect 364 132 381 149
rect 364 83 381 100
rect 508 132 525 149
rect 508 83 525 100
rect 560 78 577 95
rect 612 78 629 95
rect 660 78 677 95
rect 708 78 725 95
<< pdiffc >>
rect 512 678 529 695
rect 512 636 529 653
rect 22 589 39 606
rect 70 589 87 606
rect 118 589 135 606
rect 166 589 183 606
rect 214 589 231 606
rect 262 589 279 606
rect 310 589 327 606
rect 364 589 381 606
rect 412 589 429 606
rect 460 589 477 606
rect 512 594 529 611
rect 560 678 577 695
rect 560 636 577 653
rect 560 594 577 611
rect 612 678 629 695
rect 612 636 629 653
rect 612 594 629 611
rect 660 678 677 695
rect 660 636 677 653
rect 660 594 677 611
rect 708 678 725 695
rect 708 636 725 653
rect 708 594 725 611
<< psubdiff >>
rect 120 9 156 21
rect 120 -9 129 9
rect 147 -9 156 9
rect 120 -21 156 -9
rect 277 9 313 21
rect 277 -9 286 9
rect 304 -9 313 9
rect 277 -21 313 -9
rect 434 9 470 21
rect 434 -9 443 9
rect 461 -9 470 9
rect 434 -21 470 -9
rect 591 9 627 21
rect 591 -9 600 9
rect 618 -9 627 9
rect 591 -21 627 -9
<< nsubdiff >>
rect 120 778 156 790
rect 120 760 129 778
rect 147 760 156 778
rect 120 748 156 760
rect 277 778 313 790
rect 277 760 286 778
rect 304 760 313 778
rect 277 748 313 760
rect 434 778 470 790
rect 434 760 443 778
rect 461 760 470 778
rect 434 748 470 760
rect 591 778 627 790
rect 591 760 600 778
rect 618 760 627 778
rect 591 748 627 760
<< psubdiffcont >>
rect 129 -9 147 9
rect 286 -9 304 9
rect 443 -9 461 9
rect 600 -9 618 9
<< nsubdiffcont >>
rect 129 760 147 778
rect 286 760 304 778
rect 443 760 461 778
rect 600 760 618 778
<< poly >>
rect 537 712 552 725
rect 637 712 652 725
rect 685 712 700 725
rect 47 619 62 632
rect 95 619 110 632
rect 143 619 158 632
rect 191 619 206 632
rect 239 619 254 632
rect 287 619 302 632
rect 389 619 404 632
rect 437 619 452 632
rect 485 619 500 632
rect 47 560 62 577
rect 35 552 62 560
rect 35 535 40 552
rect 57 535 62 552
rect 35 527 62 535
rect 47 166 62 527
rect 95 517 110 577
rect 83 509 110 517
rect 83 492 88 509
rect 105 492 110 509
rect 83 484 110 492
rect 95 166 110 484
rect 143 474 158 577
rect 131 466 158 474
rect 131 449 136 466
rect 153 449 158 466
rect 131 441 158 449
rect 143 166 158 441
rect 191 431 206 577
rect 179 423 206 431
rect 179 406 184 423
rect 201 406 206 423
rect 179 398 206 406
rect 191 166 206 398
rect 239 388 254 577
rect 227 380 254 388
rect 227 363 232 380
rect 249 363 254 380
rect 227 355 254 363
rect 239 166 254 355
rect 287 345 302 577
rect 275 337 302 345
rect 275 320 280 337
rect 297 320 302 337
rect 275 312 302 320
rect 287 166 302 312
rect 389 302 404 577
rect 377 294 404 302
rect 377 277 382 294
rect 399 277 404 294
rect 377 269 404 277
rect 389 166 404 269
rect 437 259 452 577
rect 425 251 452 259
rect 425 234 430 251
rect 447 234 452 251
rect 425 226 452 234
rect 437 166 452 226
rect 485 216 500 577
rect 537 319 552 577
rect 525 311 552 319
rect 525 294 530 311
rect 547 294 552 311
rect 525 286 552 294
rect 473 208 500 216
rect 473 191 478 208
rect 495 191 500 208
rect 473 183 500 191
rect 485 166 500 183
rect 537 108 552 286
rect 637 420 652 577
rect 685 560 700 577
rect 673 552 700 560
rect 673 535 678 552
rect 695 535 700 552
rect 673 527 700 535
rect 637 412 664 420
rect 637 395 642 412
rect 659 395 664 412
rect 637 387 664 395
rect 637 108 652 387
rect 685 108 700 527
rect 47 53 62 66
rect 95 53 110 66
rect 143 53 158 66
rect 191 53 206 66
rect 239 53 254 66
rect 287 53 302 66
rect 389 53 404 66
rect 437 53 452 66
rect 485 53 500 66
rect 537 53 552 66
rect 637 53 652 66
rect 685 53 700 66
<< polycont >>
rect 40 535 57 552
rect 88 492 105 509
rect 136 449 153 466
rect 184 406 201 423
rect 232 363 249 380
rect 280 320 297 337
rect 382 277 399 294
rect 430 234 447 251
rect 530 294 547 311
rect 478 191 495 208
rect 678 535 695 552
rect 642 395 659 412
<< locali >>
rect 129 778 147 786
rect 286 778 304 786
rect 443 778 461 786
rect 600 778 618 786
rect 70 760 129 778
rect 147 760 286 778
rect 304 760 443 778
rect 461 760 600 778
rect 618 760 677 778
rect 70 619 87 760
rect 129 752 147 760
rect 166 619 183 760
rect 262 752 304 760
rect 412 752 461 760
rect 262 619 279 752
rect 412 619 429 752
rect 512 712 529 760
rect 600 752 618 760
rect 660 712 677 760
rect 508 695 532 712
rect 508 678 512 695
rect 529 678 532 695
rect 508 653 532 678
rect 508 636 512 653
rect 529 636 532 653
rect 18 606 42 619
rect 18 589 22 606
rect 39 589 42 606
rect 18 577 42 589
rect 67 606 90 619
rect 67 589 70 606
rect 87 589 90 606
rect 67 577 90 589
rect 115 606 138 619
rect 115 589 118 606
rect 135 589 138 606
rect 115 577 138 589
rect 163 606 186 619
rect 163 589 166 606
rect 183 589 186 606
rect 163 577 186 589
rect 211 606 234 619
rect 211 589 214 606
rect 231 589 234 606
rect 211 577 234 589
rect 259 606 282 619
rect 259 589 262 606
rect 279 589 282 606
rect 259 577 282 589
rect 307 606 331 619
rect 307 589 310 606
rect 327 589 331 606
rect 307 577 331 589
rect 360 606 384 619
rect 360 589 364 606
rect 381 589 384 606
rect 360 577 384 589
rect 409 606 432 619
rect 409 589 412 606
rect 429 589 432 606
rect 409 577 432 589
rect 457 606 480 619
rect 457 589 460 606
rect 477 589 480 606
rect 457 577 480 589
rect 508 611 532 636
rect 508 594 512 611
rect 529 594 532 611
rect 508 577 532 594
rect 557 695 581 712
rect 557 678 560 695
rect 577 678 581 695
rect 557 653 581 678
rect 557 636 560 653
rect 577 636 581 653
rect 557 611 581 636
rect 557 594 560 611
rect 577 594 581 611
rect 557 577 581 594
rect 40 552 57 560
rect 40 527 57 535
rect 348 538 364 555
rect 88 509 105 517
rect 88 484 105 492
rect 136 466 153 474
rect 136 441 153 449
rect 184 423 201 431
rect 184 398 201 406
rect 232 380 249 388
rect 232 355 249 363
rect 280 337 297 345
rect 280 312 297 320
rect 314 295 331 398
rect 22 278 331 295
rect 22 166 39 278
rect 348 261 365 538
rect 463 327 480 577
rect 463 311 547 327
rect 463 310 530 311
rect 382 294 399 302
rect 530 286 547 294
rect 564 304 581 577
rect 608 695 632 712
rect 608 678 612 695
rect 629 678 632 695
rect 608 653 632 678
rect 608 636 612 653
rect 629 636 632 653
rect 608 611 632 636
rect 608 594 612 611
rect 629 594 632 611
rect 608 577 632 594
rect 657 695 680 712
rect 657 678 660 695
rect 677 678 680 695
rect 657 653 680 678
rect 657 636 660 653
rect 677 636 680 653
rect 657 611 680 636
rect 657 594 660 611
rect 677 594 680 611
rect 657 577 680 594
rect 705 695 729 712
rect 705 678 708 695
rect 725 678 729 695
rect 705 653 729 678
rect 705 636 708 653
rect 725 636 729 653
rect 705 611 729 636
rect 705 594 708 611
rect 725 594 729 611
rect 705 577 729 594
rect 608 365 625 577
rect 678 552 695 560
rect 678 527 695 535
rect 712 438 729 577
rect 642 412 659 420
rect 642 387 659 395
rect 564 287 567 304
rect 382 269 399 277
rect 310 244 365 261
rect 430 251 447 259
rect 310 166 327 244
rect 430 226 447 234
rect 478 208 495 216
rect 478 183 495 191
rect 18 149 42 166
rect 18 132 22 149
rect 39 132 42 149
rect 18 100 42 132
rect 18 83 22 100
rect 39 83 42 100
rect 18 66 42 83
rect 163 149 186 166
rect 163 132 166 149
rect 183 132 186 149
rect 163 100 186 132
rect 163 83 166 100
rect 183 83 186 100
rect 163 66 186 83
rect 307 149 331 166
rect 307 132 310 149
rect 327 132 331 149
rect 307 100 331 132
rect 307 83 310 100
rect 327 83 331 100
rect 307 66 331 83
rect 360 149 384 166
rect 360 132 364 149
rect 381 132 384 149
rect 360 100 384 132
rect 360 83 364 100
rect 381 83 384 100
rect 360 66 384 83
rect 505 149 529 166
rect 505 132 508 149
rect 525 132 529 149
rect 505 100 529 132
rect 564 108 581 287
rect 505 83 508 100
rect 525 83 529 100
rect 505 66 529 83
rect 557 95 581 108
rect 557 78 560 95
rect 577 78 581 95
rect 557 66 581 78
rect 608 108 625 348
rect 712 108 729 421
rect 608 95 632 108
rect 608 78 612 95
rect 629 78 632 95
rect 608 66 632 78
rect 657 95 680 108
rect 657 78 660 95
rect 677 78 680 95
rect 657 66 680 78
rect 705 95 729 108
rect 705 78 708 95
rect 725 78 729 95
rect 705 66 729 78
rect 129 9 147 21
rect 166 9 183 66
rect 286 9 304 21
rect 443 9 461 21
rect 508 9 525 66
rect 600 9 618 21
rect 660 9 677 66
rect 70 -9 129 9
rect 147 -9 286 9
rect 304 -9 443 9
rect 461 -9 600 9
rect 618 -9 677 9
rect 129 -21 147 -9
rect 286 -21 304 -9
rect 443 -21 461 -9
rect 600 -21 618 -9
<< viali >>
rect 129 760 147 778
rect 286 760 304 778
rect 443 760 461 778
rect 600 760 618 778
rect 22 589 39 606
rect 118 589 135 606
rect 214 589 231 606
rect 310 589 327 606
rect 364 589 381 606
rect 460 589 477 606
rect 40 535 57 552
rect 364 538 381 555
rect 88 492 105 509
rect 136 449 153 466
rect 184 406 201 423
rect 314 398 331 415
rect 232 363 249 380
rect 280 320 297 337
rect 382 277 399 294
rect 530 294 547 311
rect 678 535 695 552
rect 712 421 729 438
rect 642 395 659 412
rect 608 348 625 365
rect 567 287 584 304
rect 430 234 447 251
rect 478 191 495 208
rect 364 83 381 100
rect 129 -9 147 9
rect 286 -9 304 9
rect 443 -9 461 9
rect 600 -9 618 9
<< metal1 >>
rect 0 778 747 784
rect 0 760 129 778
rect 147 760 286 778
rect 304 760 443 778
rect 461 760 600 778
rect 618 760 747 778
rect 0 754 747 760
rect 19 606 138 612
rect 19 589 22 606
rect 39 598 118 606
rect 39 589 42 598
rect 19 583 42 589
rect 115 589 118 598
rect 135 589 138 606
rect 115 583 138 589
rect 211 606 330 612
rect 211 589 214 606
rect 231 598 310 606
rect 231 589 234 598
rect 211 583 234 589
rect 307 589 310 598
rect 327 589 330 606
rect 307 583 330 589
rect 361 606 480 612
rect 361 589 364 606
rect 381 598 460 606
rect 381 589 384 598
rect 361 583 384 589
rect 457 589 460 598
rect 477 589 480 606
rect 457 583 480 589
rect 124 565 138 583
rect 36 552 63 559
rect 36 542 40 552
rect 35 535 40 542
rect 57 535 63 552
rect 124 551 253 565
rect 35 528 63 535
rect 84 509 111 516
rect 84 499 88 509
rect 83 492 88 499
rect 105 492 111 509
rect 83 485 111 492
rect 132 466 159 473
rect 132 456 136 466
rect 131 449 136 456
rect 153 449 159 466
rect 239 465 253 551
rect 316 561 330 583
rect 316 558 384 561
rect 316 555 698 558
rect 316 547 364 555
rect 361 538 364 547
rect 381 552 698 555
rect 381 544 678 552
rect 381 538 384 544
rect 361 532 384 538
rect 675 535 678 544
rect 695 535 698 552
rect 675 529 698 535
rect 239 451 321 465
rect 131 442 159 449
rect 180 423 207 430
rect 180 413 184 423
rect 179 406 184 413
rect 201 406 207 423
rect 179 399 207 406
rect 307 418 321 451
rect 709 438 732 444
rect 709 421 712 438
rect 729 424 747 438
rect 729 421 732 424
rect 307 415 662 418
rect 709 415 732 421
rect 307 398 314 415
rect 331 412 662 415
rect 331 404 642 412
rect 331 398 337 404
rect 307 393 337 398
rect 639 395 642 404
rect 659 395 662 412
rect 639 389 662 395
rect 228 380 255 387
rect 228 370 232 380
rect 227 363 232 370
rect 249 363 255 380
rect 227 356 255 363
rect 605 365 628 371
rect 605 348 608 365
rect 625 351 747 365
rect 625 348 628 351
rect 276 337 303 344
rect 605 342 628 348
rect 276 327 280 337
rect 275 320 280 327
rect 297 320 303 337
rect 275 313 303 320
rect 527 311 550 317
rect 378 294 405 301
rect 378 284 382 294
rect 377 277 382 284
rect 399 277 405 294
rect 527 294 530 311
rect 547 294 550 311
rect 527 288 550 294
rect 377 270 405 277
rect 426 251 453 258
rect 426 241 430 251
rect 425 234 430 241
rect 447 234 453 251
rect 425 227 453 234
rect 474 208 501 215
rect 474 198 478 208
rect 473 191 478 198
rect 495 191 501 208
rect 473 184 501 191
rect 536 106 550 288
rect 564 304 587 310
rect 564 287 567 304
rect 584 290 747 304
rect 584 287 587 290
rect 564 281 587 287
rect 361 100 550 106
rect 361 83 364 100
rect 381 92 550 100
rect 381 83 384 92
rect 361 77 384 83
rect 0 9 747 15
rect 0 -9 129 9
rect 147 -9 286 9
rect 304 -9 443 9
rect 461 -9 600 9
rect 618 -9 747 9
rect 0 -15 747 -9
<< labels >>
flabel metal1 736 296 736 296 0 FreeSans 80 0 0 0 OUT2
port 11 nsew
flabel metal1 348 0 348 0 0 FreeSans 80 0 0 0 gnd
port 13 nsew
flabel locali 475 375 475 375 0 FreeSans 80 0 0 0 net9
flabel metal1 742 430 742 430 0 FreeSans 80 0 0 0 OUT0
port 14 nsew
flabel metal1 740 354 740 354 0 FreeSans 80 0 0 0 OUT1
port 15 nsew
flabel metal1 355 768 355 768 0 FreeSans 80 0 0 0 vdd
port 12 nsew
flabel metal1 326 551 326 551 0 FreeSans 80 0 0 0 net6
flabel metal1 179 553 179 553 0 FreeSans 80 0 0 0 net3
flabel metal1 35 535 35 535 0 FreeSans 80 0 0 0 A0
port 0 nsew
flabel metal1 83 491 83 491 0 FreeSans 80 0 0 0 B0
port 1 nsew
flabel metal1 131 446 131 446 0 FreeSans 80 0 0 0 C0
port 2 nsew
flabel metal1 179 404 179 404 0 FreeSans 80 0 0 0 A1
port 3 nsew
flabel metal1 227 361 227 361 0 FreeSans 80 0 0 0 B1
port 4 nsew
flabel metal1 275 318 275 318 0 FreeSans 80 0 0 0 C1
port 5 nsew
flabel metal1 377 277 377 277 0 FreeSans 80 0 0 0 A2
port 6 nsew
flabel metal1 425 234 425 234 0 FreeSans 80 0 0 0 B2
port 7 nsew
flabel ndiff 217 109 217 109 0 FreeSans 80 0 0 0 net4
flabel ndiff 266 108 266 108 0 FreeSans 80 0 0 0 net5
flabel ndiff 126 108 126 108 0 FreeSans 80 0 0 0 net1
flabel ndiff 79 104 79 104 0 FreeSans 80 0 0 0 net2
flabel ndiff 466 121 466 121 0 FreeSans 80 0 0 0 net7
flabel ndiff 420 119 420 119 0 FreeSans 80 0 0 0 net8
flabel metal1 473 190 473 190 0 FreeSans 80 0 0 0 C2
port 8 nsew
<< properties >>
string FIXED_BBOX 0 0 747 769
<< end >>
