magic
tech sky130A
timestamp 1644969367
<< checkpaint >>
rect -630 -630 631 631
<< properties >>
string GDS_FILE sram_0rw2r1w_32_128_sky130A.gds
string GDS_END 2525156
string GDS_START 2524704
<< end >>
