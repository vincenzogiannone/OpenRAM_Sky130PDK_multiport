magic
tech sky130A
magscale 1 2
timestamp 1643678851
<< checkpaint >>
rect -1271 -1260 105410 56414
<< viali >>
rect 4973 4348 5007 4382
rect 4973 3426 5007 3460
rect 4973 2672 5007 2706
rect 4973 1750 5007 1784
<< metal1 >>
rect 6717 54398 6858 54426
rect 6717 54354 6745 54398
rect 6568 54326 6745 54354
rect 6717 54272 6858 54300
rect 6717 54228 6745 54272
rect 6568 54200 6745 54228
rect 6717 54046 6858 54074
rect 6717 54002 6745 54046
rect 6568 53974 6745 54002
rect 6717 52986 6858 53014
rect 6717 52962 6745 52986
rect 6568 52934 6745 52962
rect 6717 52760 6858 52788
rect 6717 52736 6745 52760
rect 6568 52708 6745 52736
rect 6717 52634 6858 52662
rect 6717 52610 6745 52634
rect 6568 52582 6745 52610
rect 6717 51318 6858 51346
rect 6717 51278 6745 51318
rect 6568 51250 6745 51278
rect 6717 51192 6858 51220
rect 6717 51152 6745 51192
rect 6568 51124 6745 51152
rect 6717 50966 6858 50994
rect 6717 50926 6745 50966
rect 6568 50898 6745 50926
rect 6717 49906 6858 49934
rect 6717 49886 6745 49906
rect 6568 49858 6745 49886
rect 6717 49680 6858 49708
rect 6717 49660 6745 49680
rect 6568 49632 6745 49660
rect 6717 49554 6858 49582
rect 6717 49534 6745 49554
rect 6568 49506 6745 49534
rect 6717 48238 6858 48266
rect 6717 48202 6745 48238
rect 6568 48174 6745 48202
rect 6717 48112 6858 48140
rect 6717 48076 6745 48112
rect 6568 48048 6745 48076
rect 6717 47886 6858 47914
rect 6717 47850 6745 47886
rect 6568 47822 6745 47850
rect 6717 46826 6858 46854
rect 6717 46810 6745 46826
rect 6568 46782 6745 46810
rect 6717 46600 6858 46628
rect 6717 46584 6745 46600
rect 6568 46556 6745 46584
rect 6717 46474 6858 46502
rect 6717 46458 6745 46474
rect 6568 46430 6745 46458
rect 6717 45158 6858 45186
rect 6717 45126 6745 45158
rect 6568 45098 6745 45126
rect 6717 45032 6858 45060
rect 6717 45000 6745 45032
rect 6568 44972 6745 45000
rect 6717 44806 6858 44834
rect 6717 44774 6745 44806
rect 6568 44746 6745 44774
rect 6717 43746 6858 43774
rect 6717 43734 6745 43746
rect 6568 43706 6745 43734
rect 6717 43520 6858 43548
rect 6717 43508 6745 43520
rect 6568 43480 6745 43508
rect 6717 43394 6858 43422
rect 6717 43382 6745 43394
rect 6568 43354 6745 43382
rect 6717 42078 6858 42106
rect 6717 42050 6745 42078
rect 6568 42022 6745 42050
rect 6717 41952 6858 41980
rect 6717 41924 6745 41952
rect 6568 41896 6745 41924
rect 6717 41726 6858 41754
rect 6717 41698 6745 41726
rect 6568 41670 6745 41698
rect 6717 40666 6858 40694
rect 6717 40658 6745 40666
rect 6568 40630 6745 40658
rect 6717 40440 6858 40468
rect 6717 40432 6745 40440
rect 6568 40404 6745 40432
rect 6717 40314 6858 40342
rect 6717 40306 6745 40314
rect 6568 40278 6745 40306
rect 6717 38998 6858 39026
rect 6717 38974 6745 38998
rect 6568 38946 6745 38974
rect 6717 38872 6858 38900
rect 6717 38848 6745 38872
rect 6568 38820 6745 38848
rect 6717 38646 6858 38674
rect 6717 38622 6745 38646
rect 6568 38594 6745 38622
rect 6717 37586 6858 37614
rect 6717 37582 6745 37586
rect 6568 37554 6745 37582
rect 6717 37360 6858 37388
rect 6717 37356 6745 37360
rect 6568 37328 6745 37356
rect 6717 37234 6858 37262
rect 6717 37230 6745 37234
rect 6568 37202 6745 37230
rect 6717 35918 6858 35946
rect 6717 35898 6745 35918
rect 6568 35870 6745 35898
rect 6717 35792 6858 35820
rect 6717 35772 6745 35792
rect 6568 35744 6745 35772
rect 6717 35566 6858 35594
rect 6717 35546 6745 35566
rect 6568 35518 6745 35546
rect 6717 34506 6858 34534
rect 6568 34478 6745 34506
rect 6717 34280 6858 34308
rect 6568 34252 6745 34280
rect 6717 34154 6858 34182
rect 6568 34126 6745 34154
rect 6717 32838 6858 32866
rect 6717 32822 6745 32838
rect 6568 32794 6745 32822
rect 6717 32712 6858 32740
rect 6717 32696 6745 32712
rect 6568 32668 6745 32696
rect 6717 32486 6858 32514
rect 6717 32470 6745 32486
rect 6568 32442 6745 32470
rect 6717 31430 6858 31454
rect 6568 31426 6858 31430
rect 6568 31402 6745 31426
rect 6717 31204 6858 31228
rect 6568 31200 6858 31204
rect 6568 31176 6745 31200
rect 6717 31078 6858 31102
rect 6568 31074 6858 31078
rect 6568 31050 6745 31074
rect 6717 29758 6858 29786
rect 6717 29746 6745 29758
rect 6568 29718 6745 29746
rect 6717 29632 6858 29660
rect 6717 29620 6745 29632
rect 6568 29592 6745 29620
rect 6717 29406 6858 29434
rect 6717 29394 6745 29406
rect 6568 29366 6745 29394
rect 6717 28354 6858 28374
rect 6568 28346 6858 28354
rect 6568 28326 6745 28346
rect 6717 28128 6858 28148
rect 6568 28120 6858 28128
rect 6568 28100 6745 28120
rect 6717 28002 6858 28022
rect 6568 27994 6858 28002
rect 6568 27974 6745 27994
rect 6717 26678 6858 26706
rect 6717 26670 6745 26678
rect 6568 26642 6745 26670
rect 6717 26552 6858 26580
rect 6717 26544 6745 26552
rect 6568 26516 6745 26544
rect 6717 26326 6858 26354
rect 6717 26318 6745 26326
rect 6568 26290 6745 26318
rect 6717 25278 6858 25294
rect 6568 25266 6858 25278
rect 6568 25250 6745 25266
rect 6717 25052 6858 25068
rect 6568 25040 6858 25052
rect 6568 25024 6745 25040
rect 6717 24926 6858 24942
rect 6568 24914 6858 24926
rect 6568 24898 6745 24914
rect 6717 23598 6858 23626
rect 6717 23594 6745 23598
rect 6568 23566 6745 23594
rect 6717 23472 6858 23500
rect 6717 23468 6745 23472
rect 6568 23440 6745 23468
rect 6717 23246 6858 23274
rect 6717 23242 6745 23246
rect 6568 23214 6745 23242
rect 6717 22202 6858 22214
rect 6568 22186 6858 22202
rect 6568 22174 6745 22186
rect 6717 21976 6858 21988
rect 6568 21960 6858 21976
rect 6568 21948 6745 21960
rect 6717 21850 6858 21862
rect 6568 21834 6858 21850
rect 6568 21822 6745 21834
rect 6717 20518 6858 20546
rect 6568 20490 6745 20518
rect 6717 20392 6858 20420
rect 6568 20364 6745 20392
rect 6717 20166 6858 20194
rect 6568 20138 6745 20166
rect 6717 19126 6858 19134
rect 6568 19106 6858 19126
rect 6568 19098 6745 19106
rect 6717 18900 6858 18908
rect 6568 18880 6858 18900
rect 6568 18872 6745 18880
rect 6717 18774 6858 18782
rect 6568 18754 6858 18774
rect 6568 18746 6745 18754
rect 6717 17442 6858 17466
rect 6568 17438 6858 17442
rect 6568 17414 6745 17438
rect 6717 17316 6858 17340
rect 6568 17312 6858 17316
rect 6568 17288 6745 17312
rect 6717 17090 6858 17114
rect 6568 17086 6858 17090
rect 6568 17062 6745 17086
rect 6717 16050 6858 16054
rect 6568 16026 6858 16050
rect 6568 16022 6745 16026
rect 6717 15824 6858 15828
rect 6568 15800 6858 15824
rect 6568 15796 6745 15800
rect 6717 15698 6858 15702
rect 6568 15674 6858 15698
rect 6568 15670 6745 15674
rect 6717 14366 6858 14386
rect 6568 14358 6858 14366
rect 6568 14338 6745 14358
rect 6717 14240 6858 14260
rect 6568 14232 6858 14240
rect 6568 14212 6745 14232
rect 6717 14014 6858 14034
rect 6568 14006 6858 14014
rect 6568 13986 6745 14006
rect 6568 12946 6858 12974
rect 6568 12720 6858 12748
rect 6568 12594 6858 12622
rect 6717 11290 6858 11306
rect 6568 11278 6858 11290
rect 6568 11262 6745 11278
rect 6717 11164 6858 11180
rect 6568 11152 6858 11164
rect 6568 11136 6745 11152
rect 6717 10938 6858 10954
rect 6568 10926 6858 10938
rect 6568 10910 6745 10926
rect 6568 9894 6745 9898
rect 6568 9870 6858 9894
rect 6717 9866 6858 9870
rect 6568 9668 6745 9672
rect 6568 9644 6858 9668
rect 6717 9640 6858 9644
rect 6568 9542 6745 9546
rect 6568 9518 6858 9542
rect 6717 9514 6858 9518
rect 6717 8214 6858 8226
rect 6568 8198 6858 8214
rect 6568 8186 6745 8198
rect 6717 8088 6858 8100
rect 6568 8072 6858 8088
rect 6568 8060 6745 8072
rect 6717 7862 6858 7874
rect 6568 7846 6858 7862
rect 6568 7834 6745 7846
rect 6568 6814 6745 6822
rect 6568 6794 6858 6814
rect 6717 6786 6858 6794
rect 6568 6588 6745 6596
rect 6568 6568 6858 6588
rect 6717 6560 6858 6568
rect 6568 6462 6745 6470
rect 6568 6442 6858 6462
rect 6717 6434 6858 6442
rect 6526 5338 30547 5366
rect 4961 4382 5019 4388
rect 4961 4379 4973 4382
rect 2644 4351 4973 4379
rect 4961 4348 4973 4351
rect 5007 4348 5019 4382
rect 4961 4342 5019 4348
rect 4961 3460 5019 3466
rect 4961 3457 4973 3460
rect 2702 3429 4973 3457
rect 4961 3426 4973 3429
rect 5007 3426 5019 3460
rect 4961 3420 5019 3426
rect 2528 3110 6872 3138
rect 2586 3052 6872 3080
rect 2702 2994 6872 3022
rect 2644 2936 6872 2964
rect 4961 2706 5019 2712
rect 4961 2703 4973 2706
rect 2586 2675 4973 2703
rect 4961 2672 4973 2675
rect 5007 2672 5019 2706
rect 4961 2666 5019 2672
rect 4961 1784 5019 1790
rect 4961 1781 4973 1784
rect 2528 1753 4973 1781
rect 4961 1750 4973 1753
rect 5007 1750 5019 1784
rect 4961 1744 5019 1750
rect 32143 1171 56948 1199
<< via1 >>
rect 6474 5326 6526 5378
rect 2592 4339 2644 4391
rect 2650 3417 2702 3469
rect 2476 3098 2528 3150
rect 2534 3040 2586 3092
rect 2650 2982 2702 3034
rect 2592 2924 2644 2976
rect 2534 2663 2586 2715
rect 2476 1741 2528 1793
rect 56948 1159 57000 1211
<< metal2 >>
rect 5364 54992 5392 55020
rect 1 5790 29 36582
rect 69 5790 97 36582
rect 137 5790 165 36582
rect 205 5790 233 36582
rect 273 5790 301 36582
rect 341 5790 369 36582
rect 409 5790 437 36582
rect 6486 5378 6514 5722
rect 7054 5422 7108 5450
rect 10166 5422 10220 5450
rect 13278 5422 13332 5450
rect 16390 5422 16444 5450
rect 19502 5422 19556 5450
rect 22614 5422 22668 5450
rect 25726 5422 25780 5450
rect 28838 5422 28892 5450
rect 31950 5422 32004 5450
rect 35062 5422 35116 5450
rect 38174 5422 38228 5450
rect 41286 5422 41340 5450
rect 44398 5422 44452 5450
rect 47510 5422 47564 5450
rect 50622 5422 50676 5450
rect 53734 5422 53788 5450
rect 2488 1793 2516 3098
rect 2546 2715 2574 3040
rect 2604 2976 2632 4339
rect 2662 3034 2690 3417
rect 3089 2674 3119 2704
rect 2965 1752 2995 1782
rect 6486 0 6514 5326
rect 7608 4326 7636 4566
rect 10720 4326 10748 4566
rect 13832 4326 13860 4566
rect 16944 4326 16972 4566
rect 20056 4326 20084 4566
rect 23168 4326 23196 4566
rect 26280 4326 26308 4566
rect 29392 4326 29420 4566
rect 32504 4326 32532 4566
rect 35616 4326 35644 4566
rect 38728 4326 38756 4566
rect 41840 4326 41868 4566
rect 44952 4326 44980 4566
rect 48064 4326 48092 4566
rect 51176 4326 51204 4566
rect 54288 4326 54316 4566
rect 56960 1211 56988 55154
rect 56960 0 56988 1159
<< metal3 >>
rect 6502 54973 6634 55039
rect 5298 54205 5430 54271
rect 6502 53435 6634 53501
rect 5298 52691 5430 52757
rect 6502 51897 6634 51963
rect 5298 51177 5430 51243
rect 6502 50359 6634 50425
rect 5298 49663 5430 49729
rect 6502 48821 6634 48887
rect 5298 48149 5430 48215
rect 6502 47283 6634 47349
rect 5298 46635 5430 46701
rect 6502 45745 6634 45811
rect 5298 45121 5430 45187
rect 6502 44207 6634 44273
rect 5298 43607 5430 43673
rect 6502 42669 6634 42735
rect 5298 42093 5430 42159
rect 6502 41131 6634 41197
rect 5298 40579 5430 40645
rect 6502 39593 6634 39659
rect 5298 39065 5430 39131
rect 6502 38055 6634 38121
rect 5298 37551 5430 37617
rect 751 36549 883 36615
rect 1646 36549 1778 36615
rect 6502 36517 6634 36583
rect 5298 36037 5430 36103
rect 751 35009 883 35075
rect 1646 35009 1778 35075
rect 6502 34979 6634 35045
rect 5298 34523 5430 34589
rect 751 33469 883 33535
rect 1646 33469 1778 33535
rect 6502 33441 6634 33507
rect 5298 33009 5430 33075
rect 751 31929 883 31995
rect 1646 31929 1778 31995
rect 6502 31903 6634 31969
rect 5298 31495 5430 31561
rect 751 30389 883 30455
rect 1646 30389 1778 30455
rect 6502 30365 6634 30431
rect 5298 29981 5430 30047
rect 751 28849 883 28915
rect 1646 28849 1778 28915
rect 6502 28827 6634 28893
rect 5298 28467 5430 28533
rect 751 27309 883 27375
rect 1646 27309 1778 27375
rect 6502 27289 6634 27355
rect 5298 26953 5430 27019
rect 751 25769 883 25835
rect 1646 25769 1778 25835
rect 6502 25751 6634 25817
rect 5298 25439 5430 25505
rect 751 24229 883 24295
rect 1646 24229 1778 24295
rect 6502 24213 6634 24279
rect 5298 23925 5430 23991
rect 6502 22675 6634 22741
rect 5298 22411 5430 22477
rect 1045 21153 1177 21219
rect 1804 21153 1936 21219
rect 6502 21137 6634 21203
rect 5298 20897 5430 20963
rect 1045 19613 1177 19679
rect 1804 19613 1936 19679
rect 6502 19599 6634 19665
rect 5298 19383 5430 19449
rect 1045 18073 1177 18139
rect 1804 18073 1936 18139
rect 6502 18061 6634 18127
rect 5298 17869 5430 17935
rect 1045 16533 1177 16599
rect 1804 16533 1936 16599
rect 6502 16523 6634 16589
rect 5298 16355 5430 16421
rect 1045 14993 1177 15059
rect 1804 14993 1936 15059
rect 6502 14985 6634 15051
rect 5298 14841 5430 14907
rect 6502 13447 6634 13513
rect 5298 13327 5430 13393
rect 1045 11917 1177 11983
rect 1804 11917 1936 11983
rect 6502 11909 6634 11975
rect 5298 11813 5430 11879
rect 1045 10377 1177 10443
rect 1804 10377 1936 10443
rect 6502 10371 6634 10437
rect 5298 10299 5430 10365
rect 1045 8837 1177 8903
rect 1804 8837 1936 8903
rect 5298 8785 5430 8851
rect 6502 8833 6634 8899
rect 1045 7297 1177 7363
rect 1804 7297 1936 7363
rect 5298 7271 5430 7337
rect 6502 7295 6634 7361
rect 1045 5757 1177 5823
rect 1804 5757 1936 5823
rect 5298 5757 5430 5823
rect 6502 5757 6634 5823
rect 7174 5614 7240 5746
rect 10286 5614 10352 5746
rect 13398 5614 13464 5746
rect 16510 5614 16576 5746
rect 19622 5614 19688 5746
rect 22734 5614 22800 5746
rect 25846 5614 25912 5746
rect 28958 5614 29024 5746
rect 32070 5614 32136 5746
rect 35182 5614 35248 5746
rect 38294 5614 38360 5746
rect 41406 5614 41472 5746
rect 44518 5614 44584 5746
rect 47630 5614 47696 5746
rect 50742 5614 50808 5746
rect 53854 5614 53920 5746
rect 7174 4782 7240 4914
rect 10286 4782 10352 4914
rect 13398 4782 13464 4914
rect 16510 4782 16576 4914
rect 19622 4782 19688 4914
rect 22734 4782 22800 4914
rect 25846 4782 25912 4914
rect 28958 4782 29024 4914
rect 32070 4782 32136 4914
rect 35182 4782 35248 4914
rect 38294 4782 38360 4914
rect 41406 4782 41472 4914
rect 44518 4782 44584 4914
rect 47630 4782 47696 4914
rect 50742 4782 50808 4914
rect 53854 4782 53920 4914
rect 3212 4709 3344 4775
rect 4307 4709 4439 4775
rect 7476 4499 7608 4565
rect 10588 4499 10720 4565
rect 13700 4499 13832 4565
rect 16812 4499 16944 4565
rect 19924 4499 20056 4565
rect 23036 4499 23168 4565
rect 26148 4499 26280 4565
rect 29260 4499 29392 4565
rect 32372 4499 32504 4565
rect 35484 4499 35616 4565
rect 38596 4499 38728 4565
rect 41708 4499 41840 4565
rect 44820 4499 44952 4565
rect 47932 4499 48064 4565
rect 51044 4499 51176 4565
rect 54156 4499 54288 4565
rect 57268 4499 57400 4565
rect 60380 4499 60512 4565
rect 63492 4499 63624 4565
rect 66604 4499 66736 4565
rect 69716 4499 69848 4565
rect 72828 4499 72960 4565
rect 75940 4499 76072 4565
rect 79052 4499 79184 4565
rect 82164 4499 82296 4565
rect 85276 4499 85408 4565
rect 88388 4499 88520 4565
rect 91500 4499 91632 4565
rect 94612 4499 94744 4565
rect 97724 4499 97856 4565
rect 100836 4499 100968 4565
rect 103948 4499 104080 4565
rect 3212 3871 3344 3937
rect 4307 3871 4439 3937
rect 7476 3553 7608 3619
rect 10588 3553 10720 3619
rect 13700 3553 13832 3619
rect 16812 3553 16944 3619
rect 19924 3553 20056 3619
rect 23036 3553 23168 3619
rect 26148 3553 26280 3619
rect 29260 3553 29392 3619
rect 32372 3553 32504 3619
rect 35484 3553 35616 3619
rect 38596 3553 38728 3619
rect 41708 3553 41840 3619
rect 44820 3553 44952 3619
rect 47932 3553 48064 3619
rect 51044 3553 51176 3619
rect 54156 3553 54288 3619
rect 57268 3553 57400 3619
rect 60380 3553 60512 3619
rect 63492 3553 63624 3619
rect 66604 3553 66736 3619
rect 69716 3553 69848 3619
rect 72828 3553 72960 3619
rect 75940 3553 76072 3619
rect 79052 3553 79184 3619
rect 82164 3553 82296 3619
rect 85276 3553 85408 3619
rect 88388 3553 88520 3619
rect 91500 3553 91632 3619
rect 94612 3553 94744 3619
rect 97724 3553 97856 3619
rect 100836 3553 100968 3619
rect 103948 3553 104080 3619
rect 3212 3033 3344 3099
rect 4307 3033 4439 3099
rect 3212 2195 3344 2261
rect 4307 2195 4439 2261
rect 7570 2114 7702 2180
rect 8348 2114 8480 2180
rect 9126 2114 9258 2180
rect 9904 2114 10036 2180
rect 10682 2114 10814 2180
rect 11460 2114 11592 2180
rect 12238 2114 12370 2180
rect 13016 2114 13148 2180
rect 13794 2114 13926 2180
rect 14572 2114 14704 2180
rect 15350 2114 15482 2180
rect 16128 2114 16260 2180
rect 16906 2114 17038 2180
rect 17684 2114 17816 2180
rect 18462 2114 18594 2180
rect 19240 2114 19372 2180
rect 20018 2114 20150 2180
rect 20796 2114 20928 2180
rect 21574 2114 21706 2180
rect 22352 2114 22484 2180
rect 23130 2114 23262 2180
rect 23908 2114 24040 2180
rect 24686 2114 24818 2180
rect 25464 2114 25596 2180
rect 26242 2114 26374 2180
rect 27020 2114 27152 2180
rect 27798 2114 27930 2180
rect 28576 2114 28708 2180
rect 29354 2114 29486 2180
rect 30132 2114 30264 2180
rect 30910 2114 31042 2180
rect 31688 2114 31820 2180
rect 32466 2114 32598 2180
rect 33244 2114 33376 2180
rect 34022 2114 34154 2180
rect 34800 2114 34932 2180
rect 35578 2114 35710 2180
rect 36356 2114 36488 2180
rect 37134 2114 37266 2180
rect 37912 2114 38044 2180
rect 38690 2114 38822 2180
rect 39468 2114 39600 2180
rect 40246 2114 40378 2180
rect 41024 2114 41156 2180
rect 41802 2114 41934 2180
rect 42580 2114 42712 2180
rect 43358 2114 43490 2180
rect 44136 2114 44268 2180
rect 44914 2114 45046 2180
rect 45692 2114 45824 2180
rect 46470 2114 46602 2180
rect 47248 2114 47380 2180
rect 48026 2114 48158 2180
rect 48804 2114 48936 2180
rect 49582 2114 49714 2180
rect 50360 2114 50492 2180
rect 51138 2114 51270 2180
rect 51916 2114 52048 2180
rect 52694 2114 52826 2180
rect 53472 2114 53604 2180
rect 54250 2114 54382 2180
rect 55028 2114 55160 2180
rect 55806 2114 55938 2180
rect 56584 2114 56716 2180
rect 3212 1357 3344 1423
rect 4307 1357 4439 1423
rect 7018 248 7084 380
rect 7796 248 7862 380
rect 8574 248 8640 380
rect 9352 248 9418 380
rect 10130 248 10196 380
rect 10908 248 10974 380
rect 11686 248 11752 380
rect 12464 248 12530 380
rect 13242 248 13308 380
rect 14020 248 14086 380
rect 14798 248 14864 380
rect 15576 248 15642 380
rect 16354 248 16420 380
rect 17132 248 17198 380
rect 17910 248 17976 380
rect 18688 248 18754 380
rect 19466 248 19532 380
rect 20244 248 20310 380
rect 21022 248 21088 380
rect 21800 248 21866 380
rect 22578 248 22644 380
rect 23356 248 23422 380
rect 24134 248 24200 380
rect 24912 248 24978 380
rect 25690 248 25756 380
rect 26468 248 26534 380
rect 27246 248 27312 380
rect 28024 248 28090 380
rect 28802 248 28868 380
rect 29580 248 29646 380
rect 30358 248 30424 380
rect 31136 248 31202 380
rect 31914 248 31980 380
rect 32692 248 32758 380
rect 33470 248 33536 380
rect 34248 248 34314 380
rect 35026 248 35092 380
rect 35804 248 35870 380
rect 36582 248 36648 380
rect 37360 248 37426 380
rect 38138 248 38204 380
rect 38916 248 38982 380
rect 39694 248 39760 380
rect 40472 248 40538 380
rect 41250 248 41316 380
rect 42028 248 42094 380
rect 42806 248 42872 380
rect 43584 248 43650 380
rect 44362 248 44428 380
rect 45140 248 45206 380
rect 45918 248 45984 380
rect 46696 248 46762 380
rect 47474 248 47540 380
rect 48252 248 48318 380
rect 49030 248 49096 380
rect 49808 248 49874 380
rect 50586 248 50652 380
rect 51364 248 51430 380
rect 52142 248 52208 380
rect 52920 248 52986 380
rect 53698 248 53764 380
rect 54476 248 54542 380
rect 55254 248 55320 380
rect 56032 248 56098 380
rect 56810 248 56876 380
use contact_17  contact_17_0
timestamp 1643678851
transform 1 0 56959 0 1 1170
box 0 0 1 1
use contact_17  contact_17_1
timestamp 1643678851
transform 1 0 6485 0 1 5337
box 0 0 1 1
use contact_17  contact_17_2
timestamp 1643678851
transform 1 0 2661 0 1 2993
box 0 0 1 1
use contact_13  contact_13_0
timestamp 1643678851
transform 1 0 4961 0 1 3420
box 0 0 1 1
use contact_17  contact_17_3
timestamp 1643678851
transform 1 0 2661 0 1 3428
box 0 0 1 1
use contact_17  contact_17_4
timestamp 1643678851
transform 1 0 2603 0 1 2935
box 0 0 1 1
use contact_13  contact_13_1
timestamp 1643678851
transform 1 0 4961 0 1 4342
box 0 0 1 1
use contact_17  contact_17_5
timestamp 1643678851
transform 1 0 2603 0 1 4350
box 0 0 1 1
use contact_17  contact_17_6
timestamp 1643678851
transform 1 0 2545 0 1 3051
box 0 0 1 1
use contact_13  contact_13_2
timestamp 1643678851
transform 1 0 4961 0 1 2666
box 0 0 1 1
use contact_17  contact_17_7
timestamp 1643678851
transform 1 0 2545 0 1 2674
box 0 0 1 1
use contact_17  contact_17_8
timestamp 1643678851
transform 1 0 2487 0 1 3109
box 0 0 1 1
use contact_13  contact_13_3
timestamp 1643678851
transform 1 0 4961 0 1 1744
box 0 0 1 1
use contact_17  contact_17_9
timestamp 1643678851
transform 1 0 2487 0 1 1752
box 0 0 1 1
use hierarchical_predecode2x4_0  hierarchical_predecode2x4_0_0
timestamp 1643678851
transform 1 0 2842 0 1 1390
box 0 -34 2356 3386
use port_address  port_address_0
timestamp 1643678851
transform 1 0 0 0 1 5790
box -11 -42 6634 49258
use port_data  port_data_0
timestamp 1643678851
transform 1 0 6858 0 1 0
box 0 190 97292 5746
use replica_bitcell_array  replica_bitcell_array_0
timestamp 1643678851
transform 1 0 6858 0 1 5790
box 0 -42 49792 49322
<< labels >>
rlabel metal2 s 6486 0 6514 5722 4 w_en
rlabel metal2 s 5364 54992 5392 55020 4 wl_en
rlabel metal2 s 56960 0 56988 55154 4 p_en_bar
rlabel metal2 s 7054 5422 7108 5450 4 din0_0
rlabel metal2 s 10166 5422 10220 5450 4 din0_1
rlabel metal2 s 13278 5422 13332 5450 4 din0_2
rlabel metal2 s 16390 5422 16444 5450 4 din0_3
rlabel metal2 s 19502 5422 19556 5450 4 din0_4
rlabel metal2 s 22614 5422 22668 5450 4 din0_5
rlabel metal2 s 25726 5422 25780 5450 4 din0_6
rlabel metal2 s 28838 5422 28892 5450 4 din0_7
rlabel metal2 s 31950 5422 32004 5450 4 din0_8
rlabel metal2 s 35062 5422 35116 5450 4 din0_9
rlabel metal2 s 38174 5422 38228 5450 4 din0_10
rlabel metal2 s 41286 5422 41340 5450 4 din0_11
rlabel metal2 s 44398 5422 44452 5450 4 din0_12
rlabel metal2 s 47510 5422 47564 5450 4 din0_13
rlabel metal2 s 50622 5422 50676 5450 4 din0_14
rlabel metal2 s 53734 5422 53788 5450 4 din0_15
rlabel metal2 s 7608 4326 7636 4566 4 dout0_0
rlabel metal2 s 7622 4446 7622 4446 4 dout1_0
rlabel metal2 s 10720 4326 10748 4566 4 dout0_1
rlabel metal2 s 10734 4446 10734 4446 4 dout1_1
rlabel metal2 s 13832 4326 13860 4566 4 dout0_2
rlabel metal2 s 13846 4446 13846 4446 4 dout1_2
rlabel metal2 s 16944 4326 16972 4566 4 dout0_3
rlabel metal2 s 16958 4446 16958 4446 4 dout1_3
rlabel metal2 s 20056 4326 20084 4566 4 dout0_4
rlabel metal2 s 20070 4446 20070 4446 4 dout1_4
rlabel metal2 s 23168 4326 23196 4566 4 dout0_5
rlabel metal2 s 23182 4446 23182 4446 4 dout1_5
rlabel metal2 s 26280 4326 26308 4566 4 dout0_6
rlabel metal2 s 26294 4446 26294 4446 4 dout1_6
rlabel metal2 s 29392 4326 29420 4566 4 dout0_7
rlabel metal2 s 29406 4446 29406 4446 4 dout1_7
rlabel metal2 s 32504 4326 32532 4566 4 dout0_8
rlabel metal2 s 32518 4446 32518 4446 4 dout1_8
rlabel metal2 s 35616 4326 35644 4566 4 dout0_9
rlabel metal2 s 35630 4446 35630 4446 4 dout1_9
rlabel metal2 s 38728 4326 38756 4566 4 dout0_10
rlabel metal2 s 38742 4446 38742 4446 4 dout1_10
rlabel metal2 s 41840 4326 41868 4566 4 dout0_11
rlabel metal2 s 41854 4446 41854 4446 4 dout1_11
rlabel metal2 s 44952 4326 44980 4566 4 dout0_12
rlabel metal2 s 44966 4446 44966 4446 4 dout1_12
rlabel metal2 s 48064 4326 48092 4566 4 dout0_13
rlabel metal2 s 48078 4446 48078 4446 4 dout1_13
rlabel metal2 s 51176 4326 51204 4566 4 dout0_14
rlabel metal2 s 51190 4446 51190 4446 4 dout1_14
rlabel metal2 s 54288 4326 54316 4566 4 dout0_15
rlabel metal2 s 54302 4446 54302 4446 4 dout1_15
rlabel metal2 s 0 5790 28 36582 4 addr2
rlabel metal2 s 68 5790 96 36582 4 addr3
rlabel metal2 s 136 5790 164 36582 4 addr4
rlabel metal2 s 204 5790 232 36582 4 addr5
rlabel metal2 s 272 5790 300 36582 4 addr6
rlabel metal2 s 340 5790 368 36582 4 addr7
rlabel metal2 s 408 5790 436 36582 4 addr8
rlabel metal2 s 2964 1752 2994 1782 4 addr0
rlabel metal2 s 3088 2674 3118 2704 4 addr1
rlabel metal3 s 1804 10376 1936 10442 4 vdd
rlabel metal3 s 38916 248 38982 380 4 vdd
rlabel metal3 s 35484 3552 35616 3618 4 vdd
rlabel metal3 s 32692 248 32758 380 4 vdd
rlabel metal3 s 54156 3552 54288 3618 4 vdd
rlabel metal3 s 47630 4782 47696 4914 4 vdd
rlabel metal3 s 6502 13446 6634 13512 4 vdd
rlabel metal3 s 10588 3552 10720 3618 4 vdd
rlabel metal3 s 23036 3552 23168 3618 4 vdd
rlabel metal3 s 35182 4782 35248 4914 4 vdd
rlabel metal3 s 5298 40578 5430 40644 4 vdd
rlabel metal3 s 49808 248 49874 380 4 vdd
rlabel metal3 s 7476 3552 7608 3618 4 vdd
rlabel metal3 s 88388 3552 88520 3618 4 vdd
rlabel metal3 s 47932 3552 48064 3618 4 vdd
rlabel metal3 s 6502 19598 6634 19664 4 vdd
rlabel metal3 s 6502 44206 6634 44272 4 vdd
rlabel metal3 s 41250 248 41316 380 4 vdd
rlabel metal3 s 24134 248 24200 380 4 vdd
rlabel metal3 s 91500 3552 91632 3618 4 vdd
rlabel metal3 s 63492 3552 63624 3618 4 vdd
rlabel metal3 s 18688 248 18754 380 4 vdd
rlabel metal3 s 13398 4782 13464 4914 4 vdd
rlabel metal3 s 56810 248 56876 380 4 vdd
rlabel metal3 s 12464 248 12530 380 4 vdd
rlabel metal3 s 10130 248 10196 380 4 vdd
rlabel metal3 s 30358 248 30424 380 4 vdd
rlabel metal3 s 40472 248 40538 380 4 vdd
rlabel metal3 s 27246 248 27312 380 4 vdd
rlabel metal3 s 6502 50358 6634 50424 4 vdd
rlabel metal3 s 19622 4782 19688 4914 4 vdd
rlabel metal3 s 5298 46634 5430 46700 4 vdd
rlabel metal3 s 42806 248 42872 380 4 vdd
rlabel metal3 s 13242 248 13308 380 4 vdd
rlabel metal3 s 44362 248 44428 380 4 vdd
rlabel metal3 s 1804 19612 1936 19678 4 vdd
rlabel metal3 s 5298 10298 5430 10364 4 vdd
rlabel metal3 s 6502 22674 6634 22740 4 vdd
rlabel metal3 s 36582 248 36648 380 4 vdd
rlabel metal3 s 25690 248 25756 380 4 vdd
rlabel metal3 s 3212 2194 3344 2260 4 vdd
rlabel metal3 s 69716 3552 69848 3618 4 vdd
rlabel metal3 s 21022 248 21088 380 4 vdd
rlabel metal3 s 51044 3552 51176 3618 4 vdd
rlabel metal3 s 6502 16522 6634 16588 4 vdd
rlabel metal3 s 37360 248 37426 380 4 vdd
rlabel metal3 s 17132 248 17198 380 4 vdd
rlabel metal3 s 14798 248 14864 380 4 vdd
rlabel metal3 s 85276 3552 85408 3618 4 vdd
rlabel metal3 s 94612 3552 94744 3618 4 vdd
rlabel metal3 s 750 25768 882 25834 4 vdd
rlabel metal3 s 26148 3552 26280 3618 4 vdd
rlabel metal3 s 6502 31902 6634 31968 4 vdd
rlabel metal3 s 10908 248 10974 380 4 vdd
rlabel metal3 s 52142 248 52208 380 4 vdd
rlabel metal3 s 21800 248 21866 380 4 vdd
rlabel metal3 s 39694 248 39760 380 4 vdd
rlabel metal3 s 1646 31928 1778 31994 4 vdd
rlabel metal3 s 38138 248 38204 380 4 vdd
rlabel metal3 s 28958 4782 29024 4914 4 vdd
rlabel metal3 s 50742 4782 50808 4914 4 vdd
rlabel metal3 s 31914 248 31980 380 4 vdd
rlabel metal3 s 57268 3552 57400 3618 4 vdd
rlabel metal3 s 29260 3552 29392 3618 4 vdd
rlabel metal3 s 45140 248 45206 380 4 vdd
rlabel metal3 s 750 28848 882 28914 4 vdd
rlabel metal3 s 43584 248 43650 380 4 vdd
rlabel metal3 s 79052 3552 79184 3618 4 vdd
rlabel metal3 s 35026 248 35092 380 4 vdd
rlabel metal3 s 26468 248 26534 380 4 vdd
rlabel metal3 s 60380 3552 60512 3618 4 vdd
rlabel metal3 s 16510 4782 16576 4914 4 vdd
rlabel metal3 s 4306 3870 4438 3936 4 vdd
rlabel metal3 s 6502 7294 6634 7360 4 vdd
rlabel metal3 s 25846 4782 25912 4914 4 vdd
rlabel metal3 s 100836 3552 100968 3618 4 vdd
rlabel metal3 s 9352 248 9418 380 4 vdd
rlabel metal3 s 44518 4782 44584 4914 4 vdd
rlabel metal3 s 55254 248 55320 380 4 vdd
rlabel metal3 s 19924 3552 20056 3618 4 vdd
rlabel metal3 s 1804 7296 1936 7362 4 vdd
rlabel metal3 s 6502 38054 6634 38120 4 vdd
rlabel metal3 s 35804 248 35870 380 4 vdd
rlabel metal3 s 34248 248 34314 380 4 vdd
rlabel metal3 s 22578 248 22644 380 4 vdd
rlabel metal3 s 8574 248 8640 380 4 vdd
rlabel metal3 s 11686 248 11752 380 4 vdd
rlabel metal3 s 5298 25438 5430 25504 4 vdd
rlabel metal3 s 1646 35008 1778 35074 4 vdd
rlabel metal3 s 66604 3552 66736 3618 4 vdd
rlabel metal3 s 54476 248 54542 380 4 vdd
rlabel metal3 s 1646 25768 1778 25834 4 vdd
rlabel metal3 s 750 35008 882 35074 4 vdd
rlabel metal3 s 41406 4782 41472 4914 4 vdd
rlabel metal3 s 1804 16532 1936 16598 4 vdd
rlabel metal3 s 15576 248 15642 380 4 vdd
rlabel metal3 s 49030 248 49096 380 4 vdd
rlabel metal3 s 7018 248 7084 380 4 vdd
rlabel metal3 s 16812 3552 16944 3618 4 vdd
rlabel metal3 s 19466 248 19532 380 4 vdd
rlabel metal3 s 6502 53434 6634 53500 4 vdd
rlabel metal3 s 51364 248 51430 380 4 vdd
rlabel metal3 s 45918 248 45984 380 4 vdd
rlabel metal3 s 97724 3552 97856 3618 4 vdd
rlabel metal3 s 24912 248 24978 380 4 vdd
rlabel metal3 s 53698 248 53764 380 4 vdd
rlabel metal3 s 16354 248 16420 380 4 vdd
rlabel metal3 s 75940 3552 76072 3618 4 vdd
rlabel metal3 s 31136 248 31202 380 4 vdd
rlabel metal3 s 38294 4782 38360 4914 4 vdd
rlabel metal3 s 47474 248 47540 380 4 vdd
rlabel metal3 s 56032 248 56098 380 4 vdd
rlabel metal3 s 48252 248 48318 380 4 vdd
rlabel metal3 s 1044 19612 1176 19678 4 vdd
rlabel metal3 s 5298 52690 5430 52756 4 vdd
rlabel metal3 s 7174 4782 7240 4914 4 vdd
rlabel metal3 s 5298 31494 5430 31560 4 vdd
rlabel metal3 s 17910 248 17976 380 4 vdd
rlabel metal3 s 5298 34522 5430 34588 4 vdd
rlabel metal3 s 750 31928 882 31994 4 vdd
rlabel metal3 s 5298 19382 5430 19448 4 vdd
rlabel metal3 s 32372 3552 32504 3618 4 vdd
rlabel metal3 s 41708 3552 41840 3618 4 vdd
rlabel metal3 s 29580 248 29646 380 4 vdd
rlabel metal3 s 32070 4782 32136 4914 4 vdd
rlabel metal3 s 6502 47282 6634 47348 4 vdd
rlabel metal3 s 1646 28848 1778 28914 4 vdd
rlabel metal3 s 3212 3870 3344 3936 4 vdd
rlabel metal3 s 6502 34978 6634 35044 4 vdd
rlabel metal3 s 1044 10376 1176 10442 4 vdd
rlabel metal3 s 20244 248 20310 380 4 vdd
rlabel metal3 s 5298 16354 5430 16420 4 vdd
rlabel metal3 s 5298 7270 5430 7336 4 vdd
rlabel metal3 s 5298 28466 5430 28532 4 vdd
rlabel metal3 s 6502 41130 6634 41196 4 vdd
rlabel metal3 s 5298 37550 5430 37616 4 vdd
rlabel metal3 s 1044 16532 1176 16598 4 vdd
rlabel metal3 s 10286 4782 10352 4914 4 vdd
rlabel metal3 s 38596 3552 38728 3618 4 vdd
rlabel metal3 s 14020 248 14086 380 4 vdd
rlabel metal3 s 6502 25750 6634 25816 4 vdd
rlabel metal3 s 23356 248 23422 380 4 vdd
rlabel metal3 s 4306 2194 4438 2260 4 vdd
rlabel metal3 s 42028 248 42094 380 4 vdd
rlabel metal3 s 52920 248 52986 380 4 vdd
rlabel metal3 s 46696 248 46762 380 4 vdd
rlabel metal3 s 5298 13326 5430 13392 4 vdd
rlabel metal3 s 1044 7296 1176 7362 4 vdd
rlabel metal3 s 6502 28826 6634 28892 4 vdd
rlabel metal3 s 22734 4782 22800 4914 4 vdd
rlabel metal3 s 13700 3552 13832 3618 4 vdd
rlabel metal3 s 72828 3552 72960 3618 4 vdd
rlabel metal3 s 33470 248 33536 380 4 vdd
rlabel metal3 s 28024 248 28090 380 4 vdd
rlabel metal3 s 53854 4782 53920 4914 4 vdd
rlabel metal3 s 5298 49662 5430 49728 4 vdd
rlabel metal3 s 103948 3552 104080 3618 4 vdd
rlabel metal3 s 6502 10370 6634 10436 4 vdd
rlabel metal3 s 28802 248 28868 380 4 vdd
rlabel metal3 s 7796 248 7862 380 4 vdd
rlabel metal3 s 82164 3552 82296 3618 4 vdd
rlabel metal3 s 44820 3552 44952 3618 4 vdd
rlabel metal3 s 50586 248 50652 380 4 vdd
rlabel metal3 s 5298 43606 5430 43672 4 vdd
rlabel metal3 s 5298 22410 5430 22476 4 vdd
rlabel metal3 s 35484 4498 35616 4564 4 gnd
rlabel metal3 s 41024 2114 41156 2180 4 gnd
rlabel metal3 s 32070 5614 32136 5746 4 gnd
rlabel metal3 s 26148 4498 26280 4564 4 gnd
rlabel metal3 s 63492 4498 63624 4564 4 gnd
rlabel metal3 s 6502 36516 6634 36582 4 gnd
rlabel metal3 s 5298 20896 5430 20962 4 gnd
rlabel metal3 s 5298 54204 5430 54270 4 gnd
rlabel metal3 s 5298 8784 5430 8850 4 gnd
rlabel metal3 s 5298 29980 5430 30046 4 gnd
rlabel metal3 s 19622 5614 19688 5746 4 gnd
rlabel metal3 s 40246 2114 40378 2180 4 gnd
rlabel metal3 s 26242 2114 26374 2180 4 gnd
rlabel metal3 s 10286 5614 10352 5746 4 gnd
rlabel metal3 s 23130 2114 23262 2180 4 gnd
rlabel metal3 s 19240 2114 19372 2180 4 gnd
rlabel metal3 s 5298 45120 5430 45186 4 gnd
rlabel metal3 s 47248 2114 47380 2180 4 gnd
rlabel metal3 s 5298 26952 5430 27018 4 gnd
rlabel metal3 s 6502 54972 6634 55038 4 gnd
rlabel metal3 s 60380 4498 60512 4564 4 gnd
rlabel metal3 s 22352 2114 22484 2180 4 gnd
rlabel metal3 s 44136 2114 44268 2180 4 gnd
rlabel metal3 s 13700 4498 13832 4564 4 gnd
rlabel metal3 s 8348 2114 8480 2180 4 gnd
rlabel metal3 s 28576 2114 28708 2180 4 gnd
rlabel metal3 s 48026 2114 48158 2180 4 gnd
rlabel metal3 s 1646 27308 1778 27374 4 gnd
rlabel metal3 s 69716 4498 69848 4564 4 gnd
rlabel metal3 s 20796 2114 20928 2180 4 gnd
rlabel metal3 s 49582 2114 49714 2180 4 gnd
rlabel metal3 s 9126 2114 9258 2180 4 gnd
rlabel metal3 s 29260 4498 29392 4564 4 gnd
rlabel metal3 s 3212 3032 3344 3098 4 gnd
rlabel metal3 s 6502 5756 6634 5822 4 gnd
rlabel metal3 s 44820 4498 44952 4564 4 gnd
rlabel metal3 s 44914 2114 45046 2180 4 gnd
rlabel metal3 s 33244 2114 33376 2180 4 gnd
rlabel metal3 s 25846 5614 25912 5746 4 gnd
rlabel metal3 s 47630 5614 47696 5746 4 gnd
rlabel metal3 s 10682 2114 10814 2180 4 gnd
rlabel metal3 s 19924 4498 20056 4564 4 gnd
rlabel metal3 s 15350 2114 15482 2180 4 gnd
rlabel metal3 s 88388 4498 88520 4564 4 gnd
rlabel metal3 s 50360 2114 50492 2180 4 gnd
rlabel metal3 s 1044 5756 1176 5822 4 gnd
rlabel metal3 s 1804 11916 1936 11982 4 gnd
rlabel metal3 s 28958 5614 29024 5746 4 gnd
rlabel metal3 s 35578 2114 35710 2180 4 gnd
rlabel metal3 s 53472 2114 53604 2180 4 gnd
rlabel metal3 s 6502 11908 6634 11974 4 gnd
rlabel metal3 s 750 33468 882 33534 4 gnd
rlabel metal3 s 6502 39592 6634 39658 4 gnd
rlabel metal3 s 3212 4708 3344 4774 4 gnd
rlabel metal3 s 31688 2114 31820 2180 4 gnd
rlabel metal3 s 6502 27288 6634 27354 4 gnd
rlabel metal3 s 42580 2114 42712 2180 4 gnd
rlabel metal3 s 1044 11916 1176 11982 4 gnd
rlabel metal3 s 82164 4498 82296 4564 4 gnd
rlabel metal3 s 7476 4498 7608 4564 4 gnd
rlabel metal3 s 45692 2114 45824 2180 4 gnd
rlabel metal3 s 91500 4498 91632 4564 4 gnd
rlabel metal3 s 22734 5614 22800 5746 4 gnd
rlabel metal3 s 1646 33468 1778 33534 4 gnd
rlabel metal3 s 24686 2114 24818 2180 4 gnd
rlabel metal3 s 12238 2114 12370 2180 4 gnd
rlabel metal3 s 4306 4708 4438 4774 4 gnd
rlabel metal3 s 16906 2114 17038 2180 4 gnd
rlabel metal3 s 32466 2114 32598 2180 4 gnd
rlabel metal3 s 54156 4498 54288 4564 4 gnd
rlabel metal3 s 6502 33440 6634 33506 4 gnd
rlabel metal3 s 1044 8836 1176 8902 4 gnd
rlabel metal3 s 1804 5756 1936 5822 4 gnd
rlabel metal3 s 55028 2114 55160 2180 4 gnd
rlabel metal3 s 20018 2114 20150 2180 4 gnd
rlabel metal3 s 5298 11812 5430 11878 4 gnd
rlabel metal3 s 9904 2114 10036 2180 4 gnd
rlabel metal3 s 13794 2114 13926 2180 4 gnd
rlabel metal3 s 7174 5614 7240 5746 4 gnd
rlabel metal3 s 38690 2114 38822 2180 4 gnd
rlabel metal3 s 1044 14992 1176 15058 4 gnd
rlabel metal3 s 6502 18060 6634 18126 4 gnd
rlabel metal3 s 6502 14984 6634 15050 4 gnd
rlabel metal3 s 56584 2114 56716 2180 4 gnd
rlabel metal3 s 29354 2114 29486 2180 4 gnd
rlabel metal3 s 4306 1356 4438 1422 4 gnd
rlabel metal3 s 34022 2114 34154 2180 4 gnd
rlabel metal3 s 6502 21136 6634 21202 4 gnd
rlabel metal3 s 18462 2114 18594 2180 4 gnd
rlabel metal3 s 1646 36548 1778 36614 4 gnd
rlabel metal3 s 6502 8832 6634 8898 4 gnd
rlabel metal3 s 3212 1356 3344 1422 4 gnd
rlabel metal3 s 43358 2114 43490 2180 4 gnd
rlabel metal3 s 5298 23924 5430 23990 4 gnd
rlabel metal3 s 51138 2114 51270 2180 4 gnd
rlabel metal3 s 41708 4498 41840 4564 4 gnd
rlabel metal3 s 57268 4498 57400 4564 4 gnd
rlabel metal3 s 21574 2114 21706 2180 4 gnd
rlabel metal3 s 1804 8836 1936 8902 4 gnd
rlabel metal3 s 94612 4498 94744 4564 4 gnd
rlabel metal3 s 13398 5614 13464 5746 4 gnd
rlabel metal3 s 37912 2114 38044 2180 4 gnd
rlabel metal3 s 5298 36036 5430 36102 4 gnd
rlabel metal3 s 5298 17868 5430 17934 4 gnd
rlabel metal3 s 53854 5614 53920 5746 4 gnd
rlabel metal3 s 38596 4498 38728 4564 4 gnd
rlabel metal3 s 103948 4498 104080 4564 4 gnd
rlabel metal3 s 5298 5756 5430 5822 4 gnd
rlabel metal3 s 35182 5614 35248 5746 4 gnd
rlabel metal3 s 23036 4498 23168 4564 4 gnd
rlabel metal3 s 36356 2114 36488 2180 4 gnd
rlabel metal3 s 37134 2114 37266 2180 4 gnd
rlabel metal3 s 16812 4498 16944 4564 4 gnd
rlabel metal3 s 23908 2114 24040 2180 4 gnd
rlabel metal3 s 17684 2114 17816 2180 4 gnd
rlabel metal3 s 79052 4498 79184 4564 4 gnd
rlabel metal3 s 32372 4498 32504 4564 4 gnd
rlabel metal3 s 5298 39064 5430 39130 4 gnd
rlabel metal3 s 47932 4498 48064 4564 4 gnd
rlabel metal3 s 85276 4498 85408 4564 4 gnd
rlabel metal3 s 1646 30388 1778 30454 4 gnd
rlabel metal3 s 97724 4498 97856 4564 4 gnd
rlabel metal3 s 14572 2114 14704 2180 4 gnd
rlabel metal3 s 1044 18072 1176 18138 4 gnd
rlabel metal3 s 750 36548 882 36614 4 gnd
rlabel metal3 s 13016 2114 13148 2180 4 gnd
rlabel metal3 s 51916 2114 52048 2180 4 gnd
rlabel metal3 s 52694 2114 52826 2180 4 gnd
rlabel metal3 s 10588 4498 10720 4564 4 gnd
rlabel metal3 s 39468 2114 39600 2180 4 gnd
rlabel metal3 s 51044 4498 51176 4564 4 gnd
rlabel metal3 s 100836 4498 100968 4564 4 gnd
rlabel metal3 s 5298 42092 5430 42158 4 gnd
rlabel metal3 s 6502 24212 6634 24278 4 gnd
rlabel metal3 s 30910 2114 31042 2180 4 gnd
rlabel metal3 s 55806 2114 55938 2180 4 gnd
rlabel metal3 s 5298 14840 5430 14906 4 gnd
rlabel metal3 s 5298 33008 5430 33074 4 gnd
rlabel metal3 s 5298 51176 5430 51242 4 gnd
rlabel metal3 s 25464 2114 25596 2180 4 gnd
rlabel metal3 s 1646 24228 1778 24294 4 gnd
rlabel metal3 s 6502 45744 6634 45810 4 gnd
rlabel metal3 s 41406 5614 41472 5746 4 gnd
rlabel metal3 s 50742 5614 50808 5746 4 gnd
rlabel metal3 s 16128 2114 16260 2180 4 gnd
rlabel metal3 s 46470 2114 46602 2180 4 gnd
rlabel metal3 s 6502 48820 6634 48886 4 gnd
rlabel metal3 s 41802 2114 41934 2180 4 gnd
rlabel metal3 s 44518 5614 44584 5746 4 gnd
rlabel metal3 s 4306 3032 4438 3098 4 gnd
rlabel metal3 s 7570 2114 7702 2180 4 gnd
rlabel metal3 s 1804 21152 1936 21218 4 gnd
rlabel metal3 s 750 27308 882 27374 4 gnd
rlabel metal3 s 11460 2114 11592 2180 4 gnd
rlabel metal3 s 16510 5614 16576 5746 4 gnd
rlabel metal3 s 6502 51896 6634 51962 4 gnd
rlabel metal3 s 34800 2114 34932 2180 4 gnd
rlabel metal3 s 72828 4498 72960 4564 4 gnd
rlabel metal3 s 1044 21152 1176 21218 4 gnd
rlabel metal3 s 38294 5614 38360 5746 4 gnd
rlabel metal3 s 27798 2114 27930 2180 4 gnd
rlabel metal3 s 30132 2114 30264 2180 4 gnd
rlabel metal3 s 750 24228 882 24294 4 gnd
rlabel metal3 s 54250 2114 54382 2180 4 gnd
rlabel metal3 s 1804 18072 1936 18138 4 gnd
rlabel metal3 s 27020 2114 27152 2180 4 gnd
rlabel metal3 s 750 30388 882 30454 4 gnd
rlabel metal3 s 48804 2114 48936 2180 4 gnd
rlabel metal3 s 5298 48148 5430 48214 4 gnd
rlabel metal3 s 1804 14992 1936 15058 4 gnd
rlabel metal3 s 75940 4498 76072 4564 4 gnd
rlabel metal3 s 6502 30364 6634 30430 4 gnd
rlabel metal3 s 6502 42668 6634 42734 4 gnd
rlabel metal3 s 66604 4498 66736 4564 4 gnd
<< properties >>
string FIXED_BBOX 0 0 104234 55154
string GDS_FILE sram_0rw2r1w_16_128_sky130A.gds
string GDS_END 339328
string GDS_START 232738
<< end >>
