magic
tech sky130A
timestamp 1643593061
<< checkpaint >>
rect -630 -630 726 720
<< metal1 >>
rect 0 0 3 90
rect 93 0 96 90
<< via1 >>
rect 3 0 93 90
<< properties >>
string FIXED_BBOX 0 0 96 90
string GDS_FILE sram_0rw2r1w_2_16_sky130A.gds
string GDS_END 582752
string GDS_START 581916
<< end >>
