magic
tech sky130A
magscale 1 2
timestamp 1644969367
<< checkpaint >>
rect -1260 -1286 1518 1400
<< scnmos >>
rect 60 0 90 84
rect 168 0 198 84
<< ndiff >>
rect 0 59 60 84
rect 0 25 8 59
rect 42 25 60 59
rect 0 0 60 25
rect 90 59 168 84
rect 90 25 112 59
rect 146 25 168 59
rect 90 0 168 25
rect 198 59 258 84
rect 198 25 216 59
rect 250 25 258 59
rect 198 0 258 25
<< ndiffc >>
rect 8 25 42 59
rect 112 25 146 59
rect 216 25 250 59
<< poly >>
rect 60 110 198 140
rect 60 84 90 110
rect 168 84 198 110
rect 60 -26 90 0
rect 168 -26 198 0
<< locali >>
rect 8 59 42 75
rect 8 9 42 25
rect 112 59 146 75
rect 112 9 146 25
rect 216 59 250 75
rect 216 9 250 25
use contact_8  contact_8_0
timestamp 1644969367
transform 1 0 208 0 1 1
box 0 0 1 1
use contact_8  contact_8_1
timestamp 1644969367
transform 1 0 104 0 1 1
box 0 0 1 1
use contact_8  contact_8_2
timestamp 1644969367
transform 1 0 0 0 1 1
box 0 0 1 1
<< labels >>
rlabel mvvaractor s 129 125 129 125 4 G
rlabel locali s 233 42 233 42 4 S
rlabel locali s 25 42 25 42 4 S
rlabel locali s 129 42 129 42 4 D
<< properties >>
string FIXED_BBOX -25 -26 283 140
string GDS_FILE sram_0rw2r1w_32_128_sky130A.gds
string GDS_END 3263002
string GDS_START 3262014
<< end >>
