magic
tech sky130A
magscale 1 2
timestamp 1644951705
<< checkpaint >>
rect -1296 -1277 3122 2155
<< locali >>
rect 0 821 1826 855
rect 196 381 262 447
rect 330 390 364 561
rect 330 356 459 390
rect 1099 356 1133 390
rect 96 257 162 323
rect 0 -17 1826 17
use pdriver_0  pdriver_0_0
timestamp 1644951705
transform 1 0 378 0 1 0
box -36 -17 1484 895
use pnand2_0  pnand2_0_0
timestamp 1644951705
transform 1 0 0 0 1 0
box -36 -17 414 895
<< labels >>
rlabel locali s 1116 373 1116 373 4 Z
rlabel locali s 129 290 129 290 4 A
rlabel locali s 229 414 229 414 4 B
rlabel locali s 913 0 913 0 4 gnd
rlabel locali s 913 838 913 838 4 vdd
<< properties >>
string FIXED_BBOX 0 0 1826 838
string GDS_FILE sram_0rw2r1w_16_128_sky130A.gds
string GDS_END 2020942
string GDS_START 2019808
<< end >>
