magic
tech sky130A
magscale 1 2
timestamp 1644951705
<< checkpaint >>
rect -1260 -1212 51118 3328
<< poly >>
rect 374 287 404 588
rect 1152 367 1182 588
rect 1930 447 1960 588
rect 2708 527 2738 588
rect 2690 511 2756 527
rect 2690 477 2706 511
rect 2740 477 2756 511
rect 2690 461 2756 477
rect 1912 431 1978 447
rect 1912 397 1928 431
rect 1962 397 1978 431
rect 1912 381 1978 397
rect 1134 351 1200 367
rect 1134 317 1150 351
rect 1184 317 1200 351
rect 1134 301 1200 317
rect 3486 287 3516 588
rect 4264 367 4294 588
rect 5042 447 5072 588
rect 5820 527 5850 588
rect 5802 511 5868 527
rect 5802 477 5818 511
rect 5852 477 5868 511
rect 5802 461 5868 477
rect 5024 431 5090 447
rect 5024 397 5040 431
rect 5074 397 5090 431
rect 5024 381 5090 397
rect 4246 351 4312 367
rect 4246 317 4262 351
rect 4296 317 4312 351
rect 4246 301 4312 317
rect 6598 287 6628 588
rect 7376 367 7406 588
rect 8154 447 8184 588
rect 8932 527 8962 588
rect 8914 511 8980 527
rect 8914 477 8930 511
rect 8964 477 8980 511
rect 8914 461 8980 477
rect 8136 431 8202 447
rect 8136 397 8152 431
rect 8186 397 8202 431
rect 8136 381 8202 397
rect 7358 351 7424 367
rect 7358 317 7374 351
rect 7408 317 7424 351
rect 7358 301 7424 317
rect 9710 287 9740 588
rect 10488 367 10518 588
rect 11266 447 11296 588
rect 12044 527 12074 588
rect 12026 511 12092 527
rect 12026 477 12042 511
rect 12076 477 12092 511
rect 12026 461 12092 477
rect 11248 431 11314 447
rect 11248 397 11264 431
rect 11298 397 11314 431
rect 11248 381 11314 397
rect 10470 351 10536 367
rect 10470 317 10486 351
rect 10520 317 10536 351
rect 10470 301 10536 317
rect 12822 287 12852 588
rect 13600 367 13630 588
rect 14378 447 14408 588
rect 15156 527 15186 588
rect 15138 511 15204 527
rect 15138 477 15154 511
rect 15188 477 15204 511
rect 15138 461 15204 477
rect 14360 431 14426 447
rect 14360 397 14376 431
rect 14410 397 14426 431
rect 14360 381 14426 397
rect 13582 351 13648 367
rect 13582 317 13598 351
rect 13632 317 13648 351
rect 13582 301 13648 317
rect 15934 287 15964 588
rect 16712 367 16742 588
rect 17490 447 17520 588
rect 18268 527 18298 588
rect 18250 511 18316 527
rect 18250 477 18266 511
rect 18300 477 18316 511
rect 18250 461 18316 477
rect 17472 431 17538 447
rect 17472 397 17488 431
rect 17522 397 17538 431
rect 17472 381 17538 397
rect 16694 351 16760 367
rect 16694 317 16710 351
rect 16744 317 16760 351
rect 16694 301 16760 317
rect 19046 287 19076 588
rect 19824 367 19854 588
rect 20602 447 20632 588
rect 21380 527 21410 588
rect 21362 511 21428 527
rect 21362 477 21378 511
rect 21412 477 21428 511
rect 21362 461 21428 477
rect 20584 431 20650 447
rect 20584 397 20600 431
rect 20634 397 20650 431
rect 20584 381 20650 397
rect 19806 351 19872 367
rect 19806 317 19822 351
rect 19856 317 19872 351
rect 19806 301 19872 317
rect 22158 287 22188 588
rect 22936 367 22966 588
rect 23714 447 23744 588
rect 24492 527 24522 588
rect 24474 511 24540 527
rect 24474 477 24490 511
rect 24524 477 24540 511
rect 24474 461 24540 477
rect 23696 431 23762 447
rect 23696 397 23712 431
rect 23746 397 23762 431
rect 23696 381 23762 397
rect 22918 351 22984 367
rect 22918 317 22934 351
rect 22968 317 22984 351
rect 22918 301 22984 317
rect 25270 287 25300 588
rect 26048 367 26078 588
rect 26826 447 26856 588
rect 27604 527 27634 588
rect 27586 511 27652 527
rect 27586 477 27602 511
rect 27636 477 27652 511
rect 27586 461 27652 477
rect 26808 431 26874 447
rect 26808 397 26824 431
rect 26858 397 26874 431
rect 26808 381 26874 397
rect 26030 351 26096 367
rect 26030 317 26046 351
rect 26080 317 26096 351
rect 26030 301 26096 317
rect 28382 287 28412 588
rect 29160 367 29190 588
rect 29938 447 29968 588
rect 30716 527 30746 588
rect 30698 511 30764 527
rect 30698 477 30714 511
rect 30748 477 30764 511
rect 30698 461 30764 477
rect 29920 431 29986 447
rect 29920 397 29936 431
rect 29970 397 29986 431
rect 29920 381 29986 397
rect 29142 351 29208 367
rect 29142 317 29158 351
rect 29192 317 29208 351
rect 29142 301 29208 317
rect 31494 287 31524 588
rect 32272 367 32302 588
rect 33050 447 33080 588
rect 33828 527 33858 588
rect 33810 511 33876 527
rect 33810 477 33826 511
rect 33860 477 33876 511
rect 33810 461 33876 477
rect 33032 431 33098 447
rect 33032 397 33048 431
rect 33082 397 33098 431
rect 33032 381 33098 397
rect 32254 351 32320 367
rect 32254 317 32270 351
rect 32304 317 32320 351
rect 32254 301 32320 317
rect 34606 287 34636 588
rect 35384 367 35414 588
rect 36162 447 36192 588
rect 36940 527 36970 588
rect 36922 511 36988 527
rect 36922 477 36938 511
rect 36972 477 36988 511
rect 36922 461 36988 477
rect 36144 431 36210 447
rect 36144 397 36160 431
rect 36194 397 36210 431
rect 36144 381 36210 397
rect 35366 351 35432 367
rect 35366 317 35382 351
rect 35416 317 35432 351
rect 35366 301 35432 317
rect 37718 287 37748 588
rect 38496 367 38526 588
rect 39274 447 39304 588
rect 40052 527 40082 588
rect 40034 511 40100 527
rect 40034 477 40050 511
rect 40084 477 40100 511
rect 40034 461 40100 477
rect 39256 431 39322 447
rect 39256 397 39272 431
rect 39306 397 39322 431
rect 39256 381 39322 397
rect 38478 351 38544 367
rect 38478 317 38494 351
rect 38528 317 38544 351
rect 38478 301 38544 317
rect 40830 287 40860 588
rect 41608 367 41638 588
rect 42386 447 42416 588
rect 43164 527 43194 588
rect 43146 511 43212 527
rect 43146 477 43162 511
rect 43196 477 43212 511
rect 43146 461 43212 477
rect 42368 431 42434 447
rect 42368 397 42384 431
rect 42418 397 42434 431
rect 42368 381 42434 397
rect 41590 351 41656 367
rect 41590 317 41606 351
rect 41640 317 41656 351
rect 41590 301 41656 317
rect 43942 287 43972 588
rect 44720 367 44750 588
rect 45498 447 45528 588
rect 46276 527 46306 588
rect 46258 511 46324 527
rect 46258 477 46274 511
rect 46308 477 46324 511
rect 46258 461 46324 477
rect 45480 431 45546 447
rect 45480 397 45496 431
rect 45530 397 45546 431
rect 45480 381 45546 397
rect 44702 351 44768 367
rect 44702 317 44718 351
rect 44752 317 44768 351
rect 44702 301 44768 317
rect 47054 287 47084 588
rect 47832 367 47862 588
rect 48610 447 48640 588
rect 49388 527 49418 588
rect 49370 511 49436 527
rect 49370 477 49386 511
rect 49420 477 49436 511
rect 49370 461 49436 477
rect 48592 431 48658 447
rect 48592 397 48608 431
rect 48642 397 48658 431
rect 48592 381 48658 397
rect 47814 351 47880 367
rect 47814 317 47830 351
rect 47864 317 47880 351
rect 47814 301 47880 317
rect 356 271 422 287
rect 356 237 372 271
rect 406 237 422 271
rect 356 221 422 237
rect 3468 271 3534 287
rect 3468 237 3484 271
rect 3518 237 3534 271
rect 3468 221 3534 237
rect 6580 271 6646 287
rect 6580 237 6596 271
rect 6630 237 6646 271
rect 6580 221 6646 237
rect 9692 271 9758 287
rect 9692 237 9708 271
rect 9742 237 9758 271
rect 9692 221 9758 237
rect 12804 271 12870 287
rect 12804 237 12820 271
rect 12854 237 12870 271
rect 12804 221 12870 237
rect 15916 271 15982 287
rect 15916 237 15932 271
rect 15966 237 15982 271
rect 15916 221 15982 237
rect 19028 271 19094 287
rect 19028 237 19044 271
rect 19078 237 19094 271
rect 19028 221 19094 237
rect 22140 271 22206 287
rect 22140 237 22156 271
rect 22190 237 22206 271
rect 22140 221 22206 237
rect 25252 271 25318 287
rect 25252 237 25268 271
rect 25302 237 25318 271
rect 25252 221 25318 237
rect 28364 271 28430 287
rect 28364 237 28380 271
rect 28414 237 28430 271
rect 28364 221 28430 237
rect 31476 271 31542 287
rect 31476 237 31492 271
rect 31526 237 31542 271
rect 31476 221 31542 237
rect 34588 271 34654 287
rect 34588 237 34604 271
rect 34638 237 34654 271
rect 34588 221 34654 237
rect 37700 271 37766 287
rect 37700 237 37716 271
rect 37750 237 37766 271
rect 37700 221 37766 237
rect 40812 271 40878 287
rect 40812 237 40828 271
rect 40862 237 40878 271
rect 40812 221 40878 237
rect 43924 271 43990 287
rect 43924 237 43940 271
rect 43974 237 43990 271
rect 43924 221 43990 237
rect 47036 271 47102 287
rect 47036 237 47052 271
rect 47086 237 47102 271
rect 47036 221 47102 237
<< polycont >>
rect 2706 477 2740 511
rect 1928 397 1962 431
rect 1150 317 1184 351
rect 5818 477 5852 511
rect 5040 397 5074 431
rect 4262 317 4296 351
rect 8930 477 8964 511
rect 8152 397 8186 431
rect 7374 317 7408 351
rect 12042 477 12076 511
rect 11264 397 11298 431
rect 10486 317 10520 351
rect 15154 477 15188 511
rect 14376 397 14410 431
rect 13598 317 13632 351
rect 18266 477 18300 511
rect 17488 397 17522 431
rect 16710 317 16744 351
rect 21378 477 21412 511
rect 20600 397 20634 431
rect 19822 317 19856 351
rect 24490 477 24524 511
rect 23712 397 23746 431
rect 22934 317 22968 351
rect 27602 477 27636 511
rect 26824 397 26858 431
rect 26046 317 26080 351
rect 30714 477 30748 511
rect 29936 397 29970 431
rect 29158 317 29192 351
rect 33826 477 33860 511
rect 33048 397 33082 431
rect 32270 317 32304 351
rect 36938 477 36972 511
rect 36160 397 36194 431
rect 35382 317 35416 351
rect 40050 477 40084 511
rect 39272 397 39306 431
rect 38494 317 38528 351
rect 43162 477 43196 511
rect 42384 397 42418 431
rect 41606 317 41640 351
rect 46274 477 46308 511
rect 45496 397 45530 431
rect 44718 317 44752 351
rect 49386 477 49420 511
rect 48608 397 48642 431
rect 47830 317 47864 351
rect 372 237 406 271
rect 3484 237 3518 271
rect 6596 237 6630 271
rect 9708 237 9742 271
rect 12820 237 12854 271
rect 15932 237 15966 271
rect 19044 237 19078 271
rect 22156 237 22190 271
rect 25268 237 25302 271
rect 28380 237 28414 271
rect 31492 237 31526 271
rect 34604 237 34638 271
rect 37716 237 37750 271
rect 40828 237 40862 271
rect 43940 237 43974 271
rect 47052 237 47086 271
<< locali >>
rect 2690 511 2756 527
rect 2690 477 2706 511
rect 2740 477 2756 511
rect 2690 461 2756 477
rect 5802 511 5868 527
rect 5802 477 5818 511
rect 5852 477 5868 511
rect 5802 461 5868 477
rect 8914 511 8980 527
rect 8914 477 8930 511
rect 8964 477 8980 511
rect 8914 461 8980 477
rect 12026 511 12092 527
rect 12026 477 12042 511
rect 12076 477 12092 511
rect 12026 461 12092 477
rect 15138 511 15204 527
rect 15138 477 15154 511
rect 15188 477 15204 511
rect 15138 461 15204 477
rect 18250 511 18316 527
rect 18250 477 18266 511
rect 18300 477 18316 511
rect 18250 461 18316 477
rect 21362 511 21428 527
rect 21362 477 21378 511
rect 21412 477 21428 511
rect 21362 461 21428 477
rect 24474 511 24540 527
rect 24474 477 24490 511
rect 24524 477 24540 511
rect 24474 461 24540 477
rect 27586 511 27652 527
rect 27586 477 27602 511
rect 27636 477 27652 511
rect 27586 461 27652 477
rect 30698 511 30764 527
rect 30698 477 30714 511
rect 30748 477 30764 511
rect 30698 461 30764 477
rect 33810 511 33876 527
rect 33810 477 33826 511
rect 33860 477 33876 511
rect 33810 461 33876 477
rect 36922 511 36988 527
rect 36922 477 36938 511
rect 36972 477 36988 511
rect 36922 461 36988 477
rect 40034 511 40100 527
rect 40034 477 40050 511
rect 40084 477 40100 511
rect 40034 461 40100 477
rect 43146 511 43212 527
rect 43146 477 43162 511
rect 43196 477 43212 511
rect 43146 461 43212 477
rect 46258 511 46324 527
rect 46258 477 46274 511
rect 46308 477 46324 511
rect 46258 461 46324 477
rect 49370 511 49436 527
rect 49370 477 49386 511
rect 49420 477 49436 511
rect 49370 461 49436 477
rect 1912 431 1978 447
rect 1912 397 1928 431
rect 1962 397 1978 431
rect 1912 381 1978 397
rect 5024 431 5090 447
rect 5024 397 5040 431
rect 5074 397 5090 431
rect 5024 381 5090 397
rect 8136 431 8202 447
rect 8136 397 8152 431
rect 8186 397 8202 431
rect 8136 381 8202 397
rect 11248 431 11314 447
rect 11248 397 11264 431
rect 11298 397 11314 431
rect 11248 381 11314 397
rect 14360 431 14426 447
rect 14360 397 14376 431
rect 14410 397 14426 431
rect 14360 381 14426 397
rect 17472 431 17538 447
rect 17472 397 17488 431
rect 17522 397 17538 431
rect 17472 381 17538 397
rect 20584 431 20650 447
rect 20584 397 20600 431
rect 20634 397 20650 431
rect 20584 381 20650 397
rect 23696 431 23762 447
rect 23696 397 23712 431
rect 23746 397 23762 431
rect 23696 381 23762 397
rect 26808 431 26874 447
rect 26808 397 26824 431
rect 26858 397 26874 431
rect 26808 381 26874 397
rect 29920 431 29986 447
rect 29920 397 29936 431
rect 29970 397 29986 431
rect 29920 381 29986 397
rect 33032 431 33098 447
rect 33032 397 33048 431
rect 33082 397 33098 431
rect 33032 381 33098 397
rect 36144 431 36210 447
rect 36144 397 36160 431
rect 36194 397 36210 431
rect 36144 381 36210 397
rect 39256 431 39322 447
rect 39256 397 39272 431
rect 39306 397 39322 431
rect 39256 381 39322 397
rect 42368 431 42434 447
rect 42368 397 42384 431
rect 42418 397 42434 431
rect 42368 381 42434 397
rect 45480 431 45546 447
rect 45480 397 45496 431
rect 45530 397 45546 431
rect 45480 381 45546 397
rect 48592 431 48658 447
rect 48592 397 48608 431
rect 48642 397 48658 431
rect 48592 381 48658 397
rect 1134 351 1200 367
rect 1134 317 1150 351
rect 1184 317 1200 351
rect 1134 301 1200 317
rect 4246 351 4312 367
rect 4246 317 4262 351
rect 4296 317 4312 351
rect 4246 301 4312 317
rect 7358 351 7424 367
rect 7358 317 7374 351
rect 7408 317 7424 351
rect 7358 301 7424 317
rect 10470 351 10536 367
rect 10470 317 10486 351
rect 10520 317 10536 351
rect 10470 301 10536 317
rect 13582 351 13648 367
rect 13582 317 13598 351
rect 13632 317 13648 351
rect 13582 301 13648 317
rect 16694 351 16760 367
rect 16694 317 16710 351
rect 16744 317 16760 351
rect 16694 301 16760 317
rect 19806 351 19872 367
rect 19806 317 19822 351
rect 19856 317 19872 351
rect 19806 301 19872 317
rect 22918 351 22984 367
rect 22918 317 22934 351
rect 22968 317 22984 351
rect 22918 301 22984 317
rect 26030 351 26096 367
rect 26030 317 26046 351
rect 26080 317 26096 351
rect 26030 301 26096 317
rect 29142 351 29208 367
rect 29142 317 29158 351
rect 29192 317 29208 351
rect 29142 301 29208 317
rect 32254 351 32320 367
rect 32254 317 32270 351
rect 32304 317 32320 351
rect 32254 301 32320 317
rect 35366 351 35432 367
rect 35366 317 35382 351
rect 35416 317 35432 351
rect 35366 301 35432 317
rect 38478 351 38544 367
rect 38478 317 38494 351
rect 38528 317 38544 351
rect 38478 301 38544 317
rect 41590 351 41656 367
rect 41590 317 41606 351
rect 41640 317 41656 351
rect 41590 301 41656 317
rect 44702 351 44768 367
rect 44702 317 44718 351
rect 44752 317 44768 351
rect 44702 301 44768 317
rect 47814 351 47880 367
rect 47814 317 47830 351
rect 47864 317 47880 351
rect 47814 301 47880 317
rect 356 271 422 287
rect 356 237 372 271
rect 406 237 422 271
rect 356 221 422 237
rect 3468 271 3534 287
rect 3468 237 3484 271
rect 3518 237 3534 271
rect 3468 221 3534 237
rect 6580 271 6646 287
rect 6580 237 6596 271
rect 6630 237 6646 271
rect 6580 221 6646 237
rect 9692 271 9758 287
rect 9692 237 9708 271
rect 9742 237 9758 271
rect 9692 221 9758 237
rect 12804 271 12870 287
rect 12804 237 12820 271
rect 12854 237 12870 271
rect 12804 221 12870 237
rect 15916 271 15982 287
rect 15916 237 15932 271
rect 15966 237 15982 271
rect 15916 221 15982 237
rect 19028 271 19094 287
rect 19028 237 19044 271
rect 19078 237 19094 271
rect 19028 221 19094 237
rect 22140 271 22206 287
rect 22140 237 22156 271
rect 22190 237 22206 271
rect 22140 221 22206 237
rect 25252 271 25318 287
rect 25252 237 25268 271
rect 25302 237 25318 271
rect 25252 221 25318 237
rect 28364 271 28430 287
rect 28364 237 28380 271
rect 28414 237 28430 271
rect 28364 221 28430 237
rect 31476 271 31542 287
rect 31476 237 31492 271
rect 31526 237 31542 271
rect 31476 221 31542 237
rect 34588 271 34654 287
rect 34588 237 34604 271
rect 34638 237 34654 271
rect 34588 221 34654 237
rect 37700 271 37766 287
rect 37700 237 37716 271
rect 37750 237 37766 271
rect 37700 221 37766 237
rect 40812 271 40878 287
rect 40812 237 40828 271
rect 40862 237 40878 271
rect 40812 221 40878 237
rect 43924 271 43990 287
rect 43924 237 43940 271
rect 43974 237 43990 271
rect 43924 221 43990 237
rect 47036 271 47102 287
rect 47036 237 47052 271
rect 47086 237 47102 271
rect 47036 221 47102 237
<< viali >>
rect 2706 477 2740 511
rect 5818 477 5852 511
rect 8930 477 8964 511
rect 12042 477 12076 511
rect 15154 477 15188 511
rect 18266 477 18300 511
rect 21378 477 21412 511
rect 24490 477 24524 511
rect 27602 477 27636 511
rect 30714 477 30748 511
rect 33826 477 33860 511
rect 36938 477 36972 511
rect 40050 477 40084 511
rect 43162 477 43196 511
rect 46274 477 46308 511
rect 49386 477 49420 511
rect 1928 397 1962 431
rect 5040 397 5074 431
rect 8152 397 8186 431
rect 11264 397 11298 431
rect 14376 397 14410 431
rect 17488 397 17522 431
rect 20600 397 20634 431
rect 23712 397 23746 431
rect 26824 397 26858 431
rect 29936 397 29970 431
rect 33048 397 33082 431
rect 36160 397 36194 431
rect 39272 397 39306 431
rect 42384 397 42418 431
rect 45496 397 45530 431
rect 48608 397 48642 431
rect 1150 317 1184 351
rect 4262 317 4296 351
rect 7374 317 7408 351
rect 10486 317 10520 351
rect 13598 317 13632 351
rect 16710 317 16744 351
rect 19822 317 19856 351
rect 22934 317 22968 351
rect 26046 317 26080 351
rect 29158 317 29192 351
rect 32270 317 32304 351
rect 35382 317 35416 351
rect 38494 317 38528 351
rect 41606 317 41640 351
rect 44718 317 44752 351
rect 47830 317 47864 351
rect 372 237 406 271
rect 3484 237 3518 271
rect 6596 237 6630 271
rect 9708 237 9742 271
rect 12820 237 12854 271
rect 15932 237 15966 271
rect 19044 237 19078 271
rect 22156 237 22190 271
rect 25268 237 25302 271
rect 28380 237 28414 271
rect 31492 237 31526 271
rect 34604 237 34638 271
rect 37716 237 37750 271
rect 40828 237 40862 271
rect 43940 237 43974 271
rect 47052 237 47086 271
<< metal1 >>
rect 2694 511 2752 517
rect 2694 508 2706 511
rect 0 480 2706 508
rect 2694 477 2706 480
rect 2740 508 2752 511
rect 5806 511 5864 517
rect 5806 508 5818 511
rect 2740 480 5818 508
rect 2740 477 2752 480
rect 2694 471 2752 477
rect 5806 477 5818 480
rect 5852 508 5864 511
rect 8918 511 8976 517
rect 8918 508 8930 511
rect 5852 480 8930 508
rect 5852 477 5864 480
rect 5806 471 5864 477
rect 8918 477 8930 480
rect 8964 508 8976 511
rect 12030 511 12088 517
rect 12030 508 12042 511
rect 8964 480 12042 508
rect 8964 477 8976 480
rect 8918 471 8976 477
rect 12030 477 12042 480
rect 12076 508 12088 511
rect 15142 511 15200 517
rect 15142 508 15154 511
rect 12076 480 15154 508
rect 12076 477 12088 480
rect 12030 471 12088 477
rect 15142 477 15154 480
rect 15188 508 15200 511
rect 18254 511 18312 517
rect 18254 508 18266 511
rect 15188 480 18266 508
rect 15188 477 15200 480
rect 15142 471 15200 477
rect 18254 477 18266 480
rect 18300 508 18312 511
rect 21366 511 21424 517
rect 21366 508 21378 511
rect 18300 480 21378 508
rect 18300 477 18312 480
rect 18254 471 18312 477
rect 21366 477 21378 480
rect 21412 508 21424 511
rect 24478 511 24536 517
rect 24478 508 24490 511
rect 21412 480 24490 508
rect 21412 477 21424 480
rect 21366 471 21424 477
rect 24478 477 24490 480
rect 24524 508 24536 511
rect 27590 511 27648 517
rect 27590 508 27602 511
rect 24524 480 27602 508
rect 24524 477 24536 480
rect 24478 471 24536 477
rect 27590 477 27602 480
rect 27636 508 27648 511
rect 30702 511 30760 517
rect 30702 508 30714 511
rect 27636 480 30714 508
rect 27636 477 27648 480
rect 27590 471 27648 477
rect 30702 477 30714 480
rect 30748 508 30760 511
rect 33814 511 33872 517
rect 33814 508 33826 511
rect 30748 480 33826 508
rect 30748 477 30760 480
rect 30702 471 30760 477
rect 33814 477 33826 480
rect 33860 508 33872 511
rect 36926 511 36984 517
rect 36926 508 36938 511
rect 33860 480 36938 508
rect 33860 477 33872 480
rect 33814 471 33872 477
rect 36926 477 36938 480
rect 36972 508 36984 511
rect 40038 511 40096 517
rect 40038 508 40050 511
rect 36972 480 40050 508
rect 36972 477 36984 480
rect 36926 471 36984 477
rect 40038 477 40050 480
rect 40084 508 40096 511
rect 43150 511 43208 517
rect 43150 508 43162 511
rect 40084 480 43162 508
rect 40084 477 40096 480
rect 40038 471 40096 477
rect 43150 477 43162 480
rect 43196 508 43208 511
rect 46262 511 46320 517
rect 46262 508 46274 511
rect 43196 480 46274 508
rect 43196 477 43208 480
rect 43150 471 43208 477
rect 46262 477 46274 480
rect 46308 508 46320 511
rect 49374 511 49432 517
rect 49374 508 49386 511
rect 46308 480 49386 508
rect 46308 477 46320 480
rect 46262 471 46320 477
rect 49374 477 49386 480
rect 49420 508 49432 511
rect 49420 480 49792 508
rect 49420 477 49432 480
rect 49374 471 49432 477
rect 1916 431 1974 437
rect 1916 428 1928 431
rect 0 400 1928 428
rect 1916 397 1928 400
rect 1962 428 1974 431
rect 5028 431 5086 437
rect 5028 428 5040 431
rect 1962 400 5040 428
rect 1962 397 1974 400
rect 1916 391 1974 397
rect 5028 397 5040 400
rect 5074 428 5086 431
rect 8140 431 8198 437
rect 8140 428 8152 431
rect 5074 400 8152 428
rect 5074 397 5086 400
rect 5028 391 5086 397
rect 8140 397 8152 400
rect 8186 428 8198 431
rect 11252 431 11310 437
rect 11252 428 11264 431
rect 8186 400 11264 428
rect 8186 397 8198 400
rect 8140 391 8198 397
rect 11252 397 11264 400
rect 11298 428 11310 431
rect 14364 431 14422 437
rect 14364 428 14376 431
rect 11298 400 14376 428
rect 11298 397 11310 400
rect 11252 391 11310 397
rect 14364 397 14376 400
rect 14410 428 14422 431
rect 17476 431 17534 437
rect 17476 428 17488 431
rect 14410 400 17488 428
rect 14410 397 14422 400
rect 14364 391 14422 397
rect 17476 397 17488 400
rect 17522 428 17534 431
rect 20588 431 20646 437
rect 20588 428 20600 431
rect 17522 400 20600 428
rect 17522 397 17534 400
rect 17476 391 17534 397
rect 20588 397 20600 400
rect 20634 428 20646 431
rect 23700 431 23758 437
rect 23700 428 23712 431
rect 20634 400 23712 428
rect 20634 397 20646 400
rect 20588 391 20646 397
rect 23700 397 23712 400
rect 23746 428 23758 431
rect 26812 431 26870 437
rect 26812 428 26824 431
rect 23746 400 26824 428
rect 23746 397 23758 400
rect 23700 391 23758 397
rect 26812 397 26824 400
rect 26858 428 26870 431
rect 29924 431 29982 437
rect 29924 428 29936 431
rect 26858 400 29936 428
rect 26858 397 26870 400
rect 26812 391 26870 397
rect 29924 397 29936 400
rect 29970 428 29982 431
rect 33036 431 33094 437
rect 33036 428 33048 431
rect 29970 400 33048 428
rect 29970 397 29982 400
rect 29924 391 29982 397
rect 33036 397 33048 400
rect 33082 428 33094 431
rect 36148 431 36206 437
rect 36148 428 36160 431
rect 33082 400 36160 428
rect 33082 397 33094 400
rect 33036 391 33094 397
rect 36148 397 36160 400
rect 36194 428 36206 431
rect 39260 431 39318 437
rect 39260 428 39272 431
rect 36194 400 39272 428
rect 36194 397 36206 400
rect 36148 391 36206 397
rect 39260 397 39272 400
rect 39306 428 39318 431
rect 42372 431 42430 437
rect 42372 428 42384 431
rect 39306 400 42384 428
rect 39306 397 39318 400
rect 39260 391 39318 397
rect 42372 397 42384 400
rect 42418 428 42430 431
rect 45484 431 45542 437
rect 45484 428 45496 431
rect 42418 400 45496 428
rect 42418 397 42430 400
rect 42372 391 42430 397
rect 45484 397 45496 400
rect 45530 428 45542 431
rect 48596 431 48654 437
rect 48596 428 48608 431
rect 45530 400 48608 428
rect 45530 397 45542 400
rect 45484 391 45542 397
rect 48596 397 48608 400
rect 48642 428 48654 431
rect 48642 400 49792 428
rect 48642 397 48654 400
rect 48596 391 48654 397
rect 1138 351 1196 357
rect 1138 348 1150 351
rect 0 320 1150 348
rect 1138 317 1150 320
rect 1184 348 1196 351
rect 4250 351 4308 357
rect 4250 348 4262 351
rect 1184 320 4262 348
rect 1184 317 1196 320
rect 1138 311 1196 317
rect 4250 317 4262 320
rect 4296 348 4308 351
rect 7362 351 7420 357
rect 7362 348 7374 351
rect 4296 320 7374 348
rect 4296 317 4308 320
rect 4250 311 4308 317
rect 7362 317 7374 320
rect 7408 348 7420 351
rect 10474 351 10532 357
rect 10474 348 10486 351
rect 7408 320 10486 348
rect 7408 317 7420 320
rect 7362 311 7420 317
rect 10474 317 10486 320
rect 10520 348 10532 351
rect 13586 351 13644 357
rect 13586 348 13598 351
rect 10520 320 13598 348
rect 10520 317 10532 320
rect 10474 311 10532 317
rect 13586 317 13598 320
rect 13632 348 13644 351
rect 16698 351 16756 357
rect 16698 348 16710 351
rect 13632 320 16710 348
rect 13632 317 13644 320
rect 13586 311 13644 317
rect 16698 317 16710 320
rect 16744 348 16756 351
rect 19810 351 19868 357
rect 19810 348 19822 351
rect 16744 320 19822 348
rect 16744 317 16756 320
rect 16698 311 16756 317
rect 19810 317 19822 320
rect 19856 348 19868 351
rect 22922 351 22980 357
rect 22922 348 22934 351
rect 19856 320 22934 348
rect 19856 317 19868 320
rect 19810 311 19868 317
rect 22922 317 22934 320
rect 22968 348 22980 351
rect 26034 351 26092 357
rect 26034 348 26046 351
rect 22968 320 26046 348
rect 22968 317 22980 320
rect 22922 311 22980 317
rect 26034 317 26046 320
rect 26080 348 26092 351
rect 29146 351 29204 357
rect 29146 348 29158 351
rect 26080 320 29158 348
rect 26080 317 26092 320
rect 26034 311 26092 317
rect 29146 317 29158 320
rect 29192 348 29204 351
rect 32258 351 32316 357
rect 32258 348 32270 351
rect 29192 320 32270 348
rect 29192 317 29204 320
rect 29146 311 29204 317
rect 32258 317 32270 320
rect 32304 348 32316 351
rect 35370 351 35428 357
rect 35370 348 35382 351
rect 32304 320 35382 348
rect 32304 317 32316 320
rect 32258 311 32316 317
rect 35370 317 35382 320
rect 35416 348 35428 351
rect 38482 351 38540 357
rect 38482 348 38494 351
rect 35416 320 38494 348
rect 35416 317 35428 320
rect 35370 311 35428 317
rect 38482 317 38494 320
rect 38528 348 38540 351
rect 41594 351 41652 357
rect 41594 348 41606 351
rect 38528 320 41606 348
rect 38528 317 38540 320
rect 38482 311 38540 317
rect 41594 317 41606 320
rect 41640 348 41652 351
rect 44706 351 44764 357
rect 44706 348 44718 351
rect 41640 320 44718 348
rect 41640 317 41652 320
rect 41594 311 41652 317
rect 44706 317 44718 320
rect 44752 348 44764 351
rect 47818 351 47876 357
rect 47818 348 47830 351
rect 44752 320 47830 348
rect 44752 317 44764 320
rect 44706 311 44764 317
rect 47818 317 47830 320
rect 47864 348 47876 351
rect 47864 320 49792 348
rect 47864 317 47876 320
rect 47818 311 47876 317
rect 360 271 418 277
rect 360 268 372 271
rect 0 240 372 268
rect 360 237 372 240
rect 406 268 418 271
rect 3472 271 3530 277
rect 3472 268 3484 271
rect 406 240 3484 268
rect 406 237 418 240
rect 360 231 418 237
rect 3472 237 3484 240
rect 3518 268 3530 271
rect 6584 271 6642 277
rect 6584 268 6596 271
rect 3518 240 6596 268
rect 3518 237 3530 240
rect 3472 231 3530 237
rect 6584 237 6596 240
rect 6630 268 6642 271
rect 9696 271 9754 277
rect 9696 268 9708 271
rect 6630 240 9708 268
rect 6630 237 6642 240
rect 6584 231 6642 237
rect 9696 237 9708 240
rect 9742 268 9754 271
rect 12808 271 12866 277
rect 12808 268 12820 271
rect 9742 240 12820 268
rect 9742 237 9754 240
rect 9696 231 9754 237
rect 12808 237 12820 240
rect 12854 268 12866 271
rect 15920 271 15978 277
rect 15920 268 15932 271
rect 12854 240 15932 268
rect 12854 237 12866 240
rect 12808 231 12866 237
rect 15920 237 15932 240
rect 15966 268 15978 271
rect 19032 271 19090 277
rect 19032 268 19044 271
rect 15966 240 19044 268
rect 15966 237 15978 240
rect 15920 231 15978 237
rect 19032 237 19044 240
rect 19078 268 19090 271
rect 22144 271 22202 277
rect 22144 268 22156 271
rect 19078 240 22156 268
rect 19078 237 19090 240
rect 19032 231 19090 237
rect 22144 237 22156 240
rect 22190 268 22202 271
rect 25256 271 25314 277
rect 25256 268 25268 271
rect 22190 240 25268 268
rect 22190 237 22202 240
rect 22144 231 22202 237
rect 25256 237 25268 240
rect 25302 268 25314 271
rect 28368 271 28426 277
rect 28368 268 28380 271
rect 25302 240 28380 268
rect 25302 237 25314 240
rect 25256 231 25314 237
rect 28368 237 28380 240
rect 28414 268 28426 271
rect 31480 271 31538 277
rect 31480 268 31492 271
rect 28414 240 31492 268
rect 28414 237 28426 240
rect 28368 231 28426 237
rect 31480 237 31492 240
rect 31526 268 31538 271
rect 34592 271 34650 277
rect 34592 268 34604 271
rect 31526 240 34604 268
rect 31526 237 31538 240
rect 31480 231 31538 237
rect 34592 237 34604 240
rect 34638 268 34650 271
rect 37704 271 37762 277
rect 37704 268 37716 271
rect 34638 240 37716 268
rect 34638 237 34650 240
rect 34592 231 34650 237
rect 37704 237 37716 240
rect 37750 268 37762 271
rect 40816 271 40874 277
rect 40816 268 40828 271
rect 37750 240 40828 268
rect 37750 237 37762 240
rect 37704 231 37762 237
rect 40816 237 40828 240
rect 40862 268 40874 271
rect 43928 271 43986 277
rect 43928 268 43940 271
rect 40862 240 43940 268
rect 40862 237 40874 240
rect 40816 231 40874 237
rect 43928 237 43940 240
rect 43974 268 43986 271
rect 47040 271 47098 277
rect 47040 268 47052 271
rect 43974 240 47052 268
rect 43974 237 43986 240
rect 43928 231 43986 237
rect 47040 237 47052 240
rect 47086 268 47098 271
rect 47086 240 49792 268
rect 47086 237 47098 240
rect 47040 231 47098 237
rect 66 134 72 186
rect 124 174 130 186
rect 844 174 850 186
rect 124 146 850 174
rect 124 134 130 146
rect 844 134 850 146
rect 902 174 908 186
rect 1622 174 1628 186
rect 902 146 1628 174
rect 902 134 908 146
rect 1622 134 1628 146
rect 1680 174 1686 186
rect 2400 174 2406 186
rect 1680 146 2406 174
rect 1680 134 1686 146
rect 2400 134 2406 146
rect 2458 134 2464 186
rect 3178 134 3184 186
rect 3236 174 3242 186
rect 3956 174 3962 186
rect 3236 146 3962 174
rect 3236 134 3242 146
rect 3956 134 3962 146
rect 4014 174 4020 186
rect 4734 174 4740 186
rect 4014 146 4740 174
rect 4014 134 4020 146
rect 4734 134 4740 146
rect 4792 174 4798 186
rect 5512 174 5518 186
rect 4792 146 5518 174
rect 4792 134 4798 146
rect 5512 134 5518 146
rect 5570 134 5576 186
rect 6290 134 6296 186
rect 6348 174 6354 186
rect 7068 174 7074 186
rect 6348 146 7074 174
rect 6348 134 6354 146
rect 7068 134 7074 146
rect 7126 174 7132 186
rect 7846 174 7852 186
rect 7126 146 7852 174
rect 7126 134 7132 146
rect 7846 134 7852 146
rect 7904 174 7910 186
rect 8624 174 8630 186
rect 7904 146 8630 174
rect 7904 134 7910 146
rect 8624 134 8630 146
rect 8682 134 8688 186
rect 9402 134 9408 186
rect 9460 174 9466 186
rect 10180 174 10186 186
rect 9460 146 10186 174
rect 9460 134 9466 146
rect 10180 134 10186 146
rect 10238 174 10244 186
rect 10958 174 10964 186
rect 10238 146 10964 174
rect 10238 134 10244 146
rect 10958 134 10964 146
rect 11016 174 11022 186
rect 11736 174 11742 186
rect 11016 146 11742 174
rect 11016 134 11022 146
rect 11736 134 11742 146
rect 11794 134 11800 186
rect 12514 134 12520 186
rect 12572 174 12578 186
rect 13292 174 13298 186
rect 12572 146 13298 174
rect 12572 134 12578 146
rect 13292 134 13298 146
rect 13350 174 13356 186
rect 14070 174 14076 186
rect 13350 146 14076 174
rect 13350 134 13356 146
rect 14070 134 14076 146
rect 14128 174 14134 186
rect 14848 174 14854 186
rect 14128 146 14854 174
rect 14128 134 14134 146
rect 14848 134 14854 146
rect 14906 134 14912 186
rect 15626 134 15632 186
rect 15684 174 15690 186
rect 16404 174 16410 186
rect 15684 146 16410 174
rect 15684 134 15690 146
rect 16404 134 16410 146
rect 16462 174 16468 186
rect 17182 174 17188 186
rect 16462 146 17188 174
rect 16462 134 16468 146
rect 17182 134 17188 146
rect 17240 174 17246 186
rect 17960 174 17966 186
rect 17240 146 17966 174
rect 17240 134 17246 146
rect 17960 134 17966 146
rect 18018 134 18024 186
rect 18738 134 18744 186
rect 18796 174 18802 186
rect 19516 174 19522 186
rect 18796 146 19522 174
rect 18796 134 18802 146
rect 19516 134 19522 146
rect 19574 174 19580 186
rect 20294 174 20300 186
rect 19574 146 20300 174
rect 19574 134 19580 146
rect 20294 134 20300 146
rect 20352 174 20358 186
rect 21072 174 21078 186
rect 20352 146 21078 174
rect 20352 134 20358 146
rect 21072 134 21078 146
rect 21130 134 21136 186
rect 21850 134 21856 186
rect 21908 174 21914 186
rect 22628 174 22634 186
rect 21908 146 22634 174
rect 21908 134 21914 146
rect 22628 134 22634 146
rect 22686 174 22692 186
rect 23406 174 23412 186
rect 22686 146 23412 174
rect 22686 134 22692 146
rect 23406 134 23412 146
rect 23464 174 23470 186
rect 24184 174 24190 186
rect 23464 146 24190 174
rect 23464 134 23470 146
rect 24184 134 24190 146
rect 24242 134 24248 186
rect 24962 134 24968 186
rect 25020 174 25026 186
rect 25740 174 25746 186
rect 25020 146 25746 174
rect 25020 134 25026 146
rect 25740 134 25746 146
rect 25798 174 25804 186
rect 26518 174 26524 186
rect 25798 146 26524 174
rect 25798 134 25804 146
rect 26518 134 26524 146
rect 26576 174 26582 186
rect 27296 174 27302 186
rect 26576 146 27302 174
rect 26576 134 26582 146
rect 27296 134 27302 146
rect 27354 134 27360 186
rect 28074 134 28080 186
rect 28132 174 28138 186
rect 28852 174 28858 186
rect 28132 146 28858 174
rect 28132 134 28138 146
rect 28852 134 28858 146
rect 28910 174 28916 186
rect 29630 174 29636 186
rect 28910 146 29636 174
rect 28910 134 28916 146
rect 29630 134 29636 146
rect 29688 174 29694 186
rect 30408 174 30414 186
rect 29688 146 30414 174
rect 29688 134 29694 146
rect 30408 134 30414 146
rect 30466 134 30472 186
rect 31186 134 31192 186
rect 31244 174 31250 186
rect 31964 174 31970 186
rect 31244 146 31970 174
rect 31244 134 31250 146
rect 31964 134 31970 146
rect 32022 174 32028 186
rect 32742 174 32748 186
rect 32022 146 32748 174
rect 32022 134 32028 146
rect 32742 134 32748 146
rect 32800 174 32806 186
rect 33520 174 33526 186
rect 32800 146 33526 174
rect 32800 134 32806 146
rect 33520 134 33526 146
rect 33578 134 33584 186
rect 34298 134 34304 186
rect 34356 174 34362 186
rect 35076 174 35082 186
rect 34356 146 35082 174
rect 34356 134 34362 146
rect 35076 134 35082 146
rect 35134 174 35140 186
rect 35854 174 35860 186
rect 35134 146 35860 174
rect 35134 134 35140 146
rect 35854 134 35860 146
rect 35912 174 35918 186
rect 36632 174 36638 186
rect 35912 146 36638 174
rect 35912 134 35918 146
rect 36632 134 36638 146
rect 36690 134 36696 186
rect 37410 134 37416 186
rect 37468 174 37474 186
rect 38188 174 38194 186
rect 37468 146 38194 174
rect 37468 134 37474 146
rect 38188 134 38194 146
rect 38246 174 38252 186
rect 38966 174 38972 186
rect 38246 146 38972 174
rect 38246 134 38252 146
rect 38966 134 38972 146
rect 39024 174 39030 186
rect 39744 174 39750 186
rect 39024 146 39750 174
rect 39024 134 39030 146
rect 39744 134 39750 146
rect 39802 134 39808 186
rect 40522 134 40528 186
rect 40580 174 40586 186
rect 41300 174 41306 186
rect 40580 146 41306 174
rect 40580 134 40586 146
rect 41300 134 41306 146
rect 41358 174 41364 186
rect 42078 174 42084 186
rect 41358 146 42084 174
rect 41358 134 41364 146
rect 42078 134 42084 146
rect 42136 174 42142 186
rect 42856 174 42862 186
rect 42136 146 42862 174
rect 42136 134 42142 146
rect 42856 134 42862 146
rect 42914 134 42920 186
rect 43634 134 43640 186
rect 43692 174 43698 186
rect 44412 174 44418 186
rect 43692 146 44418 174
rect 43692 134 43698 146
rect 44412 134 44418 146
rect 44470 174 44476 186
rect 45190 174 45196 186
rect 44470 146 45196 174
rect 44470 134 44476 146
rect 45190 134 45196 146
rect 45248 174 45254 186
rect 45968 174 45974 186
rect 45248 146 45974 174
rect 45248 134 45254 146
rect 45968 134 45974 146
rect 46026 134 46032 186
rect 46746 134 46752 186
rect 46804 174 46810 186
rect 47524 174 47530 186
rect 46804 146 47530 174
rect 46804 134 46810 146
rect 47524 134 47530 146
rect 47582 174 47588 186
rect 48302 174 48308 186
rect 47582 146 48308 174
rect 47582 134 47588 146
rect 48302 134 48308 146
rect 48360 174 48366 186
rect 49080 174 49086 186
rect 48360 146 49086 174
rect 48360 134 48366 146
rect 49080 134 49086 146
rect 49138 134 49144 186
rect 676 54 682 106
rect 734 94 740 106
rect 1454 94 1460 106
rect 734 66 1460 94
rect 734 54 740 66
rect 1454 54 1460 66
rect 1512 94 1518 106
rect 2232 94 2238 106
rect 1512 66 2238 94
rect 1512 54 1518 66
rect 2232 54 2238 66
rect 2290 94 2296 106
rect 3010 94 3016 106
rect 2290 66 3016 94
rect 2290 54 2296 66
rect 3010 54 3016 66
rect 3068 54 3074 106
rect 3788 54 3794 106
rect 3846 94 3852 106
rect 4566 94 4572 106
rect 3846 66 4572 94
rect 3846 54 3852 66
rect 4566 54 4572 66
rect 4624 94 4630 106
rect 5344 94 5350 106
rect 4624 66 5350 94
rect 4624 54 4630 66
rect 5344 54 5350 66
rect 5402 94 5408 106
rect 6122 94 6128 106
rect 5402 66 6128 94
rect 5402 54 5408 66
rect 6122 54 6128 66
rect 6180 54 6186 106
rect 6900 54 6906 106
rect 6958 94 6964 106
rect 7678 94 7684 106
rect 6958 66 7684 94
rect 6958 54 6964 66
rect 7678 54 7684 66
rect 7736 94 7742 106
rect 8456 94 8462 106
rect 7736 66 8462 94
rect 7736 54 7742 66
rect 8456 54 8462 66
rect 8514 94 8520 106
rect 9234 94 9240 106
rect 8514 66 9240 94
rect 8514 54 8520 66
rect 9234 54 9240 66
rect 9292 54 9298 106
rect 10012 54 10018 106
rect 10070 94 10076 106
rect 10790 94 10796 106
rect 10070 66 10796 94
rect 10070 54 10076 66
rect 10790 54 10796 66
rect 10848 94 10854 106
rect 11568 94 11574 106
rect 10848 66 11574 94
rect 10848 54 10854 66
rect 11568 54 11574 66
rect 11626 94 11632 106
rect 12346 94 12352 106
rect 11626 66 12352 94
rect 11626 54 11632 66
rect 12346 54 12352 66
rect 12404 54 12410 106
rect 13124 54 13130 106
rect 13182 94 13188 106
rect 13902 94 13908 106
rect 13182 66 13908 94
rect 13182 54 13188 66
rect 13902 54 13908 66
rect 13960 94 13966 106
rect 14680 94 14686 106
rect 13960 66 14686 94
rect 13960 54 13966 66
rect 14680 54 14686 66
rect 14738 94 14744 106
rect 15458 94 15464 106
rect 14738 66 15464 94
rect 14738 54 14744 66
rect 15458 54 15464 66
rect 15516 54 15522 106
rect 16236 54 16242 106
rect 16294 94 16300 106
rect 17014 94 17020 106
rect 16294 66 17020 94
rect 16294 54 16300 66
rect 17014 54 17020 66
rect 17072 94 17078 106
rect 17792 94 17798 106
rect 17072 66 17798 94
rect 17072 54 17078 66
rect 17792 54 17798 66
rect 17850 94 17856 106
rect 18570 94 18576 106
rect 17850 66 18576 94
rect 17850 54 17856 66
rect 18570 54 18576 66
rect 18628 54 18634 106
rect 19348 54 19354 106
rect 19406 94 19412 106
rect 20126 94 20132 106
rect 19406 66 20132 94
rect 19406 54 19412 66
rect 20126 54 20132 66
rect 20184 94 20190 106
rect 20904 94 20910 106
rect 20184 66 20910 94
rect 20184 54 20190 66
rect 20904 54 20910 66
rect 20962 94 20968 106
rect 21682 94 21688 106
rect 20962 66 21688 94
rect 20962 54 20968 66
rect 21682 54 21688 66
rect 21740 54 21746 106
rect 22460 54 22466 106
rect 22518 94 22524 106
rect 23238 94 23244 106
rect 22518 66 23244 94
rect 22518 54 22524 66
rect 23238 54 23244 66
rect 23296 94 23302 106
rect 24016 94 24022 106
rect 23296 66 24022 94
rect 23296 54 23302 66
rect 24016 54 24022 66
rect 24074 94 24080 106
rect 24794 94 24800 106
rect 24074 66 24800 94
rect 24074 54 24080 66
rect 24794 54 24800 66
rect 24852 54 24858 106
rect 25572 54 25578 106
rect 25630 94 25636 106
rect 26350 94 26356 106
rect 25630 66 26356 94
rect 25630 54 25636 66
rect 26350 54 26356 66
rect 26408 94 26414 106
rect 27128 94 27134 106
rect 26408 66 27134 94
rect 26408 54 26414 66
rect 27128 54 27134 66
rect 27186 94 27192 106
rect 27906 94 27912 106
rect 27186 66 27912 94
rect 27186 54 27192 66
rect 27906 54 27912 66
rect 27964 54 27970 106
rect 28684 54 28690 106
rect 28742 94 28748 106
rect 29462 94 29468 106
rect 28742 66 29468 94
rect 28742 54 28748 66
rect 29462 54 29468 66
rect 29520 94 29526 106
rect 30240 94 30246 106
rect 29520 66 30246 94
rect 29520 54 29526 66
rect 30240 54 30246 66
rect 30298 94 30304 106
rect 31018 94 31024 106
rect 30298 66 31024 94
rect 30298 54 30304 66
rect 31018 54 31024 66
rect 31076 54 31082 106
rect 31796 54 31802 106
rect 31854 94 31860 106
rect 32574 94 32580 106
rect 31854 66 32580 94
rect 31854 54 31860 66
rect 32574 54 32580 66
rect 32632 94 32638 106
rect 33352 94 33358 106
rect 32632 66 33358 94
rect 32632 54 32638 66
rect 33352 54 33358 66
rect 33410 94 33416 106
rect 34130 94 34136 106
rect 33410 66 34136 94
rect 33410 54 33416 66
rect 34130 54 34136 66
rect 34188 54 34194 106
rect 34908 54 34914 106
rect 34966 94 34972 106
rect 35686 94 35692 106
rect 34966 66 35692 94
rect 34966 54 34972 66
rect 35686 54 35692 66
rect 35744 94 35750 106
rect 36464 94 36470 106
rect 35744 66 36470 94
rect 35744 54 35750 66
rect 36464 54 36470 66
rect 36522 94 36528 106
rect 37242 94 37248 106
rect 36522 66 37248 94
rect 36522 54 36528 66
rect 37242 54 37248 66
rect 37300 54 37306 106
rect 38020 54 38026 106
rect 38078 94 38084 106
rect 38798 94 38804 106
rect 38078 66 38804 94
rect 38078 54 38084 66
rect 38798 54 38804 66
rect 38856 94 38862 106
rect 39576 94 39582 106
rect 38856 66 39582 94
rect 38856 54 38862 66
rect 39576 54 39582 66
rect 39634 94 39640 106
rect 40354 94 40360 106
rect 39634 66 40360 94
rect 39634 54 39640 66
rect 40354 54 40360 66
rect 40412 54 40418 106
rect 41132 54 41138 106
rect 41190 94 41196 106
rect 41910 94 41916 106
rect 41190 66 41916 94
rect 41190 54 41196 66
rect 41910 54 41916 66
rect 41968 94 41974 106
rect 42688 94 42694 106
rect 41968 66 42694 94
rect 41968 54 41974 66
rect 42688 54 42694 66
rect 42746 94 42752 106
rect 43466 94 43472 106
rect 42746 66 43472 94
rect 42746 54 42752 66
rect 43466 54 43472 66
rect 43524 54 43530 106
rect 44244 54 44250 106
rect 44302 94 44308 106
rect 45022 94 45028 106
rect 44302 66 45028 94
rect 44302 54 44308 66
rect 45022 54 45028 66
rect 45080 94 45086 106
rect 45800 94 45806 106
rect 45080 66 45806 94
rect 45080 54 45086 66
rect 45800 54 45806 66
rect 45858 94 45864 106
rect 46578 94 46584 106
rect 45858 66 46584 94
rect 45858 54 45864 66
rect 46578 54 46584 66
rect 46636 54 46642 106
rect 47356 54 47362 106
rect 47414 94 47420 106
rect 48134 94 48140 106
rect 47414 66 48140 94
rect 47414 54 47420 66
rect 48134 54 48140 66
rect 48192 94 48198 106
rect 48912 94 48918 106
rect 48192 66 48918 94
rect 48192 54 48198 66
rect 48912 54 48918 66
rect 48970 94 48976 106
rect 49690 94 49696 106
rect 48970 66 49696 94
rect 48970 54 48976 66
rect 49690 54 49696 66
rect 49748 54 49754 106
<< via1 >>
rect 72 134 124 186
rect 850 134 902 186
rect 1628 134 1680 186
rect 2406 134 2458 186
rect 3184 134 3236 186
rect 3962 134 4014 186
rect 4740 134 4792 186
rect 5518 134 5570 186
rect 6296 134 6348 186
rect 7074 134 7126 186
rect 7852 134 7904 186
rect 8630 134 8682 186
rect 9408 134 9460 186
rect 10186 134 10238 186
rect 10964 134 11016 186
rect 11742 134 11794 186
rect 12520 134 12572 186
rect 13298 134 13350 186
rect 14076 134 14128 186
rect 14854 134 14906 186
rect 15632 134 15684 186
rect 16410 134 16462 186
rect 17188 134 17240 186
rect 17966 134 18018 186
rect 18744 134 18796 186
rect 19522 134 19574 186
rect 20300 134 20352 186
rect 21078 134 21130 186
rect 21856 134 21908 186
rect 22634 134 22686 186
rect 23412 134 23464 186
rect 24190 134 24242 186
rect 24968 134 25020 186
rect 25746 134 25798 186
rect 26524 134 26576 186
rect 27302 134 27354 186
rect 28080 134 28132 186
rect 28858 134 28910 186
rect 29636 134 29688 186
rect 30414 134 30466 186
rect 31192 134 31244 186
rect 31970 134 32022 186
rect 32748 134 32800 186
rect 33526 134 33578 186
rect 34304 134 34356 186
rect 35082 134 35134 186
rect 35860 134 35912 186
rect 36638 134 36690 186
rect 37416 134 37468 186
rect 38194 134 38246 186
rect 38972 134 39024 186
rect 39750 134 39802 186
rect 40528 134 40580 186
rect 41306 134 41358 186
rect 42084 134 42136 186
rect 42862 134 42914 186
rect 43640 134 43692 186
rect 44418 134 44470 186
rect 45196 134 45248 186
rect 45974 134 46026 186
rect 46752 134 46804 186
rect 47530 134 47582 186
rect 48308 134 48360 186
rect 49086 134 49138 186
rect 682 54 734 106
rect 1460 54 1512 106
rect 2238 54 2290 106
rect 3016 54 3068 106
rect 3794 54 3846 106
rect 4572 54 4624 106
rect 5350 54 5402 106
rect 6128 54 6180 106
rect 6906 54 6958 106
rect 7684 54 7736 106
rect 8462 54 8514 106
rect 9240 54 9292 106
rect 10018 54 10070 106
rect 10796 54 10848 106
rect 11574 54 11626 106
rect 12352 54 12404 106
rect 13130 54 13182 106
rect 13908 54 13960 106
rect 14686 54 14738 106
rect 15464 54 15516 106
rect 16242 54 16294 106
rect 17020 54 17072 106
rect 17798 54 17850 106
rect 18576 54 18628 106
rect 19354 54 19406 106
rect 20132 54 20184 106
rect 20910 54 20962 106
rect 21688 54 21740 106
rect 22466 54 22518 106
rect 23244 54 23296 106
rect 24022 54 24074 106
rect 24800 54 24852 106
rect 25578 54 25630 106
rect 26356 54 26408 106
rect 27134 54 27186 106
rect 27912 54 27964 106
rect 28690 54 28742 106
rect 29468 54 29520 106
rect 30246 54 30298 106
rect 31024 54 31076 106
rect 31802 54 31854 106
rect 32580 54 32632 106
rect 33358 54 33410 106
rect 34136 54 34188 106
rect 34914 54 34966 106
rect 35692 54 35744 106
rect 36470 54 36522 106
rect 37248 54 37300 106
rect 38026 54 38078 106
rect 38804 54 38856 106
rect 39582 54 39634 106
rect 40360 54 40412 106
rect 41138 54 41190 106
rect 41916 54 41968 106
rect 42694 54 42746 106
rect 43472 54 43524 106
rect 44250 54 44302 106
rect 45028 54 45080 106
rect 45806 54 45858 106
rect 46584 54 46636 106
rect 47362 54 47414 106
rect 48140 54 48192 106
rect 48918 54 48970 106
rect 49696 54 49748 106
<< metal2 >>
rect 84 2012 112 2068
rect 694 2012 722 2068
rect 862 2012 890 2068
rect 1472 2012 1500 2068
rect 1640 2012 1668 2068
rect 2250 2012 2278 2068
rect 2418 2012 2446 2068
rect 3028 2012 3056 2068
rect 3196 2012 3224 2068
rect 3806 2012 3834 2068
rect 3974 2012 4002 2068
rect 4584 2012 4612 2068
rect 4752 2012 4780 2068
rect 5362 2012 5390 2068
rect 5530 2012 5558 2068
rect 6140 2012 6168 2068
rect 6308 2012 6336 2068
rect 6918 2012 6946 2068
rect 7086 2012 7114 2068
rect 7696 2012 7724 2068
rect 7864 2012 7892 2068
rect 8474 2012 8502 2068
rect 8642 2012 8670 2068
rect 9252 2012 9280 2068
rect 9420 2012 9448 2068
rect 10030 2012 10058 2068
rect 10198 2012 10226 2068
rect 10808 2012 10836 2068
rect 10976 2012 11004 2068
rect 11586 2012 11614 2068
rect 11754 2012 11782 2068
rect 12364 2012 12392 2068
rect 12532 2012 12560 2068
rect 13142 2012 13170 2068
rect 13310 2012 13338 2068
rect 13920 2012 13948 2068
rect 14088 2012 14116 2068
rect 14698 2012 14726 2068
rect 14866 2012 14894 2068
rect 15476 2012 15504 2068
rect 15644 2012 15672 2068
rect 16254 2012 16282 2068
rect 16422 2012 16450 2068
rect 17032 2012 17060 2068
rect 17200 2012 17228 2068
rect 17810 2012 17838 2068
rect 17978 2012 18006 2068
rect 18588 2012 18616 2068
rect 18756 2012 18784 2068
rect 19366 2012 19394 2068
rect 19534 2012 19562 2068
rect 20144 2012 20172 2068
rect 20312 2012 20340 2068
rect 20922 2012 20950 2068
rect 21090 2012 21118 2068
rect 21700 2012 21728 2068
rect 21868 2012 21896 2068
rect 22478 2012 22506 2068
rect 22646 2012 22674 2068
rect 23256 2012 23284 2068
rect 23424 2012 23452 2068
rect 24034 2012 24062 2068
rect 24202 2012 24230 2068
rect 24812 2012 24840 2068
rect 24980 2012 25008 2068
rect 25590 2012 25618 2068
rect 25758 2012 25786 2068
rect 26368 2012 26396 2068
rect 26536 2012 26564 2068
rect 27146 2012 27174 2068
rect 27314 2012 27342 2068
rect 27924 2012 27952 2068
rect 28092 2012 28120 2068
rect 28702 2012 28730 2068
rect 28870 2012 28898 2068
rect 29480 2012 29508 2068
rect 29648 2012 29676 2068
rect 30258 2012 30286 2068
rect 30426 2012 30454 2068
rect 31036 2012 31064 2068
rect 31204 2012 31232 2068
rect 31814 2012 31842 2068
rect 31982 2012 32010 2068
rect 32592 2012 32620 2068
rect 32760 2012 32788 2068
rect 33370 2012 33398 2068
rect 33538 2012 33566 2068
rect 34148 2012 34176 2068
rect 34316 2012 34344 2068
rect 34926 2012 34954 2068
rect 35094 2012 35122 2068
rect 35704 2012 35732 2068
rect 35872 2012 35900 2068
rect 36482 2012 36510 2068
rect 36650 2012 36678 2068
rect 37260 2012 37288 2068
rect 37428 2012 37456 2068
rect 38038 2012 38066 2068
rect 38206 2012 38234 2068
rect 38816 2012 38844 2068
rect 38984 2012 39012 2068
rect 39594 2012 39622 2068
rect 39762 2012 39790 2068
rect 40372 2012 40400 2068
rect 40540 2012 40568 2068
rect 41150 2012 41178 2068
rect 41318 2012 41346 2068
rect 41928 2012 41956 2068
rect 42096 2012 42124 2068
rect 42706 2012 42734 2068
rect 42874 2012 42902 2068
rect 43484 2012 43512 2068
rect 43652 2012 43680 2068
rect 44262 2012 44290 2068
rect 44430 2012 44458 2068
rect 45040 2012 45068 2068
rect 45208 2012 45236 2068
rect 45818 2012 45846 2068
rect 45986 2012 46014 2068
rect 46596 2012 46624 2068
rect 46764 2012 46792 2068
rect 47374 2012 47402 2068
rect 47542 2012 47570 2068
rect 48152 2012 48180 2068
rect 48320 2012 48348 2068
rect 48930 2012 48958 2068
rect 49098 2012 49126 2068
rect 49708 2012 49736 2068
rect 84 192 112 560
rect 72 186 124 192
rect 72 128 124 134
rect 694 112 722 560
rect 862 192 890 560
rect 850 186 902 192
rect 850 128 902 134
rect 1472 112 1500 560
rect 1640 192 1668 560
rect 1628 186 1680 192
rect 1628 128 1680 134
rect 2250 112 2278 560
rect 2418 192 2446 560
rect 2406 186 2458 192
rect 2406 128 2458 134
rect 3028 112 3056 560
rect 3196 192 3224 560
rect 3184 186 3236 192
rect 3184 128 3236 134
rect 3806 112 3834 560
rect 3974 192 4002 560
rect 3962 186 4014 192
rect 3962 128 4014 134
rect 4584 112 4612 560
rect 4752 192 4780 560
rect 4740 186 4792 192
rect 4740 128 4792 134
rect 5362 112 5390 560
rect 5530 192 5558 560
rect 5518 186 5570 192
rect 5518 128 5570 134
rect 6140 112 6168 560
rect 6308 192 6336 560
rect 6296 186 6348 192
rect 6296 128 6348 134
rect 6918 112 6946 560
rect 7086 192 7114 560
rect 7074 186 7126 192
rect 7074 128 7126 134
rect 7696 112 7724 560
rect 7864 192 7892 560
rect 7852 186 7904 192
rect 7852 128 7904 134
rect 8474 112 8502 560
rect 8642 192 8670 560
rect 8630 186 8682 192
rect 8630 128 8682 134
rect 9252 112 9280 560
rect 9420 192 9448 560
rect 9408 186 9460 192
rect 9408 128 9460 134
rect 10030 112 10058 560
rect 10198 192 10226 560
rect 10186 186 10238 192
rect 10186 128 10238 134
rect 10808 112 10836 560
rect 10976 192 11004 560
rect 10964 186 11016 192
rect 10964 128 11016 134
rect 11586 112 11614 560
rect 11754 192 11782 560
rect 11742 186 11794 192
rect 11742 128 11794 134
rect 12364 112 12392 560
rect 12532 192 12560 560
rect 12520 186 12572 192
rect 12520 128 12572 134
rect 13142 112 13170 560
rect 13310 192 13338 560
rect 13298 186 13350 192
rect 13298 128 13350 134
rect 13920 112 13948 560
rect 14088 192 14116 560
rect 14076 186 14128 192
rect 14076 128 14128 134
rect 14698 112 14726 560
rect 14866 192 14894 560
rect 14854 186 14906 192
rect 14854 128 14906 134
rect 15476 112 15504 560
rect 15644 192 15672 560
rect 15632 186 15684 192
rect 15632 128 15684 134
rect 16254 112 16282 560
rect 16422 192 16450 560
rect 16410 186 16462 192
rect 16410 128 16462 134
rect 17032 112 17060 560
rect 17200 192 17228 560
rect 17188 186 17240 192
rect 17188 128 17240 134
rect 17810 112 17838 560
rect 17978 192 18006 560
rect 17966 186 18018 192
rect 17966 128 18018 134
rect 18588 112 18616 560
rect 18756 192 18784 560
rect 18744 186 18796 192
rect 18744 128 18796 134
rect 19366 112 19394 560
rect 19534 192 19562 560
rect 19522 186 19574 192
rect 19522 128 19574 134
rect 20144 112 20172 560
rect 20312 192 20340 560
rect 20300 186 20352 192
rect 20300 128 20352 134
rect 20922 112 20950 560
rect 21090 192 21118 560
rect 21078 186 21130 192
rect 21078 128 21130 134
rect 21700 112 21728 560
rect 21868 192 21896 560
rect 21856 186 21908 192
rect 21856 128 21908 134
rect 22478 112 22506 560
rect 22646 192 22674 560
rect 22634 186 22686 192
rect 22634 128 22686 134
rect 23256 112 23284 560
rect 23424 192 23452 560
rect 23412 186 23464 192
rect 23412 128 23464 134
rect 24034 112 24062 560
rect 24202 192 24230 560
rect 24190 186 24242 192
rect 24190 128 24242 134
rect 24812 112 24840 560
rect 24980 192 25008 560
rect 24968 186 25020 192
rect 24968 128 25020 134
rect 25590 112 25618 560
rect 25758 192 25786 560
rect 25746 186 25798 192
rect 25746 128 25798 134
rect 26368 112 26396 560
rect 26536 192 26564 560
rect 26524 186 26576 192
rect 26524 128 26576 134
rect 27146 112 27174 560
rect 27314 192 27342 560
rect 27302 186 27354 192
rect 27302 128 27354 134
rect 27924 112 27952 560
rect 28092 192 28120 560
rect 28080 186 28132 192
rect 28080 128 28132 134
rect 28702 112 28730 560
rect 28870 192 28898 560
rect 28858 186 28910 192
rect 28858 128 28910 134
rect 29480 112 29508 560
rect 29648 192 29676 560
rect 29636 186 29688 192
rect 29636 128 29688 134
rect 30258 112 30286 560
rect 30426 192 30454 560
rect 30414 186 30466 192
rect 30414 128 30466 134
rect 31036 112 31064 560
rect 31204 192 31232 560
rect 31192 186 31244 192
rect 31192 128 31244 134
rect 31814 112 31842 560
rect 31982 192 32010 560
rect 31970 186 32022 192
rect 31970 128 32022 134
rect 32592 112 32620 560
rect 32760 192 32788 560
rect 32748 186 32800 192
rect 32748 128 32800 134
rect 33370 112 33398 560
rect 33538 192 33566 560
rect 33526 186 33578 192
rect 33526 128 33578 134
rect 34148 112 34176 560
rect 34316 192 34344 560
rect 34304 186 34356 192
rect 34304 128 34356 134
rect 34926 112 34954 560
rect 35094 192 35122 560
rect 35082 186 35134 192
rect 35082 128 35134 134
rect 35704 112 35732 560
rect 35872 192 35900 560
rect 35860 186 35912 192
rect 35860 128 35912 134
rect 36482 112 36510 560
rect 36650 192 36678 560
rect 36638 186 36690 192
rect 36638 128 36690 134
rect 37260 112 37288 560
rect 37428 192 37456 560
rect 37416 186 37468 192
rect 37416 128 37468 134
rect 38038 112 38066 560
rect 38206 192 38234 560
rect 38194 186 38246 192
rect 38194 128 38246 134
rect 38816 112 38844 560
rect 38984 192 39012 560
rect 38972 186 39024 192
rect 38972 128 39024 134
rect 39594 112 39622 560
rect 39762 192 39790 560
rect 39750 186 39802 192
rect 39750 128 39802 134
rect 40372 112 40400 560
rect 40540 192 40568 560
rect 40528 186 40580 192
rect 40528 128 40580 134
rect 41150 112 41178 560
rect 41318 192 41346 560
rect 41306 186 41358 192
rect 41306 128 41358 134
rect 41928 112 41956 560
rect 42096 192 42124 560
rect 42084 186 42136 192
rect 42084 128 42136 134
rect 42706 112 42734 560
rect 42874 192 42902 560
rect 42862 186 42914 192
rect 42862 128 42914 134
rect 43484 112 43512 560
rect 43652 192 43680 560
rect 43640 186 43692 192
rect 43640 128 43692 134
rect 44262 112 44290 560
rect 44430 192 44458 560
rect 44418 186 44470 192
rect 44418 128 44470 134
rect 45040 112 45068 560
rect 45208 192 45236 560
rect 45196 186 45248 192
rect 45196 128 45248 134
rect 45818 112 45846 560
rect 45986 192 46014 560
rect 45974 186 46026 192
rect 45974 128 46026 134
rect 46596 112 46624 560
rect 46764 192 46792 560
rect 46752 186 46804 192
rect 46752 128 46804 134
rect 47374 112 47402 560
rect 47542 192 47570 560
rect 47530 186 47582 192
rect 47530 128 47582 134
rect 48152 112 48180 560
rect 48320 192 48348 560
rect 48308 186 48360 192
rect 48308 128 48360 134
rect 48930 112 48958 560
rect 49098 192 49126 560
rect 49086 186 49138 192
rect 49086 128 49138 134
rect 49708 112 49736 560
rect 682 106 734 112
rect 682 48 734 54
rect 1460 106 1512 112
rect 1460 48 1512 54
rect 2238 106 2290 112
rect 2238 48 2290 54
rect 3016 106 3068 112
rect 3016 48 3068 54
rect 3794 106 3846 112
rect 3794 48 3846 54
rect 4572 106 4624 112
rect 4572 48 4624 54
rect 5350 106 5402 112
rect 5350 48 5402 54
rect 6128 106 6180 112
rect 6128 48 6180 54
rect 6906 106 6958 112
rect 6906 48 6958 54
rect 7684 106 7736 112
rect 7684 48 7736 54
rect 8462 106 8514 112
rect 8462 48 8514 54
rect 9240 106 9292 112
rect 9240 48 9292 54
rect 10018 106 10070 112
rect 10018 48 10070 54
rect 10796 106 10848 112
rect 10796 48 10848 54
rect 11574 106 11626 112
rect 11574 48 11626 54
rect 12352 106 12404 112
rect 12352 48 12404 54
rect 13130 106 13182 112
rect 13130 48 13182 54
rect 13908 106 13960 112
rect 13908 48 13960 54
rect 14686 106 14738 112
rect 14686 48 14738 54
rect 15464 106 15516 112
rect 15464 48 15516 54
rect 16242 106 16294 112
rect 16242 48 16294 54
rect 17020 106 17072 112
rect 17020 48 17072 54
rect 17798 106 17850 112
rect 17798 48 17850 54
rect 18576 106 18628 112
rect 18576 48 18628 54
rect 19354 106 19406 112
rect 19354 48 19406 54
rect 20132 106 20184 112
rect 20132 48 20184 54
rect 20910 106 20962 112
rect 20910 48 20962 54
rect 21688 106 21740 112
rect 21688 48 21740 54
rect 22466 106 22518 112
rect 22466 48 22518 54
rect 23244 106 23296 112
rect 23244 48 23296 54
rect 24022 106 24074 112
rect 24022 48 24074 54
rect 24800 106 24852 112
rect 24800 48 24852 54
rect 25578 106 25630 112
rect 25578 48 25630 54
rect 26356 106 26408 112
rect 26356 48 26408 54
rect 27134 106 27186 112
rect 27134 48 27186 54
rect 27912 106 27964 112
rect 27912 48 27964 54
rect 28690 106 28742 112
rect 28690 48 28742 54
rect 29468 106 29520 112
rect 29468 48 29520 54
rect 30246 106 30298 112
rect 30246 48 30298 54
rect 31024 106 31076 112
rect 31024 48 31076 54
rect 31802 106 31854 112
rect 31802 48 31854 54
rect 32580 106 32632 112
rect 32580 48 32632 54
rect 33358 106 33410 112
rect 33358 48 33410 54
rect 34136 106 34188 112
rect 34136 48 34188 54
rect 34914 106 34966 112
rect 34914 48 34966 54
rect 35692 106 35744 112
rect 35692 48 35744 54
rect 36470 106 36522 112
rect 36470 48 36522 54
rect 37248 106 37300 112
rect 37248 48 37300 54
rect 38026 106 38078 112
rect 38026 48 38078 54
rect 38804 106 38856 112
rect 38804 48 38856 54
rect 39582 106 39634 112
rect 39582 48 39634 54
rect 40360 106 40412 112
rect 40360 48 40412 54
rect 41138 106 41190 112
rect 41138 48 41190 54
rect 41916 106 41968 112
rect 41916 48 41968 54
rect 42694 106 42746 112
rect 42694 48 42746 54
rect 43472 106 43524 112
rect 43472 48 43524 54
rect 44250 106 44302 112
rect 44250 48 44302 54
rect 45028 106 45080 112
rect 45028 48 45080 54
rect 45806 106 45858 112
rect 45806 48 45858 54
rect 46584 106 46636 112
rect 46584 48 46636 54
rect 47362 106 47414 112
rect 47362 48 47414 54
rect 48140 106 48192 112
rect 48140 48 48192 54
rect 48918 106 48970 112
rect 48918 48 48970 54
rect 49696 106 49748 112
rect 49696 48 49748 54
<< metal3 >>
rect 712 1282 844 1356
rect 1490 1282 1622 1356
rect 2268 1282 2400 1356
rect 3046 1282 3178 1356
rect 3824 1282 3956 1356
rect 4602 1282 4734 1356
rect 5380 1282 5512 1356
rect 6158 1282 6290 1356
rect 6936 1282 7068 1356
rect 7714 1282 7846 1356
rect 8492 1282 8624 1356
rect 9270 1282 9402 1356
rect 10048 1282 10180 1356
rect 10826 1282 10958 1356
rect 11604 1282 11736 1356
rect 12382 1282 12514 1356
rect 13160 1282 13292 1356
rect 13938 1282 14070 1356
rect 14716 1282 14848 1356
rect 15494 1282 15626 1356
rect 16272 1282 16404 1356
rect 17050 1282 17182 1356
rect 17828 1282 17960 1356
rect 18606 1282 18738 1356
rect 19384 1282 19516 1356
rect 20162 1282 20294 1356
rect 20940 1282 21072 1356
rect 21718 1282 21850 1356
rect 22496 1282 22628 1356
rect 23274 1282 23406 1356
rect 24052 1282 24184 1356
rect 24830 1282 24962 1356
rect 25608 1282 25740 1356
rect 26386 1282 26518 1356
rect 27164 1282 27296 1356
rect 27942 1282 28074 1356
rect 28720 1282 28852 1356
rect 29498 1282 29630 1356
rect 30276 1282 30408 1356
rect 31054 1282 31186 1356
rect 31832 1282 31964 1356
rect 32610 1282 32742 1356
rect 33388 1282 33520 1356
rect 34166 1282 34298 1356
rect 34944 1282 35076 1356
rect 35722 1282 35854 1356
rect 36500 1282 36632 1356
rect 37278 1282 37410 1356
rect 38056 1282 38188 1356
rect 38834 1282 38966 1356
rect 39612 1282 39744 1356
rect 40390 1282 40522 1356
rect 41168 1282 41300 1356
rect 41946 1282 42078 1356
rect 42724 1282 42856 1356
rect 43502 1282 43634 1356
rect 44280 1282 44412 1356
rect 45058 1282 45190 1356
rect 45836 1282 45968 1356
rect 46614 1282 46746 1356
rect 47392 1282 47524 1356
rect 48170 1282 48302 1356
rect 48948 1282 49080 1356
rect 49726 1282 49858 1356
use contact_14  contact_14_0
timestamp 1644951705
transform 1 0 49690 0 1 48
box 0 0 1 1
use contact_14  contact_14_1
timestamp 1644951705
transform 1 0 49080 0 1 128
box 0 0 1 1
use contact_14  contact_14_2
timestamp 1644951705
transform 1 0 48912 0 1 48
box 0 0 1 1
use contact_14  contact_14_3
timestamp 1644951705
transform 1 0 48302 0 1 128
box 0 0 1 1
use contact_14  contact_14_4
timestamp 1644951705
transform 1 0 48134 0 1 48
box 0 0 1 1
use contact_14  contact_14_5
timestamp 1644951705
transform 1 0 47524 0 1 128
box 0 0 1 1
use contact_14  contact_14_6
timestamp 1644951705
transform 1 0 47356 0 1 48
box 0 0 1 1
use contact_14  contact_14_7
timestamp 1644951705
transform 1 0 46746 0 1 128
box 0 0 1 1
use contact_14  contact_14_8
timestamp 1644951705
transform 1 0 46578 0 1 48
box 0 0 1 1
use contact_14  contact_14_9
timestamp 1644951705
transform 1 0 45968 0 1 128
box 0 0 1 1
use contact_14  contact_14_10
timestamp 1644951705
transform 1 0 45800 0 1 48
box 0 0 1 1
use contact_14  contact_14_11
timestamp 1644951705
transform 1 0 45190 0 1 128
box 0 0 1 1
use contact_14  contact_14_12
timestamp 1644951705
transform 1 0 45022 0 1 48
box 0 0 1 1
use contact_14  contact_14_13
timestamp 1644951705
transform 1 0 44412 0 1 128
box 0 0 1 1
use contact_14  contact_14_14
timestamp 1644951705
transform 1 0 44244 0 1 48
box 0 0 1 1
use contact_14  contact_14_15
timestamp 1644951705
transform 1 0 43634 0 1 128
box 0 0 1 1
use contact_14  contact_14_16
timestamp 1644951705
transform 1 0 43466 0 1 48
box 0 0 1 1
use contact_14  contact_14_17
timestamp 1644951705
transform 1 0 42856 0 1 128
box 0 0 1 1
use contact_14  contact_14_18
timestamp 1644951705
transform 1 0 42688 0 1 48
box 0 0 1 1
use contact_14  contact_14_19
timestamp 1644951705
transform 1 0 42078 0 1 128
box 0 0 1 1
use contact_14  contact_14_20
timestamp 1644951705
transform 1 0 41910 0 1 48
box 0 0 1 1
use contact_14  contact_14_21
timestamp 1644951705
transform 1 0 41300 0 1 128
box 0 0 1 1
use contact_14  contact_14_22
timestamp 1644951705
transform 1 0 41132 0 1 48
box 0 0 1 1
use contact_14  contact_14_23
timestamp 1644951705
transform 1 0 40522 0 1 128
box 0 0 1 1
use contact_14  contact_14_24
timestamp 1644951705
transform 1 0 40354 0 1 48
box 0 0 1 1
use contact_14  contact_14_25
timestamp 1644951705
transform 1 0 39744 0 1 128
box 0 0 1 1
use contact_14  contact_14_26
timestamp 1644951705
transform 1 0 39576 0 1 48
box 0 0 1 1
use contact_14  contact_14_27
timestamp 1644951705
transform 1 0 38966 0 1 128
box 0 0 1 1
use contact_14  contact_14_28
timestamp 1644951705
transform 1 0 38798 0 1 48
box 0 0 1 1
use contact_14  contact_14_29
timestamp 1644951705
transform 1 0 38188 0 1 128
box 0 0 1 1
use contact_14  contact_14_30
timestamp 1644951705
transform 1 0 38020 0 1 48
box 0 0 1 1
use contact_14  contact_14_31
timestamp 1644951705
transform 1 0 37410 0 1 128
box 0 0 1 1
use contact_14  contact_14_32
timestamp 1644951705
transform 1 0 37242 0 1 48
box 0 0 1 1
use contact_14  contact_14_33
timestamp 1644951705
transform 1 0 36632 0 1 128
box 0 0 1 1
use contact_14  contact_14_34
timestamp 1644951705
transform 1 0 36464 0 1 48
box 0 0 1 1
use contact_14  contact_14_35
timestamp 1644951705
transform 1 0 35854 0 1 128
box 0 0 1 1
use contact_14  contact_14_36
timestamp 1644951705
transform 1 0 35686 0 1 48
box 0 0 1 1
use contact_14  contact_14_37
timestamp 1644951705
transform 1 0 35076 0 1 128
box 0 0 1 1
use contact_14  contact_14_38
timestamp 1644951705
transform 1 0 34908 0 1 48
box 0 0 1 1
use contact_14  contact_14_39
timestamp 1644951705
transform 1 0 34298 0 1 128
box 0 0 1 1
use contact_14  contact_14_40
timestamp 1644951705
transform 1 0 34130 0 1 48
box 0 0 1 1
use contact_14  contact_14_41
timestamp 1644951705
transform 1 0 33520 0 1 128
box 0 0 1 1
use contact_14  contact_14_42
timestamp 1644951705
transform 1 0 33352 0 1 48
box 0 0 1 1
use contact_14  contact_14_43
timestamp 1644951705
transform 1 0 32742 0 1 128
box 0 0 1 1
use contact_14  contact_14_44
timestamp 1644951705
transform 1 0 32574 0 1 48
box 0 0 1 1
use contact_14  contact_14_45
timestamp 1644951705
transform 1 0 31964 0 1 128
box 0 0 1 1
use contact_14  contact_14_46
timestamp 1644951705
transform 1 0 31796 0 1 48
box 0 0 1 1
use contact_14  contact_14_47
timestamp 1644951705
transform 1 0 31186 0 1 128
box 0 0 1 1
use contact_14  contact_14_48
timestamp 1644951705
transform 1 0 31018 0 1 48
box 0 0 1 1
use contact_14  contact_14_49
timestamp 1644951705
transform 1 0 30408 0 1 128
box 0 0 1 1
use contact_14  contact_14_50
timestamp 1644951705
transform 1 0 30240 0 1 48
box 0 0 1 1
use contact_14  contact_14_51
timestamp 1644951705
transform 1 0 29630 0 1 128
box 0 0 1 1
use contact_14  contact_14_52
timestamp 1644951705
transform 1 0 29462 0 1 48
box 0 0 1 1
use contact_14  contact_14_53
timestamp 1644951705
transform 1 0 28852 0 1 128
box 0 0 1 1
use contact_14  contact_14_54
timestamp 1644951705
transform 1 0 28684 0 1 48
box 0 0 1 1
use contact_14  contact_14_55
timestamp 1644951705
transform 1 0 28074 0 1 128
box 0 0 1 1
use contact_14  contact_14_56
timestamp 1644951705
transform 1 0 27906 0 1 48
box 0 0 1 1
use contact_14  contact_14_57
timestamp 1644951705
transform 1 0 27296 0 1 128
box 0 0 1 1
use contact_14  contact_14_58
timestamp 1644951705
transform 1 0 27128 0 1 48
box 0 0 1 1
use contact_14  contact_14_59
timestamp 1644951705
transform 1 0 26518 0 1 128
box 0 0 1 1
use contact_14  contact_14_60
timestamp 1644951705
transform 1 0 26350 0 1 48
box 0 0 1 1
use contact_14  contact_14_61
timestamp 1644951705
transform 1 0 25740 0 1 128
box 0 0 1 1
use contact_14  contact_14_62
timestamp 1644951705
transform 1 0 25572 0 1 48
box 0 0 1 1
use contact_14  contact_14_63
timestamp 1644951705
transform 1 0 24962 0 1 128
box 0 0 1 1
use contact_14  contact_14_64
timestamp 1644951705
transform 1 0 24794 0 1 48
box 0 0 1 1
use contact_14  contact_14_65
timestamp 1644951705
transform 1 0 24184 0 1 128
box 0 0 1 1
use contact_14  contact_14_66
timestamp 1644951705
transform 1 0 24016 0 1 48
box 0 0 1 1
use contact_14  contact_14_67
timestamp 1644951705
transform 1 0 23406 0 1 128
box 0 0 1 1
use contact_14  contact_14_68
timestamp 1644951705
transform 1 0 23238 0 1 48
box 0 0 1 1
use contact_14  contact_14_69
timestamp 1644951705
transform 1 0 22628 0 1 128
box 0 0 1 1
use contact_14  contact_14_70
timestamp 1644951705
transform 1 0 22460 0 1 48
box 0 0 1 1
use contact_14  contact_14_71
timestamp 1644951705
transform 1 0 21850 0 1 128
box 0 0 1 1
use contact_14  contact_14_72
timestamp 1644951705
transform 1 0 21682 0 1 48
box 0 0 1 1
use contact_14  contact_14_73
timestamp 1644951705
transform 1 0 21072 0 1 128
box 0 0 1 1
use contact_14  contact_14_74
timestamp 1644951705
transform 1 0 20904 0 1 48
box 0 0 1 1
use contact_14  contact_14_75
timestamp 1644951705
transform 1 0 20294 0 1 128
box 0 0 1 1
use contact_14  contact_14_76
timestamp 1644951705
transform 1 0 20126 0 1 48
box 0 0 1 1
use contact_14  contact_14_77
timestamp 1644951705
transform 1 0 19516 0 1 128
box 0 0 1 1
use contact_14  contact_14_78
timestamp 1644951705
transform 1 0 19348 0 1 48
box 0 0 1 1
use contact_14  contact_14_79
timestamp 1644951705
transform 1 0 18738 0 1 128
box 0 0 1 1
use contact_14  contact_14_80
timestamp 1644951705
transform 1 0 18570 0 1 48
box 0 0 1 1
use contact_14  contact_14_81
timestamp 1644951705
transform 1 0 17960 0 1 128
box 0 0 1 1
use contact_14  contact_14_82
timestamp 1644951705
transform 1 0 17792 0 1 48
box 0 0 1 1
use contact_14  contact_14_83
timestamp 1644951705
transform 1 0 17182 0 1 128
box 0 0 1 1
use contact_14  contact_14_84
timestamp 1644951705
transform 1 0 17014 0 1 48
box 0 0 1 1
use contact_14  contact_14_85
timestamp 1644951705
transform 1 0 16404 0 1 128
box 0 0 1 1
use contact_14  contact_14_86
timestamp 1644951705
transform 1 0 16236 0 1 48
box 0 0 1 1
use contact_14  contact_14_87
timestamp 1644951705
transform 1 0 15626 0 1 128
box 0 0 1 1
use contact_14  contact_14_88
timestamp 1644951705
transform 1 0 15458 0 1 48
box 0 0 1 1
use contact_14  contact_14_89
timestamp 1644951705
transform 1 0 14848 0 1 128
box 0 0 1 1
use contact_14  contact_14_90
timestamp 1644951705
transform 1 0 14680 0 1 48
box 0 0 1 1
use contact_14  contact_14_91
timestamp 1644951705
transform 1 0 14070 0 1 128
box 0 0 1 1
use contact_14  contact_14_92
timestamp 1644951705
transform 1 0 13902 0 1 48
box 0 0 1 1
use contact_14  contact_14_93
timestamp 1644951705
transform 1 0 13292 0 1 128
box 0 0 1 1
use contact_14  contact_14_94
timestamp 1644951705
transform 1 0 13124 0 1 48
box 0 0 1 1
use contact_14  contact_14_95
timestamp 1644951705
transform 1 0 12514 0 1 128
box 0 0 1 1
use contact_14  contact_14_96
timestamp 1644951705
transform 1 0 12346 0 1 48
box 0 0 1 1
use contact_14  contact_14_97
timestamp 1644951705
transform 1 0 11736 0 1 128
box 0 0 1 1
use contact_14  contact_14_98
timestamp 1644951705
transform 1 0 11568 0 1 48
box 0 0 1 1
use contact_14  contact_14_99
timestamp 1644951705
transform 1 0 10958 0 1 128
box 0 0 1 1
use contact_14  contact_14_100
timestamp 1644951705
transform 1 0 10790 0 1 48
box 0 0 1 1
use contact_14  contact_14_101
timestamp 1644951705
transform 1 0 10180 0 1 128
box 0 0 1 1
use contact_14  contact_14_102
timestamp 1644951705
transform 1 0 10012 0 1 48
box 0 0 1 1
use contact_14  contact_14_103
timestamp 1644951705
transform 1 0 9402 0 1 128
box 0 0 1 1
use contact_14  contact_14_104
timestamp 1644951705
transform 1 0 9234 0 1 48
box 0 0 1 1
use contact_14  contact_14_105
timestamp 1644951705
transform 1 0 8624 0 1 128
box 0 0 1 1
use contact_14  contact_14_106
timestamp 1644951705
transform 1 0 8456 0 1 48
box 0 0 1 1
use contact_14  contact_14_107
timestamp 1644951705
transform 1 0 7846 0 1 128
box 0 0 1 1
use contact_14  contact_14_108
timestamp 1644951705
transform 1 0 7678 0 1 48
box 0 0 1 1
use contact_14  contact_14_109
timestamp 1644951705
transform 1 0 7068 0 1 128
box 0 0 1 1
use contact_14  contact_14_110
timestamp 1644951705
transform 1 0 6900 0 1 48
box 0 0 1 1
use contact_14  contact_14_111
timestamp 1644951705
transform 1 0 6290 0 1 128
box 0 0 1 1
use contact_14  contact_14_112
timestamp 1644951705
transform 1 0 6122 0 1 48
box 0 0 1 1
use contact_14  contact_14_113
timestamp 1644951705
transform 1 0 5512 0 1 128
box 0 0 1 1
use contact_14  contact_14_114
timestamp 1644951705
transform 1 0 5344 0 1 48
box 0 0 1 1
use contact_14  contact_14_115
timestamp 1644951705
transform 1 0 4734 0 1 128
box 0 0 1 1
use contact_14  contact_14_116
timestamp 1644951705
transform 1 0 4566 0 1 48
box 0 0 1 1
use contact_14  contact_14_117
timestamp 1644951705
transform 1 0 3956 0 1 128
box 0 0 1 1
use contact_14  contact_14_118
timestamp 1644951705
transform 1 0 3788 0 1 48
box 0 0 1 1
use contact_14  contact_14_119
timestamp 1644951705
transform 1 0 3178 0 1 128
box 0 0 1 1
use contact_14  contact_14_120
timestamp 1644951705
transform 1 0 3010 0 1 48
box 0 0 1 1
use contact_14  contact_14_121
timestamp 1644951705
transform 1 0 2400 0 1 128
box 0 0 1 1
use contact_14  contact_14_122
timestamp 1644951705
transform 1 0 2232 0 1 48
box 0 0 1 1
use contact_14  contact_14_123
timestamp 1644951705
transform 1 0 1622 0 1 128
box 0 0 1 1
use contact_14  contact_14_124
timestamp 1644951705
transform 1 0 1454 0 1 48
box 0 0 1 1
use contact_14  contact_14_125
timestamp 1644951705
transform 1 0 844 0 1 128
box 0 0 1 1
use contact_14  contact_14_126
timestamp 1644951705
transform 1 0 676 0 1 48
box 0 0 1 1
use contact_14  contact_14_127
timestamp 1644951705
transform 1 0 66 0 1 128
box 0 0 1 1
use contact_27  contact_27_0
timestamp 1644951705
transform 1 0 49374 0 1 471
box 0 0 1 1
use contact_26  contact_26_0
timestamp 1644951705
transform 1 0 49370 0 1 461
box 0 0 1 1
use contact_27  contact_27_1
timestamp 1644951705
transform 1 0 48596 0 1 391
box 0 0 1 1
use contact_26  contact_26_1
timestamp 1644951705
transform 1 0 48592 0 1 381
box 0 0 1 1
use contact_27  contact_27_2
timestamp 1644951705
transform 1 0 47818 0 1 311
box 0 0 1 1
use contact_26  contact_26_2
timestamp 1644951705
transform 1 0 47814 0 1 301
box 0 0 1 1
use contact_27  contact_27_3
timestamp 1644951705
transform 1 0 47040 0 1 231
box 0 0 1 1
use contact_26  contact_26_3
timestamp 1644951705
transform 1 0 47036 0 1 221
box 0 0 1 1
use contact_27  contact_27_4
timestamp 1644951705
transform 1 0 46262 0 1 471
box 0 0 1 1
use contact_26  contact_26_4
timestamp 1644951705
transform 1 0 46258 0 1 461
box 0 0 1 1
use contact_27  contact_27_5
timestamp 1644951705
transform 1 0 45484 0 1 391
box 0 0 1 1
use contact_26  contact_26_5
timestamp 1644951705
transform 1 0 45480 0 1 381
box 0 0 1 1
use contact_27  contact_27_6
timestamp 1644951705
transform 1 0 44706 0 1 311
box 0 0 1 1
use contact_26  contact_26_6
timestamp 1644951705
transform 1 0 44702 0 1 301
box 0 0 1 1
use contact_27  contact_27_7
timestamp 1644951705
transform 1 0 43928 0 1 231
box 0 0 1 1
use contact_26  contact_26_7
timestamp 1644951705
transform 1 0 43924 0 1 221
box 0 0 1 1
use contact_27  contact_27_8
timestamp 1644951705
transform 1 0 43150 0 1 471
box 0 0 1 1
use contact_26  contact_26_8
timestamp 1644951705
transform 1 0 43146 0 1 461
box 0 0 1 1
use contact_27  contact_27_9
timestamp 1644951705
transform 1 0 42372 0 1 391
box 0 0 1 1
use contact_26  contact_26_9
timestamp 1644951705
transform 1 0 42368 0 1 381
box 0 0 1 1
use contact_27  contact_27_10
timestamp 1644951705
transform 1 0 41594 0 1 311
box 0 0 1 1
use contact_26  contact_26_10
timestamp 1644951705
transform 1 0 41590 0 1 301
box 0 0 1 1
use contact_27  contact_27_11
timestamp 1644951705
transform 1 0 40816 0 1 231
box 0 0 1 1
use contact_26  contact_26_11
timestamp 1644951705
transform 1 0 40812 0 1 221
box 0 0 1 1
use contact_27  contact_27_12
timestamp 1644951705
transform 1 0 40038 0 1 471
box 0 0 1 1
use contact_26  contact_26_12
timestamp 1644951705
transform 1 0 40034 0 1 461
box 0 0 1 1
use contact_27  contact_27_13
timestamp 1644951705
transform 1 0 39260 0 1 391
box 0 0 1 1
use contact_26  contact_26_13
timestamp 1644951705
transform 1 0 39256 0 1 381
box 0 0 1 1
use contact_27  contact_27_14
timestamp 1644951705
transform 1 0 38482 0 1 311
box 0 0 1 1
use contact_26  contact_26_14
timestamp 1644951705
transform 1 0 38478 0 1 301
box 0 0 1 1
use contact_27  contact_27_15
timestamp 1644951705
transform 1 0 37704 0 1 231
box 0 0 1 1
use contact_26  contact_26_15
timestamp 1644951705
transform 1 0 37700 0 1 221
box 0 0 1 1
use contact_27  contact_27_16
timestamp 1644951705
transform 1 0 36926 0 1 471
box 0 0 1 1
use contact_26  contact_26_16
timestamp 1644951705
transform 1 0 36922 0 1 461
box 0 0 1 1
use contact_27  contact_27_17
timestamp 1644951705
transform 1 0 36148 0 1 391
box 0 0 1 1
use contact_26  contact_26_17
timestamp 1644951705
transform 1 0 36144 0 1 381
box 0 0 1 1
use contact_27  contact_27_18
timestamp 1644951705
transform 1 0 35370 0 1 311
box 0 0 1 1
use contact_26  contact_26_18
timestamp 1644951705
transform 1 0 35366 0 1 301
box 0 0 1 1
use contact_27  contact_27_19
timestamp 1644951705
transform 1 0 34592 0 1 231
box 0 0 1 1
use contact_26  contact_26_19
timestamp 1644951705
transform 1 0 34588 0 1 221
box 0 0 1 1
use contact_27  contact_27_20
timestamp 1644951705
transform 1 0 33814 0 1 471
box 0 0 1 1
use contact_26  contact_26_20
timestamp 1644951705
transform 1 0 33810 0 1 461
box 0 0 1 1
use contact_27  contact_27_21
timestamp 1644951705
transform 1 0 33036 0 1 391
box 0 0 1 1
use contact_26  contact_26_21
timestamp 1644951705
transform 1 0 33032 0 1 381
box 0 0 1 1
use contact_27  contact_27_22
timestamp 1644951705
transform 1 0 32258 0 1 311
box 0 0 1 1
use contact_26  contact_26_22
timestamp 1644951705
transform 1 0 32254 0 1 301
box 0 0 1 1
use contact_27  contact_27_23
timestamp 1644951705
transform 1 0 31480 0 1 231
box 0 0 1 1
use contact_26  contact_26_23
timestamp 1644951705
transform 1 0 31476 0 1 221
box 0 0 1 1
use contact_27  contact_27_24
timestamp 1644951705
transform 1 0 30702 0 1 471
box 0 0 1 1
use contact_26  contact_26_24
timestamp 1644951705
transform 1 0 30698 0 1 461
box 0 0 1 1
use contact_27  contact_27_25
timestamp 1644951705
transform 1 0 29924 0 1 391
box 0 0 1 1
use contact_26  contact_26_25
timestamp 1644951705
transform 1 0 29920 0 1 381
box 0 0 1 1
use contact_27  contact_27_26
timestamp 1644951705
transform 1 0 29146 0 1 311
box 0 0 1 1
use contact_26  contact_26_26
timestamp 1644951705
transform 1 0 29142 0 1 301
box 0 0 1 1
use contact_27  contact_27_27
timestamp 1644951705
transform 1 0 28368 0 1 231
box 0 0 1 1
use contact_26  contact_26_27
timestamp 1644951705
transform 1 0 28364 0 1 221
box 0 0 1 1
use contact_27  contact_27_28
timestamp 1644951705
transform 1 0 27590 0 1 471
box 0 0 1 1
use contact_26  contact_26_28
timestamp 1644951705
transform 1 0 27586 0 1 461
box 0 0 1 1
use contact_27  contact_27_29
timestamp 1644951705
transform 1 0 26812 0 1 391
box 0 0 1 1
use contact_26  contact_26_29
timestamp 1644951705
transform 1 0 26808 0 1 381
box 0 0 1 1
use contact_27  contact_27_30
timestamp 1644951705
transform 1 0 26034 0 1 311
box 0 0 1 1
use contact_26  contact_26_30
timestamp 1644951705
transform 1 0 26030 0 1 301
box 0 0 1 1
use contact_27  contact_27_31
timestamp 1644951705
transform 1 0 25256 0 1 231
box 0 0 1 1
use contact_26  contact_26_31
timestamp 1644951705
transform 1 0 25252 0 1 221
box 0 0 1 1
use contact_27  contact_27_32
timestamp 1644951705
transform 1 0 24478 0 1 471
box 0 0 1 1
use contact_26  contact_26_32
timestamp 1644951705
transform 1 0 24474 0 1 461
box 0 0 1 1
use contact_27  contact_27_33
timestamp 1644951705
transform 1 0 23700 0 1 391
box 0 0 1 1
use contact_26  contact_26_33
timestamp 1644951705
transform 1 0 23696 0 1 381
box 0 0 1 1
use contact_27  contact_27_34
timestamp 1644951705
transform 1 0 22922 0 1 311
box 0 0 1 1
use contact_26  contact_26_34
timestamp 1644951705
transform 1 0 22918 0 1 301
box 0 0 1 1
use contact_27  contact_27_35
timestamp 1644951705
transform 1 0 22144 0 1 231
box 0 0 1 1
use contact_26  contact_26_35
timestamp 1644951705
transform 1 0 22140 0 1 221
box 0 0 1 1
use contact_27  contact_27_36
timestamp 1644951705
transform 1 0 21366 0 1 471
box 0 0 1 1
use contact_26  contact_26_36
timestamp 1644951705
transform 1 0 21362 0 1 461
box 0 0 1 1
use contact_27  contact_27_37
timestamp 1644951705
transform 1 0 20588 0 1 391
box 0 0 1 1
use contact_26  contact_26_37
timestamp 1644951705
transform 1 0 20584 0 1 381
box 0 0 1 1
use contact_27  contact_27_38
timestamp 1644951705
transform 1 0 19810 0 1 311
box 0 0 1 1
use contact_26  contact_26_38
timestamp 1644951705
transform 1 0 19806 0 1 301
box 0 0 1 1
use contact_27  contact_27_39
timestamp 1644951705
transform 1 0 19032 0 1 231
box 0 0 1 1
use contact_26  contact_26_39
timestamp 1644951705
transform 1 0 19028 0 1 221
box 0 0 1 1
use contact_27  contact_27_40
timestamp 1644951705
transform 1 0 18254 0 1 471
box 0 0 1 1
use contact_26  contact_26_40
timestamp 1644951705
transform 1 0 18250 0 1 461
box 0 0 1 1
use contact_27  contact_27_41
timestamp 1644951705
transform 1 0 17476 0 1 391
box 0 0 1 1
use contact_26  contact_26_41
timestamp 1644951705
transform 1 0 17472 0 1 381
box 0 0 1 1
use contact_27  contact_27_42
timestamp 1644951705
transform 1 0 16698 0 1 311
box 0 0 1 1
use contact_26  contact_26_42
timestamp 1644951705
transform 1 0 16694 0 1 301
box 0 0 1 1
use contact_27  contact_27_43
timestamp 1644951705
transform 1 0 15920 0 1 231
box 0 0 1 1
use contact_26  contact_26_43
timestamp 1644951705
transform 1 0 15916 0 1 221
box 0 0 1 1
use contact_27  contact_27_44
timestamp 1644951705
transform 1 0 15142 0 1 471
box 0 0 1 1
use contact_26  contact_26_44
timestamp 1644951705
transform 1 0 15138 0 1 461
box 0 0 1 1
use contact_27  contact_27_45
timestamp 1644951705
transform 1 0 14364 0 1 391
box 0 0 1 1
use contact_26  contact_26_45
timestamp 1644951705
transform 1 0 14360 0 1 381
box 0 0 1 1
use contact_27  contact_27_46
timestamp 1644951705
transform 1 0 13586 0 1 311
box 0 0 1 1
use contact_26  contact_26_46
timestamp 1644951705
transform 1 0 13582 0 1 301
box 0 0 1 1
use contact_27  contact_27_47
timestamp 1644951705
transform 1 0 12808 0 1 231
box 0 0 1 1
use contact_26  contact_26_47
timestamp 1644951705
transform 1 0 12804 0 1 221
box 0 0 1 1
use contact_27  contact_27_48
timestamp 1644951705
transform 1 0 12030 0 1 471
box 0 0 1 1
use contact_26  contact_26_48
timestamp 1644951705
transform 1 0 12026 0 1 461
box 0 0 1 1
use contact_27  contact_27_49
timestamp 1644951705
transform 1 0 11252 0 1 391
box 0 0 1 1
use contact_26  contact_26_49
timestamp 1644951705
transform 1 0 11248 0 1 381
box 0 0 1 1
use contact_27  contact_27_50
timestamp 1644951705
transform 1 0 10474 0 1 311
box 0 0 1 1
use contact_26  contact_26_50
timestamp 1644951705
transform 1 0 10470 0 1 301
box 0 0 1 1
use contact_27  contact_27_51
timestamp 1644951705
transform 1 0 9696 0 1 231
box 0 0 1 1
use contact_26  contact_26_51
timestamp 1644951705
transform 1 0 9692 0 1 221
box 0 0 1 1
use contact_27  contact_27_52
timestamp 1644951705
transform 1 0 8918 0 1 471
box 0 0 1 1
use contact_26  contact_26_52
timestamp 1644951705
transform 1 0 8914 0 1 461
box 0 0 1 1
use contact_27  contact_27_53
timestamp 1644951705
transform 1 0 8140 0 1 391
box 0 0 1 1
use contact_26  contact_26_53
timestamp 1644951705
transform 1 0 8136 0 1 381
box 0 0 1 1
use contact_27  contact_27_54
timestamp 1644951705
transform 1 0 7362 0 1 311
box 0 0 1 1
use contact_26  contact_26_54
timestamp 1644951705
transform 1 0 7358 0 1 301
box 0 0 1 1
use contact_27  contact_27_55
timestamp 1644951705
transform 1 0 6584 0 1 231
box 0 0 1 1
use contact_26  contact_26_55
timestamp 1644951705
transform 1 0 6580 0 1 221
box 0 0 1 1
use contact_27  contact_27_56
timestamp 1644951705
transform 1 0 5806 0 1 471
box 0 0 1 1
use contact_26  contact_26_56
timestamp 1644951705
transform 1 0 5802 0 1 461
box 0 0 1 1
use contact_27  contact_27_57
timestamp 1644951705
transform 1 0 5028 0 1 391
box 0 0 1 1
use contact_26  contact_26_57
timestamp 1644951705
transform 1 0 5024 0 1 381
box 0 0 1 1
use contact_27  contact_27_58
timestamp 1644951705
transform 1 0 4250 0 1 311
box 0 0 1 1
use contact_26  contact_26_58
timestamp 1644951705
transform 1 0 4246 0 1 301
box 0 0 1 1
use contact_27  contact_27_59
timestamp 1644951705
transform 1 0 3472 0 1 231
box 0 0 1 1
use contact_26  contact_26_59
timestamp 1644951705
transform 1 0 3468 0 1 221
box 0 0 1 1
use contact_27  contact_27_60
timestamp 1644951705
transform 1 0 2694 0 1 471
box 0 0 1 1
use contact_26  contact_26_60
timestamp 1644951705
transform 1 0 2690 0 1 461
box 0 0 1 1
use contact_27  contact_27_61
timestamp 1644951705
transform 1 0 1916 0 1 391
box 0 0 1 1
use contact_26  contact_26_61
timestamp 1644951705
transform 1 0 1912 0 1 381
box 0 0 1 1
use contact_27  contact_27_62
timestamp 1644951705
transform 1 0 1138 0 1 311
box 0 0 1 1
use contact_26  contact_26_62
timestamp 1644951705
transform 1 0 1134 0 1 301
box 0 0 1 1
use contact_27  contact_27_63
timestamp 1644951705
transform 1 0 360 0 1 231
box 0 0 1 1
use contact_26  contact_26_63
timestamp 1644951705
transform 1 0 356 0 1 221
box 0 0 1 1
use column_mux_multiport  column_mux_multiport_0
timestamp 1644951705
transform 1 0 49014 0 1 560
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_1
timestamp 1644951705
transform 1 0 48236 0 1 560
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_2
timestamp 1644951705
transform 1 0 47458 0 1 560
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_3
timestamp 1644951705
transform 1 0 46680 0 1 560
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_4
timestamp 1644951705
transform 1 0 45902 0 1 560
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_5
timestamp 1644951705
transform 1 0 45124 0 1 560
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_6
timestamp 1644951705
transform 1 0 44346 0 1 560
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_7
timestamp 1644951705
transform 1 0 43568 0 1 560
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_8
timestamp 1644951705
transform 1 0 42790 0 1 560
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_9
timestamp 1644951705
transform 1 0 42012 0 1 560
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_10
timestamp 1644951705
transform 1 0 41234 0 1 560
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_11
timestamp 1644951705
transform 1 0 40456 0 1 560
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_12
timestamp 1644951705
transform 1 0 39678 0 1 560
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_13
timestamp 1644951705
transform 1 0 38900 0 1 560
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_14
timestamp 1644951705
transform 1 0 38122 0 1 560
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_15
timestamp 1644951705
transform 1 0 37344 0 1 560
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_16
timestamp 1644951705
transform 1 0 36566 0 1 560
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_17
timestamp 1644951705
transform 1 0 35788 0 1 560
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_18
timestamp 1644951705
transform 1 0 35010 0 1 560
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_19
timestamp 1644951705
transform 1 0 34232 0 1 560
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_20
timestamp 1644951705
transform 1 0 33454 0 1 560
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_21
timestamp 1644951705
transform 1 0 32676 0 1 560
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_22
timestamp 1644951705
transform 1 0 31898 0 1 560
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_23
timestamp 1644951705
transform 1 0 31120 0 1 560
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_24
timestamp 1644951705
transform 1 0 30342 0 1 560
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_25
timestamp 1644951705
transform 1 0 29564 0 1 560
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_26
timestamp 1644951705
transform 1 0 28786 0 1 560
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_27
timestamp 1644951705
transform 1 0 28008 0 1 560
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_28
timestamp 1644951705
transform 1 0 27230 0 1 560
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_29
timestamp 1644951705
transform 1 0 26452 0 1 560
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_30
timestamp 1644951705
transform 1 0 25674 0 1 560
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_31
timestamp 1644951705
transform 1 0 24896 0 1 560
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_32
timestamp 1644951705
transform 1 0 24118 0 1 560
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_33
timestamp 1644951705
transform 1 0 23340 0 1 560
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_34
timestamp 1644951705
transform 1 0 22562 0 1 560
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_35
timestamp 1644951705
transform 1 0 21784 0 1 560
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_36
timestamp 1644951705
transform 1 0 21006 0 1 560
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_37
timestamp 1644951705
transform 1 0 20228 0 1 560
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_38
timestamp 1644951705
transform 1 0 19450 0 1 560
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_39
timestamp 1644951705
transform 1 0 18672 0 1 560
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_40
timestamp 1644951705
transform 1 0 17894 0 1 560
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_41
timestamp 1644951705
transform 1 0 17116 0 1 560
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_42
timestamp 1644951705
transform 1 0 16338 0 1 560
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_43
timestamp 1644951705
transform 1 0 15560 0 1 560
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_44
timestamp 1644951705
transform 1 0 14782 0 1 560
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_45
timestamp 1644951705
transform 1 0 14004 0 1 560
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_46
timestamp 1644951705
transform 1 0 13226 0 1 560
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_47
timestamp 1644951705
transform 1 0 12448 0 1 560
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_48
timestamp 1644951705
transform 1 0 11670 0 1 560
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_49
timestamp 1644951705
transform 1 0 10892 0 1 560
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_50
timestamp 1644951705
transform 1 0 10114 0 1 560
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_51
timestamp 1644951705
transform 1 0 9336 0 1 560
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_52
timestamp 1644951705
transform 1 0 8558 0 1 560
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_53
timestamp 1644951705
transform 1 0 7780 0 1 560
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_54
timestamp 1644951705
transform 1 0 7002 0 1 560
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_55
timestamp 1644951705
transform 1 0 6224 0 1 560
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_56
timestamp 1644951705
transform 1 0 5446 0 1 560
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_57
timestamp 1644951705
transform 1 0 4668 0 1 560
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_58
timestamp 1644951705
transform 1 0 3890 0 1 560
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_59
timestamp 1644951705
transform 1 0 3112 0 1 560
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_60
timestamp 1644951705
transform 1 0 2334 0 1 560
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_61
timestamp 1644951705
transform 1 0 1556 0 1 560
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_62
timestamp 1644951705
transform 1 0 778 0 1 560
box 49 0 844 1508
use column_mux_multiport  column_mux_multiport_63
timestamp 1644951705
transform 1 0 0 0 1 560
box 49 0 844 1508
<< labels >>
rlabel metal1 s 0 240 49792 268 4 sel_0
rlabel metal1 s 0 320 49792 348 4 sel_1
rlabel metal1 s 0 400 49792 428 4 sel_2
rlabel metal1 s 0 480 49792 508 4 sel_3
rlabel metal2 s 84 160 112 560 4 rbl0_out_0
rlabel metal2 s 694 80 722 560 4 rbl1_out_0
rlabel metal2 s 3196 160 3224 560 4 rbl0_out_1
rlabel metal2 s 3806 80 3834 560 4 rbl1_out_1
rlabel metal2 s 6308 160 6336 560 4 rbl0_out_2
rlabel metal2 s 6918 80 6946 560 4 rbl1_out_2
rlabel metal2 s 9420 160 9448 560 4 rbl0_out_3
rlabel metal2 s 10030 80 10058 560 4 rbl1_out_3
rlabel metal2 s 12532 160 12560 560 4 rbl0_out_4
rlabel metal2 s 13142 80 13170 560 4 rbl1_out_4
rlabel metal2 s 15644 160 15672 560 4 rbl0_out_5
rlabel metal2 s 16254 80 16282 560 4 rbl1_out_5
rlabel metal2 s 18756 160 18784 560 4 rbl0_out_6
rlabel metal2 s 19366 80 19394 560 4 rbl1_out_6
rlabel metal2 s 21868 160 21896 560 4 rbl0_out_7
rlabel metal2 s 22478 80 22506 560 4 rbl1_out_7
rlabel metal2 s 24980 160 25008 560 4 rbl0_out_8
rlabel metal2 s 25590 80 25618 560 4 rbl1_out_8
rlabel metal2 s 28092 160 28120 560 4 rbl0_out_9
rlabel metal2 s 28702 80 28730 560 4 rbl1_out_9
rlabel metal2 s 31204 160 31232 560 4 rbl0_out_10
rlabel metal2 s 31814 80 31842 560 4 rbl1_out_10
rlabel metal2 s 34316 160 34344 560 4 rbl0_out_11
rlabel metal2 s 34926 80 34954 560 4 rbl1_out_11
rlabel metal2 s 37428 160 37456 560 4 rbl0_out_12
rlabel metal2 s 38038 80 38066 560 4 rbl1_out_12
rlabel metal2 s 40540 160 40568 560 4 rbl0_out_13
rlabel metal2 s 41150 80 41178 560 4 rbl1_out_13
rlabel metal2 s 43652 160 43680 560 4 rbl0_out_14
rlabel metal2 s 44262 80 44290 560 4 rbl1_out_14
rlabel metal2 s 46764 160 46792 560 4 rbl0_out_15
rlabel metal2 s 47374 80 47402 560 4 rbl1_out_15
rlabel metal2 s 84 2012 112 2068 4 rbl0_0
rlabel metal2 s 694 2012 722 2068 4 rbl1_0
rlabel metal2 s 862 2012 890 2068 4 rbl0_1
rlabel metal2 s 1472 2012 1500 2068 4 rbl1_1
rlabel metal2 s 1640 2012 1668 2068 4 rbl0_2
rlabel metal2 s 2250 2012 2278 2068 4 rbl1_2
rlabel metal2 s 2418 2012 2446 2068 4 rbl0_3
rlabel metal2 s 3028 2012 3056 2068 4 rbl1_3
rlabel metal2 s 3196 2012 3224 2068 4 rbl0_4
rlabel metal2 s 3806 2012 3834 2068 4 rbl1_4
rlabel metal2 s 3974 2012 4002 2068 4 rbl0_5
rlabel metal2 s 4584 2012 4612 2068 4 rbl1_5
rlabel metal2 s 4752 2012 4780 2068 4 rbl0_6
rlabel metal2 s 5362 2012 5390 2068 4 rbl1_6
rlabel metal2 s 5530 2012 5558 2068 4 rbl0_7
rlabel metal2 s 6140 2012 6168 2068 4 rbl1_7
rlabel metal2 s 6308 2012 6336 2068 4 rbl0_8
rlabel metal2 s 6918 2012 6946 2068 4 rbl1_8
rlabel metal2 s 7086 2012 7114 2068 4 rbl0_9
rlabel metal2 s 7696 2012 7724 2068 4 rbl1_9
rlabel metal2 s 7864 2012 7892 2068 4 rbl0_10
rlabel metal2 s 8474 2012 8502 2068 4 rbl1_10
rlabel metal2 s 8642 2012 8670 2068 4 rbl0_11
rlabel metal2 s 9252 2012 9280 2068 4 rbl1_11
rlabel metal2 s 9420 2012 9448 2068 4 rbl0_12
rlabel metal2 s 10030 2012 10058 2068 4 rbl1_12
rlabel metal2 s 10198 2012 10226 2068 4 rbl0_13
rlabel metal2 s 10808 2012 10836 2068 4 rbl1_13
rlabel metal2 s 10976 2012 11004 2068 4 rbl0_14
rlabel metal2 s 11586 2012 11614 2068 4 rbl1_14
rlabel metal2 s 11754 2012 11782 2068 4 rbl0_15
rlabel metal2 s 12364 2012 12392 2068 4 rbl1_15
rlabel metal2 s 12532 2012 12560 2068 4 rbl0_16
rlabel metal2 s 13142 2012 13170 2068 4 rbl1_16
rlabel metal2 s 13310 2012 13338 2068 4 rbl0_17
rlabel metal2 s 13920 2012 13948 2068 4 rbl1_17
rlabel metal2 s 14088 2012 14116 2068 4 rbl0_18
rlabel metal2 s 14698 2012 14726 2068 4 rbl1_18
rlabel metal2 s 14866 2012 14894 2068 4 rbl0_19
rlabel metal2 s 15476 2012 15504 2068 4 rbl1_19
rlabel metal2 s 15644 2012 15672 2068 4 rbl0_20
rlabel metal2 s 16254 2012 16282 2068 4 rbl1_20
rlabel metal2 s 16422 2012 16450 2068 4 rbl0_21
rlabel metal2 s 17032 2012 17060 2068 4 rbl1_21
rlabel metal2 s 17200 2012 17228 2068 4 rbl0_22
rlabel metal2 s 17810 2012 17838 2068 4 rbl1_22
rlabel metal2 s 17978 2012 18006 2068 4 rbl0_23
rlabel metal2 s 18588 2012 18616 2068 4 rbl1_23
rlabel metal2 s 18756 2012 18784 2068 4 rbl0_24
rlabel metal2 s 19366 2012 19394 2068 4 rbl1_24
rlabel metal2 s 19534 2012 19562 2068 4 rbl0_25
rlabel metal2 s 20144 2012 20172 2068 4 rbl1_25
rlabel metal2 s 20312 2012 20340 2068 4 rbl0_26
rlabel metal2 s 20922 2012 20950 2068 4 rbl1_26
rlabel metal2 s 21090 2012 21118 2068 4 rbl0_27
rlabel metal2 s 21700 2012 21728 2068 4 rbl1_27
rlabel metal2 s 21868 2012 21896 2068 4 rbl0_28
rlabel metal2 s 22478 2012 22506 2068 4 rbl1_28
rlabel metal2 s 22646 2012 22674 2068 4 rbl0_29
rlabel metal2 s 23256 2012 23284 2068 4 rbl1_29
rlabel metal2 s 23424 2012 23452 2068 4 rbl0_30
rlabel metal2 s 24034 2012 24062 2068 4 rbl1_30
rlabel metal2 s 24202 2012 24230 2068 4 rbl0_31
rlabel metal2 s 24812 2012 24840 2068 4 rbl1_31
rlabel metal2 s 24980 2012 25008 2068 4 rbl0_32
rlabel metal2 s 25590 2012 25618 2068 4 rbl1_32
rlabel metal2 s 25758 2012 25786 2068 4 rbl0_33
rlabel metal2 s 26368 2012 26396 2068 4 rbl1_33
rlabel metal2 s 26536 2012 26564 2068 4 rbl0_34
rlabel metal2 s 27146 2012 27174 2068 4 rbl1_34
rlabel metal2 s 27314 2012 27342 2068 4 rbl0_35
rlabel metal2 s 27924 2012 27952 2068 4 rbl1_35
rlabel metal2 s 28092 2012 28120 2068 4 rbl0_36
rlabel metal2 s 28702 2012 28730 2068 4 rbl1_36
rlabel metal2 s 28870 2012 28898 2068 4 rbl0_37
rlabel metal2 s 29480 2012 29508 2068 4 rbl1_37
rlabel metal2 s 29648 2012 29676 2068 4 rbl0_38
rlabel metal2 s 30258 2012 30286 2068 4 rbl1_38
rlabel metal2 s 30426 2012 30454 2068 4 rbl0_39
rlabel metal2 s 31036 2012 31064 2068 4 rbl1_39
rlabel metal2 s 31204 2012 31232 2068 4 rbl0_40
rlabel metal2 s 31814 2012 31842 2068 4 rbl1_40
rlabel metal2 s 31982 2012 32010 2068 4 rbl0_41
rlabel metal2 s 32592 2012 32620 2068 4 rbl1_41
rlabel metal2 s 32760 2012 32788 2068 4 rbl0_42
rlabel metal2 s 33370 2012 33398 2068 4 rbl1_42
rlabel metal2 s 33538 2012 33566 2068 4 rbl0_43
rlabel metal2 s 34148 2012 34176 2068 4 rbl1_43
rlabel metal2 s 34316 2012 34344 2068 4 rbl0_44
rlabel metal2 s 34926 2012 34954 2068 4 rbl1_44
rlabel metal2 s 35094 2012 35122 2068 4 rbl0_45
rlabel metal2 s 35704 2012 35732 2068 4 rbl1_45
rlabel metal2 s 35872 2012 35900 2068 4 rbl0_46
rlabel metal2 s 36482 2012 36510 2068 4 rbl1_46
rlabel metal2 s 36650 2012 36678 2068 4 rbl0_47
rlabel metal2 s 37260 2012 37288 2068 4 rbl1_47
rlabel metal2 s 37428 2012 37456 2068 4 rbl0_48
rlabel metal2 s 38038 2012 38066 2068 4 rbl1_48
rlabel metal2 s 38206 2012 38234 2068 4 rbl0_49
rlabel metal2 s 38816 2012 38844 2068 4 rbl1_49
rlabel metal2 s 38984 2012 39012 2068 4 rbl0_50
rlabel metal2 s 39594 2012 39622 2068 4 rbl1_50
rlabel metal2 s 39762 2012 39790 2068 4 rbl0_51
rlabel metal2 s 40372 2012 40400 2068 4 rbl1_51
rlabel metal2 s 40540 2012 40568 2068 4 rbl0_52
rlabel metal2 s 41150 2012 41178 2068 4 rbl1_52
rlabel metal2 s 41318 2012 41346 2068 4 rbl0_53
rlabel metal2 s 41928 2012 41956 2068 4 rbl1_53
rlabel metal2 s 42096 2012 42124 2068 4 rbl0_54
rlabel metal2 s 42706 2012 42734 2068 4 rbl1_54
rlabel metal2 s 42874 2012 42902 2068 4 rbl0_55
rlabel metal2 s 43484 2012 43512 2068 4 rbl1_55
rlabel metal2 s 43652 2012 43680 2068 4 rbl0_56
rlabel metal2 s 44262 2012 44290 2068 4 rbl1_56
rlabel metal2 s 44430 2012 44458 2068 4 rbl0_57
rlabel metal2 s 45040 2012 45068 2068 4 rbl1_57
rlabel metal2 s 45208 2012 45236 2068 4 rbl0_58
rlabel metal2 s 45818 2012 45846 2068 4 rbl1_58
rlabel metal2 s 45986 2012 46014 2068 4 rbl0_59
rlabel metal2 s 46596 2012 46624 2068 4 rbl1_59
rlabel metal2 s 46764 2012 46792 2068 4 rbl0_60
rlabel metal2 s 47374 2012 47402 2068 4 rbl1_60
rlabel metal2 s 47542 2012 47570 2068 4 rbl0_61
rlabel metal2 s 48152 2012 48180 2068 4 rbl1_61
rlabel metal2 s 48320 2012 48348 2068 4 rbl0_62
rlabel metal2 s 48930 2012 48958 2068 4 rbl1_62
rlabel metal2 s 49098 2012 49126 2068 4 rbl0_63
rlabel metal2 s 49708 2012 49736 2068 4 rbl1_63
rlabel metal3 s 24830 1282 24962 1356 4 gnd
rlabel metal3 s 29498 1282 29630 1356 4 gnd
rlabel metal3 s 31054 1282 31186 1356 4 gnd
rlabel metal3 s 19384 1282 19516 1356 4 gnd
rlabel metal3 s 33388 1282 33520 1356 4 gnd
rlabel metal3 s 34166 1282 34298 1356 4 gnd
rlabel metal3 s 38056 1282 38188 1356 4 gnd
rlabel metal3 s 49726 1282 49858 1356 4 gnd
rlabel metal3 s 35722 1282 35854 1356 4 gnd
rlabel metal3 s 43502 1282 43634 1356 4 gnd
rlabel metal3 s 13938 1282 14070 1356 4 gnd
rlabel metal3 s 12382 1282 12514 1356 4 gnd
rlabel metal3 s 40390 1282 40522 1356 4 gnd
rlabel metal3 s 26386 1282 26518 1356 4 gnd
rlabel metal3 s 21718 1282 21850 1356 4 gnd
rlabel metal3 s 41168 1282 41300 1356 4 gnd
rlabel metal3 s 3046 1282 3178 1356 4 gnd
rlabel metal3 s 22496 1282 22628 1356 4 gnd
rlabel metal3 s 3824 1282 3956 1356 4 gnd
rlabel metal3 s 11604 1282 11736 1356 4 gnd
rlabel metal3 s 31832 1282 31964 1356 4 gnd
rlabel metal3 s 4602 1282 4734 1356 4 gnd
rlabel metal3 s 42724 1282 42856 1356 4 gnd
rlabel metal3 s 38834 1282 38966 1356 4 gnd
rlabel metal3 s 13160 1282 13292 1356 4 gnd
rlabel metal3 s 16272 1282 16404 1356 4 gnd
rlabel metal3 s 18606 1282 18738 1356 4 gnd
rlabel metal3 s 10048 1282 10180 1356 4 gnd
rlabel metal3 s 32610 1282 32742 1356 4 gnd
rlabel metal3 s 27164 1282 27296 1356 4 gnd
rlabel metal3 s 27942 1282 28074 1356 4 gnd
rlabel metal3 s 41946 1282 42078 1356 4 gnd
rlabel metal3 s 17828 1282 17960 1356 4 gnd
rlabel metal3 s 45836 1282 45968 1356 4 gnd
rlabel metal3 s 25608 1282 25740 1356 4 gnd
rlabel metal3 s 47392 1282 47524 1356 4 gnd
rlabel metal3 s 48170 1282 48302 1356 4 gnd
rlabel metal3 s 20940 1282 21072 1356 4 gnd
rlabel metal3 s 9270 1282 9402 1356 4 gnd
rlabel metal3 s 30276 1282 30408 1356 4 gnd
rlabel metal3 s 1490 1282 1622 1356 4 gnd
rlabel metal3 s 6936 1282 7068 1356 4 gnd
rlabel metal3 s 24052 1282 24184 1356 4 gnd
rlabel metal3 s 36500 1282 36632 1356 4 gnd
rlabel metal3 s 6158 1282 6290 1356 4 gnd
rlabel metal3 s 39612 1282 39744 1356 4 gnd
rlabel metal3 s 28720 1282 28852 1356 4 gnd
rlabel metal3 s 8492 1282 8624 1356 4 gnd
rlabel metal3 s 15494 1282 15626 1356 4 gnd
rlabel metal3 s 23274 1282 23406 1356 4 gnd
rlabel metal3 s 48948 1282 49080 1356 4 gnd
rlabel metal3 s 7714 1282 7846 1356 4 gnd
rlabel metal3 s 37278 1282 37410 1356 4 gnd
rlabel metal3 s 5380 1282 5512 1356 4 gnd
rlabel metal3 s 2268 1282 2400 1356 4 gnd
rlabel metal3 s 712 1282 844 1356 4 gnd
rlabel metal3 s 17050 1282 17182 1356 4 gnd
rlabel metal3 s 20162 1282 20294 1356 4 gnd
rlabel metal3 s 34944 1282 35076 1356 4 gnd
rlabel metal3 s 44280 1282 44412 1356 4 gnd
rlabel metal3 s 45058 1282 45190 1356 4 gnd
rlabel metal3 s 46614 1282 46746 1356 4 gnd
rlabel metal3 s 14716 1282 14848 1356 4 gnd
rlabel metal3 s 10826 1282 10958 1356 4 gnd
<< properties >>
string FIXED_BBOX 0 0 49792 2068
string GDS_FILE sram_0rw2r1w_16_128_sky130A.gds
string GDS_END 1591982
string GDS_START 1523018
<< end >>
