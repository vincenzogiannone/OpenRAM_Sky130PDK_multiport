magic
tech sky130A
magscale 1 2
timestamp 1643671299
<< checkpaint >>
rect -1263 -1302 2742 8006
<< via1 >>
rect 715 6678 767 6730
rect 715 5840 767 5892
rect 715 5002 767 5054
rect 715 4164 767 4216
rect 715 3326 767 3378
rect 715 2488 767 2540
rect 715 1650 767 1702
rect 715 812 767 864
rect 715 -26 767 26
<< metal2 >>
rect 721 6732 761 6738
rect 0 328 28 6704
rect 721 6670 761 6676
rect 180 6444 234 6472
rect 1260 6448 1314 6476
rect 721 5894 761 5900
rect 721 5832 761 5838
rect 180 5260 234 5288
rect 1260 5256 1314 5284
rect 721 5056 761 5062
rect 721 4994 761 5000
rect 180 4768 234 4796
rect 1260 4772 1314 4800
rect 721 4218 761 4224
rect 721 4156 761 4162
rect 180 3584 234 3612
rect 1260 3580 1314 3608
rect 721 3380 761 3386
rect 721 3318 761 3324
rect 180 3092 234 3120
rect 1260 3096 1314 3124
rect 721 2542 761 2548
rect 721 2480 761 2486
rect 180 1908 234 1936
rect 1260 1904 1314 1932
rect 721 1704 761 1710
rect 721 1642 761 1648
rect 180 1416 234 1444
rect 1260 1420 1314 1448
rect 721 866 761 872
rect 721 804 761 810
rect 0 0 28 272
rect 180 232 234 260
rect 1260 228 1314 256
rect 721 28 761 34
rect 721 -34 761 -28
<< via2 >>
rect 713 6730 769 6732
rect 713 6678 715 6730
rect 715 6678 767 6730
rect 767 6678 769 6730
rect 713 6676 769 6678
rect 713 5892 769 5894
rect 713 5840 715 5892
rect 715 5840 767 5892
rect 767 5840 769 5892
rect 713 5838 769 5840
rect 713 5054 769 5056
rect 713 5002 715 5054
rect 715 5002 767 5054
rect 767 5002 769 5054
rect 713 5000 769 5002
rect 713 4216 769 4218
rect 713 4164 715 4216
rect 715 4164 767 4216
rect 767 4164 769 4216
rect 713 4162 769 4164
rect 713 3378 769 3380
rect 713 3326 715 3378
rect 715 3326 767 3378
rect 767 3326 769 3378
rect 713 3324 769 3326
rect 713 2540 769 2542
rect 713 2488 715 2540
rect 715 2488 767 2540
rect 767 2488 769 2540
rect 713 2486 769 2488
rect 713 1702 769 1704
rect 713 1650 715 1702
rect 715 1650 767 1702
rect 767 1650 769 1702
rect 713 1648 769 1650
rect 713 864 769 866
rect 713 812 715 864
rect 715 812 767 864
rect 767 812 769 864
rect 713 810 769 812
rect -1 272 55 328
rect 713 26 769 28
rect 713 -26 715 26
rect 715 -26 767 26
rect 767 -26 769 26
rect 713 -28 769 -26
<< metal3 >>
rect 711 6732 771 6734
rect 711 6676 713 6732
rect 769 6676 771 6732
rect 711 6674 771 6676
rect 711 5894 771 5896
rect 711 5838 713 5894
rect 769 5838 771 5894
rect 711 5836 771 5838
rect 711 5056 771 5058
rect 711 5000 713 5056
rect 769 5000 771 5056
rect 711 4998 771 5000
rect 711 4218 771 4220
rect 711 4162 713 4218
rect 769 4162 771 4218
rect 711 4160 771 4162
rect 711 3380 771 3382
rect 711 3324 713 3380
rect 769 3324 771 3380
rect 711 3322 771 3324
rect 711 2542 771 2544
rect 711 2486 713 2542
rect 769 2486 771 2542
rect 711 2484 771 2486
rect 711 1704 771 1706
rect 711 1648 713 1704
rect 769 1648 771 1704
rect 711 1646 771 1648
rect 711 866 771 868
rect 711 810 713 866
rect 769 810 771 866
rect 711 808 771 810
rect -3 328 1482 330
rect -3 272 -1 328
rect 55 272 1482 328
rect -3 270 1482 272
rect 711 28 771 30
rect 711 -28 713 28
rect 769 -28 771 28
rect 711 -30 771 -28
use contact_18  contact_18_0
timestamp 1643671299
transform 1 0 -3 0 1 270
box 0 0 1 1
use contact_18  contact_18_1
timestamp 1643671299
transform 1 0 711 0 1 6674
box 0 0 1 1
use contact_17  contact_17_0
timestamp 1643671299
transform 1 0 726 0 1 6689
box 0 0 1 1
use contact_18  contact_18_2
timestamp 1643671299
transform 1 0 711 0 1 5836
box 0 0 1 1
use contact_17  contact_17_1
timestamp 1643671299
transform 1 0 726 0 1 5851
box 0 0 1 1
use contact_18  contact_18_3
timestamp 1643671299
transform 1 0 711 0 1 4998
box 0 0 1 1
use contact_17  contact_17_2
timestamp 1643671299
transform 1 0 726 0 1 5013
box 0 0 1 1
use contact_18  contact_18_4
timestamp 1643671299
transform 1 0 711 0 1 5836
box 0 0 1 1
use contact_17  contact_17_3
timestamp 1643671299
transform 1 0 726 0 1 5851
box 0 0 1 1
use contact_18  contact_18_5
timestamp 1643671299
transform 1 0 711 0 1 4998
box 0 0 1 1
use contact_17  contact_17_4
timestamp 1643671299
transform 1 0 726 0 1 5013
box 0 0 1 1
use contact_18  contact_18_6
timestamp 1643671299
transform 1 0 711 0 1 4160
box 0 0 1 1
use contact_17  contact_17_5
timestamp 1643671299
transform 1 0 726 0 1 4175
box 0 0 1 1
use contact_18  contact_18_7
timestamp 1643671299
transform 1 0 711 0 1 3322
box 0 0 1 1
use contact_17  contact_17_6
timestamp 1643671299
transform 1 0 726 0 1 3337
box 0 0 1 1
use contact_18  contact_18_8
timestamp 1643671299
transform 1 0 711 0 1 4160
box 0 0 1 1
use contact_17  contact_17_7
timestamp 1643671299
transform 1 0 726 0 1 4175
box 0 0 1 1
use contact_18  contact_18_9
timestamp 1643671299
transform 1 0 711 0 1 3322
box 0 0 1 1
use contact_17  contact_17_8
timestamp 1643671299
transform 1 0 726 0 1 3337
box 0 0 1 1
use contact_18  contact_18_10
timestamp 1643671299
transform 1 0 711 0 1 2484
box 0 0 1 1
use contact_17  contact_17_9
timestamp 1643671299
transform 1 0 726 0 1 2499
box 0 0 1 1
use contact_18  contact_18_11
timestamp 1643671299
transform 1 0 711 0 1 1646
box 0 0 1 1
use contact_17  contact_17_10
timestamp 1643671299
transform 1 0 726 0 1 1661
box 0 0 1 1
use contact_18  contact_18_12
timestamp 1643671299
transform 1 0 711 0 1 2484
box 0 0 1 1
use contact_17  contact_17_11
timestamp 1643671299
transform 1 0 726 0 1 2499
box 0 0 1 1
use contact_18  contact_18_13
timestamp 1643671299
transform 1 0 711 0 1 1646
box 0 0 1 1
use contact_17  contact_17_12
timestamp 1643671299
transform 1 0 726 0 1 1661
box 0 0 1 1
use contact_18  contact_18_14
timestamp 1643671299
transform 1 0 711 0 1 808
box 0 0 1 1
use contact_17  contact_17_13
timestamp 1643671299
transform 1 0 726 0 1 823
box 0 0 1 1
use contact_18  contact_18_15
timestamp 1643671299
transform 1 0 711 0 1 -30
box 0 0 1 1
use contact_17  contact_17_14
timestamp 1643671299
transform 1 0 726 0 1 -15
box 0 0 1 1
use contact_18  contact_18_16
timestamp 1643671299
transform 1 0 711 0 1 808
box 0 0 1 1
use contact_17  contact_17_15
timestamp 1643671299
transform 1 0 726 0 1 823
box 0 0 1 1
use dff  dff_0
timestamp 1643671299
transform 1 0 0 0 -1 6704
box 0 -42 1482 916
use dff  dff_1
timestamp 1643671299
transform 1 0 0 0 1 5028
box 0 -42 1482 916
use dff  dff_2
timestamp 1643671299
transform 1 0 0 0 -1 5028
box 0 -42 1482 916
use dff  dff_3
timestamp 1643671299
transform 1 0 0 0 1 3352
box 0 -42 1482 916
use dff  dff_4
timestamp 1643671299
transform 1 0 0 0 -1 3352
box 0 -42 1482 916
use dff  dff_5
timestamp 1643671299
transform 1 0 0 0 1 1676
box 0 -42 1482 916
use dff  dff_6
timestamp 1643671299
transform 1 0 0 0 -1 1676
box 0 -42 1482 916
use dff  dff_7
timestamp 1643671299
transform 1 0 0 0 1 0
box 0 -42 1482 916
<< labels >>
rlabel metal3 s 711 808 771 868 4 vdd
rlabel metal3 s 711 2484 771 2544 4 vdd
rlabel metal3 s 741 2514 741 2514 4 vdd
rlabel metal3 s 711 4160 771 4220 4 vdd
rlabel metal3 s 711 5836 771 5896 4 vdd
rlabel metal3 s 741 5866 741 5866 4 vdd
rlabel metal3 s 741 838 741 838 4 vdd
rlabel metal3 s 711 4998 771 5058 4 gnd
rlabel metal3 s 711 -30 771 30 4 gnd
rlabel metal3 s 711 1646 771 1706 4 gnd
rlabel metal3 s 711 3322 771 3382 4 gnd
rlabel metal3 s 711 6674 771 6734 4 gnd
rlabel metal2 s 180 232 234 260 4 din_0
rlabel metal2 s 1260 228 1314 256 4 dout_0
rlabel metal2 s 180 1416 234 1444 4 din_1
rlabel metal2 s 1260 1420 1314 1448 4 dout_1
rlabel metal2 s 180 1908 234 1936 4 din_2
rlabel metal2 s 1260 1904 1314 1932 4 dout_2
rlabel metal2 s 180 3092 234 3120 4 din_3
rlabel metal2 s 1260 3096 1314 3124 4 dout_3
rlabel metal2 s 180 3584 234 3612 4 din_4
rlabel metal2 s 1260 3580 1314 3608 4 dout_4
rlabel metal2 s 180 4768 234 4796 4 din_5
rlabel metal2 s 1260 4772 1314 4800 4 dout_5
rlabel metal2 s 180 5260 234 5288 4 din_6
rlabel metal2 s 1260 5256 1314 5284 4 dout_6
rlabel metal2 s 180 6444 234 6472 4 din_7
rlabel metal2 s 1260 6448 1314 6476 4 dout_7
rlabel metal3 s 0 270 1482 330 4 clk
<< properties >>
string FIXED_BBOX 711 -30 771 0
string GDS_FILE sram_0rw2r1w_16_32_sky130A.gds
string GDS_END 1232036
string GDS_START 1223798
<< end >>
