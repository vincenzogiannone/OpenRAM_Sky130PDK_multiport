magic
tech sky130A
magscale 1 2
timestamp 1644951705
<< checkpaint >>
rect -1319 -1314 1469 1566
<< nwell >>
rect -54 210 204 306
rect -59 42 209 210
rect -54 -54 204 42
<< scpmos >>
rect 60 0 90 252
<< pdiff >>
rect 0 143 60 252
rect 0 109 8 143
rect 42 109 60 143
rect 0 0 60 109
rect 90 143 150 252
rect 90 109 108 143
rect 142 109 150 143
rect 90 0 150 109
<< pdiffc >>
rect 8 109 42 143
rect 108 109 142 143
<< poly >>
rect 60 252 90 278
rect 60 -26 90 0
<< locali >>
rect 8 143 42 159
rect 8 93 42 109
rect 108 143 142 159
rect 108 93 142 109
use contact_9  contact_9_0
timestamp 1644951705
transform 1 0 100 0 1 85
box 0 0 2 2
use contact_9  contact_9_1
timestamp 1644951705
transform 1 0 0 0 1 85
box 0 0 2 2
<< labels >>
rlabel mvvaractor s 75 126 75 126 4 G
rlabel locali s 25 126 25 126 4 S
rlabel locali s 125 126 125 126 4 D
<< properties >>
string FIXED_BBOX -54 -54 204 42
string GDS_FILE sram_0rw2r1w_16_128_sky130A.gds
string GDS_END 1785046
string GDS_START 1784218
<< end >>
