magic
tech sky130A
magscale 1 2
timestamp 1644951705
<< checkpaint >>
rect -1260 -1297 3650 4649
<< locali >>
rect 0 3335 419 3369
rect 453 3335 1531 3369
rect 1565 3335 2354 3369
rect 2165 2958 2199 2992
rect 0 2497 419 2531
rect 453 2497 1531 2531
rect 1565 2497 2354 2531
rect 2165 2036 2199 2070
rect 0 1659 419 1693
rect 453 1659 1531 1693
rect 1565 1659 2354 1693
rect 2165 1282 2199 1316
rect 0 821 419 855
rect 453 821 1531 855
rect 1565 821 2354 855
rect 2165 360 2199 394
rect 0 -17 419 17
rect 453 -17 1531 17
rect 1565 -17 2354 17
<< viali >>
rect 419 3335 453 3369
rect 1531 3335 1565 3369
rect 1720 3045 1754 3079
rect 1820 2921 1854 2955
rect 419 2497 453 2531
rect 1531 2497 1565 2531
rect 1820 2073 1854 2107
rect 1720 1949 1754 1983
rect 419 1659 453 1693
rect 1531 1659 1565 1693
rect 1720 1369 1754 1403
rect 560 1282 594 1316
rect 692 1282 726 1316
rect 1820 1245 1854 1279
rect 419 821 453 855
rect 1531 821 1565 855
rect 1820 397 1854 431
rect 560 360 594 394
rect 692 360 726 394
rect 1720 273 1754 307
rect 419 -17 453 17
rect 1531 -17 1565 17
<< metal1 >>
rect 404 3326 410 3378
rect 462 3326 468 3378
rect 1516 3326 1522 3378
rect 1574 3326 1580 3378
rect 106 3036 112 3088
rect 164 3076 170 3088
rect 1218 3076 1224 3088
rect 164 3048 1224 3076
rect 164 3036 170 3048
rect 1218 3036 1224 3048
rect 1276 3076 1282 3088
rect 1708 3079 1766 3085
rect 1708 3076 1720 3079
rect 1276 3048 1720 3076
rect 1276 3036 1282 3048
rect 1708 3045 1720 3048
rect 1754 3045 1766 3079
rect 1708 3039 1766 3045
rect 230 2912 236 2964
rect 288 2952 294 2964
rect 1342 2952 1348 2964
rect 288 2924 1348 2952
rect 288 2912 294 2924
rect 1342 2912 1348 2924
rect 1400 2952 1406 2964
rect 1808 2955 1866 2961
rect 1808 2952 1820 2955
rect 1400 2924 1820 2952
rect 1400 2912 1406 2924
rect 1808 2921 1820 2924
rect 1854 2921 1866 2955
rect 1808 2915 1866 2921
rect 404 2488 410 2540
rect 462 2488 468 2540
rect 1516 2488 1522 2540
rect 1574 2488 1580 2540
rect 1342 2064 1348 2116
rect 1400 2104 1406 2116
rect 1808 2107 1866 2113
rect 1808 2104 1820 2107
rect 1400 2076 1820 2104
rect 1400 2064 1406 2076
rect 1808 2073 1820 2076
rect 1854 2073 1866 2107
rect 1808 2067 1866 2073
rect 970 1940 976 1992
rect 1028 1980 1034 1992
rect 1708 1983 1766 1989
rect 1708 1980 1720 1983
rect 1028 1952 1720 1980
rect 1028 1940 1034 1952
rect 1708 1949 1720 1952
rect 1754 1949 1766 1983
rect 1708 1943 1766 1949
rect 404 1650 410 1702
rect 462 1650 468 1702
rect 1516 1650 1522 1702
rect 1574 1650 1580 1702
rect 1094 1610 1100 1622
rect 850 1582 1100 1610
rect 230 1273 236 1325
rect 288 1313 294 1325
rect 548 1316 606 1322
rect 548 1313 560 1316
rect 288 1285 560 1313
rect 288 1273 294 1285
rect 548 1282 560 1285
rect 594 1282 606 1316
rect 548 1276 606 1282
rect 680 1316 738 1322
rect 680 1282 692 1316
rect 726 1313 738 1316
rect 850 1313 878 1582
rect 1094 1570 1100 1582
rect 1152 1570 1158 1622
rect 1218 1360 1224 1412
rect 1276 1400 1282 1412
rect 1708 1403 1766 1409
rect 1708 1400 1720 1403
rect 1276 1372 1720 1400
rect 1276 1360 1282 1372
rect 1708 1369 1720 1372
rect 1754 1369 1766 1403
rect 1708 1363 1766 1369
rect 726 1285 878 1313
rect 726 1282 738 1285
rect 680 1276 738 1282
rect 1094 1236 1100 1288
rect 1152 1276 1158 1288
rect 1808 1279 1866 1285
rect 1808 1276 1820 1279
rect 1152 1248 1820 1276
rect 1152 1236 1158 1248
rect 1808 1245 1820 1248
rect 1854 1245 1866 1279
rect 1808 1239 1866 1245
rect 404 812 410 864
rect 462 812 468 864
rect 1516 812 1522 864
rect 1574 812 1580 864
rect 970 772 976 784
rect 850 744 976 772
rect 106 351 112 403
rect 164 391 170 403
rect 548 394 606 400
rect 548 391 560 394
rect 164 363 560 391
rect 164 351 170 363
rect 548 360 560 363
rect 594 360 606 394
rect 548 354 606 360
rect 680 394 738 400
rect 680 360 692 394
rect 726 391 738 394
rect 850 391 878 744
rect 970 732 976 744
rect 1028 732 1034 784
rect 726 363 878 391
rect 1094 388 1100 440
rect 1152 428 1158 440
rect 1808 431 1866 437
rect 1808 428 1820 431
rect 1152 400 1820 428
rect 1152 388 1158 400
rect 1808 397 1820 400
rect 1854 397 1866 431
rect 1808 391 1866 397
rect 726 360 738 363
rect 680 354 738 360
rect 970 264 976 316
rect 1028 304 1034 316
rect 1708 307 1766 313
rect 1708 304 1720 307
rect 1028 276 1720 304
rect 1028 264 1034 276
rect 1708 273 1720 276
rect 1754 273 1766 307
rect 1708 267 1766 273
rect 404 -26 410 26
rect 462 -26 468 26
rect 1516 -26 1522 26
rect 1574 -26 1580 26
<< via1 >>
rect 410 3369 462 3378
rect 410 3335 419 3369
rect 419 3335 453 3369
rect 453 3335 462 3369
rect 410 3326 462 3335
rect 1522 3369 1574 3378
rect 1522 3335 1531 3369
rect 1531 3335 1565 3369
rect 1565 3335 1574 3369
rect 1522 3326 1574 3335
rect 112 3036 164 3088
rect 1224 3036 1276 3088
rect 236 2912 288 2964
rect 1348 2912 1400 2964
rect 410 2531 462 2540
rect 410 2497 419 2531
rect 419 2497 453 2531
rect 453 2497 462 2531
rect 410 2488 462 2497
rect 1522 2531 1574 2540
rect 1522 2497 1531 2531
rect 1531 2497 1565 2531
rect 1565 2497 1574 2531
rect 1522 2488 1574 2497
rect 1348 2064 1400 2116
rect 976 1940 1028 1992
rect 410 1693 462 1702
rect 410 1659 419 1693
rect 419 1659 453 1693
rect 453 1659 462 1693
rect 410 1650 462 1659
rect 1522 1693 1574 1702
rect 1522 1659 1531 1693
rect 1531 1659 1565 1693
rect 1565 1659 1574 1693
rect 1522 1650 1574 1659
rect 236 1273 288 1325
rect 1100 1570 1152 1622
rect 1224 1360 1276 1412
rect 1100 1236 1152 1288
rect 410 855 462 864
rect 410 821 419 855
rect 419 821 453 855
rect 453 821 462 855
rect 410 812 462 821
rect 1522 855 1574 864
rect 1522 821 1531 855
rect 1531 821 1565 855
rect 1565 821 1574 855
rect 1522 812 1574 821
rect 112 351 164 403
rect 976 732 1028 784
rect 1100 388 1152 440
rect 976 264 1028 316
rect 410 17 462 26
rect 410 -17 419 17
rect 419 -17 453 17
rect 453 -17 462 17
rect 410 -26 462 -17
rect 1522 17 1574 26
rect 1522 -17 1531 17
rect 1531 -17 1565 17
rect 1565 -17 1574 17
rect 1522 -26 1574 -17
<< metal2 >>
rect 408 3380 464 3389
rect 124 3094 152 3352
rect 112 3088 164 3094
rect 112 3030 164 3036
rect 124 409 152 3030
rect 248 2970 276 3352
rect 1520 3380 1576 3389
rect 408 3315 464 3324
rect 236 2964 288 2970
rect 236 2906 288 2912
rect 248 1331 276 2906
rect 408 2542 464 2551
rect 408 2477 464 2486
rect 988 1998 1016 3352
rect 976 1992 1028 1998
rect 976 1934 1028 1940
rect 408 1704 464 1713
rect 408 1639 464 1648
rect 236 1325 288 1331
rect 236 1267 288 1273
rect 112 403 164 409
rect 112 345 164 351
rect 124 124 152 345
rect 248 124 276 1267
rect 408 866 464 875
rect 408 801 464 810
rect 988 790 1016 1934
rect 1112 1628 1140 3352
rect 1236 3094 1264 3352
rect 1224 3088 1276 3094
rect 1224 3030 1276 3036
rect 1100 1622 1152 1628
rect 1100 1564 1152 1570
rect 1112 1294 1140 1564
rect 1236 1418 1264 3030
rect 1360 2970 1388 3352
rect 1520 3315 1576 3324
rect 1348 2964 1400 2970
rect 1348 2906 1400 2912
rect 1360 2122 1388 2906
rect 1520 2542 1576 2551
rect 1520 2477 1576 2486
rect 1348 2116 1400 2122
rect 1348 2058 1400 2064
rect 1224 1412 1276 1418
rect 1224 1354 1276 1360
rect 1100 1288 1152 1294
rect 1100 1230 1152 1236
rect 976 784 1028 790
rect 976 726 1028 732
rect 988 322 1016 726
rect 1112 446 1140 1230
rect 1100 440 1152 446
rect 1100 382 1152 388
rect 976 316 1028 322
rect 976 258 1028 264
rect 988 124 1016 258
rect 1112 124 1140 382
rect 1236 124 1264 1354
rect 1360 124 1388 2058
rect 1520 1704 1576 1713
rect 1520 1639 1576 1648
rect 1520 866 1576 875
rect 1520 801 1576 810
rect 408 28 464 37
rect 408 -37 464 -28
rect 1520 28 1576 37
rect 1520 -37 1576 -28
<< via2 >>
rect 408 3378 464 3380
rect 408 3326 410 3378
rect 410 3326 462 3378
rect 462 3326 464 3378
rect 1520 3378 1576 3380
rect 408 3324 464 3326
rect 408 2540 464 2542
rect 408 2488 410 2540
rect 410 2488 462 2540
rect 462 2488 464 2540
rect 408 2486 464 2488
rect 408 1702 464 1704
rect 408 1650 410 1702
rect 410 1650 462 1702
rect 462 1650 464 1702
rect 408 1648 464 1650
rect 408 864 464 866
rect 408 812 410 864
rect 410 812 462 864
rect 462 812 464 864
rect 408 810 464 812
rect 1520 3326 1522 3378
rect 1522 3326 1574 3378
rect 1574 3326 1576 3378
rect 1520 3324 1576 3326
rect 1520 2540 1576 2542
rect 1520 2488 1522 2540
rect 1522 2488 1574 2540
rect 1574 2488 1576 2540
rect 1520 2486 1576 2488
rect 1520 1702 1576 1704
rect 1520 1650 1522 1702
rect 1522 1650 1574 1702
rect 1574 1650 1576 1702
rect 1520 1648 1576 1650
rect 1520 864 1576 866
rect 1520 812 1522 864
rect 1522 812 1574 864
rect 1574 812 1576 864
rect 1520 810 1576 812
rect 408 26 464 28
rect 408 -26 410 26
rect 410 -26 462 26
rect 462 -26 464 26
rect 408 -28 464 -26
rect 1520 26 1576 28
rect 1520 -26 1522 26
rect 1522 -26 1574 26
rect 1574 -26 1576 26
rect 1520 -28 1576 -26
<< metal3 >>
rect 370 3380 502 3389
rect 370 3324 408 3380
rect 464 3324 502 3380
rect 370 3315 502 3324
rect 1482 3380 1614 3389
rect 1482 3324 1520 3380
rect 1576 3324 1614 3380
rect 1482 3315 1614 3324
rect 370 2542 502 2551
rect 370 2486 408 2542
rect 464 2486 502 2542
rect 370 2477 502 2486
rect 1482 2542 1614 2551
rect 1482 2486 1520 2542
rect 1576 2486 1614 2542
rect 1482 2477 1614 2486
rect 370 1704 502 1713
rect 370 1648 408 1704
rect 464 1648 502 1704
rect 370 1639 502 1648
rect 1482 1704 1614 1713
rect 1482 1648 1520 1704
rect 1576 1648 1614 1704
rect 1482 1639 1614 1648
rect 370 866 502 875
rect 370 810 408 866
rect 464 810 502 866
rect 370 801 502 810
rect 1482 866 1614 875
rect 1482 810 1520 866
rect 1576 810 1614 866
rect 1482 801 1614 810
rect 370 28 502 37
rect 370 -28 408 28
rect 464 -28 502 28
rect 370 -37 502 -28
rect 1482 28 1614 37
rect 1482 -28 1520 28
rect 1576 -28 1614 28
rect 1482 -37 1614 -28
use contact_18  contact_18_0
timestamp 1644951705
transform 1 0 1482 0 1 3315
box 0 0 1 1
use contact_17  contact_17_0
timestamp 1644951705
transform 1 0 1516 0 1 3320
box 0 0 1 1
use contact_13  contact_13_0
timestamp 1644951705
transform 1 0 1519 0 1 3329
box 0 0 1 1
use contact_18  contact_18_1
timestamp 1644951705
transform 1 0 370 0 1 3315
box 0 0 1 1
use contact_17  contact_17_1
timestamp 1644951705
transform 1 0 404 0 1 3320
box 0 0 1 1
use contact_13  contact_13_1
timestamp 1644951705
transform 1 0 407 0 1 3329
box 0 0 1 1
use contact_18  contact_18_2
timestamp 1644951705
transform 1 0 1482 0 1 2477
box 0 0 1 1
use contact_17  contact_17_2
timestamp 1644951705
transform 1 0 1516 0 1 2482
box 0 0 1 1
use contact_13  contact_13_2
timestamp 1644951705
transform 1 0 1519 0 1 2491
box 0 0 1 1
use contact_18  contact_18_3
timestamp 1644951705
transform 1 0 370 0 1 2477
box 0 0 1 1
use contact_17  contact_17_3
timestamp 1644951705
transform 1 0 404 0 1 2482
box 0 0 1 1
use contact_13  contact_13_3
timestamp 1644951705
transform 1 0 407 0 1 2491
box 0 0 1 1
use contact_18  contact_18_4
timestamp 1644951705
transform 1 0 1482 0 1 1639
box 0 0 1 1
use contact_17  contact_17_4
timestamp 1644951705
transform 1 0 1516 0 1 1644
box 0 0 1 1
use contact_13  contact_13_4
timestamp 1644951705
transform 1 0 1519 0 1 1653
box 0 0 1 1
use contact_18  contact_18_5
timestamp 1644951705
transform 1 0 370 0 1 1639
box 0 0 1 1
use contact_17  contact_17_5
timestamp 1644951705
transform 1 0 404 0 1 1644
box 0 0 1 1
use contact_13  contact_13_5
timestamp 1644951705
transform 1 0 407 0 1 1653
box 0 0 1 1
use contact_18  contact_18_6
timestamp 1644951705
transform 1 0 1482 0 1 2477
box 0 0 1 1
use contact_17  contact_17_6
timestamp 1644951705
transform 1 0 1516 0 1 2482
box 0 0 1 1
use contact_13  contact_13_6
timestamp 1644951705
transform 1 0 1519 0 1 2491
box 0 0 1 1
use contact_18  contact_18_7
timestamp 1644951705
transform 1 0 370 0 1 2477
box 0 0 1 1
use contact_17  contact_17_7
timestamp 1644951705
transform 1 0 404 0 1 2482
box 0 0 1 1
use contact_13  contact_13_7
timestamp 1644951705
transform 1 0 407 0 1 2491
box 0 0 1 1
use contact_18  contact_18_8
timestamp 1644951705
transform 1 0 1482 0 1 1639
box 0 0 1 1
use contact_17  contact_17_8
timestamp 1644951705
transform 1 0 1516 0 1 1644
box 0 0 1 1
use contact_13  contact_13_8
timestamp 1644951705
transform 1 0 1519 0 1 1653
box 0 0 1 1
use contact_18  contact_18_9
timestamp 1644951705
transform 1 0 370 0 1 1639
box 0 0 1 1
use contact_17  contact_17_9
timestamp 1644951705
transform 1 0 404 0 1 1644
box 0 0 1 1
use contact_13  contact_13_9
timestamp 1644951705
transform 1 0 407 0 1 1653
box 0 0 1 1
use contact_18  contact_18_10
timestamp 1644951705
transform 1 0 1482 0 1 801
box 0 0 1 1
use contact_17  contact_17_10
timestamp 1644951705
transform 1 0 1516 0 1 806
box 0 0 1 1
use contact_13  contact_13_10
timestamp 1644951705
transform 1 0 1519 0 1 815
box 0 0 1 1
use contact_18  contact_18_11
timestamp 1644951705
transform 1 0 370 0 1 801
box 0 0 1 1
use contact_17  contact_17_11
timestamp 1644951705
transform 1 0 404 0 1 806
box 0 0 1 1
use contact_13  contact_13_11
timestamp 1644951705
transform 1 0 407 0 1 815
box 0 0 1 1
use contact_18  contact_18_12
timestamp 1644951705
transform 1 0 1482 0 1 -37
box 0 0 1 1
use contact_17  contact_17_12
timestamp 1644951705
transform 1 0 1516 0 1 -32
box 0 0 1 1
use contact_13  contact_13_12
timestamp 1644951705
transform 1 0 1519 0 1 -23
box 0 0 1 1
use contact_18  contact_18_13
timestamp 1644951705
transform 1 0 370 0 1 -37
box 0 0 1 1
use contact_17  contact_17_13
timestamp 1644951705
transform 1 0 404 0 1 -32
box 0 0 1 1
use contact_13  contact_13_13
timestamp 1644951705
transform 1 0 407 0 1 -23
box 0 0 1 1
use contact_18  contact_18_14
timestamp 1644951705
transform 1 0 1482 0 1 801
box 0 0 1 1
use contact_17  contact_17_14
timestamp 1644951705
transform 1 0 1516 0 1 806
box 0 0 1 1
use contact_13  contact_13_14
timestamp 1644951705
transform 1 0 1519 0 1 815
box 0 0 1 1
use contact_18  contact_18_15
timestamp 1644951705
transform 1 0 370 0 1 801
box 0 0 1 1
use contact_17  contact_17_15
timestamp 1644951705
transform 1 0 404 0 1 806
box 0 0 1 1
use contact_13  contact_13_15
timestamp 1644951705
transform 1 0 407 0 1 815
box 0 0 1 1
use contact_17  contact_17_16
timestamp 1644951705
transform 1 0 1342 0 1 2906
box 0 0 1 1
use contact_17  contact_17_17
timestamp 1644951705
transform 1 0 230 0 1 2906
box 0 0 1 1
use contact_17  contact_17_18
timestamp 1644951705
transform 1 0 1218 0 1 3030
box 0 0 1 1
use contact_17  contact_17_19
timestamp 1644951705
transform 1 0 106 0 1 3030
box 0 0 1 1
use contact_14  contact_14_0
timestamp 1644951705
transform 1 0 1094 0 1 1564
box 0 0 1 1
use contact_13  contact_13_16
timestamp 1644951705
transform 1 0 680 0 1 1276
box 0 0 1 1
use contact_14  contact_14_1
timestamp 1644951705
transform 1 0 970 0 1 726
box 0 0 1 1
use contact_13  contact_13_17
timestamp 1644951705
transform 1 0 680 0 1 354
box 0 0 1 1
use contact_15  contact_15_0
timestamp 1644951705
transform 1 0 1808 0 1 2915
box 0 0 1 1
use contact_14  contact_14_2
timestamp 1644951705
transform 1 0 1342 0 1 2906
box 0 0 1 1
use contact_13  contact_13_18
timestamp 1644951705
transform 1 0 1708 0 1 3039
box 0 0 1 1
use contact_14  contact_14_3
timestamp 1644951705
transform 1 0 1218 0 1 3030
box 0 0 1 1
use contact_15  contact_15_1
timestamp 1644951705
transform 1 0 1808 0 1 2067
box 0 0 1 1
use contact_14  contact_14_4
timestamp 1644951705
transform 1 0 1342 0 1 2058
box 0 0 1 1
use contact_13  contact_13_19
timestamp 1644951705
transform 1 0 1708 0 1 1943
box 0 0 1 1
use contact_14  contact_14_5
timestamp 1644951705
transform 1 0 970 0 1 1934
box 0 0 1 1
use contact_15  contact_15_2
timestamp 1644951705
transform 1 0 1808 0 1 1239
box 0 0 1 1
use contact_14  contact_14_6
timestamp 1644951705
transform 1 0 1094 0 1 1230
box 0 0 1 1
use contact_13  contact_13_20
timestamp 1644951705
transform 1 0 1708 0 1 1363
box 0 0 1 1
use contact_14  contact_14_7
timestamp 1644951705
transform 1 0 1218 0 1 1354
box 0 0 1 1
use contact_15  contact_15_3
timestamp 1644951705
transform 1 0 1808 0 1 391
box 0 0 1 1
use contact_14  contact_14_8
timestamp 1644951705
transform 1 0 1094 0 1 382
box 0 0 1 1
use contact_13  contact_13_21
timestamp 1644951705
transform 1 0 1708 0 1 267
box 0 0 1 1
use contact_14  contact_14_9
timestamp 1644951705
transform 1 0 970 0 1 258
box 0 0 1 1
use contact_14  contact_14_10
timestamp 1644951705
transform 1 0 230 0 1 1267
box 0 0 1 1
use contact_13  contact_13_22
timestamp 1644951705
transform 1 0 548 0 1 1276
box 0 0 1 1
use contact_14  contact_14_11
timestamp 1644951705
transform 1 0 106 0 1 345
box 0 0 1 1
use contact_13  contact_13_23
timestamp 1644951705
transform 1 0 548 0 1 354
box 0 0 1 1
use pand2  pand2_0
timestamp 1644951705
transform 1 0 1608 0 -1 3352
box -36 -17 782 895
use pand2  pand2_1
timestamp 1644951705
transform 1 0 1608 0 1 1676
box -36 -17 782 895
use pand2  pand2_2
timestamp 1644951705
transform 1 0 1608 0 -1 1676
box -36 -17 782 895
use pand2  pand2_3
timestamp 1644951705
transform 1 0 1608 0 1 0
box -36 -17 782 895
use pinv_1  pinv_1_0
timestamp 1644951705
transform 1 0 496 0 -1 1676
box -36 -17 404 895
use pinv_1  pinv_1_1
timestamp 1644951705
transform 1 0 496 0 1 0
box -36 -17 404 895
<< labels >>
rlabel metal2 s 112 345 164 409 4 in_0
rlabel metal2 s 236 1267 288 1331 4 in_1
rlabel locali s 2182 377 2182 377 4 out_0
rlabel locali s 2182 1299 2182 1299 4 out_1
rlabel locali s 2182 2053 2182 2053 4 out_2
rlabel locali s 2182 2975 2182 2975 4 out_3
rlabel metal3 s 1482 2477 1614 2551 4 vdd
rlabel metal3 s 1482 801 1614 875 4 vdd
rlabel metal3 s 370 2477 502 2551 4 vdd
rlabel metal3 s 370 801 502 875 4 vdd
rlabel metal3 s 1482 1639 1614 1713 4 gnd
rlabel metal3 s 1482 -37 1614 37 4 gnd
rlabel metal3 s 370 -37 502 37 4 gnd
rlabel metal3 s 370 1639 502 1713 4 gnd
rlabel metal3 s 370 3315 502 3389 4 gnd
rlabel metal3 s 1482 3315 1614 3389 4 gnd
<< properties >>
string FIXED_BBOX 1482 -37 1614 0
string GDS_FILE sram_0rw2r1w_16_128_sky130A.gds
string GDS_END 1928824
string GDS_START 1918356
<< end >>
