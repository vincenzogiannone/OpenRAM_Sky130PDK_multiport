magic
tech sky130A
magscale 1 2
timestamp 1644969367
<< checkpaint >>
rect -1260 -1297 3340 7457
<< locali >>
rect 0 6143 291 6177
rect 325 6143 1163 6177
rect 1197 6143 2044 6177
rect 1855 5415 1889 5449
rect 0 4603 291 4637
rect 325 4603 1163 4637
rect 1197 4603 2044 4637
rect 1855 3791 1889 3825
rect 0 3063 291 3097
rect 325 3063 1163 3097
rect 1197 3063 2044 3097
rect 1855 2335 1889 2369
rect 0 1523 291 1557
rect 325 1523 1163 1557
rect 1197 1523 2044 1557
rect 1855 711 1889 745
rect 0 -17 291 17
rect 325 -17 1163 17
rect 1197 -17 2044 17
<< viali >>
rect 291 6143 325 6177
rect 1163 6143 1197 6177
rect 1320 5853 1354 5887
rect 1420 5729 1454 5763
rect 291 4603 325 4637
rect 1163 4603 1197 4637
rect 1420 3477 1454 3511
rect 1320 3353 1354 3387
rect 291 3063 325 3097
rect 1163 3063 1197 3097
rect 1320 2773 1354 2807
rect 1420 2649 1454 2683
rect 400 2335 434 2369
rect 532 2335 566 2369
rect 291 1523 325 1557
rect 1163 1523 1197 1557
rect 400 711 434 745
rect 532 711 566 745
rect 1420 397 1454 431
rect 1320 273 1354 307
rect 291 -17 325 17
rect 1163 -17 1197 17
<< metal1 >>
rect 276 6134 282 6186
rect 334 6134 340 6186
rect 1148 6134 1154 6186
rect 1206 6134 1212 6186
rect 66 5844 72 5896
rect 124 5884 130 5896
rect 938 5884 944 5896
rect 124 5856 944 5884
rect 124 5844 130 5856
rect 938 5844 944 5856
rect 996 5884 1002 5896
rect 1308 5887 1366 5893
rect 1308 5884 1320 5887
rect 996 5856 1320 5884
rect 996 5844 1002 5856
rect 1308 5853 1320 5856
rect 1354 5853 1366 5887
rect 1308 5847 1366 5853
rect 150 5720 156 5772
rect 208 5760 214 5772
rect 1022 5760 1028 5772
rect 208 5732 1028 5760
rect 208 5720 214 5732
rect 1022 5720 1028 5732
rect 1080 5760 1086 5772
rect 1408 5763 1466 5769
rect 1408 5760 1420 5763
rect 1080 5732 1420 5760
rect 1080 5720 1086 5732
rect 1408 5729 1420 5732
rect 1454 5729 1466 5763
rect 1408 5723 1466 5729
rect 276 4594 282 4646
rect 334 4594 340 4646
rect 1148 4594 1154 4646
rect 1206 4594 1212 4646
rect 1022 3468 1028 3520
rect 1080 3508 1086 3520
rect 1408 3511 1466 3517
rect 1408 3508 1420 3511
rect 1080 3480 1420 3508
rect 1080 3468 1086 3480
rect 1408 3477 1420 3480
rect 1454 3477 1466 3511
rect 1408 3471 1466 3477
rect 770 3344 776 3396
rect 828 3384 834 3396
rect 1308 3387 1366 3393
rect 1308 3384 1320 3387
rect 828 3356 1320 3384
rect 828 3344 834 3356
rect 1308 3353 1320 3356
rect 1354 3353 1366 3387
rect 1308 3347 1366 3353
rect 276 3054 282 3106
rect 334 3054 340 3106
rect 1148 3054 1154 3106
rect 1206 3054 1212 3106
rect 854 3014 860 3026
rect 690 2986 860 3014
rect 150 2326 156 2378
rect 208 2366 214 2378
rect 388 2369 446 2375
rect 388 2366 400 2369
rect 208 2338 400 2366
rect 208 2326 214 2338
rect 388 2335 400 2338
rect 434 2335 446 2369
rect 388 2329 446 2335
rect 520 2369 578 2375
rect 520 2335 532 2369
rect 566 2366 578 2369
rect 690 2366 718 2986
rect 854 2974 860 2986
rect 912 2974 918 3026
rect 938 2764 944 2816
rect 996 2804 1002 2816
rect 1308 2807 1366 2813
rect 1308 2804 1320 2807
rect 996 2776 1320 2804
rect 996 2764 1002 2776
rect 1308 2773 1320 2776
rect 1354 2773 1366 2807
rect 1308 2767 1366 2773
rect 854 2640 860 2692
rect 912 2680 918 2692
rect 1408 2683 1466 2689
rect 1408 2680 1420 2683
rect 912 2652 1420 2680
rect 912 2640 918 2652
rect 1408 2649 1420 2652
rect 1454 2649 1466 2683
rect 1408 2643 1466 2649
rect 566 2338 718 2366
rect 566 2335 578 2338
rect 520 2329 578 2335
rect 276 1514 282 1566
rect 334 1514 340 1566
rect 1148 1514 1154 1566
rect 1206 1514 1212 1566
rect 770 1474 776 1486
rect 690 1446 776 1474
rect 66 702 72 754
rect 124 742 130 754
rect 388 745 446 751
rect 388 742 400 745
rect 124 714 400 742
rect 124 702 130 714
rect 388 711 400 714
rect 434 711 446 745
rect 388 705 446 711
rect 520 745 578 751
rect 520 711 532 745
rect 566 742 578 745
rect 690 742 718 1446
rect 770 1434 776 1446
rect 828 1434 834 1486
rect 566 714 718 742
rect 566 711 578 714
rect 520 705 578 711
rect 854 388 860 440
rect 912 428 918 440
rect 1408 431 1466 437
rect 1408 428 1420 431
rect 912 400 1420 428
rect 912 388 918 400
rect 1408 397 1420 400
rect 1454 397 1466 431
rect 1408 391 1466 397
rect 770 264 776 316
rect 828 304 834 316
rect 1308 307 1366 313
rect 1308 304 1320 307
rect 828 276 1320 304
rect 828 264 834 276
rect 1308 273 1320 276
rect 1354 273 1366 307
rect 1308 267 1366 273
rect 276 -26 282 26
rect 334 -26 340 26
rect 1148 -26 1154 26
rect 1206 -26 1212 26
<< via1 >>
rect 282 6177 334 6186
rect 282 6143 291 6177
rect 291 6143 325 6177
rect 325 6143 334 6177
rect 282 6134 334 6143
rect 1154 6177 1206 6186
rect 1154 6143 1163 6177
rect 1163 6143 1197 6177
rect 1197 6143 1206 6177
rect 1154 6134 1206 6143
rect 72 5844 124 5896
rect 944 5844 996 5896
rect 156 5720 208 5772
rect 1028 5720 1080 5772
rect 282 4637 334 4646
rect 282 4603 291 4637
rect 291 4603 325 4637
rect 325 4603 334 4637
rect 282 4594 334 4603
rect 1154 4637 1206 4646
rect 1154 4603 1163 4637
rect 1163 4603 1197 4637
rect 1197 4603 1206 4637
rect 1154 4594 1206 4603
rect 1028 3468 1080 3520
rect 776 3344 828 3396
rect 282 3097 334 3106
rect 282 3063 291 3097
rect 291 3063 325 3097
rect 325 3063 334 3097
rect 282 3054 334 3063
rect 1154 3097 1206 3106
rect 1154 3063 1163 3097
rect 1163 3063 1197 3097
rect 1197 3063 1206 3097
rect 1154 3054 1206 3063
rect 156 2326 208 2378
rect 860 2974 912 3026
rect 944 2764 996 2816
rect 860 2640 912 2692
rect 282 1557 334 1566
rect 282 1523 291 1557
rect 291 1523 325 1557
rect 325 1523 334 1557
rect 282 1514 334 1523
rect 1154 1557 1206 1566
rect 1154 1523 1163 1557
rect 1163 1523 1197 1557
rect 1197 1523 1206 1557
rect 1154 1514 1206 1523
rect 72 702 124 754
rect 776 1434 828 1486
rect 860 388 912 440
rect 776 264 828 316
rect 282 17 334 26
rect 282 -17 291 17
rect 291 -17 325 17
rect 325 -17 334 17
rect 282 -26 334 -17
rect 1154 17 1206 26
rect 1154 -17 1163 17
rect 1163 -17 1197 17
rect 1197 -17 1206 17
rect 1154 -26 1206 -17
<< metal2 >>
rect 280 6188 336 6197
rect 84 5902 112 6160
rect 72 5896 124 5902
rect 72 5838 124 5844
rect 84 760 112 5838
rect 168 5778 196 6160
rect 1152 6188 1208 6197
rect 280 6123 336 6132
rect 156 5772 208 5778
rect 156 5714 208 5720
rect 168 2384 196 5714
rect 280 4648 336 4657
rect 280 4583 336 4592
rect 788 3402 816 6160
rect 776 3396 828 3402
rect 776 3338 828 3344
rect 280 3108 336 3117
rect 280 3043 336 3052
rect 156 2378 208 2384
rect 156 2320 208 2326
rect 72 754 124 760
rect 72 696 124 702
rect 84 84 112 696
rect 168 84 196 2320
rect 280 1568 336 1577
rect 280 1503 336 1512
rect 788 1492 816 3338
rect 872 3032 900 6160
rect 956 5902 984 6160
rect 944 5896 996 5902
rect 944 5838 996 5844
rect 860 3026 912 3032
rect 860 2968 912 2974
rect 872 2698 900 2968
rect 956 2822 984 5838
rect 1040 5778 1068 6160
rect 1152 6123 1208 6132
rect 1028 5772 1080 5778
rect 1028 5714 1080 5720
rect 1040 3526 1068 5714
rect 1152 4648 1208 4657
rect 1152 4583 1208 4592
rect 1028 3520 1080 3526
rect 1028 3462 1080 3468
rect 944 2816 996 2822
rect 944 2758 996 2764
rect 860 2692 912 2698
rect 860 2634 912 2640
rect 776 1486 828 1492
rect 776 1428 828 1434
rect 788 322 816 1428
rect 872 446 900 2634
rect 860 440 912 446
rect 860 382 912 388
rect 776 316 828 322
rect 776 258 828 264
rect 788 84 816 258
rect 872 84 900 382
rect 956 84 984 2758
rect 1040 84 1068 3462
rect 1152 3108 1208 3117
rect 1152 3043 1208 3052
rect 1152 1568 1208 1577
rect 1152 1503 1208 1512
rect 280 28 336 37
rect 280 -37 336 -28
rect 1152 28 1208 37
rect 1152 -37 1208 -28
<< via2 >>
rect 280 6186 336 6188
rect 280 6134 282 6186
rect 282 6134 334 6186
rect 334 6134 336 6186
rect 1152 6186 1208 6188
rect 280 6132 336 6134
rect 280 4646 336 4648
rect 280 4594 282 4646
rect 282 4594 334 4646
rect 334 4594 336 4646
rect 280 4592 336 4594
rect 280 3106 336 3108
rect 280 3054 282 3106
rect 282 3054 334 3106
rect 334 3054 336 3106
rect 280 3052 336 3054
rect 280 1566 336 1568
rect 280 1514 282 1566
rect 282 1514 334 1566
rect 334 1514 336 1566
rect 280 1512 336 1514
rect 1152 6134 1154 6186
rect 1154 6134 1206 6186
rect 1206 6134 1208 6186
rect 1152 6132 1208 6134
rect 1152 4646 1208 4648
rect 1152 4594 1154 4646
rect 1154 4594 1206 4646
rect 1206 4594 1208 4646
rect 1152 4592 1208 4594
rect 1152 3106 1208 3108
rect 1152 3054 1154 3106
rect 1154 3054 1206 3106
rect 1206 3054 1208 3106
rect 1152 3052 1208 3054
rect 1152 1566 1208 1568
rect 1152 1514 1154 1566
rect 1154 1514 1206 1566
rect 1206 1514 1208 1566
rect 1152 1512 1208 1514
rect 280 26 336 28
rect 280 -26 282 26
rect 282 -26 334 26
rect 334 -26 336 26
rect 280 -28 336 -26
rect 1152 26 1208 28
rect 1152 -26 1154 26
rect 1154 -26 1206 26
rect 1206 -26 1208 26
rect 1152 -28 1208 -26
<< metal3 >>
rect 242 6188 374 6197
rect 242 6132 280 6188
rect 336 6132 374 6188
rect 242 6123 374 6132
rect 1114 6188 1246 6197
rect 1114 6132 1152 6188
rect 1208 6132 1246 6188
rect 1114 6123 1246 6132
rect 242 4648 374 4657
rect 242 4592 280 4648
rect 336 4592 374 4648
rect 242 4583 374 4592
rect 1114 4648 1246 4657
rect 1114 4592 1152 4648
rect 1208 4592 1246 4648
rect 1114 4583 1246 4592
rect 242 3108 374 3117
rect 242 3052 280 3108
rect 336 3052 374 3108
rect 242 3043 374 3052
rect 1114 3108 1246 3117
rect 1114 3052 1152 3108
rect 1208 3052 1246 3108
rect 1114 3043 1246 3052
rect 242 1568 374 1577
rect 242 1512 280 1568
rect 336 1512 374 1568
rect 242 1503 374 1512
rect 1114 1568 1246 1577
rect 1114 1512 1152 1568
rect 1208 1512 1246 1568
rect 1114 1503 1246 1512
rect 242 28 374 37
rect 242 -28 280 28
rect 336 -28 374 28
rect 242 -37 374 -28
rect 1114 28 1246 37
rect 1114 -28 1152 28
rect 1208 -28 1246 28
rect 1114 -37 1246 -28
use contact_18  contact_18_0
timestamp 1644969367
transform 1 0 1114 0 1 6123
box 0 0 1 1
use contact_17  contact_17_0
timestamp 1644969367
transform 1 0 1148 0 1 6128
box 0 0 1 1
use contact_13  contact_13_0
timestamp 1644969367
transform 1 0 1151 0 1 6137
box 0 0 1 1
use contact_18  contact_18_1
timestamp 1644969367
transform 1 0 242 0 1 6123
box 0 0 1 1
use contact_17  contact_17_1
timestamp 1644969367
transform 1 0 276 0 1 6128
box 0 0 1 1
use contact_13  contact_13_1
timestamp 1644969367
transform 1 0 279 0 1 6137
box 0 0 1 1
use contact_18  contact_18_2
timestamp 1644969367
transform 1 0 1114 0 1 4583
box 0 0 1 1
use contact_17  contact_17_2
timestamp 1644969367
transform 1 0 1148 0 1 4588
box 0 0 1 1
use contact_13  contact_13_2
timestamp 1644969367
transform 1 0 1151 0 1 4597
box 0 0 1 1
use contact_18  contact_18_3
timestamp 1644969367
transform 1 0 242 0 1 4583
box 0 0 1 1
use contact_17  contact_17_3
timestamp 1644969367
transform 1 0 276 0 1 4588
box 0 0 1 1
use contact_13  contact_13_3
timestamp 1644969367
transform 1 0 279 0 1 4597
box 0 0 1 1
use contact_18  contact_18_4
timestamp 1644969367
transform 1 0 1114 0 1 3043
box 0 0 1 1
use contact_17  contact_17_4
timestamp 1644969367
transform 1 0 1148 0 1 3048
box 0 0 1 1
use contact_13  contact_13_4
timestamp 1644969367
transform 1 0 1151 0 1 3057
box 0 0 1 1
use contact_18  contact_18_5
timestamp 1644969367
transform 1 0 242 0 1 3043
box 0 0 1 1
use contact_17  contact_17_5
timestamp 1644969367
transform 1 0 276 0 1 3048
box 0 0 1 1
use contact_13  contact_13_5
timestamp 1644969367
transform 1 0 279 0 1 3057
box 0 0 1 1
use contact_18  contact_18_6
timestamp 1644969367
transform 1 0 1114 0 1 4583
box 0 0 1 1
use contact_17  contact_17_6
timestamp 1644969367
transform 1 0 1148 0 1 4588
box 0 0 1 1
use contact_13  contact_13_6
timestamp 1644969367
transform 1 0 1151 0 1 4597
box 0 0 1 1
use contact_18  contact_18_7
timestamp 1644969367
transform 1 0 242 0 1 4583
box 0 0 1 1
use contact_17  contact_17_7
timestamp 1644969367
transform 1 0 276 0 1 4588
box 0 0 1 1
use contact_13  contact_13_7
timestamp 1644969367
transform 1 0 279 0 1 4597
box 0 0 1 1
use contact_18  contact_18_8
timestamp 1644969367
transform 1 0 1114 0 1 3043
box 0 0 1 1
use contact_17  contact_17_8
timestamp 1644969367
transform 1 0 1148 0 1 3048
box 0 0 1 1
use contact_13  contact_13_8
timestamp 1644969367
transform 1 0 1151 0 1 3057
box 0 0 1 1
use contact_18  contact_18_9
timestamp 1644969367
transform 1 0 242 0 1 3043
box 0 0 1 1
use contact_17  contact_17_9
timestamp 1644969367
transform 1 0 276 0 1 3048
box 0 0 1 1
use contact_13  contact_13_9
timestamp 1644969367
transform 1 0 279 0 1 3057
box 0 0 1 1
use contact_18  contact_18_10
timestamp 1644969367
transform 1 0 1114 0 1 1503
box 0 0 1 1
use contact_17  contact_17_10
timestamp 1644969367
transform 1 0 1148 0 1 1508
box 0 0 1 1
use contact_13  contact_13_10
timestamp 1644969367
transform 1 0 1151 0 1 1517
box 0 0 1 1
use contact_18  contact_18_11
timestamp 1644969367
transform 1 0 242 0 1 1503
box 0 0 1 1
use contact_17  contact_17_11
timestamp 1644969367
transform 1 0 276 0 1 1508
box 0 0 1 1
use contact_13  contact_13_11
timestamp 1644969367
transform 1 0 279 0 1 1517
box 0 0 1 1
use contact_18  contact_18_12
timestamp 1644969367
transform 1 0 1114 0 1 -37
box 0 0 1 1
use contact_17  contact_17_12
timestamp 1644969367
transform 1 0 1148 0 1 -32
box 0 0 1 1
use contact_13  contact_13_12
timestamp 1644969367
transform 1 0 1151 0 1 -23
box 0 0 1 1
use contact_18  contact_18_13
timestamp 1644969367
transform 1 0 242 0 1 -37
box 0 0 1 1
use contact_17  contact_17_13
timestamp 1644969367
transform 1 0 276 0 1 -32
box 0 0 1 1
use contact_13  contact_13_13
timestamp 1644969367
transform 1 0 279 0 1 -23
box 0 0 1 1
use contact_18  contact_18_14
timestamp 1644969367
transform 1 0 1114 0 1 1503
box 0 0 1 1
use contact_17  contact_17_14
timestamp 1644969367
transform 1 0 1148 0 1 1508
box 0 0 1 1
use contact_13  contact_13_14
timestamp 1644969367
transform 1 0 1151 0 1 1517
box 0 0 1 1
use contact_18  contact_18_15
timestamp 1644969367
transform 1 0 242 0 1 1503
box 0 0 1 1
use contact_17  contact_17_15
timestamp 1644969367
transform 1 0 276 0 1 1508
box 0 0 1 1
use contact_13  contact_13_15
timestamp 1644969367
transform 1 0 279 0 1 1517
box 0 0 1 1
use contact_17  contact_17_16
timestamp 1644969367
transform 1 0 1022 0 1 5714
box 0 0 1 1
use contact_17  contact_17_17
timestamp 1644969367
transform 1 0 150 0 1 5714
box 0 0 1 1
use contact_17  contact_17_18
timestamp 1644969367
transform 1 0 938 0 1 5838
box 0 0 1 1
use contact_17  contact_17_19
timestamp 1644969367
transform 1 0 66 0 1 5838
box 0 0 1 1
use contact_14  contact_14_0
timestamp 1644969367
transform 1 0 854 0 1 2968
box 0 0 1 1
use contact_13  contact_13_16
timestamp 1644969367
transform 1 0 520 0 1 2329
box 0 0 1 1
use contact_14  contact_14_1
timestamp 1644969367
transform 1 0 770 0 1 1428
box 0 0 1 1
use contact_13  contact_13_17
timestamp 1644969367
transform 1 0 520 0 1 705
box 0 0 1 1
use contact_15  contact_15_0
timestamp 1644969367
transform 1 0 1408 0 1 5723
box 0 0 1 1
use contact_14  contact_14_2
timestamp 1644969367
transform 1 0 1022 0 1 5714
box 0 0 1 1
use contact_13  contact_13_18
timestamp 1644969367
transform 1 0 1308 0 1 5847
box 0 0 1 1
use contact_14  contact_14_3
timestamp 1644969367
transform 1 0 938 0 1 5838
box 0 0 1 1
use contact_15  contact_15_1
timestamp 1644969367
transform 1 0 1408 0 1 3471
box 0 0 1 1
use contact_14  contact_14_4
timestamp 1644969367
transform 1 0 1022 0 1 3462
box 0 0 1 1
use contact_13  contact_13_19
timestamp 1644969367
transform 1 0 1308 0 1 3347
box 0 0 1 1
use contact_14  contact_14_5
timestamp 1644969367
transform 1 0 770 0 1 3338
box 0 0 1 1
use contact_15  contact_15_2
timestamp 1644969367
transform 1 0 1408 0 1 2643
box 0 0 1 1
use contact_14  contact_14_6
timestamp 1644969367
transform 1 0 854 0 1 2634
box 0 0 1 1
use contact_13  contact_13_20
timestamp 1644969367
transform 1 0 1308 0 1 2767
box 0 0 1 1
use contact_14  contact_14_7
timestamp 1644969367
transform 1 0 938 0 1 2758
box 0 0 1 1
use contact_15  contact_15_3
timestamp 1644969367
transform 1 0 1408 0 1 391
box 0 0 1 1
use contact_14  contact_14_8
timestamp 1644969367
transform 1 0 854 0 1 382
box 0 0 1 1
use contact_13  contact_13_21
timestamp 1644969367
transform 1 0 1308 0 1 267
box 0 0 1 1
use contact_14  contact_14_9
timestamp 1644969367
transform 1 0 770 0 1 258
box 0 0 1 1
use contact_14  contact_14_10
timestamp 1644969367
transform 1 0 150 0 1 2320
box 0 0 1 1
use contact_13  contact_13_22
timestamp 1644969367
transform 1 0 388 0 1 2329
box 0 0 1 1
use contact_14  contact_14_11
timestamp 1644969367
transform 1 0 66 0 1 696
box 0 0 1 1
use contact_13  contact_13_23
timestamp 1644969367
transform 1 0 388 0 1 705
box 0 0 1 1
use and2_dec  and2_dec_0
timestamp 1644969367
transform 1 0 1208 0 -1 6160
box -36 -17 872 1597
use and2_dec  and2_dec_1
timestamp 1644969367
transform 1 0 1208 0 1 3080
box -36 -17 872 1597
use and2_dec  and2_dec_2
timestamp 1644969367
transform 1 0 1208 0 -1 3080
box -36 -17 872 1597
use and2_dec  and2_dec_3
timestamp 1644969367
transform 1 0 1208 0 1 0
box -36 -17 872 1597
use pinv  pinv_0
timestamp 1644969367
transform 1 0 336 0 -1 3080
box -36 -17 404 1597
use pinv  pinv_1
timestamp 1644969367
transform 1 0 336 0 1 0
box -36 -17 404 1597
<< labels >>
rlabel metal2 s 72 696 124 760 4 in_0
rlabel metal2 s 156 2320 208 2384 4 in_1
rlabel locali s 1872 728 1872 728 4 out_0
rlabel locali s 1872 2352 1872 2352 4 out_1
rlabel locali s 1872 3808 1872 3808 4 out_2
rlabel locali s 1872 5432 1872 5432 4 out_3
rlabel metal3 s 242 1503 374 1577 4 vdd
rlabel metal3 s 1114 1503 1246 1577 4 vdd
rlabel metal3 s 242 4583 374 4657 4 vdd
rlabel metal3 s 1114 4583 1246 4657 4 vdd
rlabel metal3 s 1114 3043 1246 3117 4 gnd
rlabel metal3 s 242 -37 374 37 4 gnd
rlabel metal3 s 242 6123 374 6197 4 gnd
rlabel metal3 s 1114 -37 1246 37 4 gnd
rlabel metal3 s 1114 6123 1246 6197 4 gnd
rlabel metal3 s 242 3043 374 3117 4 gnd
<< properties >>
string FIXED_BBOX 1114 -37 1246 0
string GDS_FILE sram_0rw2r1w_32_128_sky130A.gds
string GDS_END 3064692
string GDS_START 3054220
<< end >>
