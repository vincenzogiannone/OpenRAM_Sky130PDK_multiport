magic
tech sky130A
timestamp 1644949024
<< checkpaint >>
rect -630 -651 2186 12971
<< metal1 >>
rect 0 11984 1556 11998
rect 0 11921 1556 11935
rect 0 11808 1556 11822
rect 0 11278 1556 11292
rect 0 11165 1556 11179
rect 0 11102 1556 11116
rect 0 10444 1556 10458
rect 0 10381 1556 10395
rect 0 10268 1556 10282
rect 0 9738 1556 9752
rect 0 9625 1556 9639
rect 0 9562 1556 9576
rect 0 8904 1556 8918
rect 0 8841 1556 8855
rect 0 8728 1556 8742
rect 0 8198 1556 8212
rect 0 8085 1556 8099
rect 0 8022 1556 8036
rect 0 7364 1556 7378
rect 0 7301 1556 7315
rect 0 7188 1556 7202
rect 0 6658 1556 6672
rect 0 6545 1556 6559
rect 0 6482 1556 6496
rect 0 5824 1556 5838
rect 0 5761 1556 5775
rect 0 5648 1556 5662
rect 0 5118 1556 5132
rect 0 5005 1556 5019
rect 0 4942 1556 4956
rect 0 4284 1556 4298
rect 0 4221 1556 4235
rect 0 4108 1556 4122
rect 0 3578 1556 3592
rect 0 3465 1556 3479
rect 0 3402 1556 3416
rect 0 2744 1556 2758
rect 0 2681 1556 2695
rect 0 2568 1556 2582
rect 0 2038 1556 2052
rect 0 1925 1556 1939
rect 0 1862 1556 1876
rect 0 1204 1556 1218
rect 0 1141 1556 1155
rect 0 1028 1556 1042
rect 0 498 1556 512
rect 0 385 1556 399
rect 0 322 1556 336
<< metal2 >>
rect 96 0 110 12320
rect 222 0 236 12320
rect 313 0 327 12320
rect 485 0 499 12320
rect 611 0 625 12320
rect 702 0 716 12320
rect 874 0 888 12320
rect 1000 0 1014 12320
rect 1091 0 1105 12320
rect 1263 0 1277 12320
rect 1389 0 1403 12320
rect 1480 0 1494 12320
use bitcell_array  bitcell_array_0
timestamp 1644949024
transform 1 0 0 0 1 0
box 0 -21 1556 12341
<< labels >>
rlabel metal1 s 0 385 1556 399 4 rwl_0_0
rlabel metal1 s 0 498 1556 512 4 rwl_1_0
rlabel metal1 s 0 322 1556 336 4 wwl_0_0
rlabel metal1 s 0 1141 1556 1155 4 rwl_0_1
rlabel metal1 s 0 1028 1556 1042 4 rwl_1_1
rlabel metal1 s 0 1204 1556 1218 4 wwl_0_1
rlabel metal1 s 0 1925 1556 1939 4 rwl_0_2
rlabel metal1 s 0 2038 1556 2052 4 rwl_1_2
rlabel metal1 s 0 1862 1556 1876 4 wwl_0_2
rlabel metal1 s 0 2681 1556 2695 4 rwl_0_3
rlabel metal1 s 0 2568 1556 2582 4 rwl_1_3
rlabel metal1 s 0 2744 1556 2758 4 wwl_0_3
rlabel metal1 s 0 3465 1556 3479 4 rwl_0_4
rlabel metal1 s 0 3578 1556 3592 4 rwl_1_4
rlabel metal1 s 0 3402 1556 3416 4 wwl_0_4
rlabel metal1 s 0 4221 1556 4235 4 rwl_0_5
rlabel metal1 s 0 4108 1556 4122 4 rwl_1_5
rlabel metal1 s 0 4284 1556 4298 4 wwl_0_5
rlabel metal1 s 0 5005 1556 5019 4 rwl_0_6
rlabel metal1 s 0 5118 1556 5132 4 rwl_1_6
rlabel metal1 s 0 4942 1556 4956 4 wwl_0_6
rlabel metal1 s 0 5761 1556 5775 4 rwl_0_7
rlabel metal1 s 0 5648 1556 5662 4 rwl_1_7
rlabel metal1 s 0 5824 1556 5838 4 wwl_0_7
rlabel metal1 s 0 6545 1556 6559 4 rwl_0_8
rlabel metal1 s 0 6658 1556 6672 4 rwl_1_8
rlabel metal1 s 0 6482 1556 6496 4 wwl_0_8
rlabel metal1 s 0 7301 1556 7315 4 rwl_0_9
rlabel metal1 s 0 7188 1556 7202 4 rwl_1_9
rlabel metal1 s 0 7364 1556 7378 4 wwl_0_9
rlabel metal1 s 0 8085 1556 8099 4 rwl_0_10
rlabel metal1 s 0 8198 1556 8212 4 rwl_1_10
rlabel metal1 s 0 8022 1556 8036 4 wwl_0_10
rlabel metal1 s 0 8841 1556 8855 4 rwl_0_11
rlabel metal1 s 0 8728 1556 8742 4 rwl_1_11
rlabel metal1 s 0 8904 1556 8918 4 wwl_0_11
rlabel metal1 s 0 9625 1556 9639 4 rwl_0_12
rlabel metal1 s 0 9738 1556 9752 4 rwl_1_12
rlabel metal1 s 0 9562 1556 9576 4 wwl_0_12
rlabel metal1 s 0 10381 1556 10395 4 rwl_0_13
rlabel metal1 s 0 10268 1556 10282 4 rwl_1_13
rlabel metal1 s 0 10444 1556 10458 4 wwl_0_13
rlabel metal1 s 0 11165 1556 11179 4 rwl_0_14
rlabel metal1 s 0 11278 1556 11292 4 rwl_1_14
rlabel metal1 s 0 11102 1556 11116 4 wwl_0_14
rlabel metal1 s 0 11921 1556 11935 4 rwl_0_15
rlabel metal1 s 0 11808 1556 11822 4 rwl_1_15
rlabel metal1 s 0 11984 1556 11998 4 wwl_0_15
rlabel metal2 s 96 0 110 12320 4 read_bl_0_0
rlabel metal2 s 485 0 499 12320 4 read_bl_0_1
rlabel metal2 s 874 0 888 12320 4 read_bl_0_2
rlabel metal2 s 1263 0 1277 12320 4 read_bl_0_3
rlabel metal2 s 222 0 236 12320 4 read_bl_1_0
rlabel metal2 s 611 0 625 12320 4 read_bl_1_1
rlabel metal2 s 1000 0 1014 12320 4 read_bl_1_2
rlabel metal2 s 1389 0 1403 12320 4 read_bl_1_3
rlabel metal2 s 313 0 327 12320 4 write_bl_0_0
rlabel metal2 s 702 0 716 12320 4 write_bl_0_1
rlabel metal2 s 1091 0 1105 12320 4 write_bl_0_2
rlabel metal2 s 1480 0 1494 12320 4 write_bl_0_3
<< properties >>
string FIXED_BBOX 0 0 3112 24640
string GDS_FILE sram_0rw2r1w_4_16_sky130A.gds
string GDS_END 121414
string GDS_START 109790
<< end >>
