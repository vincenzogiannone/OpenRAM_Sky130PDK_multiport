magic
tech sky130A
timestamp 1643678851
<< checkpaint >>
rect -630 -630 631 631
<< properties >>
string GDS_FILE sram_0rw2r1w_16_128_sky130A.gds
string GDS_END 1483052
string GDS_START 1482600
<< end >>
