magic
tech sky130A
magscale 1 2
timestamp 1643678851
<< checkpaint >>
rect -1319 -1316 2873 1602
<< nwell >>
rect -54 228 1608 342
rect -59 60 1613 228
rect -54 -54 1608 60
<< scpmos >>
rect 60 0 90 288
rect 168 0 198 288
rect 276 0 306 288
rect 384 0 414 288
rect 492 0 522 288
rect 600 0 630 288
rect 708 0 738 288
rect 816 0 846 288
rect 924 0 954 288
rect 1032 0 1062 288
rect 1140 0 1170 288
rect 1248 0 1278 288
rect 1356 0 1386 288
rect 1464 0 1494 288
<< pdiff >>
rect 0 161 60 288
rect 0 127 8 161
rect 42 127 60 161
rect 0 0 60 127
rect 90 161 168 288
rect 90 127 112 161
rect 146 127 168 161
rect 90 0 168 127
rect 198 161 276 288
rect 198 127 220 161
rect 254 127 276 161
rect 198 0 276 127
rect 306 161 384 288
rect 306 127 328 161
rect 362 127 384 161
rect 306 0 384 127
rect 414 161 492 288
rect 414 127 436 161
rect 470 127 492 161
rect 414 0 492 127
rect 522 161 600 288
rect 522 127 544 161
rect 578 127 600 161
rect 522 0 600 127
rect 630 161 708 288
rect 630 127 652 161
rect 686 127 708 161
rect 630 0 708 127
rect 738 161 816 288
rect 738 127 760 161
rect 794 127 816 161
rect 738 0 816 127
rect 846 161 924 288
rect 846 127 868 161
rect 902 127 924 161
rect 846 0 924 127
rect 954 161 1032 288
rect 954 127 976 161
rect 1010 127 1032 161
rect 954 0 1032 127
rect 1062 161 1140 288
rect 1062 127 1084 161
rect 1118 127 1140 161
rect 1062 0 1140 127
rect 1170 161 1248 288
rect 1170 127 1192 161
rect 1226 127 1248 161
rect 1170 0 1248 127
rect 1278 161 1356 288
rect 1278 127 1300 161
rect 1334 127 1356 161
rect 1278 0 1356 127
rect 1386 161 1464 288
rect 1386 127 1408 161
rect 1442 127 1464 161
rect 1386 0 1464 127
rect 1494 161 1554 288
rect 1494 127 1512 161
rect 1546 127 1554 161
rect 1494 0 1554 127
<< pdiffc >>
rect 8 127 42 161
rect 112 127 146 161
rect 220 127 254 161
rect 328 127 362 161
rect 436 127 470 161
rect 544 127 578 161
rect 652 127 686 161
rect 760 127 794 161
rect 868 127 902 161
rect 976 127 1010 161
rect 1084 127 1118 161
rect 1192 127 1226 161
rect 1300 127 1334 161
rect 1408 127 1442 161
rect 1512 127 1546 161
<< poly >>
rect 60 288 90 314
rect 168 288 198 314
rect 276 288 306 314
rect 384 288 414 314
rect 492 288 522 314
rect 600 288 630 314
rect 708 288 738 314
rect 816 288 846 314
rect 924 288 954 314
rect 1032 288 1062 314
rect 1140 288 1170 314
rect 1248 288 1278 314
rect 1356 288 1386 314
rect 1464 288 1494 314
rect 60 -26 90 0
rect 168 -26 198 0
rect 276 -26 306 0
rect 384 -26 414 0
rect 492 -26 522 0
rect 600 -26 630 0
rect 708 -26 738 0
rect 816 -26 846 0
rect 924 -26 954 0
rect 1032 -26 1062 0
rect 1140 -26 1170 0
rect 1248 -26 1278 0
rect 1356 -26 1386 0
rect 1464 -26 1494 0
rect 60 -56 1494 -26
<< locali >>
rect 8 161 42 177
rect 8 111 42 127
rect 112 161 146 177
rect 112 77 146 127
rect 220 161 254 177
rect 220 111 254 127
rect 328 161 362 177
rect 328 77 362 127
rect 436 161 470 177
rect 436 111 470 127
rect 544 161 578 177
rect 544 77 578 127
rect 652 161 686 177
rect 652 111 686 127
rect 760 161 794 177
rect 760 77 794 127
rect 868 161 902 177
rect 868 111 902 127
rect 976 161 1010 177
rect 976 77 1010 127
rect 1084 161 1118 177
rect 1084 111 1118 127
rect 1192 161 1226 177
rect 1192 77 1226 127
rect 1300 161 1334 177
rect 1300 111 1334 127
rect 1408 161 1442 177
rect 1408 77 1442 127
rect 1512 161 1546 177
rect 1512 111 1546 127
rect 112 43 1442 77
use contact_9  contact_9_0
timestamp 1643678851
transform 1 0 1504 0 1 103
box 0 0 2 2
use contact_9  contact_9_1
timestamp 1643678851
transform 1 0 1400 0 1 103
box 0 0 2 2
use contact_9  contact_9_2
timestamp 1643678851
transform 1 0 1292 0 1 103
box 0 0 2 2
use contact_9  contact_9_3
timestamp 1643678851
transform 1 0 1184 0 1 103
box 0 0 2 2
use contact_9  contact_9_4
timestamp 1643678851
transform 1 0 1076 0 1 103
box 0 0 2 2
use contact_9  contact_9_5
timestamp 1643678851
transform 1 0 968 0 1 103
box 0 0 2 2
use contact_9  contact_9_6
timestamp 1643678851
transform 1 0 860 0 1 103
box 0 0 2 2
use contact_9  contact_9_7
timestamp 1643678851
transform 1 0 752 0 1 103
box 0 0 2 2
use contact_9  contact_9_8
timestamp 1643678851
transform 1 0 644 0 1 103
box 0 0 2 2
use contact_9  contact_9_9
timestamp 1643678851
transform 1 0 536 0 1 103
box 0 0 2 2
use contact_9  contact_9_10
timestamp 1643678851
transform 1 0 428 0 1 103
box 0 0 2 2
use contact_9  contact_9_11
timestamp 1643678851
transform 1 0 320 0 1 103
box 0 0 2 2
use contact_9  contact_9_12
timestamp 1643678851
transform 1 0 212 0 1 103
box 0 0 2 2
use contact_9  contact_9_13
timestamp 1643678851
transform 1 0 104 0 1 103
box 0 0 2 2
use contact_9  contact_9_14
timestamp 1643678851
transform 1 0 0 0 1 103
box 0 0 2 2
<< labels >>
rlabel mvvaractor s 777 -41 777 -41 4 G
rlabel locali s 1317 144 1317 144 4 S
rlabel locali s 453 144 453 144 4 S
rlabel locali s 885 144 885 144 4 S
rlabel locali s 669 144 669 144 4 S
rlabel locali s 237 144 237 144 4 S
rlabel locali s 1101 144 1101 144 4 S
rlabel locali s 1529 144 1529 144 4 S
rlabel locali s 25 144 25 144 4 S
rlabel locali s 777 60 777 60 4 D
<< properties >>
string FIXED_BBOX -54 -56 1608 60
string GDS_FILE sram_0rw2r1w_16_128_sky130A.gds
string GDS_END 2060054
string GDS_START 2056586
<< end >>
