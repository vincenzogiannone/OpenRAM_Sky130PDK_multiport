magic
tech sky130A
timestamp 1643280717
<< nwell >>
rect 0 158 136 525
<< nmos >>
rect 61 61 76 103
<< pmos >>
rect 61 176 76 446
<< ndiff >>
rect 19 91 61 103
rect 19 74 25 91
rect 43 74 61 91
rect 19 61 61 74
rect 76 91 118 103
rect 76 74 94 91
rect 112 74 118 91
rect 76 61 118 74
<< pdiff >>
rect 19 415 61 446
rect 19 398 25 415
rect 42 398 61 415
rect 19 367 61 398
rect 19 350 25 367
rect 42 350 61 367
rect 19 319 61 350
rect 19 302 25 319
rect 42 302 61 319
rect 19 271 61 302
rect 19 254 25 271
rect 42 254 61 271
rect 19 223 61 254
rect 19 206 25 223
rect 42 206 61 223
rect 19 176 61 206
rect 76 415 118 446
rect 76 398 95 415
rect 112 398 118 415
rect 76 367 118 398
rect 76 350 95 367
rect 112 350 118 367
rect 76 319 118 350
rect 76 302 95 319
rect 112 302 118 319
rect 76 271 118 302
rect 76 254 95 271
rect 112 254 118 271
rect 76 223 118 254
rect 76 206 95 223
rect 112 206 118 223
rect 76 176 118 206
<< ndiffc >>
rect 25 74 43 91
rect 94 74 112 91
<< pdiffc >>
rect 25 398 42 415
rect 25 350 42 367
rect 25 302 42 319
rect 25 254 42 271
rect 25 206 42 223
rect 95 398 112 415
rect 95 350 112 367
rect 95 302 112 319
rect 95 254 112 271
rect 95 206 112 223
<< psubdiff >>
rect 47 26 89 34
rect 47 8 59 26
rect 77 8 89 26
rect 47 0 89 8
<< nsubdiff >>
rect 47 499 89 507
rect 47 481 59 499
rect 77 481 89 499
rect 47 473 89 481
<< psubdiffcont >>
rect 59 8 77 26
<< nsubdiffcont >>
rect 59 481 77 499
<< poly >>
rect 61 446 76 466
rect 61 153 76 176
rect 1 145 76 153
rect 1 128 6 145
rect 23 128 76 145
rect 1 120 76 128
rect 61 103 76 120
rect 61 48 76 61
<< polycont >>
rect 6 128 23 145
<< locali >>
rect 59 499 77 507
rect 31 481 59 490
rect 31 473 77 481
rect 31 446 49 473
rect 19 415 49 446
rect 19 398 25 415
rect 42 398 49 415
rect 19 367 49 398
rect 19 350 25 367
rect 42 350 49 367
rect 19 319 49 350
rect 19 302 25 319
rect 42 302 49 319
rect 19 271 49 302
rect 19 254 25 271
rect 42 254 49 271
rect 19 223 49 254
rect 19 206 25 223
rect 42 206 49 223
rect 19 176 49 206
rect 88 415 118 446
rect 88 398 95 415
rect 112 398 118 415
rect 88 367 118 398
rect 88 350 95 367
rect 112 350 118 367
rect 88 319 118 350
rect 88 302 95 319
rect 112 302 118 319
rect 88 271 118 302
rect 88 254 95 271
rect 112 254 118 271
rect 88 223 118 254
rect 88 206 95 223
rect 112 206 118 223
rect 88 176 118 206
rect 6 145 23 153
rect 6 120 23 128
rect 101 145 118 176
rect 101 103 118 128
rect 19 91 49 103
rect 19 74 25 91
rect 43 74 49 91
rect 19 61 49 74
rect 88 91 118 103
rect 88 74 94 91
rect 112 74 118 91
rect 88 61 118 74
rect 32 34 49 61
rect 32 26 77 34
rect 32 17 59 26
rect 59 0 77 8
<< viali >>
rect 59 481 77 499
rect 6 128 23 145
rect 101 128 118 145
rect 59 8 77 26
<< metal1 >>
rect 0 499 136 505
rect 0 481 59 499
rect 77 481 136 499
rect 0 475 136 481
rect 1 150 28 153
rect 1 124 2 150
rect 1 120 28 124
rect 96 149 123 152
rect 96 123 97 149
rect 96 120 123 123
rect 0 26 136 32
rect 0 8 59 26
rect 77 8 136 26
rect 0 2 136 8
<< via1 >>
rect 2 145 28 150
rect 2 128 6 145
rect 6 128 23 145
rect 23 128 28 145
rect 2 124 28 128
rect 97 145 123 149
rect 97 128 101 145
rect 101 128 118 145
rect 118 128 123 145
rect 97 123 123 128
<< metal2 >>
rect 7 153 21 525
rect 2 150 28 153
rect 101 152 115 525
rect 2 120 28 124
rect 96 149 123 152
rect 96 123 97 149
rect 96 120 123 123
rect 7 0 21 120
rect 101 0 115 120
<< labels >>
flabel metal1 16 491 16 491 0 FreeSans 80 0 0 0 vdd
port 6 nsew
flabel metal1 20 17 20 17 0 FreeSans 80 0 0 0 gnd
port 7 nsew
flabel metal2 14 116 14 116 0 FreeSans 80 0 0 0 rbl
port 10 nsew
flabel metal2 107 49 107 49 0 FreeSans 80 0 0 0 dout
port 11 nsew
<< properties >>
string FIXED_BBOX 0 0 136 525
<< end >>
