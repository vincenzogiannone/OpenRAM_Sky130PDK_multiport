magic
tech sky130A
magscale 1 2
timestamp 1644969367
<< checkpaint >>
rect -1260 -1260 1532 2310
<< nwell >>
rect 0 316 272 1050
<< pwell >>
rect 94 0 178 68
<< nmos >>
rect 122 122 152 206
<< pmos >>
rect 122 352 152 892
<< ndiff >>
rect 38 182 122 206
rect 38 148 51 182
rect 85 148 122 182
rect 38 122 122 148
rect 152 182 236 206
rect 152 148 189 182
rect 223 148 236 182
rect 152 122 236 148
<< pdiff >>
rect 38 830 122 892
rect 38 796 50 830
rect 84 796 122 830
rect 38 734 122 796
rect 38 700 50 734
rect 84 700 122 734
rect 38 638 122 700
rect 38 604 50 638
rect 84 604 122 638
rect 38 542 122 604
rect 38 508 50 542
rect 84 508 122 542
rect 38 446 122 508
rect 38 412 50 446
rect 84 412 122 446
rect 38 352 122 412
rect 152 830 236 892
rect 152 796 190 830
rect 224 796 236 830
rect 152 734 236 796
rect 152 700 190 734
rect 224 700 236 734
rect 152 638 236 700
rect 152 604 190 638
rect 224 604 236 638
rect 152 542 236 604
rect 152 508 190 542
rect 224 508 236 542
rect 152 446 236 508
rect 152 412 190 446
rect 224 412 236 446
rect 152 352 236 412
<< ndiffc >>
rect 51 148 85 182
rect 189 148 223 182
<< pdiffc >>
rect 50 796 84 830
rect 50 700 84 734
rect 50 604 84 638
rect 50 508 84 542
rect 50 412 84 446
rect 190 796 224 830
rect 190 700 224 734
rect 190 604 224 638
rect 190 508 224 542
rect 190 412 224 446
<< psubdiff >>
rect 94 51 178 68
rect 94 17 119 51
rect 153 17 178 51
rect 94 0 178 17
<< nsubdiff >>
rect 94 997 178 1014
rect 94 963 119 997
rect 153 963 178 997
rect 94 946 178 963
<< psubdiffcont >>
rect 119 17 153 51
<< nsubdiffcont >>
rect 119 963 153 997
<< poly >>
rect 122 892 152 932
rect 122 306 152 352
rect 2 290 152 306
rect 2 256 12 290
rect 46 256 152 290
rect 2 240 152 256
rect 122 206 152 240
rect 122 96 152 122
<< polycont >>
rect 12 256 46 290
<< locali >>
rect 118 997 154 1014
rect 118 980 119 997
rect 62 963 119 980
rect 153 963 154 997
rect 62 946 154 963
rect 62 892 98 946
rect 38 830 98 892
rect 38 796 50 830
rect 84 796 98 830
rect 38 734 98 796
rect 38 700 50 734
rect 84 700 98 734
rect 38 638 98 700
rect 38 604 50 638
rect 84 604 98 638
rect 38 542 98 604
rect 38 508 50 542
rect 84 508 98 542
rect 38 446 98 508
rect 38 412 50 446
rect 84 412 98 446
rect 38 352 98 412
rect 176 830 236 892
rect 176 796 190 830
rect 224 796 236 830
rect 176 734 236 796
rect 176 700 190 734
rect 224 700 236 734
rect 176 638 236 700
rect 176 604 190 638
rect 224 604 236 638
rect 176 542 236 604
rect 176 508 190 542
rect 224 508 236 542
rect 176 446 236 508
rect 176 412 190 446
rect 224 412 236 446
rect 176 352 236 412
rect 12 290 46 306
rect 12 240 46 256
rect 202 290 236 352
rect 202 206 236 256
rect 38 182 98 206
rect 38 148 51 182
rect 85 148 98 182
rect 38 122 98 148
rect 176 182 236 206
rect 176 148 189 182
rect 223 148 236 182
rect 176 122 236 148
rect 64 68 98 122
rect 64 51 154 68
rect 64 34 119 51
rect 118 17 119 34
rect 153 17 154 51
rect 118 0 154 17
<< viali >>
rect 119 963 153 997
rect 12 256 46 290
rect 202 256 236 290
rect 119 17 153 51
<< metal1 >>
rect 0 997 272 1010
rect 0 963 119 997
rect 153 963 272 997
rect 0 950 272 963
rect 2 300 56 306
rect 2 248 4 300
rect 2 240 56 248
rect 192 298 246 304
rect 192 246 194 298
rect 192 240 246 246
rect 0 51 272 64
rect 0 17 119 51
rect 153 17 272 51
rect 0 4 272 17
<< via1 >>
rect 4 290 56 300
rect 4 256 12 290
rect 12 256 46 290
rect 46 256 56 290
rect 4 248 56 256
rect 194 290 246 298
rect 194 256 202 290
rect 202 256 236 290
rect 236 256 246 290
rect 194 246 246 256
<< metal2 >>
rect 14 306 42 1050
rect 4 300 56 306
rect 202 304 230 1050
rect 4 240 56 248
rect 192 298 246 304
rect 192 246 194 298
rect 192 240 246 246
rect 14 0 42 240
rect 202 0 230 240
<< labels >>
rlabel metal1 s 0 950 272 1010 4 vdd
port 1 nsew
rlabel metal1 s 0 4 272 64 4 gnd
port 2 nsew
rlabel metal2 s 14 0 42 240 4 rbl
port 3 nsew
rlabel metal2 s 202 0 230 240 4 dout
port 4 nsew
rlabel metal2 s 28 120 28 120 4 rbl
rlabel metal2 s 216 120 216 120 4 dout
rlabel metal1 s 136 980 136 980 4 vdd
rlabel metal1 s 136 34 136 34 4 gnd
<< properties >>
string FIXED_BBOX 0 0 272 1050
string GDS_FILE sram_0rw2r1w_32_128_sky130A.gds
string GDS_END 2602382
string GDS_START 2597754
<< end >>
