magic
tech sky130A
magscale 1 2
timestamp 1643593061
<< checkpaint >>
rect -1296 -1277 4604 2155
<< nwell >>
rect -36 402 3344 895
<< locali >>
rect 0 821 3308 855
rect 48 344 114 410
rect 196 360 449 394
rect 568 360 925 394
rect 1241 354 1725 388
rect 2473 354 2507 388
rect 0 -17 3308 17
use pinv_8  pinv_8_0
timestamp 1643593061
transform 1 0 1644 0 1 0
box -36 -17 1700 895
use pinv_7  pinv_7_0
timestamp 1643593061
transform 1 0 844 0 1 0
box -36 -17 836 895
use pinv_6  pinv_6_0
timestamp 1643593061
transform 1 0 368 0 1 0
box -36 -17 512 895
use pinv_5  pinv_5_0
timestamp 1643593061
transform 1 0 0 0 1 0
box -36 -17 404 895
<< labels >>
rlabel locali s 2490 371 2490 371 4 Z
rlabel locali s 81 377 81 377 4 A
rlabel locali s 1654 0 1654 0 4 gnd
rlabel locali s 1654 838 1654 838 4 vdd
<< properties >>
string FIXED_BBOX 0 0 3308 838
string GDS_FILE sram_0rw2r1w_2_16_sky130A.gds
string GDS_END 525876
string GDS_START 524604
<< end >>
