magic
tech sky130A
magscale 1 2
timestamp 1644949024
<< checkpaint >>
rect -1260 -1284 4352 2212
<< metal1 >>
rect 323 900 375 906
rect 323 842 375 848
rect 1121 900 1173 906
rect 1121 842 1173 848
rect 1919 900 1971 906
rect 1919 842 1971 848
rect 2717 900 2769 906
rect 2717 842 2769 848
rect 0 356 3092 384
rect 323 68 375 74
rect 323 10 375 16
rect 1121 68 1173 74
rect 1121 10 1173 16
rect 1919 68 1971 74
rect 1919 10 1971 16
rect 2717 68 2769 74
rect 2717 10 2769 16
<< via1 >>
rect 323 848 375 900
rect 1121 848 1173 900
rect 1919 848 1971 900
rect 2717 848 2769 900
rect 323 16 375 68
rect 1121 16 1173 68
rect 1919 16 1971 68
rect 2717 16 2769 68
<< metal2 >>
rect 321 902 377 911
rect 321 837 377 846
rect 630 322 658 952
rect 1119 902 1175 911
rect 1119 837 1175 846
rect 1428 322 1456 952
rect 1917 902 1973 911
rect 1917 837 1973 846
rect 2226 322 2254 952
rect 2715 902 2771 911
rect 2715 837 2771 846
rect 3024 322 3052 952
rect 196 272 250 300
rect 994 272 1048 300
rect 1792 272 1846 300
rect 2590 272 2644 300
rect 321 70 377 79
rect 321 5 377 14
rect 1119 70 1175 79
rect 1119 5 1175 14
rect 1917 70 1973 79
rect 1917 5 1973 14
rect 2715 70 2771 79
rect 2715 5 2771 14
<< via2 >>
rect 321 900 377 902
rect 321 848 323 900
rect 323 848 375 900
rect 375 848 377 900
rect 321 846 377 848
rect 1119 900 1175 902
rect 1119 848 1121 900
rect 1121 848 1173 900
rect 1173 848 1175 900
rect 1119 846 1175 848
rect 1917 900 1973 902
rect 1917 848 1919 900
rect 1919 848 1971 900
rect 1971 848 1973 900
rect 1917 846 1973 848
rect 2715 900 2771 902
rect 2715 848 2717 900
rect 2717 848 2769 900
rect 2769 848 2771 900
rect 2715 846 2771 848
rect 321 68 377 70
rect 321 16 323 68
rect 323 16 375 68
rect 375 16 377 68
rect 321 14 377 16
rect 1119 68 1175 70
rect 1119 16 1121 68
rect 1121 16 1173 68
rect 1173 16 1175 68
rect 1119 14 1175 16
rect 1917 68 1973 70
rect 1917 16 1919 68
rect 1919 16 1971 68
rect 1971 16 1973 68
rect 1917 14 1973 16
rect 2715 68 2771 70
rect 2715 16 2717 68
rect 2717 16 2769 68
rect 2769 16 2771 68
rect 2715 14 2771 16
<< metal3 >>
rect 316 902 382 940
rect 316 846 321 902
rect 377 846 382 902
rect 316 808 382 846
rect 1114 902 1180 940
rect 1114 846 1119 902
rect 1175 846 1180 902
rect 1114 808 1180 846
rect 1912 902 1978 940
rect 1912 846 1917 902
rect 1973 846 1978 902
rect 1912 808 1978 846
rect 2710 902 2776 940
rect 2710 846 2715 902
rect 2771 846 2776 902
rect 2710 808 2776 846
rect 316 70 382 108
rect 316 14 321 70
rect 377 14 382 70
rect 316 -24 382 14
rect 1114 70 1180 108
rect 1114 14 1119 70
rect 1175 14 1180 70
rect 1114 -24 1180 14
rect 1912 70 1978 108
rect 1912 14 1917 70
rect 1973 14 1978 70
rect 1912 -24 1978 14
rect 2710 70 2776 108
rect 2710 14 2715 70
rect 2771 14 2776 70
rect 2710 -24 2776 14
use contact_23  contact_23_0
timestamp 1644949024
transform 1 0 2710 0 1 -24
box 0 0 1 1
use contact_22  contact_22_0
timestamp 1644949024
transform 1 0 2717 0 1 10
box 0 0 1 1
use contact_23  contact_23_1
timestamp 1644949024
transform 1 0 2710 0 1 808
box 0 0 1 1
use contact_22  contact_22_1
timestamp 1644949024
transform 1 0 2717 0 1 842
box 0 0 1 1
use contact_23  contact_23_2
timestamp 1644949024
transform 1 0 1912 0 1 -24
box 0 0 1 1
use contact_22  contact_22_2
timestamp 1644949024
transform 1 0 1919 0 1 10
box 0 0 1 1
use contact_23  contact_23_3
timestamp 1644949024
transform 1 0 1912 0 1 808
box 0 0 1 1
use contact_22  contact_22_3
timestamp 1644949024
transform 1 0 1919 0 1 842
box 0 0 1 1
use contact_23  contact_23_4
timestamp 1644949024
transform 1 0 1114 0 1 -24
box 0 0 1 1
use contact_22  contact_22_4
timestamp 1644949024
transform 1 0 1121 0 1 10
box 0 0 1 1
use contact_23  contact_23_5
timestamp 1644949024
transform 1 0 1114 0 1 808
box 0 0 1 1
use contact_22  contact_22_5
timestamp 1644949024
transform 1 0 1121 0 1 842
box 0 0 1 1
use contact_23  contact_23_6
timestamp 1644949024
transform 1 0 316 0 1 -24
box 0 0 1 1
use contact_22  contact_22_6
timestamp 1644949024
transform 1 0 323 0 1 10
box 0 0 1 1
use contact_23  contact_23_7
timestamp 1644949024
transform 1 0 316 0 1 808
box 0 0 1 1
use contact_22  contact_22_7
timestamp 1644949024
transform 1 0 323 0 1 842
box 0 0 1 1
use write_driver_multiport  write_driver_multiport_0
timestamp 1644949024
transform 1 0 2394 0 1 0
box 0 0 698 952
use write_driver_multiport  write_driver_multiport_1
timestamp 1644949024
transform 1 0 1596 0 1 0
box 0 0 698 952
use write_driver_multiport  write_driver_multiport_2
timestamp 1644949024
transform 1 0 798 0 1 0
box 0 0 698 952
use write_driver_multiport  write_driver_multiport_3
timestamp 1644949024
transform 1 0 0 0 1 0
box 0 0 698 952
<< labels >>
rlabel metal2 s 196 272 250 300 4 din_0
rlabel metal2 s 630 322 658 952 4 wbl0_0
rlabel metal3 s 1114 808 1180 940 4 vdd
rlabel metal3 s 2710 808 2776 940 4 vdd
rlabel metal3 s 1912 808 1978 940 4 vdd
rlabel metal3 s 316 808 382 940 4 vdd
rlabel metal3 s 316 -24 382 108 4 gnd
rlabel metal3 s 1114 -24 1180 108 4 gnd
rlabel metal3 s 1912 -24 1978 108 4 gnd
rlabel metal3 s 2710 -24 2776 108 4 gnd
rlabel metal2 s 994 272 1048 300 4 din_1
rlabel metal2 s 1428 322 1456 952 4 wbl0_1
rlabel metal2 s 1792 272 1846 300 4 din_2
rlabel metal2 s 2226 322 2254 952 4 wbl0_2
rlabel metal2 s 2590 272 2644 300 4 din_3
rlabel metal2 s 3024 322 3052 952 4 wbl0_3
rlabel metal1 s 0 356 3092 384 4 en
<< properties >>
string FIXED_BBOX 2710 -24 2776 0
string GDS_FILE sram_0rw2r1w_4_16_sky130A.gds
string GDS_END 219850
string GDS_START 215182
<< end >>
