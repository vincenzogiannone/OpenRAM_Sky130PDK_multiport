magic
tech sky130A
magscale 1 2
timestamp 1643678851
<< checkpaint >>
rect -1299 -1302 24972 2176
<< via1 >>
rect 715 812 767 864
rect 2197 812 2249 864
rect 3679 812 3731 864
rect 5161 812 5213 864
rect 6643 812 6695 864
rect 8125 812 8177 864
rect 9607 812 9659 864
rect 11089 812 11141 864
rect 12571 812 12623 864
rect 14053 812 14105 864
rect 15535 812 15587 864
rect 17017 812 17069 864
rect 18499 812 18551 864
rect 19981 812 20033 864
rect 21463 812 21515 864
rect 22945 812 22997 864
rect 715 -26 767 26
rect 2197 -26 2249 26
rect 3679 -26 3731 26
rect 5161 -26 5213 26
rect 6643 -26 6695 26
rect 8125 -26 8177 26
rect 9607 -26 9659 26
rect 11089 -26 11141 26
rect 12571 -26 12623 26
rect 14053 -26 14105 26
rect 15535 -26 15587 26
rect 17017 -26 17069 26
rect 18499 -26 18551 26
rect 19981 -26 20033 26
rect 21463 -26 21515 26
rect 22945 -26 22997 26
<< metal2 >>
rect 721 866 761 872
rect 2203 866 2243 872
rect 3685 866 3725 872
rect 5167 866 5207 872
rect 6649 866 6689 872
rect 8131 866 8171 872
rect 9613 866 9653 872
rect 11095 866 11135 872
rect 12577 866 12617 872
rect 14059 866 14099 872
rect 15541 866 15581 872
rect 17023 866 17063 872
rect 18505 866 18545 872
rect 19987 866 20027 872
rect 21469 866 21509 872
rect 22951 866 22991 872
rect 0 336 28 838
rect 721 804 761 810
rect 1482 336 1510 838
rect 2203 804 2243 810
rect 2964 336 2992 838
rect 3685 804 3725 810
rect 4446 336 4474 838
rect 5167 804 5207 810
rect 5928 336 5956 838
rect 6649 804 6689 810
rect 7410 336 7438 838
rect 8131 804 8171 810
rect 8892 336 8920 838
rect 9613 804 9653 810
rect 10374 336 10402 838
rect 11095 804 11135 810
rect 11856 336 11884 838
rect 12577 804 12617 810
rect 13338 336 13366 838
rect 14059 804 14099 810
rect 14820 336 14848 838
rect 15541 804 15581 810
rect 16302 336 16330 838
rect 17023 804 17063 810
rect 17784 336 17812 838
rect 18505 804 18545 810
rect 19266 336 19294 838
rect 19987 804 20027 810
rect 20748 336 20776 838
rect 21469 804 21509 810
rect 22230 336 22258 838
rect 22951 804 22991 810
rect 0 0 28 280
rect 180 232 234 260
rect 1260 228 1314 256
rect 721 28 761 34
rect 1482 0 1510 280
rect 1662 232 1716 260
rect 2742 228 2796 256
rect 2203 28 2243 34
rect 2964 0 2992 280
rect 3144 232 3198 260
rect 4224 228 4278 256
rect 3685 28 3725 34
rect 4446 0 4474 280
rect 4626 232 4680 260
rect 5706 228 5760 256
rect 5167 28 5207 34
rect 5928 0 5956 280
rect 6108 232 6162 260
rect 7188 228 7242 256
rect 6649 28 6689 34
rect 7410 0 7438 280
rect 7590 232 7644 260
rect 8670 228 8724 256
rect 8131 28 8171 34
rect 8892 0 8920 280
rect 9072 232 9126 260
rect 10152 228 10206 256
rect 9613 28 9653 34
rect 10374 0 10402 280
rect 10554 232 10608 260
rect 11634 228 11688 256
rect 11095 28 11135 34
rect 11856 0 11884 280
rect 12036 232 12090 260
rect 13116 228 13170 256
rect 12577 28 12617 34
rect 13338 0 13366 280
rect 13518 232 13572 260
rect 14598 228 14652 256
rect 14059 28 14099 34
rect 14820 0 14848 280
rect 15000 232 15054 260
rect 16080 228 16134 256
rect 15541 28 15581 34
rect 16302 0 16330 280
rect 16482 232 16536 260
rect 17562 228 17616 256
rect 17023 28 17063 34
rect 17784 0 17812 280
rect 17964 232 18018 260
rect 19044 228 19098 256
rect 18505 28 18545 34
rect 19266 0 19294 280
rect 19446 232 19500 260
rect 20526 228 20580 256
rect 19987 28 20027 34
rect 20748 0 20776 280
rect 20928 232 20982 260
rect 22008 228 22062 256
rect 21469 28 21509 34
rect 22230 0 22258 280
rect 22410 232 22464 260
rect 23490 228 23544 256
rect 22951 28 22991 34
rect 721 -34 761 -28
rect 2203 -34 2243 -28
rect 3685 -34 3725 -28
rect 5167 -34 5207 -28
rect 6649 -34 6689 -28
rect 8131 -34 8171 -28
rect 9613 -34 9653 -28
rect 11095 -34 11135 -28
rect 12577 -34 12617 -28
rect 14059 -34 14099 -28
rect 15541 -34 15581 -28
rect 17023 -34 17063 -28
rect 18505 -34 18545 -28
rect 19987 -34 20027 -28
rect 21469 -34 21509 -28
rect 22951 -34 22991 -28
<< via2 >>
rect 713 864 769 866
rect 713 812 715 864
rect 715 812 767 864
rect 767 812 769 864
rect 2195 864 2251 866
rect 713 810 769 812
rect 2195 812 2197 864
rect 2197 812 2249 864
rect 2249 812 2251 864
rect 3677 864 3733 866
rect 2195 810 2251 812
rect 3677 812 3679 864
rect 3679 812 3731 864
rect 3731 812 3733 864
rect 5159 864 5215 866
rect 3677 810 3733 812
rect 5159 812 5161 864
rect 5161 812 5213 864
rect 5213 812 5215 864
rect 6641 864 6697 866
rect 5159 810 5215 812
rect 6641 812 6643 864
rect 6643 812 6695 864
rect 6695 812 6697 864
rect 8123 864 8179 866
rect 6641 810 6697 812
rect 8123 812 8125 864
rect 8125 812 8177 864
rect 8177 812 8179 864
rect 9605 864 9661 866
rect 8123 810 8179 812
rect 9605 812 9607 864
rect 9607 812 9659 864
rect 9659 812 9661 864
rect 11087 864 11143 866
rect 9605 810 9661 812
rect 11087 812 11089 864
rect 11089 812 11141 864
rect 11141 812 11143 864
rect 12569 864 12625 866
rect 11087 810 11143 812
rect 12569 812 12571 864
rect 12571 812 12623 864
rect 12623 812 12625 864
rect 14051 864 14107 866
rect 12569 810 12625 812
rect 14051 812 14053 864
rect 14053 812 14105 864
rect 14105 812 14107 864
rect 15533 864 15589 866
rect 14051 810 14107 812
rect 15533 812 15535 864
rect 15535 812 15587 864
rect 15587 812 15589 864
rect 17015 864 17071 866
rect 15533 810 15589 812
rect 17015 812 17017 864
rect 17017 812 17069 864
rect 17069 812 17071 864
rect 18497 864 18553 866
rect 17015 810 17071 812
rect 18497 812 18499 864
rect 18499 812 18551 864
rect 18551 812 18553 864
rect 19979 864 20035 866
rect 18497 810 18553 812
rect 19979 812 19981 864
rect 19981 812 20033 864
rect 20033 812 20035 864
rect 21461 864 21517 866
rect 19979 810 20035 812
rect 21461 812 21463 864
rect 21463 812 21515 864
rect 21515 812 21517 864
rect 22943 864 22999 866
rect 21461 810 21517 812
rect 22943 812 22945 864
rect 22945 812 22997 864
rect 22997 812 22999 864
rect 22943 810 22999 812
rect -1 280 55 336
rect 1481 280 1537 336
rect 2963 280 3019 336
rect 4445 280 4501 336
rect 5927 280 5983 336
rect 7409 280 7465 336
rect 8891 280 8947 336
rect 10373 280 10429 336
rect 11855 280 11911 336
rect 13337 280 13393 336
rect 14819 280 14875 336
rect 16301 280 16357 336
rect 17783 280 17839 336
rect 19265 280 19321 336
rect 20747 280 20803 336
rect 22229 280 22285 336
rect 713 26 769 28
rect 713 -26 715 26
rect 715 -26 767 26
rect 767 -26 769 26
rect 2195 26 2251 28
rect 713 -28 769 -26
rect 2195 -26 2197 26
rect 2197 -26 2249 26
rect 2249 -26 2251 26
rect 3677 26 3733 28
rect 2195 -28 2251 -26
rect 3677 -26 3679 26
rect 3679 -26 3731 26
rect 3731 -26 3733 26
rect 5159 26 5215 28
rect 3677 -28 3733 -26
rect 5159 -26 5161 26
rect 5161 -26 5213 26
rect 5213 -26 5215 26
rect 6641 26 6697 28
rect 5159 -28 5215 -26
rect 6641 -26 6643 26
rect 6643 -26 6695 26
rect 6695 -26 6697 26
rect 8123 26 8179 28
rect 6641 -28 6697 -26
rect 8123 -26 8125 26
rect 8125 -26 8177 26
rect 8177 -26 8179 26
rect 9605 26 9661 28
rect 8123 -28 8179 -26
rect 9605 -26 9607 26
rect 9607 -26 9659 26
rect 9659 -26 9661 26
rect 11087 26 11143 28
rect 9605 -28 9661 -26
rect 11087 -26 11089 26
rect 11089 -26 11141 26
rect 11141 -26 11143 26
rect 12569 26 12625 28
rect 11087 -28 11143 -26
rect 12569 -26 12571 26
rect 12571 -26 12623 26
rect 12623 -26 12625 26
rect 14051 26 14107 28
rect 12569 -28 12625 -26
rect 14051 -26 14053 26
rect 14053 -26 14105 26
rect 14105 -26 14107 26
rect 15533 26 15589 28
rect 14051 -28 14107 -26
rect 15533 -26 15535 26
rect 15535 -26 15587 26
rect 15587 -26 15589 26
rect 17015 26 17071 28
rect 15533 -28 15589 -26
rect 17015 -26 17017 26
rect 17017 -26 17069 26
rect 17069 -26 17071 26
rect 18497 26 18553 28
rect 17015 -28 17071 -26
rect 18497 -26 18499 26
rect 18499 -26 18551 26
rect 18551 -26 18553 26
rect 19979 26 20035 28
rect 18497 -28 18553 -26
rect 19979 -26 19981 26
rect 19981 -26 20033 26
rect 20033 -26 20035 26
rect 21461 26 21517 28
rect 19979 -28 20035 -26
rect 21461 -26 21463 26
rect 21463 -26 21515 26
rect 21515 -26 21517 26
rect 22943 26 22999 28
rect 21461 -28 21517 -26
rect 22943 -26 22945 26
rect 22945 -26 22997 26
rect 22997 -26 22999 26
rect 22943 -28 22999 -26
<< metal3 >>
rect 675 866 807 871
rect 675 810 713 866
rect 769 810 807 866
rect 675 805 807 810
rect 2157 866 2289 871
rect 2157 810 2195 866
rect 2251 810 2289 866
rect 2157 805 2289 810
rect 3639 866 3771 871
rect 3639 810 3677 866
rect 3733 810 3771 866
rect 3639 805 3771 810
rect 5121 866 5253 871
rect 5121 810 5159 866
rect 5215 810 5253 866
rect 5121 805 5253 810
rect 6603 866 6735 871
rect 6603 810 6641 866
rect 6697 810 6735 866
rect 6603 805 6735 810
rect 8085 866 8217 871
rect 8085 810 8123 866
rect 8179 810 8217 866
rect 8085 805 8217 810
rect 9567 866 9699 871
rect 9567 810 9605 866
rect 9661 810 9699 866
rect 9567 805 9699 810
rect 11049 866 11181 871
rect 11049 810 11087 866
rect 11143 810 11181 866
rect 11049 805 11181 810
rect 12531 866 12663 871
rect 12531 810 12569 866
rect 12625 810 12663 866
rect 12531 805 12663 810
rect 14013 866 14145 871
rect 14013 810 14051 866
rect 14107 810 14145 866
rect 14013 805 14145 810
rect 15495 866 15627 871
rect 15495 810 15533 866
rect 15589 810 15627 866
rect 15495 805 15627 810
rect 16977 866 17109 871
rect 16977 810 17015 866
rect 17071 810 17109 866
rect 16977 805 17109 810
rect 18459 866 18591 871
rect 18459 810 18497 866
rect 18553 810 18591 866
rect 18459 805 18591 810
rect 19941 866 20073 871
rect 19941 810 19979 866
rect 20035 810 20073 866
rect 19941 805 20073 810
rect 21423 866 21555 871
rect 21423 810 21461 866
rect 21517 810 21555 866
rect 21423 805 21555 810
rect 22905 866 23037 871
rect 22905 810 22943 866
rect 22999 810 23037 866
rect 22905 805 23037 810
rect -39 338 93 341
rect 1443 338 1575 341
rect 2925 338 3057 341
rect 4407 338 4539 341
rect 5889 338 6021 341
rect 7371 338 7503 341
rect 8853 338 8985 341
rect 10335 338 10467 341
rect 11817 338 11949 341
rect 13299 338 13431 341
rect 14781 338 14913 341
rect 16263 338 16395 341
rect 17745 338 17877 341
rect 19227 338 19359 341
rect 20709 338 20841 341
rect 22191 338 22323 341
rect -39 336 23712 338
rect -39 280 -1 336
rect 55 280 1481 336
rect 1537 280 2963 336
rect 3019 280 4445 336
rect 4501 280 5927 336
rect 5983 280 7409 336
rect 7465 280 8891 336
rect 8947 280 10373 336
rect 10429 280 11855 336
rect 11911 280 13337 336
rect 13393 280 14819 336
rect 14875 280 16301 336
rect 16357 280 17783 336
rect 17839 280 19265 336
rect 19321 280 20747 336
rect 20803 280 22229 336
rect 22285 280 23712 336
rect -39 278 23712 280
rect -39 275 93 278
rect 1443 275 1575 278
rect 2925 275 3057 278
rect 4407 275 4539 278
rect 5889 275 6021 278
rect 7371 275 7503 278
rect 8853 275 8985 278
rect 10335 275 10467 278
rect 11817 275 11949 278
rect 13299 275 13431 278
rect 14781 275 14913 278
rect 16263 275 16395 278
rect 17745 275 17877 278
rect 19227 275 19359 278
rect 20709 275 20841 278
rect 22191 275 22323 278
rect 675 28 807 33
rect 675 -28 713 28
rect 769 -28 807 28
rect 675 -33 807 -28
rect 2157 28 2289 33
rect 2157 -28 2195 28
rect 2251 -28 2289 28
rect 2157 -33 2289 -28
rect 3639 28 3771 33
rect 3639 -28 3677 28
rect 3733 -28 3771 28
rect 3639 -33 3771 -28
rect 5121 28 5253 33
rect 5121 -28 5159 28
rect 5215 -28 5253 28
rect 5121 -33 5253 -28
rect 6603 28 6735 33
rect 6603 -28 6641 28
rect 6697 -28 6735 28
rect 6603 -33 6735 -28
rect 8085 28 8217 33
rect 8085 -28 8123 28
rect 8179 -28 8217 28
rect 8085 -33 8217 -28
rect 9567 28 9699 33
rect 9567 -28 9605 28
rect 9661 -28 9699 28
rect 9567 -33 9699 -28
rect 11049 28 11181 33
rect 11049 -28 11087 28
rect 11143 -28 11181 28
rect 11049 -33 11181 -28
rect 12531 28 12663 33
rect 12531 -28 12569 28
rect 12625 -28 12663 28
rect 12531 -33 12663 -28
rect 14013 28 14145 33
rect 14013 -28 14051 28
rect 14107 -28 14145 28
rect 14013 -33 14145 -28
rect 15495 28 15627 33
rect 15495 -28 15533 28
rect 15589 -28 15627 28
rect 15495 -33 15627 -28
rect 16977 28 17109 33
rect 16977 -28 17015 28
rect 17071 -28 17109 28
rect 16977 -33 17109 -28
rect 18459 28 18591 33
rect 18459 -28 18497 28
rect 18553 -28 18591 28
rect 18459 -33 18591 -28
rect 19941 28 20073 33
rect 19941 -28 19979 28
rect 20035 -28 20073 28
rect 19941 -33 20073 -28
rect 21423 28 21555 33
rect 21423 -28 21461 28
rect 21517 -28 21555 28
rect 21423 -33 21555 -28
rect 22905 28 23037 33
rect 22905 -28 22943 28
rect 22999 -28 23037 28
rect 22905 -33 23037 -28
use contact_18  contact_18_0
timestamp 1643678851
transform 1 0 22191 0 1 275
box 0 0 1 1
use contact_18  contact_18_1
timestamp 1643678851
transform 1 0 20709 0 1 275
box 0 0 1 1
use contact_18  contact_18_2
timestamp 1643678851
transform 1 0 19227 0 1 275
box 0 0 1 1
use contact_18  contact_18_3
timestamp 1643678851
transform 1 0 17745 0 1 275
box 0 0 1 1
use contact_18  contact_18_4
timestamp 1643678851
transform 1 0 16263 0 1 275
box 0 0 1 1
use contact_18  contact_18_5
timestamp 1643678851
transform 1 0 14781 0 1 275
box 0 0 1 1
use contact_18  contact_18_6
timestamp 1643678851
transform 1 0 13299 0 1 275
box 0 0 1 1
use contact_18  contact_18_7
timestamp 1643678851
transform 1 0 11817 0 1 275
box 0 0 1 1
use contact_18  contact_18_8
timestamp 1643678851
transform 1 0 10335 0 1 275
box 0 0 1 1
use contact_18  contact_18_9
timestamp 1643678851
transform 1 0 8853 0 1 275
box 0 0 1 1
use contact_18  contact_18_10
timestamp 1643678851
transform 1 0 7371 0 1 275
box 0 0 1 1
use contact_18  contact_18_11
timestamp 1643678851
transform 1 0 5889 0 1 275
box 0 0 1 1
use contact_18  contact_18_12
timestamp 1643678851
transform 1 0 4407 0 1 275
box 0 0 1 1
use contact_18  contact_18_13
timestamp 1643678851
transform 1 0 2925 0 1 275
box 0 0 1 1
use contact_18  contact_18_14
timestamp 1643678851
transform 1 0 1443 0 1 275
box 0 0 1 1
use contact_18  contact_18_15
timestamp 1643678851
transform 1 0 -39 0 1 275
box 0 0 1 1
use contact_18  contact_18_16
timestamp 1643678851
transform 1 0 22905 0 1 -33
box 0 0 1 1
use contact_17  contact_17_0
timestamp 1643678851
transform 1 0 22956 0 1 -15
box 0 0 1 1
use contact_18  contact_18_17
timestamp 1643678851
transform 1 0 22905 0 1 805
box 0 0 1 1
use contact_17  contact_17_1
timestamp 1643678851
transform 1 0 22956 0 1 823
box 0 0 1 1
use contact_18  contact_18_18
timestamp 1643678851
transform 1 0 21423 0 1 -33
box 0 0 1 1
use contact_17  contact_17_2
timestamp 1643678851
transform 1 0 21474 0 1 -15
box 0 0 1 1
use contact_18  contact_18_19
timestamp 1643678851
transform 1 0 21423 0 1 805
box 0 0 1 1
use contact_17  contact_17_3
timestamp 1643678851
transform 1 0 21474 0 1 823
box 0 0 1 1
use contact_18  contact_18_20
timestamp 1643678851
transform 1 0 19941 0 1 -33
box 0 0 1 1
use contact_17  contact_17_4
timestamp 1643678851
transform 1 0 19992 0 1 -15
box 0 0 1 1
use contact_18  contact_18_21
timestamp 1643678851
transform 1 0 19941 0 1 805
box 0 0 1 1
use contact_17  contact_17_5
timestamp 1643678851
transform 1 0 19992 0 1 823
box 0 0 1 1
use contact_18  contact_18_22
timestamp 1643678851
transform 1 0 18459 0 1 -33
box 0 0 1 1
use contact_17  contact_17_6
timestamp 1643678851
transform 1 0 18510 0 1 -15
box 0 0 1 1
use contact_18  contact_18_23
timestamp 1643678851
transform 1 0 18459 0 1 805
box 0 0 1 1
use contact_17  contact_17_7
timestamp 1643678851
transform 1 0 18510 0 1 823
box 0 0 1 1
use contact_18  contact_18_24
timestamp 1643678851
transform 1 0 16977 0 1 -33
box 0 0 1 1
use contact_17  contact_17_8
timestamp 1643678851
transform 1 0 17028 0 1 -15
box 0 0 1 1
use contact_18  contact_18_25
timestamp 1643678851
transform 1 0 16977 0 1 805
box 0 0 1 1
use contact_17  contact_17_9
timestamp 1643678851
transform 1 0 17028 0 1 823
box 0 0 1 1
use contact_18  contact_18_26
timestamp 1643678851
transform 1 0 15495 0 1 -33
box 0 0 1 1
use contact_17  contact_17_10
timestamp 1643678851
transform 1 0 15546 0 1 -15
box 0 0 1 1
use contact_18  contact_18_27
timestamp 1643678851
transform 1 0 15495 0 1 805
box 0 0 1 1
use contact_17  contact_17_11
timestamp 1643678851
transform 1 0 15546 0 1 823
box 0 0 1 1
use contact_18  contact_18_28
timestamp 1643678851
transform 1 0 14013 0 1 -33
box 0 0 1 1
use contact_17  contact_17_12
timestamp 1643678851
transform 1 0 14064 0 1 -15
box 0 0 1 1
use contact_18  contact_18_29
timestamp 1643678851
transform 1 0 14013 0 1 805
box 0 0 1 1
use contact_17  contact_17_13
timestamp 1643678851
transform 1 0 14064 0 1 823
box 0 0 1 1
use contact_18  contact_18_30
timestamp 1643678851
transform 1 0 12531 0 1 -33
box 0 0 1 1
use contact_17  contact_17_14
timestamp 1643678851
transform 1 0 12582 0 1 -15
box 0 0 1 1
use contact_18  contact_18_31
timestamp 1643678851
transform 1 0 12531 0 1 805
box 0 0 1 1
use contact_17  contact_17_15
timestamp 1643678851
transform 1 0 12582 0 1 823
box 0 0 1 1
use contact_18  contact_18_32
timestamp 1643678851
transform 1 0 11049 0 1 -33
box 0 0 1 1
use contact_17  contact_17_16
timestamp 1643678851
transform 1 0 11100 0 1 -15
box 0 0 1 1
use contact_18  contact_18_33
timestamp 1643678851
transform 1 0 11049 0 1 805
box 0 0 1 1
use contact_17  contact_17_17
timestamp 1643678851
transform 1 0 11100 0 1 823
box 0 0 1 1
use contact_18  contact_18_34
timestamp 1643678851
transform 1 0 9567 0 1 -33
box 0 0 1 1
use contact_17  contact_17_18
timestamp 1643678851
transform 1 0 9618 0 1 -15
box 0 0 1 1
use contact_18  contact_18_35
timestamp 1643678851
transform 1 0 9567 0 1 805
box 0 0 1 1
use contact_17  contact_17_19
timestamp 1643678851
transform 1 0 9618 0 1 823
box 0 0 1 1
use contact_18  contact_18_36
timestamp 1643678851
transform 1 0 8085 0 1 -33
box 0 0 1 1
use contact_17  contact_17_20
timestamp 1643678851
transform 1 0 8136 0 1 -15
box 0 0 1 1
use contact_18  contact_18_37
timestamp 1643678851
transform 1 0 8085 0 1 805
box 0 0 1 1
use contact_17  contact_17_21
timestamp 1643678851
transform 1 0 8136 0 1 823
box 0 0 1 1
use contact_18  contact_18_38
timestamp 1643678851
transform 1 0 6603 0 1 -33
box 0 0 1 1
use contact_17  contact_17_22
timestamp 1643678851
transform 1 0 6654 0 1 -15
box 0 0 1 1
use contact_18  contact_18_39
timestamp 1643678851
transform 1 0 6603 0 1 805
box 0 0 1 1
use contact_17  contact_17_23
timestamp 1643678851
transform 1 0 6654 0 1 823
box 0 0 1 1
use contact_18  contact_18_40
timestamp 1643678851
transform 1 0 5121 0 1 -33
box 0 0 1 1
use contact_17  contact_17_24
timestamp 1643678851
transform 1 0 5172 0 1 -15
box 0 0 1 1
use contact_18  contact_18_41
timestamp 1643678851
transform 1 0 5121 0 1 805
box 0 0 1 1
use contact_17  contact_17_25
timestamp 1643678851
transform 1 0 5172 0 1 823
box 0 0 1 1
use contact_18  contact_18_42
timestamp 1643678851
transform 1 0 3639 0 1 -33
box 0 0 1 1
use contact_17  contact_17_26
timestamp 1643678851
transform 1 0 3690 0 1 -15
box 0 0 1 1
use contact_18  contact_18_43
timestamp 1643678851
transform 1 0 3639 0 1 805
box 0 0 1 1
use contact_17  contact_17_27
timestamp 1643678851
transform 1 0 3690 0 1 823
box 0 0 1 1
use contact_18  contact_18_44
timestamp 1643678851
transform 1 0 2157 0 1 -33
box 0 0 1 1
use contact_17  contact_17_28
timestamp 1643678851
transform 1 0 2208 0 1 -15
box 0 0 1 1
use contact_18  contact_18_45
timestamp 1643678851
transform 1 0 2157 0 1 805
box 0 0 1 1
use contact_17  contact_17_29
timestamp 1643678851
transform 1 0 2208 0 1 823
box 0 0 1 1
use contact_18  contact_18_46
timestamp 1643678851
transform 1 0 675 0 1 -33
box 0 0 1 1
use contact_17  contact_17_30
timestamp 1643678851
transform 1 0 726 0 1 -15
box 0 0 1 1
use contact_18  contact_18_47
timestamp 1643678851
transform 1 0 675 0 1 805
box 0 0 1 1
use contact_17  contact_17_31
timestamp 1643678851
transform 1 0 726 0 1 823
box 0 0 1 1
use dff  dff_0
timestamp 1643678851
transform 1 0 22230 0 1 0
box 0 -42 1482 916
use dff  dff_1
timestamp 1643678851
transform 1 0 20748 0 1 0
box 0 -42 1482 916
use dff  dff_2
timestamp 1643678851
transform 1 0 19266 0 1 0
box 0 -42 1482 916
use dff  dff_3
timestamp 1643678851
transform 1 0 17784 0 1 0
box 0 -42 1482 916
use dff  dff_4
timestamp 1643678851
transform 1 0 16302 0 1 0
box 0 -42 1482 916
use dff  dff_5
timestamp 1643678851
transform 1 0 14820 0 1 0
box 0 -42 1482 916
use dff  dff_6
timestamp 1643678851
transform 1 0 13338 0 1 0
box 0 -42 1482 916
use dff  dff_7
timestamp 1643678851
transform 1 0 11856 0 1 0
box 0 -42 1482 916
use dff  dff_8
timestamp 1643678851
transform 1 0 10374 0 1 0
box 0 -42 1482 916
use dff  dff_9
timestamp 1643678851
transform 1 0 8892 0 1 0
box 0 -42 1482 916
use dff  dff_10
timestamp 1643678851
transform 1 0 7410 0 1 0
box 0 -42 1482 916
use dff  dff_11
timestamp 1643678851
transform 1 0 5928 0 1 0
box 0 -42 1482 916
use dff  dff_12
timestamp 1643678851
transform 1 0 4446 0 1 0
box 0 -42 1482 916
use dff  dff_13
timestamp 1643678851
transform 1 0 2964 0 1 0
box 0 -42 1482 916
use dff  dff_14
timestamp 1643678851
transform 1 0 1482 0 1 0
box 0 -42 1482 916
use dff  dff_15
timestamp 1643678851
transform 1 0 0 0 1 0
box 0 -42 1482 916
<< labels >>
rlabel metal3 s 15495 805 15627 871 4 vdd
rlabel metal3 s 675 805 807 871 4 vdd
rlabel metal3 s 3639 805 3771 871 4 vdd
rlabel metal3 s 19941 805 20073 871 4 vdd
rlabel metal3 s 22905 805 23037 871 4 vdd
rlabel metal3 s 6603 805 6735 871 4 vdd
rlabel metal3 s 5121 805 5253 871 4 vdd
rlabel metal3 s 8085 805 8217 871 4 vdd
rlabel metal3 s 9567 805 9699 871 4 vdd
rlabel metal3 s 16977 805 17109 871 4 vdd
rlabel metal3 s 11049 805 11181 871 4 vdd
rlabel metal3 s 2157 805 2289 871 4 vdd
rlabel metal3 s 21423 805 21555 871 4 vdd
rlabel metal3 s 12531 805 12663 871 4 vdd
rlabel metal3 s 14013 805 14145 871 4 vdd
rlabel metal3 s 18459 805 18591 871 4 vdd
rlabel metal3 s 22905 -33 23037 33 4 gnd
rlabel metal3 s 2157 -33 2289 33 4 gnd
rlabel metal3 s 675 -33 807 33 4 gnd
rlabel metal3 s 8085 -33 8217 33 4 gnd
rlabel metal3 s 12531 -33 12663 33 4 gnd
rlabel metal3 s 9567 -33 9699 33 4 gnd
rlabel metal3 s 18459 -33 18591 33 4 gnd
rlabel metal3 s 14013 -33 14145 33 4 gnd
rlabel metal3 s 19941 -33 20073 33 4 gnd
rlabel metal3 s 5121 -33 5253 33 4 gnd
rlabel metal3 s 6603 -33 6735 33 4 gnd
rlabel metal3 s 11049 -33 11181 33 4 gnd
rlabel metal3 s 16977 -33 17109 33 4 gnd
rlabel metal3 s 21423 -33 21555 33 4 gnd
rlabel metal3 s 3639 -33 3771 33 4 gnd
rlabel metal3 s 15495 -33 15627 33 4 gnd
rlabel metal2 s 180 232 234 260 4 din_0
rlabel metal2 s 1260 228 1314 256 4 dout_0
rlabel metal2 s 1662 232 1716 260 4 din_1
rlabel metal2 s 2742 228 2796 256 4 dout_1
rlabel metal2 s 3144 232 3198 260 4 din_2
rlabel metal2 s 4224 228 4278 256 4 dout_2
rlabel metal2 s 4626 232 4680 260 4 din_3
rlabel metal2 s 5706 228 5760 256 4 dout_3
rlabel metal2 s 6108 232 6162 260 4 din_4
rlabel metal2 s 7188 228 7242 256 4 dout_4
rlabel metal2 s 7590 232 7644 260 4 din_5
rlabel metal2 s 8670 228 8724 256 4 dout_5
rlabel metal2 s 9072 232 9126 260 4 din_6
rlabel metal2 s 10152 228 10206 256 4 dout_6
rlabel metal2 s 10554 232 10608 260 4 din_7
rlabel metal2 s 11634 228 11688 256 4 dout_7
rlabel metal2 s 12036 232 12090 260 4 din_8
rlabel metal2 s 13116 228 13170 256 4 dout_8
rlabel metal2 s 13518 232 13572 260 4 din_9
rlabel metal2 s 14598 228 14652 256 4 dout_9
rlabel metal2 s 15000 232 15054 260 4 din_10
rlabel metal2 s 16080 228 16134 256 4 dout_10
rlabel metal2 s 16482 232 16536 260 4 din_11
rlabel metal2 s 17562 228 17616 256 4 dout_11
rlabel metal2 s 17964 232 18018 260 4 din_12
rlabel metal2 s 19044 228 19098 256 4 dout_12
rlabel metal2 s 19446 232 19500 260 4 din_13
rlabel metal2 s 20526 228 20580 256 4 dout_13
rlabel metal2 s 20928 232 20982 260 4 din_14
rlabel metal2 s 22008 228 22062 256 4 dout_14
rlabel metal2 s 22410 232 22464 260 4 din_15
rlabel metal2 s 23490 228 23544 256 4 dout_15
rlabel metal3 s 0 278 23712 338 4 clk
<< properties >>
string FIXED_BBOX 22905 -33 23037 0
string GDS_FILE sram_0rw2r1w_16_128_sky130A.gds
string GDS_END 2172202
string GDS_START 2153088
<< end >>
