magic
tech sky130A
magscale 1 2
timestamp 1644951705
<< checkpaint >>
rect -1296 -1277 2312 2857
<< locali >>
rect 0 1523 1016 1557
rect 430 745 464 1279
rect 430 711 729 745
rect 827 711 861 745
rect 329 505 395 571
rect 196 381 262 447
rect 63 257 129 323
rect 0 -17 1016 17
use pinv  pinv_0
timestamp 1644951705
transform 1 0 648 0 1 0
box -36 -17 404 1597
use pnand3  pnand3_0
timestamp 1644951705
transform 1 0 0 0 1 0
box -36 -17 684 1597
<< labels >>
rlabel locali s 844 728 844 728 4 Z
rlabel locali s 96 290 96 290 4 A
rlabel locali s 229 414 229 414 4 B
rlabel locali s 362 538 362 538 4 C
rlabel locali s 508 0 508 0 4 gnd
rlabel locali s 508 1540 508 1540 4 vdd
<< properties >>
string FIXED_BBOX 0 0 1016 1540
string GDS_FILE sram_0rw2r1w_16_128_sky130A.gds
string GDS_END 1814272
string GDS_START 1813154
<< end >>
