magic
tech sky130A
magscale 1 2
timestamp 1644969367
<< checkpaint >>
rect -1143 -1263 50157 2310
<< metal1 >>
rect 221 954 227 1006
rect 279 954 285 1006
rect 493 954 499 1006
rect 551 954 557 1006
rect 1777 954 1783 1006
rect 1835 954 1841 1006
rect 2049 954 2055 1006
rect 2107 954 2113 1006
rect 3333 954 3339 1006
rect 3391 954 3397 1006
rect 3605 954 3611 1006
rect 3663 954 3669 1006
rect 4889 954 4895 1006
rect 4947 954 4953 1006
rect 5161 954 5167 1006
rect 5219 954 5225 1006
rect 6445 954 6451 1006
rect 6503 954 6509 1006
rect 6717 954 6723 1006
rect 6775 954 6781 1006
rect 8001 954 8007 1006
rect 8059 954 8065 1006
rect 8273 954 8279 1006
rect 8331 954 8337 1006
rect 9557 954 9563 1006
rect 9615 954 9621 1006
rect 9829 954 9835 1006
rect 9887 954 9893 1006
rect 11113 954 11119 1006
rect 11171 954 11177 1006
rect 11385 954 11391 1006
rect 11443 954 11449 1006
rect 12669 954 12675 1006
rect 12727 954 12733 1006
rect 12941 954 12947 1006
rect 12999 954 13005 1006
rect 14225 954 14231 1006
rect 14283 954 14289 1006
rect 14497 954 14503 1006
rect 14555 954 14561 1006
rect 15781 954 15787 1006
rect 15839 954 15845 1006
rect 16053 954 16059 1006
rect 16111 954 16117 1006
rect 17337 954 17343 1006
rect 17395 954 17401 1006
rect 17609 954 17615 1006
rect 17667 954 17673 1006
rect 18893 954 18899 1006
rect 18951 954 18957 1006
rect 19165 954 19171 1006
rect 19223 954 19229 1006
rect 20449 954 20455 1006
rect 20507 954 20513 1006
rect 20721 954 20727 1006
rect 20779 954 20785 1006
rect 22005 954 22011 1006
rect 22063 954 22069 1006
rect 22277 954 22283 1006
rect 22335 954 22341 1006
rect 23561 954 23567 1006
rect 23619 954 23625 1006
rect 23833 954 23839 1006
rect 23891 954 23897 1006
rect 25117 954 25123 1006
rect 25175 954 25181 1006
rect 25389 954 25395 1006
rect 25447 954 25453 1006
rect 26673 954 26679 1006
rect 26731 954 26737 1006
rect 26945 954 26951 1006
rect 27003 954 27009 1006
rect 28229 954 28235 1006
rect 28287 954 28293 1006
rect 28501 954 28507 1006
rect 28559 954 28565 1006
rect 29785 954 29791 1006
rect 29843 954 29849 1006
rect 30057 954 30063 1006
rect 30115 954 30121 1006
rect 31341 954 31347 1006
rect 31399 954 31405 1006
rect 31613 954 31619 1006
rect 31671 954 31677 1006
rect 32897 954 32903 1006
rect 32955 954 32961 1006
rect 33169 954 33175 1006
rect 33227 954 33233 1006
rect 34453 954 34459 1006
rect 34511 954 34517 1006
rect 34725 954 34731 1006
rect 34783 954 34789 1006
rect 36009 954 36015 1006
rect 36067 954 36073 1006
rect 36281 954 36287 1006
rect 36339 954 36345 1006
rect 37565 954 37571 1006
rect 37623 954 37629 1006
rect 37837 954 37843 1006
rect 37895 954 37901 1006
rect 39121 954 39127 1006
rect 39179 954 39185 1006
rect 39393 954 39399 1006
rect 39451 954 39457 1006
rect 40677 954 40683 1006
rect 40735 954 40741 1006
rect 40949 954 40955 1006
rect 41007 954 41013 1006
rect 42233 954 42239 1006
rect 42291 954 42297 1006
rect 42505 954 42511 1006
rect 42563 954 42569 1006
rect 43789 954 43795 1006
rect 43847 954 43853 1006
rect 44061 954 44067 1006
rect 44119 954 44125 1006
rect 45345 954 45351 1006
rect 45403 954 45409 1006
rect 45617 954 45623 1006
rect 45675 954 45681 1006
rect 46901 954 46907 1006
rect 46959 954 46965 1006
rect 47173 954 47179 1006
rect 47231 954 47237 1006
rect 48457 954 48463 1006
rect 48515 954 48521 1006
rect 48729 954 48735 1006
rect 48787 954 48793 1006
rect 221 8 227 60
rect 279 8 285 60
rect 493 8 499 60
rect 551 8 557 60
rect 1777 8 1783 60
rect 1835 8 1841 60
rect 2049 8 2055 60
rect 2107 8 2113 60
rect 3333 8 3339 60
rect 3391 8 3397 60
rect 3605 8 3611 60
rect 3663 8 3669 60
rect 4889 8 4895 60
rect 4947 8 4953 60
rect 5161 8 5167 60
rect 5219 8 5225 60
rect 6445 8 6451 60
rect 6503 8 6509 60
rect 6717 8 6723 60
rect 6775 8 6781 60
rect 8001 8 8007 60
rect 8059 8 8065 60
rect 8273 8 8279 60
rect 8331 8 8337 60
rect 9557 8 9563 60
rect 9615 8 9621 60
rect 9829 8 9835 60
rect 9887 8 9893 60
rect 11113 8 11119 60
rect 11171 8 11177 60
rect 11385 8 11391 60
rect 11443 8 11449 60
rect 12669 8 12675 60
rect 12727 8 12733 60
rect 12941 8 12947 60
rect 12999 8 13005 60
rect 14225 8 14231 60
rect 14283 8 14289 60
rect 14497 8 14503 60
rect 14555 8 14561 60
rect 15781 8 15787 60
rect 15839 8 15845 60
rect 16053 8 16059 60
rect 16111 8 16117 60
rect 17337 8 17343 60
rect 17395 8 17401 60
rect 17609 8 17615 60
rect 17667 8 17673 60
rect 18893 8 18899 60
rect 18951 8 18957 60
rect 19165 8 19171 60
rect 19223 8 19229 60
rect 20449 8 20455 60
rect 20507 8 20513 60
rect 20721 8 20727 60
rect 20779 8 20785 60
rect 22005 8 22011 60
rect 22063 8 22069 60
rect 22277 8 22283 60
rect 22335 8 22341 60
rect 23561 8 23567 60
rect 23619 8 23625 60
rect 23833 8 23839 60
rect 23891 8 23897 60
rect 25117 8 25123 60
rect 25175 8 25181 60
rect 25389 8 25395 60
rect 25447 8 25453 60
rect 26673 8 26679 60
rect 26731 8 26737 60
rect 26945 8 26951 60
rect 27003 8 27009 60
rect 28229 8 28235 60
rect 28287 8 28293 60
rect 28501 8 28507 60
rect 28559 8 28565 60
rect 29785 8 29791 60
rect 29843 8 29849 60
rect 30057 8 30063 60
rect 30115 8 30121 60
rect 31341 8 31347 60
rect 31399 8 31405 60
rect 31613 8 31619 60
rect 31671 8 31677 60
rect 32897 8 32903 60
rect 32955 8 32961 60
rect 33169 8 33175 60
rect 33227 8 33233 60
rect 34453 8 34459 60
rect 34511 8 34517 60
rect 34725 8 34731 60
rect 34783 8 34789 60
rect 36009 8 36015 60
rect 36067 8 36073 60
rect 36281 8 36287 60
rect 36339 8 36345 60
rect 37565 8 37571 60
rect 37623 8 37629 60
rect 37837 8 37843 60
rect 37895 8 37901 60
rect 39121 8 39127 60
rect 39179 8 39185 60
rect 39393 8 39399 60
rect 39451 8 39457 60
rect 40677 8 40683 60
rect 40735 8 40741 60
rect 40949 8 40955 60
rect 41007 8 41013 60
rect 42233 8 42239 60
rect 42291 8 42297 60
rect 42505 8 42511 60
rect 42563 8 42569 60
rect 43789 8 43795 60
rect 43847 8 43853 60
rect 44061 8 44067 60
rect 44119 8 44125 60
rect 45345 8 45351 60
rect 45403 8 45409 60
rect 45617 8 45623 60
rect 45675 8 45681 60
rect 46901 8 46907 60
rect 46959 8 46965 60
rect 47173 8 47179 60
rect 47231 8 47237 60
rect 48457 8 48463 60
rect 48515 8 48521 60
rect 48729 8 48735 60
rect 48787 8 48793 60
<< via1 >>
rect 227 954 279 1006
rect 499 954 551 1006
rect 1783 954 1835 1006
rect 2055 954 2107 1006
rect 3339 954 3391 1006
rect 3611 954 3663 1006
rect 4895 954 4947 1006
rect 5167 954 5219 1006
rect 6451 954 6503 1006
rect 6723 954 6775 1006
rect 8007 954 8059 1006
rect 8279 954 8331 1006
rect 9563 954 9615 1006
rect 9835 954 9887 1006
rect 11119 954 11171 1006
rect 11391 954 11443 1006
rect 12675 954 12727 1006
rect 12947 954 12999 1006
rect 14231 954 14283 1006
rect 14503 954 14555 1006
rect 15787 954 15839 1006
rect 16059 954 16111 1006
rect 17343 954 17395 1006
rect 17615 954 17667 1006
rect 18899 954 18951 1006
rect 19171 954 19223 1006
rect 20455 954 20507 1006
rect 20727 954 20779 1006
rect 22011 954 22063 1006
rect 22283 954 22335 1006
rect 23567 954 23619 1006
rect 23839 954 23891 1006
rect 25123 954 25175 1006
rect 25395 954 25447 1006
rect 26679 954 26731 1006
rect 26951 954 27003 1006
rect 28235 954 28287 1006
rect 28507 954 28559 1006
rect 29791 954 29843 1006
rect 30063 954 30115 1006
rect 31347 954 31399 1006
rect 31619 954 31671 1006
rect 32903 954 32955 1006
rect 33175 954 33227 1006
rect 34459 954 34511 1006
rect 34731 954 34783 1006
rect 36015 954 36067 1006
rect 36287 954 36339 1006
rect 37571 954 37623 1006
rect 37843 954 37895 1006
rect 39127 954 39179 1006
rect 39399 954 39451 1006
rect 40683 954 40735 1006
rect 40955 954 41007 1006
rect 42239 954 42291 1006
rect 42511 954 42563 1006
rect 43795 954 43847 1006
rect 44067 954 44119 1006
rect 45351 954 45403 1006
rect 45623 954 45675 1006
rect 46907 954 46959 1006
rect 47179 954 47231 1006
rect 48463 954 48515 1006
rect 48735 954 48787 1006
rect 227 8 279 60
rect 499 8 551 60
rect 1783 8 1835 60
rect 2055 8 2107 60
rect 3339 8 3391 60
rect 3611 8 3663 60
rect 4895 8 4947 60
rect 5167 8 5219 60
rect 6451 8 6503 60
rect 6723 8 6775 60
rect 8007 8 8059 60
rect 8279 8 8331 60
rect 9563 8 9615 60
rect 9835 8 9887 60
rect 11119 8 11171 60
rect 11391 8 11443 60
rect 12675 8 12727 60
rect 12947 8 12999 60
rect 14231 8 14283 60
rect 14503 8 14555 60
rect 15787 8 15839 60
rect 16059 8 16111 60
rect 17343 8 17395 60
rect 17615 8 17667 60
rect 18899 8 18951 60
rect 19171 8 19223 60
rect 20455 8 20507 60
rect 20727 8 20779 60
rect 22011 8 22063 60
rect 22283 8 22335 60
rect 23567 8 23619 60
rect 23839 8 23891 60
rect 25123 8 25175 60
rect 25395 8 25447 60
rect 26679 8 26731 60
rect 26951 8 27003 60
rect 28235 8 28287 60
rect 28507 8 28559 60
rect 29791 8 29843 60
rect 30063 8 30115 60
rect 31347 8 31399 60
rect 31619 8 31671 60
rect 32903 8 32955 60
rect 33175 8 33227 60
rect 34459 8 34511 60
rect 34731 8 34783 60
rect 36015 8 36067 60
rect 36287 8 36339 60
rect 37571 8 37623 60
rect 37843 8 37895 60
rect 39127 8 39179 60
rect 39399 8 39451 60
rect 40683 8 40735 60
rect 40955 8 41007 60
rect 42239 8 42291 60
rect 42511 8 42563 60
rect 43795 8 43847 60
rect 44067 8 44119 60
rect 45351 8 45403 60
rect 45623 8 45675 60
rect 46907 8 46959 60
rect 47179 8 47231 60
rect 48463 8 48515 60
rect 48735 8 48787 60
<< metal2 >>
rect 225 1008 281 1017
rect 225 943 281 952
rect 497 1008 553 1017
rect 497 943 553 952
rect 1781 1008 1837 1017
rect 1781 943 1837 952
rect 2053 1008 2109 1017
rect 2053 943 2109 952
rect 3337 1008 3393 1017
rect 3337 943 3393 952
rect 3609 1008 3665 1017
rect 3609 943 3665 952
rect 4893 1008 4949 1017
rect 4893 943 4949 952
rect 5165 1008 5221 1017
rect 5165 943 5221 952
rect 6449 1008 6505 1017
rect 6449 943 6505 952
rect 6721 1008 6777 1017
rect 6721 943 6777 952
rect 8005 1008 8061 1017
rect 8005 943 8061 952
rect 8277 1008 8333 1017
rect 8277 943 8333 952
rect 9561 1008 9617 1017
rect 9561 943 9617 952
rect 9833 1008 9889 1017
rect 9833 943 9889 952
rect 11117 1008 11173 1017
rect 11117 943 11173 952
rect 11389 1008 11445 1017
rect 11389 943 11445 952
rect 12673 1008 12729 1017
rect 12673 943 12729 952
rect 12945 1008 13001 1017
rect 12945 943 13001 952
rect 14229 1008 14285 1017
rect 14229 943 14285 952
rect 14501 1008 14557 1017
rect 14501 943 14557 952
rect 15785 1008 15841 1017
rect 15785 943 15841 952
rect 16057 1008 16113 1017
rect 16057 943 16113 952
rect 17341 1008 17397 1017
rect 17341 943 17397 952
rect 17613 1008 17669 1017
rect 17613 943 17669 952
rect 18897 1008 18953 1017
rect 18897 943 18953 952
rect 19169 1008 19225 1017
rect 19169 943 19225 952
rect 20453 1008 20509 1017
rect 20453 943 20509 952
rect 20725 1008 20781 1017
rect 20725 943 20781 952
rect 22009 1008 22065 1017
rect 22009 943 22065 952
rect 22281 1008 22337 1017
rect 22281 943 22337 952
rect 23565 1008 23621 1017
rect 23565 943 23621 952
rect 23837 1008 23893 1017
rect 23837 943 23893 952
rect 25121 1008 25177 1017
rect 25121 943 25177 952
rect 25393 1008 25449 1017
rect 25393 943 25449 952
rect 26677 1008 26733 1017
rect 26677 943 26733 952
rect 26949 1008 27005 1017
rect 26949 943 27005 952
rect 28233 1008 28289 1017
rect 28233 943 28289 952
rect 28505 1008 28561 1017
rect 28505 943 28561 952
rect 29789 1008 29845 1017
rect 29789 943 29845 952
rect 30061 1008 30117 1017
rect 30061 943 30117 952
rect 31345 1008 31401 1017
rect 31345 943 31401 952
rect 31617 1008 31673 1017
rect 31617 943 31673 952
rect 32901 1008 32957 1017
rect 32901 943 32957 952
rect 33173 1008 33229 1017
rect 33173 943 33229 952
rect 34457 1008 34513 1017
rect 34457 943 34513 952
rect 34729 1008 34785 1017
rect 34729 943 34785 952
rect 36013 1008 36069 1017
rect 36013 943 36069 952
rect 36285 1008 36341 1017
rect 36285 943 36341 952
rect 37569 1008 37625 1017
rect 37569 943 37625 952
rect 37841 1008 37897 1017
rect 37841 943 37897 952
rect 39125 1008 39181 1017
rect 39125 943 39181 952
rect 39397 1008 39453 1017
rect 39397 943 39453 952
rect 40681 1008 40737 1017
rect 40681 943 40737 952
rect 40953 1008 41009 1017
rect 40953 943 41009 952
rect 42237 1008 42293 1017
rect 42237 943 42293 952
rect 42509 1008 42565 1017
rect 42509 943 42565 952
rect 43793 1008 43849 1017
rect 43793 943 43849 952
rect 44065 1008 44121 1017
rect 44065 943 44121 952
rect 45349 1008 45405 1017
rect 45349 943 45405 952
rect 45621 1008 45677 1017
rect 45621 943 45677 952
rect 46905 1008 46961 1017
rect 46905 943 46961 952
rect 47177 1008 47233 1017
rect 47177 943 47233 952
rect 48461 1008 48517 1017
rect 48461 943 48517 952
rect 48733 1008 48789 1017
rect 48733 943 48789 952
rect 131 0 159 240
rect 225 62 281 71
rect 225 -3 281 6
rect 319 0 347 240
rect 403 0 431 240
rect 497 62 553 71
rect 497 -3 553 6
rect 591 0 619 240
rect 1687 0 1715 240
rect 1781 62 1837 71
rect 1781 -3 1837 6
rect 1875 0 1903 240
rect 1959 0 1987 240
rect 2053 62 2109 71
rect 2053 -3 2109 6
rect 2147 0 2175 240
rect 3243 0 3271 240
rect 3337 62 3393 71
rect 3337 -3 3393 6
rect 3431 0 3459 240
rect 3515 0 3543 240
rect 3609 62 3665 71
rect 3609 -3 3665 6
rect 3703 0 3731 240
rect 4799 0 4827 240
rect 4893 62 4949 71
rect 4893 -3 4949 6
rect 4987 0 5015 240
rect 5071 0 5099 240
rect 5165 62 5221 71
rect 5165 -3 5221 6
rect 5259 0 5287 240
rect 6355 0 6383 240
rect 6449 62 6505 71
rect 6449 -3 6505 6
rect 6543 0 6571 240
rect 6627 0 6655 240
rect 6721 62 6777 71
rect 6721 -3 6777 6
rect 6815 0 6843 240
rect 7911 0 7939 240
rect 8005 62 8061 71
rect 8005 -3 8061 6
rect 8099 0 8127 240
rect 8183 0 8211 240
rect 8277 62 8333 71
rect 8277 -3 8333 6
rect 8371 0 8399 240
rect 9467 0 9495 240
rect 9561 62 9617 71
rect 9561 -3 9617 6
rect 9655 0 9683 240
rect 9739 0 9767 240
rect 9833 62 9889 71
rect 9833 -3 9889 6
rect 9927 0 9955 240
rect 11023 0 11051 240
rect 11117 62 11173 71
rect 11117 -3 11173 6
rect 11211 0 11239 240
rect 11295 0 11323 240
rect 11389 62 11445 71
rect 11389 -3 11445 6
rect 11483 0 11511 240
rect 12579 0 12607 240
rect 12673 62 12729 71
rect 12673 -3 12729 6
rect 12767 0 12795 240
rect 12851 0 12879 240
rect 12945 62 13001 71
rect 12945 -3 13001 6
rect 13039 0 13067 240
rect 14135 0 14163 240
rect 14229 62 14285 71
rect 14229 -3 14285 6
rect 14323 0 14351 240
rect 14407 0 14435 240
rect 14501 62 14557 71
rect 14501 -3 14557 6
rect 14595 0 14623 240
rect 15691 0 15719 240
rect 15785 62 15841 71
rect 15785 -3 15841 6
rect 15879 0 15907 240
rect 15963 0 15991 240
rect 16057 62 16113 71
rect 16057 -3 16113 6
rect 16151 0 16179 240
rect 17247 0 17275 240
rect 17341 62 17397 71
rect 17341 -3 17397 6
rect 17435 0 17463 240
rect 17519 0 17547 240
rect 17613 62 17669 71
rect 17613 -3 17669 6
rect 17707 0 17735 240
rect 18803 0 18831 240
rect 18897 62 18953 71
rect 18897 -3 18953 6
rect 18991 0 19019 240
rect 19075 0 19103 240
rect 19169 62 19225 71
rect 19169 -3 19225 6
rect 19263 0 19291 240
rect 20359 0 20387 240
rect 20453 62 20509 71
rect 20453 -3 20509 6
rect 20547 0 20575 240
rect 20631 0 20659 240
rect 20725 62 20781 71
rect 20725 -3 20781 6
rect 20819 0 20847 240
rect 21915 0 21943 240
rect 22009 62 22065 71
rect 22009 -3 22065 6
rect 22103 0 22131 240
rect 22187 0 22215 240
rect 22281 62 22337 71
rect 22281 -3 22337 6
rect 22375 0 22403 240
rect 23471 0 23499 240
rect 23565 62 23621 71
rect 23565 -3 23621 6
rect 23659 0 23687 240
rect 23743 0 23771 240
rect 23837 62 23893 71
rect 23837 -3 23893 6
rect 23931 0 23959 240
rect 25027 0 25055 240
rect 25121 62 25177 71
rect 25121 -3 25177 6
rect 25215 0 25243 240
rect 25299 0 25327 240
rect 25393 62 25449 71
rect 25393 -3 25449 6
rect 25487 0 25515 240
rect 26583 0 26611 240
rect 26677 62 26733 71
rect 26677 -3 26733 6
rect 26771 0 26799 240
rect 26855 0 26883 240
rect 26949 62 27005 71
rect 26949 -3 27005 6
rect 27043 0 27071 240
rect 28139 0 28167 240
rect 28233 62 28289 71
rect 28233 -3 28289 6
rect 28327 0 28355 240
rect 28411 0 28439 240
rect 28505 62 28561 71
rect 28505 -3 28561 6
rect 28599 0 28627 240
rect 29695 0 29723 240
rect 29789 62 29845 71
rect 29789 -3 29845 6
rect 29883 0 29911 240
rect 29967 0 29995 240
rect 30061 62 30117 71
rect 30061 -3 30117 6
rect 30155 0 30183 240
rect 31251 0 31279 240
rect 31345 62 31401 71
rect 31345 -3 31401 6
rect 31439 0 31467 240
rect 31523 0 31551 240
rect 31617 62 31673 71
rect 31617 -3 31673 6
rect 31711 0 31739 240
rect 32807 0 32835 240
rect 32901 62 32957 71
rect 32901 -3 32957 6
rect 32995 0 33023 240
rect 33079 0 33107 240
rect 33173 62 33229 71
rect 33173 -3 33229 6
rect 33267 0 33295 240
rect 34363 0 34391 240
rect 34457 62 34513 71
rect 34457 -3 34513 6
rect 34551 0 34579 240
rect 34635 0 34663 240
rect 34729 62 34785 71
rect 34729 -3 34785 6
rect 34823 0 34851 240
rect 35919 0 35947 240
rect 36013 62 36069 71
rect 36013 -3 36069 6
rect 36107 0 36135 240
rect 36191 0 36219 240
rect 36285 62 36341 71
rect 36285 -3 36341 6
rect 36379 0 36407 240
rect 37475 0 37503 240
rect 37569 62 37625 71
rect 37569 -3 37625 6
rect 37663 0 37691 240
rect 37747 0 37775 240
rect 37841 62 37897 71
rect 37841 -3 37897 6
rect 37935 0 37963 240
rect 39031 0 39059 240
rect 39125 62 39181 71
rect 39125 -3 39181 6
rect 39219 0 39247 240
rect 39303 0 39331 240
rect 39397 62 39453 71
rect 39397 -3 39453 6
rect 39491 0 39519 240
rect 40587 0 40615 240
rect 40681 62 40737 71
rect 40681 -3 40737 6
rect 40775 0 40803 240
rect 40859 0 40887 240
rect 40953 62 41009 71
rect 40953 -3 41009 6
rect 41047 0 41075 240
rect 42143 0 42171 240
rect 42237 62 42293 71
rect 42237 -3 42293 6
rect 42331 0 42359 240
rect 42415 0 42443 240
rect 42509 62 42565 71
rect 42509 -3 42565 6
rect 42603 0 42631 240
rect 43699 0 43727 240
rect 43793 62 43849 71
rect 43793 -3 43849 6
rect 43887 0 43915 240
rect 43971 0 43999 240
rect 44065 62 44121 71
rect 44065 -3 44121 6
rect 44159 0 44187 240
rect 45255 0 45283 240
rect 45349 62 45405 71
rect 45349 -3 45405 6
rect 45443 0 45471 240
rect 45527 0 45555 240
rect 45621 62 45677 71
rect 45621 -3 45677 6
rect 45715 0 45743 240
rect 46811 0 46839 240
rect 46905 62 46961 71
rect 46905 -3 46961 6
rect 46999 0 47027 240
rect 47083 0 47111 240
rect 47177 62 47233 71
rect 47177 -3 47233 6
rect 47271 0 47299 240
rect 48367 0 48395 240
rect 48461 62 48517 71
rect 48461 -3 48517 6
rect 48555 0 48583 240
rect 48639 0 48667 240
rect 48733 62 48789 71
rect 48733 -3 48789 6
rect 48827 0 48855 240
<< via2 >>
rect 225 1006 281 1008
rect 225 954 227 1006
rect 227 954 279 1006
rect 279 954 281 1006
rect 225 952 281 954
rect 497 1006 553 1008
rect 497 954 499 1006
rect 499 954 551 1006
rect 551 954 553 1006
rect 497 952 553 954
rect 1781 1006 1837 1008
rect 1781 954 1783 1006
rect 1783 954 1835 1006
rect 1835 954 1837 1006
rect 1781 952 1837 954
rect 2053 1006 2109 1008
rect 2053 954 2055 1006
rect 2055 954 2107 1006
rect 2107 954 2109 1006
rect 2053 952 2109 954
rect 3337 1006 3393 1008
rect 3337 954 3339 1006
rect 3339 954 3391 1006
rect 3391 954 3393 1006
rect 3337 952 3393 954
rect 3609 1006 3665 1008
rect 3609 954 3611 1006
rect 3611 954 3663 1006
rect 3663 954 3665 1006
rect 3609 952 3665 954
rect 4893 1006 4949 1008
rect 4893 954 4895 1006
rect 4895 954 4947 1006
rect 4947 954 4949 1006
rect 4893 952 4949 954
rect 5165 1006 5221 1008
rect 5165 954 5167 1006
rect 5167 954 5219 1006
rect 5219 954 5221 1006
rect 5165 952 5221 954
rect 6449 1006 6505 1008
rect 6449 954 6451 1006
rect 6451 954 6503 1006
rect 6503 954 6505 1006
rect 6449 952 6505 954
rect 6721 1006 6777 1008
rect 6721 954 6723 1006
rect 6723 954 6775 1006
rect 6775 954 6777 1006
rect 6721 952 6777 954
rect 8005 1006 8061 1008
rect 8005 954 8007 1006
rect 8007 954 8059 1006
rect 8059 954 8061 1006
rect 8005 952 8061 954
rect 8277 1006 8333 1008
rect 8277 954 8279 1006
rect 8279 954 8331 1006
rect 8331 954 8333 1006
rect 8277 952 8333 954
rect 9561 1006 9617 1008
rect 9561 954 9563 1006
rect 9563 954 9615 1006
rect 9615 954 9617 1006
rect 9561 952 9617 954
rect 9833 1006 9889 1008
rect 9833 954 9835 1006
rect 9835 954 9887 1006
rect 9887 954 9889 1006
rect 9833 952 9889 954
rect 11117 1006 11173 1008
rect 11117 954 11119 1006
rect 11119 954 11171 1006
rect 11171 954 11173 1006
rect 11117 952 11173 954
rect 11389 1006 11445 1008
rect 11389 954 11391 1006
rect 11391 954 11443 1006
rect 11443 954 11445 1006
rect 11389 952 11445 954
rect 12673 1006 12729 1008
rect 12673 954 12675 1006
rect 12675 954 12727 1006
rect 12727 954 12729 1006
rect 12673 952 12729 954
rect 12945 1006 13001 1008
rect 12945 954 12947 1006
rect 12947 954 12999 1006
rect 12999 954 13001 1006
rect 12945 952 13001 954
rect 14229 1006 14285 1008
rect 14229 954 14231 1006
rect 14231 954 14283 1006
rect 14283 954 14285 1006
rect 14229 952 14285 954
rect 14501 1006 14557 1008
rect 14501 954 14503 1006
rect 14503 954 14555 1006
rect 14555 954 14557 1006
rect 14501 952 14557 954
rect 15785 1006 15841 1008
rect 15785 954 15787 1006
rect 15787 954 15839 1006
rect 15839 954 15841 1006
rect 15785 952 15841 954
rect 16057 1006 16113 1008
rect 16057 954 16059 1006
rect 16059 954 16111 1006
rect 16111 954 16113 1006
rect 16057 952 16113 954
rect 17341 1006 17397 1008
rect 17341 954 17343 1006
rect 17343 954 17395 1006
rect 17395 954 17397 1006
rect 17341 952 17397 954
rect 17613 1006 17669 1008
rect 17613 954 17615 1006
rect 17615 954 17667 1006
rect 17667 954 17669 1006
rect 17613 952 17669 954
rect 18897 1006 18953 1008
rect 18897 954 18899 1006
rect 18899 954 18951 1006
rect 18951 954 18953 1006
rect 18897 952 18953 954
rect 19169 1006 19225 1008
rect 19169 954 19171 1006
rect 19171 954 19223 1006
rect 19223 954 19225 1006
rect 19169 952 19225 954
rect 20453 1006 20509 1008
rect 20453 954 20455 1006
rect 20455 954 20507 1006
rect 20507 954 20509 1006
rect 20453 952 20509 954
rect 20725 1006 20781 1008
rect 20725 954 20727 1006
rect 20727 954 20779 1006
rect 20779 954 20781 1006
rect 20725 952 20781 954
rect 22009 1006 22065 1008
rect 22009 954 22011 1006
rect 22011 954 22063 1006
rect 22063 954 22065 1006
rect 22009 952 22065 954
rect 22281 1006 22337 1008
rect 22281 954 22283 1006
rect 22283 954 22335 1006
rect 22335 954 22337 1006
rect 22281 952 22337 954
rect 23565 1006 23621 1008
rect 23565 954 23567 1006
rect 23567 954 23619 1006
rect 23619 954 23621 1006
rect 23565 952 23621 954
rect 23837 1006 23893 1008
rect 23837 954 23839 1006
rect 23839 954 23891 1006
rect 23891 954 23893 1006
rect 23837 952 23893 954
rect 25121 1006 25177 1008
rect 25121 954 25123 1006
rect 25123 954 25175 1006
rect 25175 954 25177 1006
rect 25121 952 25177 954
rect 25393 1006 25449 1008
rect 25393 954 25395 1006
rect 25395 954 25447 1006
rect 25447 954 25449 1006
rect 25393 952 25449 954
rect 26677 1006 26733 1008
rect 26677 954 26679 1006
rect 26679 954 26731 1006
rect 26731 954 26733 1006
rect 26677 952 26733 954
rect 26949 1006 27005 1008
rect 26949 954 26951 1006
rect 26951 954 27003 1006
rect 27003 954 27005 1006
rect 26949 952 27005 954
rect 28233 1006 28289 1008
rect 28233 954 28235 1006
rect 28235 954 28287 1006
rect 28287 954 28289 1006
rect 28233 952 28289 954
rect 28505 1006 28561 1008
rect 28505 954 28507 1006
rect 28507 954 28559 1006
rect 28559 954 28561 1006
rect 28505 952 28561 954
rect 29789 1006 29845 1008
rect 29789 954 29791 1006
rect 29791 954 29843 1006
rect 29843 954 29845 1006
rect 29789 952 29845 954
rect 30061 1006 30117 1008
rect 30061 954 30063 1006
rect 30063 954 30115 1006
rect 30115 954 30117 1006
rect 30061 952 30117 954
rect 31345 1006 31401 1008
rect 31345 954 31347 1006
rect 31347 954 31399 1006
rect 31399 954 31401 1006
rect 31345 952 31401 954
rect 31617 1006 31673 1008
rect 31617 954 31619 1006
rect 31619 954 31671 1006
rect 31671 954 31673 1006
rect 31617 952 31673 954
rect 32901 1006 32957 1008
rect 32901 954 32903 1006
rect 32903 954 32955 1006
rect 32955 954 32957 1006
rect 32901 952 32957 954
rect 33173 1006 33229 1008
rect 33173 954 33175 1006
rect 33175 954 33227 1006
rect 33227 954 33229 1006
rect 33173 952 33229 954
rect 34457 1006 34513 1008
rect 34457 954 34459 1006
rect 34459 954 34511 1006
rect 34511 954 34513 1006
rect 34457 952 34513 954
rect 34729 1006 34785 1008
rect 34729 954 34731 1006
rect 34731 954 34783 1006
rect 34783 954 34785 1006
rect 34729 952 34785 954
rect 36013 1006 36069 1008
rect 36013 954 36015 1006
rect 36015 954 36067 1006
rect 36067 954 36069 1006
rect 36013 952 36069 954
rect 36285 1006 36341 1008
rect 36285 954 36287 1006
rect 36287 954 36339 1006
rect 36339 954 36341 1006
rect 36285 952 36341 954
rect 37569 1006 37625 1008
rect 37569 954 37571 1006
rect 37571 954 37623 1006
rect 37623 954 37625 1006
rect 37569 952 37625 954
rect 37841 1006 37897 1008
rect 37841 954 37843 1006
rect 37843 954 37895 1006
rect 37895 954 37897 1006
rect 37841 952 37897 954
rect 39125 1006 39181 1008
rect 39125 954 39127 1006
rect 39127 954 39179 1006
rect 39179 954 39181 1006
rect 39125 952 39181 954
rect 39397 1006 39453 1008
rect 39397 954 39399 1006
rect 39399 954 39451 1006
rect 39451 954 39453 1006
rect 39397 952 39453 954
rect 40681 1006 40737 1008
rect 40681 954 40683 1006
rect 40683 954 40735 1006
rect 40735 954 40737 1006
rect 40681 952 40737 954
rect 40953 1006 41009 1008
rect 40953 954 40955 1006
rect 40955 954 41007 1006
rect 41007 954 41009 1006
rect 40953 952 41009 954
rect 42237 1006 42293 1008
rect 42237 954 42239 1006
rect 42239 954 42291 1006
rect 42291 954 42293 1006
rect 42237 952 42293 954
rect 42509 1006 42565 1008
rect 42509 954 42511 1006
rect 42511 954 42563 1006
rect 42563 954 42565 1006
rect 42509 952 42565 954
rect 43793 1006 43849 1008
rect 43793 954 43795 1006
rect 43795 954 43847 1006
rect 43847 954 43849 1006
rect 43793 952 43849 954
rect 44065 1006 44121 1008
rect 44065 954 44067 1006
rect 44067 954 44119 1006
rect 44119 954 44121 1006
rect 44065 952 44121 954
rect 45349 1006 45405 1008
rect 45349 954 45351 1006
rect 45351 954 45403 1006
rect 45403 954 45405 1006
rect 45349 952 45405 954
rect 45621 1006 45677 1008
rect 45621 954 45623 1006
rect 45623 954 45675 1006
rect 45675 954 45677 1006
rect 45621 952 45677 954
rect 46905 1006 46961 1008
rect 46905 954 46907 1006
rect 46907 954 46959 1006
rect 46959 954 46961 1006
rect 46905 952 46961 954
rect 47177 1006 47233 1008
rect 47177 954 47179 1006
rect 47179 954 47231 1006
rect 47231 954 47233 1006
rect 47177 952 47233 954
rect 48461 1006 48517 1008
rect 48461 954 48463 1006
rect 48463 954 48515 1006
rect 48515 954 48517 1006
rect 48461 952 48517 954
rect 48733 1006 48789 1008
rect 48733 954 48735 1006
rect 48735 954 48787 1006
rect 48787 954 48789 1006
rect 48733 952 48789 954
rect 225 60 281 62
rect 225 8 227 60
rect 227 8 279 60
rect 279 8 281 60
rect 225 6 281 8
rect 497 60 553 62
rect 497 8 499 60
rect 499 8 551 60
rect 551 8 553 60
rect 497 6 553 8
rect 1781 60 1837 62
rect 1781 8 1783 60
rect 1783 8 1835 60
rect 1835 8 1837 60
rect 1781 6 1837 8
rect 2053 60 2109 62
rect 2053 8 2055 60
rect 2055 8 2107 60
rect 2107 8 2109 60
rect 2053 6 2109 8
rect 3337 60 3393 62
rect 3337 8 3339 60
rect 3339 8 3391 60
rect 3391 8 3393 60
rect 3337 6 3393 8
rect 3609 60 3665 62
rect 3609 8 3611 60
rect 3611 8 3663 60
rect 3663 8 3665 60
rect 3609 6 3665 8
rect 4893 60 4949 62
rect 4893 8 4895 60
rect 4895 8 4947 60
rect 4947 8 4949 60
rect 4893 6 4949 8
rect 5165 60 5221 62
rect 5165 8 5167 60
rect 5167 8 5219 60
rect 5219 8 5221 60
rect 5165 6 5221 8
rect 6449 60 6505 62
rect 6449 8 6451 60
rect 6451 8 6503 60
rect 6503 8 6505 60
rect 6449 6 6505 8
rect 6721 60 6777 62
rect 6721 8 6723 60
rect 6723 8 6775 60
rect 6775 8 6777 60
rect 6721 6 6777 8
rect 8005 60 8061 62
rect 8005 8 8007 60
rect 8007 8 8059 60
rect 8059 8 8061 60
rect 8005 6 8061 8
rect 8277 60 8333 62
rect 8277 8 8279 60
rect 8279 8 8331 60
rect 8331 8 8333 60
rect 8277 6 8333 8
rect 9561 60 9617 62
rect 9561 8 9563 60
rect 9563 8 9615 60
rect 9615 8 9617 60
rect 9561 6 9617 8
rect 9833 60 9889 62
rect 9833 8 9835 60
rect 9835 8 9887 60
rect 9887 8 9889 60
rect 9833 6 9889 8
rect 11117 60 11173 62
rect 11117 8 11119 60
rect 11119 8 11171 60
rect 11171 8 11173 60
rect 11117 6 11173 8
rect 11389 60 11445 62
rect 11389 8 11391 60
rect 11391 8 11443 60
rect 11443 8 11445 60
rect 11389 6 11445 8
rect 12673 60 12729 62
rect 12673 8 12675 60
rect 12675 8 12727 60
rect 12727 8 12729 60
rect 12673 6 12729 8
rect 12945 60 13001 62
rect 12945 8 12947 60
rect 12947 8 12999 60
rect 12999 8 13001 60
rect 12945 6 13001 8
rect 14229 60 14285 62
rect 14229 8 14231 60
rect 14231 8 14283 60
rect 14283 8 14285 60
rect 14229 6 14285 8
rect 14501 60 14557 62
rect 14501 8 14503 60
rect 14503 8 14555 60
rect 14555 8 14557 60
rect 14501 6 14557 8
rect 15785 60 15841 62
rect 15785 8 15787 60
rect 15787 8 15839 60
rect 15839 8 15841 60
rect 15785 6 15841 8
rect 16057 60 16113 62
rect 16057 8 16059 60
rect 16059 8 16111 60
rect 16111 8 16113 60
rect 16057 6 16113 8
rect 17341 60 17397 62
rect 17341 8 17343 60
rect 17343 8 17395 60
rect 17395 8 17397 60
rect 17341 6 17397 8
rect 17613 60 17669 62
rect 17613 8 17615 60
rect 17615 8 17667 60
rect 17667 8 17669 60
rect 17613 6 17669 8
rect 18897 60 18953 62
rect 18897 8 18899 60
rect 18899 8 18951 60
rect 18951 8 18953 60
rect 18897 6 18953 8
rect 19169 60 19225 62
rect 19169 8 19171 60
rect 19171 8 19223 60
rect 19223 8 19225 60
rect 19169 6 19225 8
rect 20453 60 20509 62
rect 20453 8 20455 60
rect 20455 8 20507 60
rect 20507 8 20509 60
rect 20453 6 20509 8
rect 20725 60 20781 62
rect 20725 8 20727 60
rect 20727 8 20779 60
rect 20779 8 20781 60
rect 20725 6 20781 8
rect 22009 60 22065 62
rect 22009 8 22011 60
rect 22011 8 22063 60
rect 22063 8 22065 60
rect 22009 6 22065 8
rect 22281 60 22337 62
rect 22281 8 22283 60
rect 22283 8 22335 60
rect 22335 8 22337 60
rect 22281 6 22337 8
rect 23565 60 23621 62
rect 23565 8 23567 60
rect 23567 8 23619 60
rect 23619 8 23621 60
rect 23565 6 23621 8
rect 23837 60 23893 62
rect 23837 8 23839 60
rect 23839 8 23891 60
rect 23891 8 23893 60
rect 23837 6 23893 8
rect 25121 60 25177 62
rect 25121 8 25123 60
rect 25123 8 25175 60
rect 25175 8 25177 60
rect 25121 6 25177 8
rect 25393 60 25449 62
rect 25393 8 25395 60
rect 25395 8 25447 60
rect 25447 8 25449 60
rect 25393 6 25449 8
rect 26677 60 26733 62
rect 26677 8 26679 60
rect 26679 8 26731 60
rect 26731 8 26733 60
rect 26677 6 26733 8
rect 26949 60 27005 62
rect 26949 8 26951 60
rect 26951 8 27003 60
rect 27003 8 27005 60
rect 26949 6 27005 8
rect 28233 60 28289 62
rect 28233 8 28235 60
rect 28235 8 28287 60
rect 28287 8 28289 60
rect 28233 6 28289 8
rect 28505 60 28561 62
rect 28505 8 28507 60
rect 28507 8 28559 60
rect 28559 8 28561 60
rect 28505 6 28561 8
rect 29789 60 29845 62
rect 29789 8 29791 60
rect 29791 8 29843 60
rect 29843 8 29845 60
rect 29789 6 29845 8
rect 30061 60 30117 62
rect 30061 8 30063 60
rect 30063 8 30115 60
rect 30115 8 30117 60
rect 30061 6 30117 8
rect 31345 60 31401 62
rect 31345 8 31347 60
rect 31347 8 31399 60
rect 31399 8 31401 60
rect 31345 6 31401 8
rect 31617 60 31673 62
rect 31617 8 31619 60
rect 31619 8 31671 60
rect 31671 8 31673 60
rect 31617 6 31673 8
rect 32901 60 32957 62
rect 32901 8 32903 60
rect 32903 8 32955 60
rect 32955 8 32957 60
rect 32901 6 32957 8
rect 33173 60 33229 62
rect 33173 8 33175 60
rect 33175 8 33227 60
rect 33227 8 33229 60
rect 33173 6 33229 8
rect 34457 60 34513 62
rect 34457 8 34459 60
rect 34459 8 34511 60
rect 34511 8 34513 60
rect 34457 6 34513 8
rect 34729 60 34785 62
rect 34729 8 34731 60
rect 34731 8 34783 60
rect 34783 8 34785 60
rect 34729 6 34785 8
rect 36013 60 36069 62
rect 36013 8 36015 60
rect 36015 8 36067 60
rect 36067 8 36069 60
rect 36013 6 36069 8
rect 36285 60 36341 62
rect 36285 8 36287 60
rect 36287 8 36339 60
rect 36339 8 36341 60
rect 36285 6 36341 8
rect 37569 60 37625 62
rect 37569 8 37571 60
rect 37571 8 37623 60
rect 37623 8 37625 60
rect 37569 6 37625 8
rect 37841 60 37897 62
rect 37841 8 37843 60
rect 37843 8 37895 60
rect 37895 8 37897 60
rect 37841 6 37897 8
rect 39125 60 39181 62
rect 39125 8 39127 60
rect 39127 8 39179 60
rect 39179 8 39181 60
rect 39125 6 39181 8
rect 39397 60 39453 62
rect 39397 8 39399 60
rect 39399 8 39451 60
rect 39451 8 39453 60
rect 39397 6 39453 8
rect 40681 60 40737 62
rect 40681 8 40683 60
rect 40683 8 40735 60
rect 40735 8 40737 60
rect 40681 6 40737 8
rect 40953 60 41009 62
rect 40953 8 40955 60
rect 40955 8 41007 60
rect 41007 8 41009 60
rect 40953 6 41009 8
rect 42237 60 42293 62
rect 42237 8 42239 60
rect 42239 8 42291 60
rect 42291 8 42293 60
rect 42237 6 42293 8
rect 42509 60 42565 62
rect 42509 8 42511 60
rect 42511 8 42563 60
rect 42563 8 42565 60
rect 42509 6 42565 8
rect 43793 60 43849 62
rect 43793 8 43795 60
rect 43795 8 43847 60
rect 43847 8 43849 60
rect 43793 6 43849 8
rect 44065 60 44121 62
rect 44065 8 44067 60
rect 44067 8 44119 60
rect 44119 8 44121 60
rect 44065 6 44121 8
rect 45349 60 45405 62
rect 45349 8 45351 60
rect 45351 8 45403 60
rect 45403 8 45405 60
rect 45349 6 45405 8
rect 45621 60 45677 62
rect 45621 8 45623 60
rect 45623 8 45675 60
rect 45675 8 45677 60
rect 45621 6 45677 8
rect 46905 60 46961 62
rect 46905 8 46907 60
rect 46907 8 46959 60
rect 46959 8 46961 60
rect 46905 6 46961 8
rect 47177 60 47233 62
rect 47177 8 47179 60
rect 47179 8 47231 60
rect 47231 8 47233 60
rect 47177 6 47233 8
rect 48461 60 48517 62
rect 48461 8 48463 60
rect 48463 8 48515 60
rect 48515 8 48517 60
rect 48461 6 48517 8
rect 48733 60 48789 62
rect 48733 8 48735 60
rect 48735 8 48787 60
rect 48787 8 48789 60
rect 48733 6 48789 8
<< metal3 >>
rect 187 1008 319 1017
rect 187 952 225 1008
rect 281 952 319 1008
rect 187 943 319 952
rect 459 1008 591 1017
rect 459 952 497 1008
rect 553 952 591 1008
rect 459 943 591 952
rect 1743 1008 1875 1017
rect 1743 952 1781 1008
rect 1837 952 1875 1008
rect 1743 943 1875 952
rect 2015 1008 2147 1017
rect 2015 952 2053 1008
rect 2109 952 2147 1008
rect 2015 943 2147 952
rect 3299 1008 3431 1017
rect 3299 952 3337 1008
rect 3393 952 3431 1008
rect 3299 943 3431 952
rect 3571 1008 3703 1017
rect 3571 952 3609 1008
rect 3665 952 3703 1008
rect 3571 943 3703 952
rect 4855 1008 4987 1017
rect 4855 952 4893 1008
rect 4949 952 4987 1008
rect 4855 943 4987 952
rect 5127 1008 5259 1017
rect 5127 952 5165 1008
rect 5221 952 5259 1008
rect 5127 943 5259 952
rect 6411 1008 6543 1017
rect 6411 952 6449 1008
rect 6505 952 6543 1008
rect 6411 943 6543 952
rect 6683 1008 6815 1017
rect 6683 952 6721 1008
rect 6777 952 6815 1008
rect 6683 943 6815 952
rect 7967 1008 8099 1017
rect 7967 952 8005 1008
rect 8061 952 8099 1008
rect 7967 943 8099 952
rect 8239 1008 8371 1017
rect 8239 952 8277 1008
rect 8333 952 8371 1008
rect 8239 943 8371 952
rect 9523 1008 9655 1017
rect 9523 952 9561 1008
rect 9617 952 9655 1008
rect 9523 943 9655 952
rect 9795 1008 9927 1017
rect 9795 952 9833 1008
rect 9889 952 9927 1008
rect 9795 943 9927 952
rect 11079 1008 11211 1017
rect 11079 952 11117 1008
rect 11173 952 11211 1008
rect 11079 943 11211 952
rect 11351 1008 11483 1017
rect 11351 952 11389 1008
rect 11445 952 11483 1008
rect 11351 943 11483 952
rect 12635 1008 12767 1017
rect 12635 952 12673 1008
rect 12729 952 12767 1008
rect 12635 943 12767 952
rect 12907 1008 13039 1017
rect 12907 952 12945 1008
rect 13001 952 13039 1008
rect 12907 943 13039 952
rect 14191 1008 14323 1017
rect 14191 952 14229 1008
rect 14285 952 14323 1008
rect 14191 943 14323 952
rect 14463 1008 14595 1017
rect 14463 952 14501 1008
rect 14557 952 14595 1008
rect 14463 943 14595 952
rect 15747 1008 15879 1017
rect 15747 952 15785 1008
rect 15841 952 15879 1008
rect 15747 943 15879 952
rect 16019 1008 16151 1017
rect 16019 952 16057 1008
rect 16113 952 16151 1008
rect 16019 943 16151 952
rect 17303 1008 17435 1017
rect 17303 952 17341 1008
rect 17397 952 17435 1008
rect 17303 943 17435 952
rect 17575 1008 17707 1017
rect 17575 952 17613 1008
rect 17669 952 17707 1008
rect 17575 943 17707 952
rect 18859 1008 18991 1017
rect 18859 952 18897 1008
rect 18953 952 18991 1008
rect 18859 943 18991 952
rect 19131 1008 19263 1017
rect 19131 952 19169 1008
rect 19225 952 19263 1008
rect 19131 943 19263 952
rect 20415 1008 20547 1017
rect 20415 952 20453 1008
rect 20509 952 20547 1008
rect 20415 943 20547 952
rect 20687 1008 20819 1017
rect 20687 952 20725 1008
rect 20781 952 20819 1008
rect 20687 943 20819 952
rect 21971 1008 22103 1017
rect 21971 952 22009 1008
rect 22065 952 22103 1008
rect 21971 943 22103 952
rect 22243 1008 22375 1017
rect 22243 952 22281 1008
rect 22337 952 22375 1008
rect 22243 943 22375 952
rect 23527 1008 23659 1017
rect 23527 952 23565 1008
rect 23621 952 23659 1008
rect 23527 943 23659 952
rect 23799 1008 23931 1017
rect 23799 952 23837 1008
rect 23893 952 23931 1008
rect 23799 943 23931 952
rect 25083 1008 25215 1017
rect 25083 952 25121 1008
rect 25177 952 25215 1008
rect 25083 943 25215 952
rect 25355 1008 25487 1017
rect 25355 952 25393 1008
rect 25449 952 25487 1008
rect 25355 943 25487 952
rect 26639 1008 26771 1017
rect 26639 952 26677 1008
rect 26733 952 26771 1008
rect 26639 943 26771 952
rect 26911 1008 27043 1017
rect 26911 952 26949 1008
rect 27005 952 27043 1008
rect 26911 943 27043 952
rect 28195 1008 28327 1017
rect 28195 952 28233 1008
rect 28289 952 28327 1008
rect 28195 943 28327 952
rect 28467 1008 28599 1017
rect 28467 952 28505 1008
rect 28561 952 28599 1008
rect 28467 943 28599 952
rect 29751 1008 29883 1017
rect 29751 952 29789 1008
rect 29845 952 29883 1008
rect 29751 943 29883 952
rect 30023 1008 30155 1017
rect 30023 952 30061 1008
rect 30117 952 30155 1008
rect 30023 943 30155 952
rect 31307 1008 31439 1017
rect 31307 952 31345 1008
rect 31401 952 31439 1008
rect 31307 943 31439 952
rect 31579 1008 31711 1017
rect 31579 952 31617 1008
rect 31673 952 31711 1008
rect 31579 943 31711 952
rect 32863 1008 32995 1017
rect 32863 952 32901 1008
rect 32957 952 32995 1008
rect 32863 943 32995 952
rect 33135 1008 33267 1017
rect 33135 952 33173 1008
rect 33229 952 33267 1008
rect 33135 943 33267 952
rect 34419 1008 34551 1017
rect 34419 952 34457 1008
rect 34513 952 34551 1008
rect 34419 943 34551 952
rect 34691 1008 34823 1017
rect 34691 952 34729 1008
rect 34785 952 34823 1008
rect 34691 943 34823 952
rect 35975 1008 36107 1017
rect 35975 952 36013 1008
rect 36069 952 36107 1008
rect 35975 943 36107 952
rect 36247 1008 36379 1017
rect 36247 952 36285 1008
rect 36341 952 36379 1008
rect 36247 943 36379 952
rect 37531 1008 37663 1017
rect 37531 952 37569 1008
rect 37625 952 37663 1008
rect 37531 943 37663 952
rect 37803 1008 37935 1017
rect 37803 952 37841 1008
rect 37897 952 37935 1008
rect 37803 943 37935 952
rect 39087 1008 39219 1017
rect 39087 952 39125 1008
rect 39181 952 39219 1008
rect 39087 943 39219 952
rect 39359 1008 39491 1017
rect 39359 952 39397 1008
rect 39453 952 39491 1008
rect 39359 943 39491 952
rect 40643 1008 40775 1017
rect 40643 952 40681 1008
rect 40737 952 40775 1008
rect 40643 943 40775 952
rect 40915 1008 41047 1017
rect 40915 952 40953 1008
rect 41009 952 41047 1008
rect 40915 943 41047 952
rect 42199 1008 42331 1017
rect 42199 952 42237 1008
rect 42293 952 42331 1008
rect 42199 943 42331 952
rect 42471 1008 42603 1017
rect 42471 952 42509 1008
rect 42565 952 42603 1008
rect 42471 943 42603 952
rect 43755 1008 43887 1017
rect 43755 952 43793 1008
rect 43849 952 43887 1008
rect 43755 943 43887 952
rect 44027 1008 44159 1017
rect 44027 952 44065 1008
rect 44121 952 44159 1008
rect 44027 943 44159 952
rect 45311 1008 45443 1017
rect 45311 952 45349 1008
rect 45405 952 45443 1008
rect 45311 943 45443 952
rect 45583 1008 45715 1017
rect 45583 952 45621 1008
rect 45677 952 45715 1008
rect 45583 943 45715 952
rect 46867 1008 46999 1017
rect 46867 952 46905 1008
rect 46961 952 46999 1008
rect 46867 943 46999 952
rect 47139 1008 47271 1017
rect 47139 952 47177 1008
rect 47233 952 47271 1008
rect 47139 943 47271 952
rect 48423 1008 48555 1017
rect 48423 952 48461 1008
rect 48517 952 48555 1008
rect 48423 943 48555 952
rect 48695 1008 48827 1017
rect 48695 952 48733 1008
rect 48789 952 48827 1008
rect 48695 943 48827 952
rect 187 62 319 71
rect 187 6 225 62
rect 281 6 319 62
rect 187 -3 319 6
rect 459 62 591 71
rect 459 6 497 62
rect 553 6 591 62
rect 459 -3 591 6
rect 1743 62 1875 71
rect 1743 6 1781 62
rect 1837 6 1875 62
rect 1743 -3 1875 6
rect 2015 62 2147 71
rect 2015 6 2053 62
rect 2109 6 2147 62
rect 2015 -3 2147 6
rect 3299 62 3431 71
rect 3299 6 3337 62
rect 3393 6 3431 62
rect 3299 -3 3431 6
rect 3571 62 3703 71
rect 3571 6 3609 62
rect 3665 6 3703 62
rect 3571 -3 3703 6
rect 4855 62 4987 71
rect 4855 6 4893 62
rect 4949 6 4987 62
rect 4855 -3 4987 6
rect 5127 62 5259 71
rect 5127 6 5165 62
rect 5221 6 5259 62
rect 5127 -3 5259 6
rect 6411 62 6543 71
rect 6411 6 6449 62
rect 6505 6 6543 62
rect 6411 -3 6543 6
rect 6683 62 6815 71
rect 6683 6 6721 62
rect 6777 6 6815 62
rect 6683 -3 6815 6
rect 7967 62 8099 71
rect 7967 6 8005 62
rect 8061 6 8099 62
rect 7967 -3 8099 6
rect 8239 62 8371 71
rect 8239 6 8277 62
rect 8333 6 8371 62
rect 8239 -3 8371 6
rect 9523 62 9655 71
rect 9523 6 9561 62
rect 9617 6 9655 62
rect 9523 -3 9655 6
rect 9795 62 9927 71
rect 9795 6 9833 62
rect 9889 6 9927 62
rect 9795 -3 9927 6
rect 11079 62 11211 71
rect 11079 6 11117 62
rect 11173 6 11211 62
rect 11079 -3 11211 6
rect 11351 62 11483 71
rect 11351 6 11389 62
rect 11445 6 11483 62
rect 11351 -3 11483 6
rect 12635 62 12767 71
rect 12635 6 12673 62
rect 12729 6 12767 62
rect 12635 -3 12767 6
rect 12907 62 13039 71
rect 12907 6 12945 62
rect 13001 6 13039 62
rect 12907 -3 13039 6
rect 14191 62 14323 71
rect 14191 6 14229 62
rect 14285 6 14323 62
rect 14191 -3 14323 6
rect 14463 62 14595 71
rect 14463 6 14501 62
rect 14557 6 14595 62
rect 14463 -3 14595 6
rect 15747 62 15879 71
rect 15747 6 15785 62
rect 15841 6 15879 62
rect 15747 -3 15879 6
rect 16019 62 16151 71
rect 16019 6 16057 62
rect 16113 6 16151 62
rect 16019 -3 16151 6
rect 17303 62 17435 71
rect 17303 6 17341 62
rect 17397 6 17435 62
rect 17303 -3 17435 6
rect 17575 62 17707 71
rect 17575 6 17613 62
rect 17669 6 17707 62
rect 17575 -3 17707 6
rect 18859 62 18991 71
rect 18859 6 18897 62
rect 18953 6 18991 62
rect 18859 -3 18991 6
rect 19131 62 19263 71
rect 19131 6 19169 62
rect 19225 6 19263 62
rect 19131 -3 19263 6
rect 20415 62 20547 71
rect 20415 6 20453 62
rect 20509 6 20547 62
rect 20415 -3 20547 6
rect 20687 62 20819 71
rect 20687 6 20725 62
rect 20781 6 20819 62
rect 20687 -3 20819 6
rect 21971 62 22103 71
rect 21971 6 22009 62
rect 22065 6 22103 62
rect 21971 -3 22103 6
rect 22243 62 22375 71
rect 22243 6 22281 62
rect 22337 6 22375 62
rect 22243 -3 22375 6
rect 23527 62 23659 71
rect 23527 6 23565 62
rect 23621 6 23659 62
rect 23527 -3 23659 6
rect 23799 62 23931 71
rect 23799 6 23837 62
rect 23893 6 23931 62
rect 23799 -3 23931 6
rect 25083 62 25215 71
rect 25083 6 25121 62
rect 25177 6 25215 62
rect 25083 -3 25215 6
rect 25355 62 25487 71
rect 25355 6 25393 62
rect 25449 6 25487 62
rect 25355 -3 25487 6
rect 26639 62 26771 71
rect 26639 6 26677 62
rect 26733 6 26771 62
rect 26639 -3 26771 6
rect 26911 62 27043 71
rect 26911 6 26949 62
rect 27005 6 27043 62
rect 26911 -3 27043 6
rect 28195 62 28327 71
rect 28195 6 28233 62
rect 28289 6 28327 62
rect 28195 -3 28327 6
rect 28467 62 28599 71
rect 28467 6 28505 62
rect 28561 6 28599 62
rect 28467 -3 28599 6
rect 29751 62 29883 71
rect 29751 6 29789 62
rect 29845 6 29883 62
rect 29751 -3 29883 6
rect 30023 62 30155 71
rect 30023 6 30061 62
rect 30117 6 30155 62
rect 30023 -3 30155 6
rect 31307 62 31439 71
rect 31307 6 31345 62
rect 31401 6 31439 62
rect 31307 -3 31439 6
rect 31579 62 31711 71
rect 31579 6 31617 62
rect 31673 6 31711 62
rect 31579 -3 31711 6
rect 32863 62 32995 71
rect 32863 6 32901 62
rect 32957 6 32995 62
rect 32863 -3 32995 6
rect 33135 62 33267 71
rect 33135 6 33173 62
rect 33229 6 33267 62
rect 33135 -3 33267 6
rect 34419 62 34551 71
rect 34419 6 34457 62
rect 34513 6 34551 62
rect 34419 -3 34551 6
rect 34691 62 34823 71
rect 34691 6 34729 62
rect 34785 6 34823 62
rect 34691 -3 34823 6
rect 35975 62 36107 71
rect 35975 6 36013 62
rect 36069 6 36107 62
rect 35975 -3 36107 6
rect 36247 62 36379 71
rect 36247 6 36285 62
rect 36341 6 36379 62
rect 36247 -3 36379 6
rect 37531 62 37663 71
rect 37531 6 37569 62
rect 37625 6 37663 62
rect 37531 -3 37663 6
rect 37803 62 37935 71
rect 37803 6 37841 62
rect 37897 6 37935 62
rect 37803 -3 37935 6
rect 39087 62 39219 71
rect 39087 6 39125 62
rect 39181 6 39219 62
rect 39087 -3 39219 6
rect 39359 62 39491 71
rect 39359 6 39397 62
rect 39453 6 39491 62
rect 39359 -3 39491 6
rect 40643 62 40775 71
rect 40643 6 40681 62
rect 40737 6 40775 62
rect 40643 -3 40775 6
rect 40915 62 41047 71
rect 40915 6 40953 62
rect 41009 6 41047 62
rect 40915 -3 41047 6
rect 42199 62 42331 71
rect 42199 6 42237 62
rect 42293 6 42331 62
rect 42199 -3 42331 6
rect 42471 62 42603 71
rect 42471 6 42509 62
rect 42565 6 42603 62
rect 42471 -3 42603 6
rect 43755 62 43887 71
rect 43755 6 43793 62
rect 43849 6 43887 62
rect 43755 -3 43887 6
rect 44027 62 44159 71
rect 44027 6 44065 62
rect 44121 6 44159 62
rect 44027 -3 44159 6
rect 45311 62 45443 71
rect 45311 6 45349 62
rect 45405 6 45443 62
rect 45311 -3 45443 6
rect 45583 62 45715 71
rect 45583 6 45621 62
rect 45677 6 45715 62
rect 45583 -3 45715 6
rect 46867 62 46999 71
rect 46867 6 46905 62
rect 46961 6 46999 62
rect 46867 -3 46999 6
rect 47139 62 47271 71
rect 47139 6 47177 62
rect 47233 6 47271 62
rect 47139 -3 47271 6
rect 48423 62 48555 71
rect 48423 6 48461 62
rect 48517 6 48555 62
rect 48423 -3 48555 6
rect 48695 62 48827 71
rect 48695 6 48733 62
rect 48789 6 48827 62
rect 48695 -3 48827 6
use contact_18  contact_18_0
timestamp 1644969367
transform 1 0 48695 0 1 943
box 0 0 1 1
use contact_17  contact_17_0
timestamp 1644969367
transform 1 0 48729 0 1 948
box 0 0 1 1
use contact_18  contact_18_1
timestamp 1644969367
transform 1 0 48695 0 1 -3
box 0 0 1 1
use contact_17  contact_17_1
timestamp 1644969367
transform 1 0 48729 0 1 2
box 0 0 1 1
use contact_18  contact_18_2
timestamp 1644969367
transform 1 0 48423 0 1 943
box 0 0 1 1
use contact_17  contact_17_2
timestamp 1644969367
transform 1 0 48457 0 1 948
box 0 0 1 1
use contact_18  contact_18_3
timestamp 1644969367
transform 1 0 48423 0 1 -3
box 0 0 1 1
use contact_17  contact_17_3
timestamp 1644969367
transform 1 0 48457 0 1 2
box 0 0 1 1
use contact_18  contact_18_4
timestamp 1644969367
transform 1 0 47139 0 1 943
box 0 0 1 1
use contact_17  contact_17_4
timestamp 1644969367
transform 1 0 47173 0 1 948
box 0 0 1 1
use contact_18  contact_18_5
timestamp 1644969367
transform 1 0 47139 0 1 -3
box 0 0 1 1
use contact_17  contact_17_5
timestamp 1644969367
transform 1 0 47173 0 1 2
box 0 0 1 1
use contact_18  contact_18_6
timestamp 1644969367
transform 1 0 46867 0 1 943
box 0 0 1 1
use contact_17  contact_17_6
timestamp 1644969367
transform 1 0 46901 0 1 948
box 0 0 1 1
use contact_18  contact_18_7
timestamp 1644969367
transform 1 0 46867 0 1 -3
box 0 0 1 1
use contact_17  contact_17_7
timestamp 1644969367
transform 1 0 46901 0 1 2
box 0 0 1 1
use contact_18  contact_18_8
timestamp 1644969367
transform 1 0 45583 0 1 943
box 0 0 1 1
use contact_17  contact_17_8
timestamp 1644969367
transform 1 0 45617 0 1 948
box 0 0 1 1
use contact_18  contact_18_9
timestamp 1644969367
transform 1 0 45583 0 1 -3
box 0 0 1 1
use contact_17  contact_17_9
timestamp 1644969367
transform 1 0 45617 0 1 2
box 0 0 1 1
use contact_18  contact_18_10
timestamp 1644969367
transform 1 0 45311 0 1 943
box 0 0 1 1
use contact_17  contact_17_10
timestamp 1644969367
transform 1 0 45345 0 1 948
box 0 0 1 1
use contact_18  contact_18_11
timestamp 1644969367
transform 1 0 45311 0 1 -3
box 0 0 1 1
use contact_17  contact_17_11
timestamp 1644969367
transform 1 0 45345 0 1 2
box 0 0 1 1
use contact_18  contact_18_12
timestamp 1644969367
transform 1 0 44027 0 1 943
box 0 0 1 1
use contact_17  contact_17_12
timestamp 1644969367
transform 1 0 44061 0 1 948
box 0 0 1 1
use contact_18  contact_18_13
timestamp 1644969367
transform 1 0 44027 0 1 -3
box 0 0 1 1
use contact_17  contact_17_13
timestamp 1644969367
transform 1 0 44061 0 1 2
box 0 0 1 1
use contact_18  contact_18_14
timestamp 1644969367
transform 1 0 43755 0 1 943
box 0 0 1 1
use contact_17  contact_17_14
timestamp 1644969367
transform 1 0 43789 0 1 948
box 0 0 1 1
use contact_18  contact_18_15
timestamp 1644969367
transform 1 0 43755 0 1 -3
box 0 0 1 1
use contact_17  contact_17_15
timestamp 1644969367
transform 1 0 43789 0 1 2
box 0 0 1 1
use contact_18  contact_18_16
timestamp 1644969367
transform 1 0 42471 0 1 943
box 0 0 1 1
use contact_17  contact_17_16
timestamp 1644969367
transform 1 0 42505 0 1 948
box 0 0 1 1
use contact_18  contact_18_17
timestamp 1644969367
transform 1 0 42471 0 1 -3
box 0 0 1 1
use contact_17  contact_17_17
timestamp 1644969367
transform 1 0 42505 0 1 2
box 0 0 1 1
use contact_18  contact_18_18
timestamp 1644969367
transform 1 0 42199 0 1 943
box 0 0 1 1
use contact_17  contact_17_18
timestamp 1644969367
transform 1 0 42233 0 1 948
box 0 0 1 1
use contact_18  contact_18_19
timestamp 1644969367
transform 1 0 42199 0 1 -3
box 0 0 1 1
use contact_17  contact_17_19
timestamp 1644969367
transform 1 0 42233 0 1 2
box 0 0 1 1
use contact_18  contact_18_20
timestamp 1644969367
transform 1 0 40915 0 1 943
box 0 0 1 1
use contact_17  contact_17_20
timestamp 1644969367
transform 1 0 40949 0 1 948
box 0 0 1 1
use contact_18  contact_18_21
timestamp 1644969367
transform 1 0 40915 0 1 -3
box 0 0 1 1
use contact_17  contact_17_21
timestamp 1644969367
transform 1 0 40949 0 1 2
box 0 0 1 1
use contact_18  contact_18_22
timestamp 1644969367
transform 1 0 40643 0 1 943
box 0 0 1 1
use contact_17  contact_17_22
timestamp 1644969367
transform 1 0 40677 0 1 948
box 0 0 1 1
use contact_18  contact_18_23
timestamp 1644969367
transform 1 0 40643 0 1 -3
box 0 0 1 1
use contact_17  contact_17_23
timestamp 1644969367
transform 1 0 40677 0 1 2
box 0 0 1 1
use contact_18  contact_18_24
timestamp 1644969367
transform 1 0 39359 0 1 943
box 0 0 1 1
use contact_17  contact_17_24
timestamp 1644969367
transform 1 0 39393 0 1 948
box 0 0 1 1
use contact_18  contact_18_25
timestamp 1644969367
transform 1 0 39359 0 1 -3
box 0 0 1 1
use contact_17  contact_17_25
timestamp 1644969367
transform 1 0 39393 0 1 2
box 0 0 1 1
use contact_18  contact_18_26
timestamp 1644969367
transform 1 0 39087 0 1 943
box 0 0 1 1
use contact_17  contact_17_26
timestamp 1644969367
transform 1 0 39121 0 1 948
box 0 0 1 1
use contact_18  contact_18_27
timestamp 1644969367
transform 1 0 39087 0 1 -3
box 0 0 1 1
use contact_17  contact_17_27
timestamp 1644969367
transform 1 0 39121 0 1 2
box 0 0 1 1
use contact_18  contact_18_28
timestamp 1644969367
transform 1 0 37803 0 1 943
box 0 0 1 1
use contact_17  contact_17_28
timestamp 1644969367
transform 1 0 37837 0 1 948
box 0 0 1 1
use contact_18  contact_18_29
timestamp 1644969367
transform 1 0 37803 0 1 -3
box 0 0 1 1
use contact_17  contact_17_29
timestamp 1644969367
transform 1 0 37837 0 1 2
box 0 0 1 1
use contact_18  contact_18_30
timestamp 1644969367
transform 1 0 37531 0 1 943
box 0 0 1 1
use contact_17  contact_17_30
timestamp 1644969367
transform 1 0 37565 0 1 948
box 0 0 1 1
use contact_18  contact_18_31
timestamp 1644969367
transform 1 0 37531 0 1 -3
box 0 0 1 1
use contact_17  contact_17_31
timestamp 1644969367
transform 1 0 37565 0 1 2
box 0 0 1 1
use contact_18  contact_18_32
timestamp 1644969367
transform 1 0 36247 0 1 943
box 0 0 1 1
use contact_17  contact_17_32
timestamp 1644969367
transform 1 0 36281 0 1 948
box 0 0 1 1
use contact_18  contact_18_33
timestamp 1644969367
transform 1 0 36247 0 1 -3
box 0 0 1 1
use contact_17  contact_17_33
timestamp 1644969367
transform 1 0 36281 0 1 2
box 0 0 1 1
use contact_18  contact_18_34
timestamp 1644969367
transform 1 0 35975 0 1 943
box 0 0 1 1
use contact_17  contact_17_34
timestamp 1644969367
transform 1 0 36009 0 1 948
box 0 0 1 1
use contact_18  contact_18_35
timestamp 1644969367
transform 1 0 35975 0 1 -3
box 0 0 1 1
use contact_17  contact_17_35
timestamp 1644969367
transform 1 0 36009 0 1 2
box 0 0 1 1
use contact_18  contact_18_36
timestamp 1644969367
transform 1 0 34691 0 1 943
box 0 0 1 1
use contact_17  contact_17_36
timestamp 1644969367
transform 1 0 34725 0 1 948
box 0 0 1 1
use contact_18  contact_18_37
timestamp 1644969367
transform 1 0 34691 0 1 -3
box 0 0 1 1
use contact_17  contact_17_37
timestamp 1644969367
transform 1 0 34725 0 1 2
box 0 0 1 1
use contact_18  contact_18_38
timestamp 1644969367
transform 1 0 34419 0 1 943
box 0 0 1 1
use contact_17  contact_17_38
timestamp 1644969367
transform 1 0 34453 0 1 948
box 0 0 1 1
use contact_18  contact_18_39
timestamp 1644969367
transform 1 0 34419 0 1 -3
box 0 0 1 1
use contact_17  contact_17_39
timestamp 1644969367
transform 1 0 34453 0 1 2
box 0 0 1 1
use contact_18  contact_18_40
timestamp 1644969367
transform 1 0 33135 0 1 943
box 0 0 1 1
use contact_17  contact_17_40
timestamp 1644969367
transform 1 0 33169 0 1 948
box 0 0 1 1
use contact_18  contact_18_41
timestamp 1644969367
transform 1 0 33135 0 1 -3
box 0 0 1 1
use contact_17  contact_17_41
timestamp 1644969367
transform 1 0 33169 0 1 2
box 0 0 1 1
use contact_18  contact_18_42
timestamp 1644969367
transform 1 0 32863 0 1 943
box 0 0 1 1
use contact_17  contact_17_42
timestamp 1644969367
transform 1 0 32897 0 1 948
box 0 0 1 1
use contact_18  contact_18_43
timestamp 1644969367
transform 1 0 32863 0 1 -3
box 0 0 1 1
use contact_17  contact_17_43
timestamp 1644969367
transform 1 0 32897 0 1 2
box 0 0 1 1
use contact_18  contact_18_44
timestamp 1644969367
transform 1 0 31579 0 1 943
box 0 0 1 1
use contact_17  contact_17_44
timestamp 1644969367
transform 1 0 31613 0 1 948
box 0 0 1 1
use contact_18  contact_18_45
timestamp 1644969367
transform 1 0 31579 0 1 -3
box 0 0 1 1
use contact_17  contact_17_45
timestamp 1644969367
transform 1 0 31613 0 1 2
box 0 0 1 1
use contact_18  contact_18_46
timestamp 1644969367
transform 1 0 31307 0 1 943
box 0 0 1 1
use contact_17  contact_17_46
timestamp 1644969367
transform 1 0 31341 0 1 948
box 0 0 1 1
use contact_18  contact_18_47
timestamp 1644969367
transform 1 0 31307 0 1 -3
box 0 0 1 1
use contact_17  contact_17_47
timestamp 1644969367
transform 1 0 31341 0 1 2
box 0 0 1 1
use contact_18  contact_18_48
timestamp 1644969367
transform 1 0 30023 0 1 943
box 0 0 1 1
use contact_17  contact_17_48
timestamp 1644969367
transform 1 0 30057 0 1 948
box 0 0 1 1
use contact_18  contact_18_49
timestamp 1644969367
transform 1 0 30023 0 1 -3
box 0 0 1 1
use contact_17  contact_17_49
timestamp 1644969367
transform 1 0 30057 0 1 2
box 0 0 1 1
use contact_18  contact_18_50
timestamp 1644969367
transform 1 0 29751 0 1 943
box 0 0 1 1
use contact_17  contact_17_50
timestamp 1644969367
transform 1 0 29785 0 1 948
box 0 0 1 1
use contact_18  contact_18_51
timestamp 1644969367
transform 1 0 29751 0 1 -3
box 0 0 1 1
use contact_17  contact_17_51
timestamp 1644969367
transform 1 0 29785 0 1 2
box 0 0 1 1
use contact_18  contact_18_52
timestamp 1644969367
transform 1 0 28467 0 1 943
box 0 0 1 1
use contact_17  contact_17_52
timestamp 1644969367
transform 1 0 28501 0 1 948
box 0 0 1 1
use contact_18  contact_18_53
timestamp 1644969367
transform 1 0 28467 0 1 -3
box 0 0 1 1
use contact_17  contact_17_53
timestamp 1644969367
transform 1 0 28501 0 1 2
box 0 0 1 1
use contact_18  contact_18_54
timestamp 1644969367
transform 1 0 28195 0 1 943
box 0 0 1 1
use contact_17  contact_17_54
timestamp 1644969367
transform 1 0 28229 0 1 948
box 0 0 1 1
use contact_18  contact_18_55
timestamp 1644969367
transform 1 0 28195 0 1 -3
box 0 0 1 1
use contact_17  contact_17_55
timestamp 1644969367
transform 1 0 28229 0 1 2
box 0 0 1 1
use contact_18  contact_18_56
timestamp 1644969367
transform 1 0 26911 0 1 943
box 0 0 1 1
use contact_17  contact_17_56
timestamp 1644969367
transform 1 0 26945 0 1 948
box 0 0 1 1
use contact_18  contact_18_57
timestamp 1644969367
transform 1 0 26911 0 1 -3
box 0 0 1 1
use contact_17  contact_17_57
timestamp 1644969367
transform 1 0 26945 0 1 2
box 0 0 1 1
use contact_18  contact_18_58
timestamp 1644969367
transform 1 0 26639 0 1 943
box 0 0 1 1
use contact_17  contact_17_58
timestamp 1644969367
transform 1 0 26673 0 1 948
box 0 0 1 1
use contact_18  contact_18_59
timestamp 1644969367
transform 1 0 26639 0 1 -3
box 0 0 1 1
use contact_17  contact_17_59
timestamp 1644969367
transform 1 0 26673 0 1 2
box 0 0 1 1
use contact_18  contact_18_60
timestamp 1644969367
transform 1 0 25355 0 1 943
box 0 0 1 1
use contact_17  contact_17_60
timestamp 1644969367
transform 1 0 25389 0 1 948
box 0 0 1 1
use contact_18  contact_18_61
timestamp 1644969367
transform 1 0 25355 0 1 -3
box 0 0 1 1
use contact_17  contact_17_61
timestamp 1644969367
transform 1 0 25389 0 1 2
box 0 0 1 1
use contact_18  contact_18_62
timestamp 1644969367
transform 1 0 25083 0 1 943
box 0 0 1 1
use contact_17  contact_17_62
timestamp 1644969367
transform 1 0 25117 0 1 948
box 0 0 1 1
use contact_18  contact_18_63
timestamp 1644969367
transform 1 0 25083 0 1 -3
box 0 0 1 1
use contact_17  contact_17_63
timestamp 1644969367
transform 1 0 25117 0 1 2
box 0 0 1 1
use contact_18  contact_18_64
timestamp 1644969367
transform 1 0 23799 0 1 943
box 0 0 1 1
use contact_17  contact_17_64
timestamp 1644969367
transform 1 0 23833 0 1 948
box 0 0 1 1
use contact_18  contact_18_65
timestamp 1644969367
transform 1 0 23799 0 1 -3
box 0 0 1 1
use contact_17  contact_17_65
timestamp 1644969367
transform 1 0 23833 0 1 2
box 0 0 1 1
use contact_18  contact_18_66
timestamp 1644969367
transform 1 0 23527 0 1 943
box 0 0 1 1
use contact_17  contact_17_66
timestamp 1644969367
transform 1 0 23561 0 1 948
box 0 0 1 1
use contact_18  contact_18_67
timestamp 1644969367
transform 1 0 23527 0 1 -3
box 0 0 1 1
use contact_17  contact_17_67
timestamp 1644969367
transform 1 0 23561 0 1 2
box 0 0 1 1
use contact_18  contact_18_68
timestamp 1644969367
transform 1 0 22243 0 1 943
box 0 0 1 1
use contact_17  contact_17_68
timestamp 1644969367
transform 1 0 22277 0 1 948
box 0 0 1 1
use contact_18  contact_18_69
timestamp 1644969367
transform 1 0 22243 0 1 -3
box 0 0 1 1
use contact_17  contact_17_69
timestamp 1644969367
transform 1 0 22277 0 1 2
box 0 0 1 1
use contact_18  contact_18_70
timestamp 1644969367
transform 1 0 21971 0 1 943
box 0 0 1 1
use contact_17  contact_17_70
timestamp 1644969367
transform 1 0 22005 0 1 948
box 0 0 1 1
use contact_18  contact_18_71
timestamp 1644969367
transform 1 0 21971 0 1 -3
box 0 0 1 1
use contact_17  contact_17_71
timestamp 1644969367
transform 1 0 22005 0 1 2
box 0 0 1 1
use contact_18  contact_18_72
timestamp 1644969367
transform 1 0 20687 0 1 943
box 0 0 1 1
use contact_17  contact_17_72
timestamp 1644969367
transform 1 0 20721 0 1 948
box 0 0 1 1
use contact_18  contact_18_73
timestamp 1644969367
transform 1 0 20687 0 1 -3
box 0 0 1 1
use contact_17  contact_17_73
timestamp 1644969367
transform 1 0 20721 0 1 2
box 0 0 1 1
use contact_18  contact_18_74
timestamp 1644969367
transform 1 0 20415 0 1 943
box 0 0 1 1
use contact_17  contact_17_74
timestamp 1644969367
transform 1 0 20449 0 1 948
box 0 0 1 1
use contact_18  contact_18_75
timestamp 1644969367
transform 1 0 20415 0 1 -3
box 0 0 1 1
use contact_17  contact_17_75
timestamp 1644969367
transform 1 0 20449 0 1 2
box 0 0 1 1
use contact_18  contact_18_76
timestamp 1644969367
transform 1 0 19131 0 1 943
box 0 0 1 1
use contact_17  contact_17_76
timestamp 1644969367
transform 1 0 19165 0 1 948
box 0 0 1 1
use contact_18  contact_18_77
timestamp 1644969367
transform 1 0 19131 0 1 -3
box 0 0 1 1
use contact_17  contact_17_77
timestamp 1644969367
transform 1 0 19165 0 1 2
box 0 0 1 1
use contact_18  contact_18_78
timestamp 1644969367
transform 1 0 18859 0 1 943
box 0 0 1 1
use contact_17  contact_17_78
timestamp 1644969367
transform 1 0 18893 0 1 948
box 0 0 1 1
use contact_18  contact_18_79
timestamp 1644969367
transform 1 0 18859 0 1 -3
box 0 0 1 1
use contact_17  contact_17_79
timestamp 1644969367
transform 1 0 18893 0 1 2
box 0 0 1 1
use contact_18  contact_18_80
timestamp 1644969367
transform 1 0 17575 0 1 943
box 0 0 1 1
use contact_17  contact_17_80
timestamp 1644969367
transform 1 0 17609 0 1 948
box 0 0 1 1
use contact_18  contact_18_81
timestamp 1644969367
transform 1 0 17575 0 1 -3
box 0 0 1 1
use contact_17  contact_17_81
timestamp 1644969367
transform 1 0 17609 0 1 2
box 0 0 1 1
use contact_18  contact_18_82
timestamp 1644969367
transform 1 0 17303 0 1 943
box 0 0 1 1
use contact_17  contact_17_82
timestamp 1644969367
transform 1 0 17337 0 1 948
box 0 0 1 1
use contact_18  contact_18_83
timestamp 1644969367
transform 1 0 17303 0 1 -3
box 0 0 1 1
use contact_17  contact_17_83
timestamp 1644969367
transform 1 0 17337 0 1 2
box 0 0 1 1
use contact_18  contact_18_84
timestamp 1644969367
transform 1 0 16019 0 1 943
box 0 0 1 1
use contact_17  contact_17_84
timestamp 1644969367
transform 1 0 16053 0 1 948
box 0 0 1 1
use contact_18  contact_18_85
timestamp 1644969367
transform 1 0 16019 0 1 -3
box 0 0 1 1
use contact_17  contact_17_85
timestamp 1644969367
transform 1 0 16053 0 1 2
box 0 0 1 1
use contact_18  contact_18_86
timestamp 1644969367
transform 1 0 15747 0 1 943
box 0 0 1 1
use contact_17  contact_17_86
timestamp 1644969367
transform 1 0 15781 0 1 948
box 0 0 1 1
use contact_18  contact_18_87
timestamp 1644969367
transform 1 0 15747 0 1 -3
box 0 0 1 1
use contact_17  contact_17_87
timestamp 1644969367
transform 1 0 15781 0 1 2
box 0 0 1 1
use contact_18  contact_18_88
timestamp 1644969367
transform 1 0 14463 0 1 943
box 0 0 1 1
use contact_17  contact_17_88
timestamp 1644969367
transform 1 0 14497 0 1 948
box 0 0 1 1
use contact_18  contact_18_89
timestamp 1644969367
transform 1 0 14463 0 1 -3
box 0 0 1 1
use contact_17  contact_17_89
timestamp 1644969367
transform 1 0 14497 0 1 2
box 0 0 1 1
use contact_18  contact_18_90
timestamp 1644969367
transform 1 0 14191 0 1 943
box 0 0 1 1
use contact_17  contact_17_90
timestamp 1644969367
transform 1 0 14225 0 1 948
box 0 0 1 1
use contact_18  contact_18_91
timestamp 1644969367
transform 1 0 14191 0 1 -3
box 0 0 1 1
use contact_17  contact_17_91
timestamp 1644969367
transform 1 0 14225 0 1 2
box 0 0 1 1
use contact_18  contact_18_92
timestamp 1644969367
transform 1 0 12907 0 1 943
box 0 0 1 1
use contact_17  contact_17_92
timestamp 1644969367
transform 1 0 12941 0 1 948
box 0 0 1 1
use contact_18  contact_18_93
timestamp 1644969367
transform 1 0 12907 0 1 -3
box 0 0 1 1
use contact_17  contact_17_93
timestamp 1644969367
transform 1 0 12941 0 1 2
box 0 0 1 1
use contact_18  contact_18_94
timestamp 1644969367
transform 1 0 12635 0 1 943
box 0 0 1 1
use contact_17  contact_17_94
timestamp 1644969367
transform 1 0 12669 0 1 948
box 0 0 1 1
use contact_18  contact_18_95
timestamp 1644969367
transform 1 0 12635 0 1 -3
box 0 0 1 1
use contact_17  contact_17_95
timestamp 1644969367
transform 1 0 12669 0 1 2
box 0 0 1 1
use contact_18  contact_18_96
timestamp 1644969367
transform 1 0 11351 0 1 943
box 0 0 1 1
use contact_17  contact_17_96
timestamp 1644969367
transform 1 0 11385 0 1 948
box 0 0 1 1
use contact_18  contact_18_97
timestamp 1644969367
transform 1 0 11351 0 1 -3
box 0 0 1 1
use contact_17  contact_17_97
timestamp 1644969367
transform 1 0 11385 0 1 2
box 0 0 1 1
use contact_18  contact_18_98
timestamp 1644969367
transform 1 0 11079 0 1 943
box 0 0 1 1
use contact_17  contact_17_98
timestamp 1644969367
transform 1 0 11113 0 1 948
box 0 0 1 1
use contact_18  contact_18_99
timestamp 1644969367
transform 1 0 11079 0 1 -3
box 0 0 1 1
use contact_17  contact_17_99
timestamp 1644969367
transform 1 0 11113 0 1 2
box 0 0 1 1
use contact_18  contact_18_100
timestamp 1644969367
transform 1 0 9795 0 1 943
box 0 0 1 1
use contact_17  contact_17_100
timestamp 1644969367
transform 1 0 9829 0 1 948
box 0 0 1 1
use contact_18  contact_18_101
timestamp 1644969367
transform 1 0 9795 0 1 -3
box 0 0 1 1
use contact_17  contact_17_101
timestamp 1644969367
transform 1 0 9829 0 1 2
box 0 0 1 1
use contact_18  contact_18_102
timestamp 1644969367
transform 1 0 9523 0 1 943
box 0 0 1 1
use contact_17  contact_17_102
timestamp 1644969367
transform 1 0 9557 0 1 948
box 0 0 1 1
use contact_18  contact_18_103
timestamp 1644969367
transform 1 0 9523 0 1 -3
box 0 0 1 1
use contact_17  contact_17_103
timestamp 1644969367
transform 1 0 9557 0 1 2
box 0 0 1 1
use contact_18  contact_18_104
timestamp 1644969367
transform 1 0 8239 0 1 943
box 0 0 1 1
use contact_17  contact_17_104
timestamp 1644969367
transform 1 0 8273 0 1 948
box 0 0 1 1
use contact_18  contact_18_105
timestamp 1644969367
transform 1 0 8239 0 1 -3
box 0 0 1 1
use contact_17  contact_17_105
timestamp 1644969367
transform 1 0 8273 0 1 2
box 0 0 1 1
use contact_18  contact_18_106
timestamp 1644969367
transform 1 0 7967 0 1 943
box 0 0 1 1
use contact_17  contact_17_106
timestamp 1644969367
transform 1 0 8001 0 1 948
box 0 0 1 1
use contact_18  contact_18_107
timestamp 1644969367
transform 1 0 7967 0 1 -3
box 0 0 1 1
use contact_17  contact_17_107
timestamp 1644969367
transform 1 0 8001 0 1 2
box 0 0 1 1
use contact_18  contact_18_108
timestamp 1644969367
transform 1 0 6683 0 1 943
box 0 0 1 1
use contact_17  contact_17_108
timestamp 1644969367
transform 1 0 6717 0 1 948
box 0 0 1 1
use contact_18  contact_18_109
timestamp 1644969367
transform 1 0 6683 0 1 -3
box 0 0 1 1
use contact_17  contact_17_109
timestamp 1644969367
transform 1 0 6717 0 1 2
box 0 0 1 1
use contact_18  contact_18_110
timestamp 1644969367
transform 1 0 6411 0 1 943
box 0 0 1 1
use contact_17  contact_17_110
timestamp 1644969367
transform 1 0 6445 0 1 948
box 0 0 1 1
use contact_18  contact_18_111
timestamp 1644969367
transform 1 0 6411 0 1 -3
box 0 0 1 1
use contact_17  contact_17_111
timestamp 1644969367
transform 1 0 6445 0 1 2
box 0 0 1 1
use contact_18  contact_18_112
timestamp 1644969367
transform 1 0 5127 0 1 943
box 0 0 1 1
use contact_17  contact_17_112
timestamp 1644969367
transform 1 0 5161 0 1 948
box 0 0 1 1
use contact_18  contact_18_113
timestamp 1644969367
transform 1 0 5127 0 1 -3
box 0 0 1 1
use contact_17  contact_17_113
timestamp 1644969367
transform 1 0 5161 0 1 2
box 0 0 1 1
use contact_18  contact_18_114
timestamp 1644969367
transform 1 0 4855 0 1 943
box 0 0 1 1
use contact_17  contact_17_114
timestamp 1644969367
transform 1 0 4889 0 1 948
box 0 0 1 1
use contact_18  contact_18_115
timestamp 1644969367
transform 1 0 4855 0 1 -3
box 0 0 1 1
use contact_17  contact_17_115
timestamp 1644969367
transform 1 0 4889 0 1 2
box 0 0 1 1
use contact_18  contact_18_116
timestamp 1644969367
transform 1 0 3571 0 1 943
box 0 0 1 1
use contact_17  contact_17_116
timestamp 1644969367
transform 1 0 3605 0 1 948
box 0 0 1 1
use contact_18  contact_18_117
timestamp 1644969367
transform 1 0 3571 0 1 -3
box 0 0 1 1
use contact_17  contact_17_117
timestamp 1644969367
transform 1 0 3605 0 1 2
box 0 0 1 1
use contact_18  contact_18_118
timestamp 1644969367
transform 1 0 3299 0 1 943
box 0 0 1 1
use contact_17  contact_17_118
timestamp 1644969367
transform 1 0 3333 0 1 948
box 0 0 1 1
use contact_18  contact_18_119
timestamp 1644969367
transform 1 0 3299 0 1 -3
box 0 0 1 1
use contact_17  contact_17_119
timestamp 1644969367
transform 1 0 3333 0 1 2
box 0 0 1 1
use contact_18  contact_18_120
timestamp 1644969367
transform 1 0 2015 0 1 943
box 0 0 1 1
use contact_17  contact_17_120
timestamp 1644969367
transform 1 0 2049 0 1 948
box 0 0 1 1
use contact_18  contact_18_121
timestamp 1644969367
transform 1 0 2015 0 1 -3
box 0 0 1 1
use contact_17  contact_17_121
timestamp 1644969367
transform 1 0 2049 0 1 2
box 0 0 1 1
use contact_18  contact_18_122
timestamp 1644969367
transform 1 0 1743 0 1 943
box 0 0 1 1
use contact_17  contact_17_122
timestamp 1644969367
transform 1 0 1777 0 1 948
box 0 0 1 1
use contact_18  contact_18_123
timestamp 1644969367
transform 1 0 1743 0 1 -3
box 0 0 1 1
use contact_17  contact_17_123
timestamp 1644969367
transform 1 0 1777 0 1 2
box 0 0 1 1
use contact_18  contact_18_124
timestamp 1644969367
transform 1 0 459 0 1 943
box 0 0 1 1
use contact_17  contact_17_124
timestamp 1644969367
transform 1 0 493 0 1 948
box 0 0 1 1
use contact_18  contact_18_125
timestamp 1644969367
transform 1 0 459 0 1 -3
box 0 0 1 1
use contact_17  contact_17_125
timestamp 1644969367
transform 1 0 493 0 1 2
box 0 0 1 1
use contact_18  contact_18_126
timestamp 1644969367
transform 1 0 187 0 1 943
box 0 0 1 1
use contact_17  contact_17_126
timestamp 1644969367
transform 1 0 221 0 1 948
box 0 0 1 1
use contact_18  contact_18_127
timestamp 1644969367
transform 1 0 187 0 1 -3
box 0 0 1 1
use contact_17  contact_17_127
timestamp 1644969367
transform 1 0 221 0 1 2
box 0 0 1 1
use sense_amp_multiport  sense_amp_multiport_0
timestamp 1644969367
transform 1 0 48625 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_1
timestamp 1644969367
transform 1 0 48353 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_2
timestamp 1644969367
transform 1 0 47069 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_3
timestamp 1644969367
transform 1 0 46797 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_4
timestamp 1644969367
transform 1 0 45513 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_5
timestamp 1644969367
transform 1 0 45241 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_6
timestamp 1644969367
transform 1 0 43957 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_7
timestamp 1644969367
transform 1 0 43685 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_8
timestamp 1644969367
transform 1 0 42401 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_9
timestamp 1644969367
transform 1 0 42129 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_10
timestamp 1644969367
transform 1 0 40845 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_11
timestamp 1644969367
transform 1 0 40573 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_12
timestamp 1644969367
transform 1 0 39289 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_13
timestamp 1644969367
transform 1 0 39017 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_14
timestamp 1644969367
transform 1 0 37733 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_15
timestamp 1644969367
transform 1 0 37461 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_16
timestamp 1644969367
transform 1 0 36177 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_17
timestamp 1644969367
transform 1 0 35905 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_18
timestamp 1644969367
transform 1 0 34621 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_19
timestamp 1644969367
transform 1 0 34349 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_20
timestamp 1644969367
transform 1 0 33065 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_21
timestamp 1644969367
transform 1 0 32793 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_22
timestamp 1644969367
transform 1 0 31509 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_23
timestamp 1644969367
transform 1 0 31237 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_24
timestamp 1644969367
transform 1 0 29953 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_25
timestamp 1644969367
transform 1 0 29681 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_26
timestamp 1644969367
transform 1 0 28397 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_27
timestamp 1644969367
transform 1 0 28125 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_28
timestamp 1644969367
transform 1 0 26841 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_29
timestamp 1644969367
transform 1 0 26569 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_30
timestamp 1644969367
transform 1 0 25285 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_31
timestamp 1644969367
transform 1 0 25013 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_32
timestamp 1644969367
transform 1 0 23729 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_33
timestamp 1644969367
transform 1 0 23457 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_34
timestamp 1644969367
transform 1 0 22173 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_35
timestamp 1644969367
transform 1 0 21901 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_36
timestamp 1644969367
transform 1 0 20617 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_37
timestamp 1644969367
transform 1 0 20345 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_38
timestamp 1644969367
transform 1 0 19061 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_39
timestamp 1644969367
transform 1 0 18789 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_40
timestamp 1644969367
transform 1 0 17505 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_41
timestamp 1644969367
transform 1 0 17233 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_42
timestamp 1644969367
transform 1 0 15949 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_43
timestamp 1644969367
transform 1 0 15677 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_44
timestamp 1644969367
transform 1 0 14393 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_45
timestamp 1644969367
transform 1 0 14121 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_46
timestamp 1644969367
transform 1 0 12837 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_47
timestamp 1644969367
transform 1 0 12565 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_48
timestamp 1644969367
transform 1 0 11281 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_49
timestamp 1644969367
transform 1 0 11009 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_50
timestamp 1644969367
transform 1 0 9725 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_51
timestamp 1644969367
transform 1 0 9453 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_52
timestamp 1644969367
transform 1 0 8169 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_53
timestamp 1644969367
transform 1 0 7897 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_54
timestamp 1644969367
transform 1 0 6613 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_55
timestamp 1644969367
transform 1 0 6341 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_56
timestamp 1644969367
transform 1 0 5057 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_57
timestamp 1644969367
transform 1 0 4785 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_58
timestamp 1644969367
transform 1 0 3501 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_59
timestamp 1644969367
transform 1 0 3229 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_60
timestamp 1644969367
transform 1 0 1945 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_61
timestamp 1644969367
transform 1 0 1673 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_62
timestamp 1644969367
transform 1 0 389 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_63
timestamp 1644969367
transform 1 0 117 0 1 0
box 0 0 272 1050
<< labels >>
rlabel metal3 s 3571 -3 3703 71 4 gnd
rlabel metal3 s 12907 -3 13039 71 4 gnd
rlabel metal3 s 42199 -3 42331 71 4 gnd
rlabel metal3 s 8239 -3 8371 71 4 gnd
rlabel metal3 s 32863 -3 32995 71 4 gnd
rlabel metal3 s 45311 -3 45443 71 4 gnd
rlabel metal3 s 44027 -3 44159 71 4 gnd
rlabel metal3 s 17575 -3 17707 71 4 gnd
rlabel metal3 s 43755 -3 43887 71 4 gnd
rlabel metal3 s 26639 -3 26771 71 4 gnd
rlabel metal3 s 34691 -3 34823 71 4 gnd
rlabel metal3 s 37531 -3 37663 71 4 gnd
rlabel metal3 s 48695 -3 48827 71 4 gnd
rlabel metal3 s 33135 -3 33267 71 4 gnd
rlabel metal3 s 22243 -3 22375 71 4 gnd
rlabel metal3 s 3299 -3 3431 71 4 gnd
rlabel metal3 s 14191 -3 14323 71 4 gnd
rlabel metal3 s 19131 -3 19263 71 4 gnd
rlabel metal3 s 20415 -3 20547 71 4 gnd
rlabel metal3 s 4855 -3 4987 71 4 gnd
rlabel metal3 s 17303 -3 17435 71 4 gnd
rlabel metal3 s 23527 -3 23659 71 4 gnd
rlabel metal3 s 25355 -3 25487 71 4 gnd
rlabel metal3 s 187 -3 319 71 4 gnd
rlabel metal3 s 40915 -3 41047 71 4 gnd
rlabel metal3 s 39359 -3 39491 71 4 gnd
rlabel metal3 s 23799 -3 23931 71 4 gnd
rlabel metal3 s 31579 -3 31711 71 4 gnd
rlabel metal3 s 34419 -3 34551 71 4 gnd
rlabel metal3 s 28195 -3 28327 71 4 gnd
rlabel metal3 s 35975 -3 36107 71 4 gnd
rlabel metal3 s 15747 -3 15879 71 4 gnd
rlabel metal3 s 16019 -3 16151 71 4 gnd
rlabel metal3 s 26911 -3 27043 71 4 gnd
rlabel metal3 s 9795 -3 9927 71 4 gnd
rlabel metal3 s 2015 -3 2147 71 4 gnd
rlabel metal3 s 459 -3 591 71 4 gnd
rlabel metal3 s 47139 -3 47271 71 4 gnd
rlabel metal3 s 5127 -3 5259 71 4 gnd
rlabel metal3 s 11351 -3 11483 71 4 gnd
rlabel metal3 s 30023 -3 30155 71 4 gnd
rlabel metal3 s 1743 -3 1875 71 4 gnd
rlabel metal3 s 7967 -3 8099 71 4 gnd
rlabel metal3 s 9523 -3 9655 71 4 gnd
rlabel metal3 s 12635 -3 12767 71 4 gnd
rlabel metal3 s 39087 -3 39219 71 4 gnd
rlabel metal3 s 42471 -3 42603 71 4 gnd
rlabel metal3 s 46867 -3 46999 71 4 gnd
rlabel metal3 s 37803 -3 37935 71 4 gnd
rlabel metal3 s 48423 -3 48555 71 4 gnd
rlabel metal3 s 21971 -3 22103 71 4 gnd
rlabel metal3 s 40643 -3 40775 71 4 gnd
rlabel metal3 s 25083 -3 25215 71 4 gnd
rlabel metal3 s 14463 -3 14595 71 4 gnd
rlabel metal3 s 20687 -3 20819 71 4 gnd
rlabel metal3 s 36247 -3 36379 71 4 gnd
rlabel metal3 s 28467 -3 28599 71 4 gnd
rlabel metal3 s 45583 -3 45715 71 4 gnd
rlabel metal3 s 31307 -3 31439 71 4 gnd
rlabel metal3 s 11079 -3 11211 71 4 gnd
rlabel metal3 s 18859 -3 18991 71 4 gnd
rlabel metal3 s 6411 -3 6543 71 4 gnd
rlabel metal3 s 29751 -3 29883 71 4 gnd
rlabel metal3 s 6683 -3 6815 71 4 gnd
rlabel metal3 s 17303 943 17435 1017 4 vdd
rlabel metal3 s 28195 943 28327 1017 4 vdd
rlabel metal3 s 37531 943 37663 1017 4 vdd
rlabel metal3 s 22243 943 22375 1017 4 vdd
rlabel metal3 s 6411 943 6543 1017 4 vdd
rlabel metal3 s 11079 943 11211 1017 4 vdd
rlabel metal3 s 16019 943 16151 1017 4 vdd
rlabel metal3 s 3571 943 3703 1017 4 vdd
rlabel metal3 s 34691 943 34823 1017 4 vdd
rlabel metal3 s 39087 943 39219 1017 4 vdd
rlabel metal3 s 9795 943 9927 1017 4 vdd
rlabel metal3 s 17575 943 17707 1017 4 vdd
rlabel metal3 s 29751 943 29883 1017 4 vdd
rlabel metal3 s 3299 943 3431 1017 4 vdd
rlabel metal3 s 19131 943 19263 1017 4 vdd
rlabel metal3 s 48423 943 48555 1017 4 vdd
rlabel metal3 s 40643 943 40775 1017 4 vdd
rlabel metal3 s 14191 943 14323 1017 4 vdd
rlabel metal3 s 14463 943 14595 1017 4 vdd
rlabel metal3 s 44027 943 44159 1017 4 vdd
rlabel metal3 s 187 943 319 1017 4 vdd
rlabel metal3 s 8239 943 8371 1017 4 vdd
rlabel metal3 s 1743 943 1875 1017 4 vdd
rlabel metal3 s 42471 943 42603 1017 4 vdd
rlabel metal3 s 47139 943 47271 1017 4 vdd
rlabel metal3 s 12907 943 13039 1017 4 vdd
rlabel metal3 s 25355 943 25487 1017 4 vdd
rlabel metal3 s 46867 943 46999 1017 4 vdd
rlabel metal3 s 40915 943 41047 1017 4 vdd
rlabel metal3 s 31307 943 31439 1017 4 vdd
rlabel metal3 s 23527 943 23659 1017 4 vdd
rlabel metal3 s 28467 943 28599 1017 4 vdd
rlabel metal3 s 459 943 591 1017 4 vdd
rlabel metal3 s 32863 943 32995 1017 4 vdd
rlabel metal3 s 25083 943 25215 1017 4 vdd
rlabel metal3 s 35975 943 36107 1017 4 vdd
rlabel metal3 s 7967 943 8099 1017 4 vdd
rlabel metal3 s 12635 943 12767 1017 4 vdd
rlabel metal3 s 15747 943 15879 1017 4 vdd
rlabel metal3 s 23799 943 23931 1017 4 vdd
rlabel metal3 s 45583 943 45715 1017 4 vdd
rlabel metal3 s 2015 943 2147 1017 4 vdd
rlabel metal3 s 26911 943 27043 1017 4 vdd
rlabel metal3 s 48695 943 48827 1017 4 vdd
rlabel metal3 s 45311 943 45443 1017 4 vdd
rlabel metal3 s 30023 943 30155 1017 4 vdd
rlabel metal3 s 33135 943 33267 1017 4 vdd
rlabel metal3 s 37803 943 37935 1017 4 vdd
rlabel metal3 s 43755 943 43887 1017 4 vdd
rlabel metal3 s 6683 943 6815 1017 4 vdd
rlabel metal3 s 31579 943 31711 1017 4 vdd
rlabel metal3 s 39359 943 39491 1017 4 vdd
rlabel metal3 s 5127 943 5259 1017 4 vdd
rlabel metal3 s 18859 943 18991 1017 4 vdd
rlabel metal3 s 20415 943 20547 1017 4 vdd
rlabel metal3 s 26639 943 26771 1017 4 vdd
rlabel metal3 s 42199 943 42331 1017 4 vdd
rlabel metal3 s 9523 943 9655 1017 4 vdd
rlabel metal3 s 34419 943 34551 1017 4 vdd
rlabel metal3 s 20687 943 20819 1017 4 vdd
rlabel metal3 s 21971 943 22103 1017 4 vdd
rlabel metal3 s 36247 943 36379 1017 4 vdd
rlabel metal3 s 4855 943 4987 1017 4 vdd
rlabel metal3 s 11351 943 11483 1017 4 vdd
rlabel metal2 s 131 0 159 240 4 rbl_0
rlabel metal2 s 319 0 347 240 4 data_0
rlabel metal2 s 403 0 431 240 4 rbl_1
rlabel metal2 s 591 0 619 240 4 data_1
rlabel metal2 s 1687 0 1715 240 4 rbl_2
rlabel metal2 s 1875 0 1903 240 4 data_2
rlabel metal2 s 1959 0 1987 240 4 rbl_3
rlabel metal2 s 2147 0 2175 240 4 data_3
rlabel metal2 s 3243 0 3271 240 4 rbl_4
rlabel metal2 s 3431 0 3459 240 4 data_4
rlabel metal2 s 3515 0 3543 240 4 rbl_5
rlabel metal2 s 3703 0 3731 240 4 data_5
rlabel metal2 s 4799 0 4827 240 4 rbl_6
rlabel metal2 s 4987 0 5015 240 4 data_6
rlabel metal2 s 5071 0 5099 240 4 rbl_7
rlabel metal2 s 5259 0 5287 240 4 data_7
rlabel metal2 s 6355 0 6383 240 4 rbl_8
rlabel metal2 s 6543 0 6571 240 4 data_8
rlabel metal2 s 6627 0 6655 240 4 rbl_9
rlabel metal2 s 6815 0 6843 240 4 data_9
rlabel metal2 s 7911 0 7939 240 4 rbl_10
rlabel metal2 s 8099 0 8127 240 4 data_10
rlabel metal2 s 8183 0 8211 240 4 rbl_11
rlabel metal2 s 8371 0 8399 240 4 data_11
rlabel metal2 s 9467 0 9495 240 4 rbl_12
rlabel metal2 s 9655 0 9683 240 4 data_12
rlabel metal2 s 9739 0 9767 240 4 rbl_13
rlabel metal2 s 9927 0 9955 240 4 data_13
rlabel metal2 s 11023 0 11051 240 4 rbl_14
rlabel metal2 s 11211 0 11239 240 4 data_14
rlabel metal2 s 11295 0 11323 240 4 rbl_15
rlabel metal2 s 11483 0 11511 240 4 data_15
rlabel metal2 s 12579 0 12607 240 4 rbl_16
rlabel metal2 s 12767 0 12795 240 4 data_16
rlabel metal2 s 12851 0 12879 240 4 rbl_17
rlabel metal2 s 13039 0 13067 240 4 data_17
rlabel metal2 s 14135 0 14163 240 4 rbl_18
rlabel metal2 s 14323 0 14351 240 4 data_18
rlabel metal2 s 14407 0 14435 240 4 rbl_19
rlabel metal2 s 14595 0 14623 240 4 data_19
rlabel metal2 s 15691 0 15719 240 4 rbl_20
rlabel metal2 s 15879 0 15907 240 4 data_20
rlabel metal2 s 15963 0 15991 240 4 rbl_21
rlabel metal2 s 16151 0 16179 240 4 data_21
rlabel metal2 s 17247 0 17275 240 4 rbl_22
rlabel metal2 s 17435 0 17463 240 4 data_22
rlabel metal2 s 17519 0 17547 240 4 rbl_23
rlabel metal2 s 17707 0 17735 240 4 data_23
rlabel metal2 s 18803 0 18831 240 4 rbl_24
rlabel metal2 s 18991 0 19019 240 4 data_24
rlabel metal2 s 19075 0 19103 240 4 rbl_25
rlabel metal2 s 19263 0 19291 240 4 data_25
rlabel metal2 s 20359 0 20387 240 4 rbl_26
rlabel metal2 s 20547 0 20575 240 4 data_26
rlabel metal2 s 20631 0 20659 240 4 rbl_27
rlabel metal2 s 20819 0 20847 240 4 data_27
rlabel metal2 s 21915 0 21943 240 4 rbl_28
rlabel metal2 s 22103 0 22131 240 4 data_28
rlabel metal2 s 22187 0 22215 240 4 rbl_29
rlabel metal2 s 22375 0 22403 240 4 data_29
rlabel metal2 s 23471 0 23499 240 4 rbl_30
rlabel metal2 s 23659 0 23687 240 4 data_30
rlabel metal2 s 23743 0 23771 240 4 rbl_31
rlabel metal2 s 23931 0 23959 240 4 data_31
rlabel metal2 s 25027 0 25055 240 4 rbl_32
rlabel metal2 s 25215 0 25243 240 4 data_32
rlabel metal2 s 25299 0 25327 240 4 rbl_33
rlabel metal2 s 25487 0 25515 240 4 data_33
rlabel metal2 s 26583 0 26611 240 4 rbl_34
rlabel metal2 s 26771 0 26799 240 4 data_34
rlabel metal2 s 26855 0 26883 240 4 rbl_35
rlabel metal2 s 27043 0 27071 240 4 data_35
rlabel metal2 s 28139 0 28167 240 4 rbl_36
rlabel metal2 s 28327 0 28355 240 4 data_36
rlabel metal2 s 28411 0 28439 240 4 rbl_37
rlabel metal2 s 28599 0 28627 240 4 data_37
rlabel metal2 s 29695 0 29723 240 4 rbl_38
rlabel metal2 s 29883 0 29911 240 4 data_38
rlabel metal2 s 29967 0 29995 240 4 rbl_39
rlabel metal2 s 30155 0 30183 240 4 data_39
rlabel metal2 s 31251 0 31279 240 4 rbl_40
rlabel metal2 s 31439 0 31467 240 4 data_40
rlabel metal2 s 31523 0 31551 240 4 rbl_41
rlabel metal2 s 31711 0 31739 240 4 data_41
rlabel metal2 s 32807 0 32835 240 4 rbl_42
rlabel metal2 s 32995 0 33023 240 4 data_42
rlabel metal2 s 33079 0 33107 240 4 rbl_43
rlabel metal2 s 33267 0 33295 240 4 data_43
rlabel metal2 s 34363 0 34391 240 4 rbl_44
rlabel metal2 s 34551 0 34579 240 4 data_44
rlabel metal2 s 34635 0 34663 240 4 rbl_45
rlabel metal2 s 34823 0 34851 240 4 data_45
rlabel metal2 s 35919 0 35947 240 4 rbl_46
rlabel metal2 s 36107 0 36135 240 4 data_46
rlabel metal2 s 36191 0 36219 240 4 rbl_47
rlabel metal2 s 36379 0 36407 240 4 data_47
rlabel metal2 s 37475 0 37503 240 4 rbl_48
rlabel metal2 s 37663 0 37691 240 4 data_48
rlabel metal2 s 37747 0 37775 240 4 rbl_49
rlabel metal2 s 37935 0 37963 240 4 data_49
rlabel metal2 s 39031 0 39059 240 4 rbl_50
rlabel metal2 s 39219 0 39247 240 4 data_50
rlabel metal2 s 39303 0 39331 240 4 rbl_51
rlabel metal2 s 39491 0 39519 240 4 data_51
rlabel metal2 s 40587 0 40615 240 4 rbl_52
rlabel metal2 s 40775 0 40803 240 4 data_52
rlabel metal2 s 40859 0 40887 240 4 rbl_53
rlabel metal2 s 41047 0 41075 240 4 data_53
rlabel metal2 s 42143 0 42171 240 4 rbl_54
rlabel metal2 s 42331 0 42359 240 4 data_54
rlabel metal2 s 42415 0 42443 240 4 rbl_55
rlabel metal2 s 42603 0 42631 240 4 data_55
rlabel metal2 s 43699 0 43727 240 4 rbl_56
rlabel metal2 s 43887 0 43915 240 4 data_56
rlabel metal2 s 43971 0 43999 240 4 rbl_57
rlabel metal2 s 44159 0 44187 240 4 data_57
rlabel metal2 s 45255 0 45283 240 4 rbl_58
rlabel metal2 s 45443 0 45471 240 4 data_58
rlabel metal2 s 45527 0 45555 240 4 rbl_59
rlabel metal2 s 45715 0 45743 240 4 data_59
rlabel metal2 s 46811 0 46839 240 4 rbl_60
rlabel metal2 s 46999 0 47027 240 4 data_60
rlabel metal2 s 47083 0 47111 240 4 rbl_61
rlabel metal2 s 47271 0 47299 240 4 data_61
rlabel metal2 s 48367 0 48395 240 4 rbl_62
rlabel metal2 s 48555 0 48583 240 4 data_62
rlabel metal2 s 48639 0 48667 240 4 rbl_63
rlabel metal2 s 48827 0 48855 240 4 data_63
<< properties >>
string FIXED_BBOX 48695 -3 48827 0
string GDS_FILE sram_0rw2r1w_32_128_sky130A.gds
string GDS_END 2597702
string GDS_START 2527958
<< end >>
