magic
tech sky130A
magscale 1 2
timestamp 1644969367
<< checkpaint >>
rect -1296 -1277 2132 2857
<< locali >>
rect 0 1523 836 1557
rect 330 745 364 1263
rect 330 711 549 745
rect 647 711 681 745
rect 196 381 262 447
rect 96 257 162 323
rect 0 -17 836 17
use pinv  pinv_0
timestamp 1644969367
transform 1 0 468 0 1 0
box -36 -17 404 1597
use pnand2  pnand2_0
timestamp 1644969367
transform 1 0 0 0 1 0
box -36 -17 504 1597
<< labels >>
rlabel locali s 664 728 664 728 4 Z
rlabel locali s 129 290 129 290 4 A
rlabel locali s 229 414 229 414 4 B
rlabel locali s 418 0 418 0 4 gnd
rlabel locali s 418 1540 418 1540 4 vdd
<< properties >>
string FIXED_BBOX 0 0 836 1540
string GDS_FILE sram_0rw2r1w_32_128_sky130A.gds
string GDS_END 3069894
string GDS_START 3068896
<< end >>
