magic
tech sky130A
magscale 1 2
timestamp 1644969367
<< checkpaint >>
rect -1260 -1302 9332 99734
<< metal1 >>
rect 6438 97850 6732 97852
rect 6438 97824 7352 97850
rect 6704 97822 7352 97824
rect 7978 97752 8006 97780
rect 6438 97702 7050 97730
rect 7978 97626 8006 97654
rect 6438 97556 6872 97584
rect 7978 97400 8006 97428
rect 7978 96360 8006 96388
rect 6438 96204 6872 96232
rect 7978 96134 8006 96162
rect 6438 96058 7050 96086
rect 7978 96008 8006 96036
rect 6704 95964 7352 95966
rect 6438 95938 7352 95964
rect 6438 95936 6732 95938
rect 6438 94774 6732 94776
rect 6438 94748 7352 94774
rect 6704 94746 7352 94748
rect 7978 94676 8006 94704
rect 6438 94626 7050 94654
rect 7978 94550 8006 94578
rect 6438 94480 6872 94508
rect 7978 94324 8006 94352
rect 7978 93284 8006 93312
rect 6438 93128 6872 93156
rect 7978 93058 8006 93086
rect 6438 92982 7050 93010
rect 7978 92932 8006 92960
rect 6704 92888 7352 92890
rect 6438 92862 7352 92888
rect 6438 92860 6732 92862
rect 6438 91698 6732 91700
rect 6438 91672 7352 91698
rect 6704 91670 7352 91672
rect 7978 91600 8006 91628
rect 6438 91550 7050 91578
rect 7978 91474 8006 91502
rect 6438 91404 6872 91432
rect 7978 91248 8006 91276
rect 7978 90208 8006 90236
rect 6438 90052 6872 90080
rect 7978 89982 8006 90010
rect 6438 89906 7050 89934
rect 7978 89856 8006 89884
rect 6704 89812 7352 89814
rect 6438 89786 7352 89812
rect 6438 89784 6732 89786
rect 6438 88622 6732 88624
rect 6438 88596 7352 88622
rect 6704 88594 7352 88596
rect 7978 88524 8006 88552
rect 6438 88474 7050 88502
rect 7978 88398 8006 88426
rect 6438 88328 6872 88356
rect 7978 88172 8006 88200
rect 7978 87132 8006 87160
rect 6438 86976 6872 87004
rect 7978 86906 8006 86934
rect 6438 86830 7050 86858
rect 7978 86780 8006 86808
rect 6704 86736 7352 86738
rect 6438 86710 7352 86736
rect 6438 86708 6732 86710
rect 6438 85546 6732 85548
rect 6438 85520 7352 85546
rect 6704 85518 7352 85520
rect 7978 85448 8006 85476
rect 6438 85398 7050 85426
rect 7978 85322 8006 85350
rect 6438 85252 6872 85280
rect 7978 85096 8006 85124
rect 7978 84056 8006 84084
rect 6438 83900 6872 83928
rect 7978 83830 8006 83858
rect 6438 83754 7050 83782
rect 7978 83704 8006 83732
rect 6704 83660 7352 83662
rect 6438 83634 7352 83660
rect 6438 83632 6732 83634
rect 6438 82470 6732 82472
rect 6438 82444 7352 82470
rect 6704 82442 7352 82444
rect 7978 82372 8006 82400
rect 6438 82322 7050 82350
rect 7978 82246 8006 82274
rect 6438 82176 6872 82204
rect 7978 82020 8006 82048
rect 7978 80980 8006 81008
rect 6438 80824 6872 80852
rect 7978 80754 8006 80782
rect 6438 80678 7050 80706
rect 7978 80628 8006 80656
rect 6704 80584 7352 80586
rect 6438 80558 7352 80584
rect 6438 80556 6732 80558
rect 6438 79394 6732 79396
rect 6438 79368 7352 79394
rect 6704 79366 7352 79368
rect 7978 79296 8006 79324
rect 6438 79246 7050 79274
rect 7978 79170 8006 79198
rect 6438 79100 6872 79128
rect 7978 78944 8006 78972
rect 7978 77904 8006 77932
rect 6438 77748 6872 77776
rect 7978 77678 8006 77706
rect 6438 77602 7050 77630
rect 7978 77552 8006 77580
rect 6704 77508 7352 77510
rect 6438 77482 7352 77508
rect 6438 77480 6732 77482
rect 6438 76318 6732 76320
rect 6438 76292 7352 76318
rect 6704 76290 7352 76292
rect 7978 76220 8006 76248
rect 6438 76170 7050 76198
rect 7978 76094 8006 76122
rect 6438 76024 6872 76052
rect 7978 75868 8006 75896
rect 7978 74828 8006 74856
rect 6438 74672 6872 74700
rect 7978 74602 8006 74630
rect 6438 74526 7050 74554
rect 7978 74476 8006 74504
rect 6704 74432 7352 74434
rect 6438 74406 7352 74432
rect 6438 74404 6732 74406
rect 6438 73242 6732 73244
rect 6438 73216 7352 73242
rect 6704 73214 7352 73216
rect 7978 73144 8006 73172
rect 6438 73094 7050 73122
rect 7978 73018 8006 73046
rect 6438 72948 6872 72976
rect 7978 72792 8006 72820
rect 7978 71752 8006 71780
rect 6438 71596 6872 71624
rect 7978 71526 8006 71554
rect 6438 71450 7050 71478
rect 7978 71400 8006 71428
rect 6704 71356 7352 71358
rect 6438 71330 7352 71356
rect 6438 71328 6732 71330
rect 6438 70166 6732 70168
rect 6438 70140 7352 70166
rect 6704 70138 7352 70140
rect 7978 70068 8006 70096
rect 6438 70018 7050 70046
rect 7978 69942 8006 69970
rect 6438 69872 6872 69900
rect 7978 69716 8006 69744
rect 7978 68676 8006 68704
rect 6438 68520 6872 68548
rect 7978 68450 8006 68478
rect 6438 68374 7050 68402
rect 7978 68324 8006 68352
rect 6704 68280 7352 68282
rect 6438 68254 7352 68280
rect 6438 68252 6732 68254
rect 6438 67090 6732 67092
rect 6438 67064 7352 67090
rect 6704 67062 7352 67064
rect 7978 66992 8006 67020
rect 6438 66942 7050 66970
rect 7978 66866 8006 66894
rect 6438 66796 6872 66824
rect 7978 66640 8006 66668
rect 7978 65600 8006 65628
rect 6438 65444 6872 65472
rect 7978 65374 8006 65402
rect 6438 65298 7050 65326
rect 7978 65248 8006 65276
rect 6704 65204 7352 65206
rect 6438 65178 7352 65204
rect 6438 65176 6732 65178
rect 6438 64014 6732 64016
rect 6438 63988 7352 64014
rect 6704 63986 7352 63988
rect 7978 63916 8006 63944
rect 6438 63866 7050 63894
rect 7978 63790 8006 63818
rect 6438 63720 6872 63748
rect 7978 63564 8006 63592
rect 7978 62524 8006 62552
rect 6438 62368 6872 62396
rect 7978 62298 8006 62326
rect 6438 62222 7050 62250
rect 7978 62172 8006 62200
rect 6704 62128 7352 62130
rect 6438 62102 7352 62128
rect 6438 62100 6732 62102
rect 6438 60938 6732 60940
rect 6438 60912 7352 60938
rect 6704 60910 7352 60912
rect 7978 60840 8006 60868
rect 6438 60790 7050 60818
rect 7978 60714 8006 60742
rect 6438 60644 6872 60672
rect 7978 60488 8006 60516
rect 7978 59448 8006 59476
rect 6438 59292 6872 59320
rect 7978 59222 8006 59250
rect 6438 59146 7050 59174
rect 7978 59096 8006 59124
rect 6704 59052 7352 59054
rect 6438 59026 7352 59052
rect 6438 59024 6732 59026
rect 6438 57862 6732 57864
rect 6438 57836 7352 57862
rect 6704 57834 7352 57836
rect 7978 57764 8006 57792
rect 6438 57714 7050 57742
rect 7978 57638 8006 57666
rect 6438 57568 6872 57596
rect 7978 57412 8006 57440
rect 7978 56372 8006 56400
rect 6438 56216 6872 56244
rect 7978 56146 8006 56174
rect 6438 56070 7050 56098
rect 7978 56020 8006 56048
rect 6704 55976 7352 55978
rect 6438 55950 7352 55976
rect 6438 55948 6732 55950
rect 6438 54786 6732 54788
rect 6438 54760 7352 54786
rect 6704 54758 7352 54760
rect 7978 54688 8006 54716
rect 6438 54638 7050 54666
rect 7978 54562 8006 54590
rect 6438 54492 6872 54520
rect 7978 54336 8006 54364
rect 7978 53296 8006 53324
rect 6438 53140 6872 53168
rect 7978 53070 8006 53098
rect 6438 52994 7050 53022
rect 7978 52944 8006 52972
rect 6704 52900 7352 52902
rect 6438 52874 7352 52900
rect 6438 52872 6732 52874
rect 6438 51710 6732 51712
rect 6438 51684 7352 51710
rect 6704 51682 7352 51684
rect 7978 51612 8006 51640
rect 6438 51562 7050 51590
rect 7978 51486 8006 51514
rect 6438 51416 6872 51444
rect 7978 51260 8006 51288
rect 7978 50220 8006 50248
rect 6438 50064 6872 50092
rect 7978 49994 8006 50022
rect 6438 49918 7050 49946
rect 7978 49868 8006 49896
rect 6704 49824 7352 49826
rect 6438 49798 7352 49824
rect 6438 49796 6732 49798
rect 6438 48634 6732 48636
rect 6438 48608 7352 48634
rect 6704 48606 7352 48608
rect 7978 48536 8006 48564
rect 6438 48486 7050 48514
rect 7978 48410 8006 48438
rect 6438 48340 6872 48368
rect 7978 48184 8006 48212
rect 7978 47144 8006 47172
rect 6438 46988 6872 47016
rect 7978 46918 8006 46946
rect 6438 46842 7050 46870
rect 7978 46792 8006 46820
rect 6704 46748 7352 46750
rect 6438 46722 7352 46748
rect 6438 46720 6732 46722
rect 6438 45558 6732 45560
rect 6438 45532 7352 45558
rect 6704 45530 7352 45532
rect 7978 45460 8006 45488
rect 6438 45410 7050 45438
rect 7978 45334 8006 45362
rect 6438 45264 6872 45292
rect 7978 45108 8006 45136
rect 7978 44068 8006 44096
rect 6438 43912 6872 43940
rect 7978 43842 8006 43870
rect 6438 43766 7050 43794
rect 7978 43716 8006 43744
rect 6704 43672 7352 43674
rect 6438 43646 7352 43672
rect 6438 43644 6732 43646
rect 6438 42482 6732 42484
rect 6438 42456 7352 42482
rect 6704 42454 7352 42456
rect 7978 42384 8006 42412
rect 6438 42334 7050 42362
rect 7978 42258 8006 42286
rect 6438 42188 6872 42216
rect 7978 42032 8006 42060
rect 7978 40992 8006 41020
rect 6438 40836 6872 40864
rect 7978 40766 8006 40794
rect 6438 40690 7050 40718
rect 7978 40640 8006 40668
rect 6704 40596 7352 40598
rect 6438 40570 7352 40596
rect 6438 40568 6732 40570
rect 6438 39406 6732 39408
rect 6438 39380 7352 39406
rect 6704 39378 7352 39380
rect 7978 39308 8006 39336
rect 6438 39258 7050 39286
rect 7978 39182 8006 39210
rect 6438 39112 6872 39140
rect 7978 38956 8006 38984
rect 7978 37916 8006 37944
rect 6438 37760 6872 37788
rect 7978 37690 8006 37718
rect 6438 37614 7050 37642
rect 7978 37564 8006 37592
rect 6704 37520 7352 37522
rect 6438 37494 7352 37520
rect 6438 37492 6732 37494
rect 6438 36330 6732 36332
rect 6438 36304 7352 36330
rect 6704 36302 7352 36304
rect 7978 36232 8006 36260
rect 6438 36182 7050 36210
rect 7978 36106 8006 36134
rect 6438 36036 6872 36064
rect 7978 35880 8006 35908
rect 7978 34840 8006 34868
rect 6438 34684 6872 34712
rect 7978 34614 8006 34642
rect 6438 34538 7050 34566
rect 7978 34488 8006 34516
rect 6704 34444 7352 34446
rect 6438 34418 7352 34444
rect 6438 34416 6732 34418
rect 6438 33254 6732 33256
rect 6438 33228 7352 33254
rect 6704 33226 7352 33228
rect 7978 33156 8006 33184
rect 6438 33106 7050 33134
rect 7978 33030 8006 33058
rect 6438 32960 6872 32988
rect 7978 32804 8006 32832
rect 7978 31764 8006 31792
rect 6438 31608 6872 31636
rect 7978 31538 8006 31566
rect 6438 31462 7050 31490
rect 7978 31412 8006 31440
rect 6704 31368 7352 31370
rect 6438 31342 7352 31368
rect 6438 31340 6732 31342
rect 6438 30178 6732 30180
rect 6438 30152 7352 30178
rect 6704 30150 7352 30152
rect 7978 30080 8006 30108
rect 6438 30030 7050 30058
rect 7978 29954 8006 29982
rect 6438 29884 6872 29912
rect 7978 29728 8006 29756
rect 7978 28688 8006 28716
rect 6438 28532 6872 28560
rect 7978 28462 8006 28490
rect 6438 28386 7050 28414
rect 7978 28336 8006 28364
rect 6704 28292 7352 28294
rect 6438 28266 7352 28292
rect 6438 28264 6732 28266
rect 6438 27102 6732 27104
rect 6438 27076 7352 27102
rect 6704 27074 7352 27076
rect 7978 27004 8006 27032
rect 6438 26954 7050 26982
rect 7978 26878 8006 26906
rect 6438 26808 6872 26836
rect 7978 26652 8006 26680
rect 7978 25612 8006 25640
rect 6438 25456 6872 25484
rect 7978 25386 8006 25414
rect 6438 25310 7050 25338
rect 7978 25260 8006 25288
rect 6704 25216 7352 25218
rect 6438 25190 7352 25216
rect 6438 25188 6732 25190
rect 6438 24026 6732 24028
rect 6438 24000 7352 24026
rect 6704 23998 7352 24000
rect 7978 23928 8006 23956
rect 6438 23878 7050 23906
rect 7978 23802 8006 23830
rect 6438 23732 6872 23760
rect 7978 23576 8006 23604
rect 7978 22536 8006 22564
rect 6438 22380 6872 22408
rect 7978 22310 8006 22338
rect 6438 22234 7050 22262
rect 7978 22184 8006 22212
rect 6704 22140 7352 22142
rect 6438 22114 7352 22140
rect 6438 22112 6732 22114
rect 6438 20950 6732 20952
rect 6438 20924 7352 20950
rect 6704 20922 7352 20924
rect 7978 20852 8006 20880
rect 6438 20802 7050 20830
rect 7978 20726 8006 20754
rect 6438 20656 6872 20684
rect 7978 20500 8006 20528
rect 7978 19460 8006 19488
rect 6438 19304 6872 19332
rect 7978 19234 8006 19262
rect 6438 19158 7050 19186
rect 7978 19108 8006 19136
rect 6704 19064 7352 19066
rect 6438 19038 7352 19064
rect 6438 19036 6732 19038
rect 6438 17874 6732 17876
rect 6438 17848 7352 17874
rect 6704 17846 7352 17848
rect 7978 17776 8006 17804
rect 6438 17726 7050 17754
rect 7978 17650 8006 17678
rect 6438 17580 6872 17608
rect 7978 17424 8006 17452
rect 7978 16384 8006 16412
rect 6438 16228 6872 16256
rect 7978 16158 8006 16186
rect 6438 16082 7050 16110
rect 7978 16032 8006 16060
rect 6704 15988 7352 15990
rect 6438 15962 7352 15988
rect 6438 15960 6732 15962
rect 6438 14798 6732 14800
rect 6438 14772 7352 14798
rect 6704 14770 7352 14772
rect 7978 14700 8006 14728
rect 6438 14650 7050 14678
rect 7978 14574 8006 14602
rect 6438 14504 6872 14532
rect 7978 14348 8006 14376
rect 7978 13308 8006 13336
rect 6438 13152 6872 13180
rect 7978 13082 8006 13110
rect 6438 13006 7050 13034
rect 7978 12956 8006 12984
rect 6704 12912 7352 12914
rect 6438 12886 7352 12912
rect 6438 12884 6732 12886
rect 6438 11722 6732 11724
rect 6438 11696 7352 11722
rect 6704 11694 7352 11696
rect 7978 11624 8006 11652
rect 6438 11574 7050 11602
rect 7978 11498 8006 11526
rect 6438 11428 6872 11456
rect 7978 11272 8006 11300
rect 7978 10232 8006 10260
rect 6438 10076 6872 10104
rect 7978 10006 8006 10034
rect 6438 9930 7050 9958
rect 7978 9880 8006 9908
rect 6704 9836 7352 9838
rect 6438 9810 7352 9836
rect 6438 9808 6732 9810
rect 6438 8646 6732 8648
rect 6438 8620 7352 8646
rect 6704 8618 7352 8620
rect 7978 8548 8006 8576
rect 6438 8498 7050 8526
rect 7978 8422 8006 8450
rect 6438 8352 6872 8380
rect 7978 8196 8006 8224
rect 7978 7156 8006 7184
rect 6438 7000 6872 7028
rect 7978 6930 8006 6958
rect 6438 6854 7050 6882
rect 7978 6804 8006 6832
rect 6704 6760 7352 6762
rect 6438 6734 7352 6760
rect 6438 6732 6732 6734
rect 6438 5570 6732 5572
rect 6438 5544 7352 5570
rect 6704 5542 7352 5544
rect 7978 5472 8006 5500
rect 6438 5422 7050 5450
rect 7978 5346 8006 5374
rect 6438 5276 6872 5304
rect 7978 5120 8006 5148
rect 7978 4080 8006 4108
rect 6438 3924 6872 3952
rect 7978 3854 8006 3882
rect 6438 3778 7050 3806
rect 7978 3728 8006 3756
rect 6704 3684 7352 3686
rect 6438 3658 7352 3684
rect 6438 3656 6732 3658
rect 6438 2494 6732 2496
rect 6438 2468 7352 2494
rect 6704 2466 7352 2468
rect 7978 2396 8006 2424
rect 6438 2346 7050 2374
rect 7978 2270 8006 2298
rect 6438 2200 6872 2228
rect 7978 2044 8006 2072
rect 7978 1004 8006 1032
rect 6438 848 6872 876
rect 7978 778 8006 806
rect 6438 702 7050 730
rect 7978 652 8006 680
rect 6704 608 7352 610
rect 6438 582 7352 608
rect 6438 580 6732 582
<< metal2 >>
rect 6616 98418 6830 98446
rect 18 0 46 36952
rect 102 0 130 36952
rect 186 0 214 36952
rect 270 0 298 36952
rect 354 0 382 36952
rect 438 0 466 36952
rect 522 0 550 36952
rect 606 0 634 36952
<< metal3 >>
rect 6400 98395 6532 98469
rect 7940 98395 8072 98469
rect 6400 96857 6532 96931
rect 7940 96857 8072 96931
rect 6400 95319 6532 95393
rect 7940 95319 8072 95393
rect 6400 93781 6532 93855
rect 7940 93781 8072 93855
rect 6400 92243 6532 92317
rect 7940 92243 8072 92317
rect 6400 90705 6532 90779
rect 7940 90705 8072 90779
rect 6400 89167 6532 89241
rect 7940 89167 8072 89241
rect 6400 87629 6532 87703
rect 7940 87629 8072 87703
rect 6400 86091 6532 86165
rect 7940 86091 8072 86165
rect 6400 84553 6532 84627
rect 7940 84553 8072 84627
rect 6400 83015 6532 83089
rect 7940 83015 8072 83089
rect 6400 81477 6532 81551
rect 7940 81477 8072 81551
rect 6400 79939 6532 80013
rect 7940 79939 8072 80013
rect 6400 78401 6532 78475
rect 7940 78401 8072 78475
rect 6400 76863 6532 76937
rect 7940 76863 8072 76937
rect 6400 75325 6532 75399
rect 7940 75325 8072 75399
rect 6400 73787 6532 73861
rect 7940 73787 8072 73861
rect 6400 72249 6532 72323
rect 7940 72249 8072 72323
rect 6400 70711 6532 70785
rect 7940 70711 8072 70785
rect 6400 69173 6532 69247
rect 7940 69173 8072 69247
rect 6400 67635 6532 67709
rect 7940 67635 8072 67709
rect 6400 66097 6532 66171
rect 7940 66097 8072 66171
rect 6400 64559 6532 64633
rect 7940 64559 8072 64633
rect 6400 63021 6532 63095
rect 7940 63021 8072 63095
rect 6400 61483 6532 61557
rect 7940 61483 8072 61557
rect 6400 59945 6532 60019
rect 7940 59945 8072 60019
rect 6400 58407 6532 58481
rect 7940 58407 8072 58481
rect 6400 56869 6532 56943
rect 7940 56869 8072 56943
rect 6400 55331 6532 55405
rect 7940 55331 8072 55405
rect 6400 53793 6532 53867
rect 7940 53793 8072 53867
rect 6400 52255 6532 52329
rect 7940 52255 8072 52329
rect 6400 50717 6532 50791
rect 7940 50717 8072 50791
rect 6400 49179 6532 49253
rect 7940 49179 8072 49253
rect 6400 47641 6532 47715
rect 7940 47641 8072 47715
rect 6400 46103 6532 46177
rect 7940 46103 8072 46177
rect 6400 44565 6532 44639
rect 7940 44565 8072 44639
rect 6400 43027 6532 43101
rect 7940 43027 8072 43101
rect 6400 41489 6532 41563
rect 7940 41489 8072 41563
rect 6400 39951 6532 40025
rect 7940 39951 8072 40025
rect 6400 38413 6532 38487
rect 7940 38413 8072 38487
rect 1044 36915 1176 36989
rect 2084 36915 2216 36989
rect 6400 36875 6532 36949
rect 7940 36875 8072 36949
rect 1044 35375 1176 35449
rect 2084 35375 2216 35449
rect 6400 35337 6532 35411
rect 7940 35337 8072 35411
rect 1044 33835 1176 33909
rect 2084 33835 2216 33909
rect 6400 33799 6532 33873
rect 7940 33799 8072 33873
rect 1044 32295 1176 32369
rect 2084 32295 2216 32369
rect 6400 32261 6532 32335
rect 7940 32261 8072 32335
rect 1044 30755 1176 30829
rect 2084 30755 2216 30829
rect 6400 30723 6532 30797
rect 7940 30723 8072 30797
rect 1044 29215 1176 29289
rect 2084 29215 2216 29289
rect 6400 29185 6532 29259
rect 7940 29185 8072 29259
rect 1044 27675 1176 27749
rect 2084 27675 2216 27749
rect 6400 27647 6532 27721
rect 7940 27647 8072 27721
rect 1044 26135 1176 26209
rect 2084 26135 2216 26209
rect 6400 26109 6532 26183
rect 7940 26109 8072 26183
rect 1044 24595 1176 24669
rect 2084 24595 2216 24669
rect 6400 24571 6532 24645
rect 7940 24571 8072 24645
rect 6400 23033 6532 23107
rect 7940 23033 8072 23107
rect 1044 21519 1176 21593
rect 2084 21519 2216 21593
rect 6400 21495 6532 21569
rect 7940 21495 8072 21569
rect 1044 19979 1176 20053
rect 2084 19979 2216 20053
rect 6400 19957 6532 20031
rect 7940 19957 8072 20031
rect 1044 18439 1176 18513
rect 2084 18439 2216 18513
rect 6400 18419 6532 18493
rect 7940 18419 8072 18493
rect 1044 16899 1176 16973
rect 2084 16899 2216 16973
rect 6400 16881 6532 16955
rect 7940 16881 8072 16955
rect 1044 15359 1176 15433
rect 2084 15359 2216 15433
rect 6400 15343 6532 15417
rect 7940 15343 8072 15417
rect 1044 13819 1176 13893
rect 2084 13819 2216 13893
rect 6400 13805 6532 13879
rect 7940 13805 8072 13879
rect 1044 12279 1176 12353
rect 2084 12279 2216 12353
rect 6400 12267 6532 12341
rect 7940 12267 8072 12341
rect 1044 10739 1176 10813
rect 2084 10739 2216 10813
rect 6400 10729 6532 10803
rect 7940 10729 8072 10803
rect 1044 9199 1176 9273
rect 2084 9199 2216 9273
rect 6400 9191 6532 9265
rect 7940 9191 8072 9265
rect 6400 7653 6532 7727
rect 7940 7653 8072 7727
rect 1392 6123 1524 6197
rect 2264 6123 2396 6197
rect 6400 6115 6532 6189
rect 7940 6115 8072 6189
rect 1392 4583 1524 4657
rect 2264 4583 2396 4657
rect 6400 4577 6532 4651
rect 7940 4577 8072 4651
rect 1392 3043 1524 3117
rect 2264 3043 2396 3117
rect 6400 3039 6532 3113
rect 7940 3039 8072 3113
rect 1392 1503 1524 1577
rect 2264 1503 2396 1577
rect 6400 1501 6532 1575
rect 7940 1501 8072 1575
rect 1392 -37 1524 37
rect 2264 -37 2396 37
rect 6400 -37 6532 37
rect 7940 -37 8072 37
use wordline_driver_array  wordline_driver_array_0
timestamp 1644969367
transform 1 0 6802 0 1 0
box 0 -42 1270 98474
use hierarchical_decoder  hierarchical_decoder_0
timestamp 1644969367
transform 1 0 0 0 1 0
box 0 -42 6532 98474
<< labels >>
rlabel metal2 s 18 0 46 36952 4 addr0
rlabel metal2 s 102 0 130 36952 4 addr1
rlabel metal2 s 186 0 214 36952 4 addr2
rlabel metal2 s 270 0 298 36952 4 addr3
rlabel metal2 s 354 0 382 36952 4 addr4
rlabel metal2 s 438 0 466 36952 4 addr5
rlabel metal2 s 522 0 550 36952 4 addr6
rlabel metal2 s 606 0 634 36952 4 addr7
rlabel metal1 s 7978 778 8006 806 4 rwl0_0
rlabel metal1 s 7978 1004 8006 1032 4 rwl1_0
rlabel metal1 s 7978 652 8006 680 4 wwl0_0
rlabel metal1 s 7978 2270 8006 2298 4 rwl0_1
rlabel metal1 s 7978 2044 8006 2072 4 rwl1_1
rlabel metal1 s 7978 2396 8006 2424 4 wwl0_1
rlabel metal1 s 7978 3854 8006 3882 4 rwl0_2
rlabel metal1 s 7978 4080 8006 4108 4 rwl1_2
rlabel metal1 s 7978 3728 8006 3756 4 wwl0_2
rlabel metal1 s 7978 5346 8006 5374 4 rwl0_3
rlabel metal1 s 7978 5120 8006 5148 4 rwl1_3
rlabel metal1 s 7978 5472 8006 5500 4 wwl0_3
rlabel metal1 s 7978 6930 8006 6958 4 rwl0_4
rlabel metal1 s 7978 7156 8006 7184 4 rwl1_4
rlabel metal1 s 7978 6804 8006 6832 4 wwl0_4
rlabel metal1 s 7978 8422 8006 8450 4 rwl0_5
rlabel metal1 s 7978 8196 8006 8224 4 rwl1_5
rlabel metal1 s 7978 8548 8006 8576 4 wwl0_5
rlabel metal1 s 7978 10006 8006 10034 4 rwl0_6
rlabel metal1 s 7978 10232 8006 10260 4 rwl1_6
rlabel metal1 s 7978 9880 8006 9908 4 wwl0_6
rlabel metal1 s 7978 11498 8006 11526 4 rwl0_7
rlabel metal1 s 7978 11272 8006 11300 4 rwl1_7
rlabel metal1 s 7978 11624 8006 11652 4 wwl0_7
rlabel metal1 s 7978 13082 8006 13110 4 rwl0_8
rlabel metal1 s 7978 13308 8006 13336 4 rwl1_8
rlabel metal1 s 7978 12956 8006 12984 4 wwl0_8
rlabel metal1 s 7978 14574 8006 14602 4 rwl0_9
rlabel metal1 s 7978 14348 8006 14376 4 rwl1_9
rlabel metal1 s 7978 14700 8006 14728 4 wwl0_9
rlabel metal1 s 7978 16158 8006 16186 4 rwl0_10
rlabel metal1 s 7978 16384 8006 16412 4 rwl1_10
rlabel metal1 s 7978 16032 8006 16060 4 wwl0_10
rlabel metal1 s 7978 17650 8006 17678 4 rwl0_11
rlabel metal1 s 7978 17424 8006 17452 4 rwl1_11
rlabel metal1 s 7978 17776 8006 17804 4 wwl0_11
rlabel metal1 s 7978 19234 8006 19262 4 rwl0_12
rlabel metal1 s 7978 19460 8006 19488 4 rwl1_12
rlabel metal1 s 7978 19108 8006 19136 4 wwl0_12
rlabel metal1 s 7978 20726 8006 20754 4 rwl0_13
rlabel metal1 s 7978 20500 8006 20528 4 rwl1_13
rlabel metal1 s 7978 20852 8006 20880 4 wwl0_13
rlabel metal1 s 7978 22310 8006 22338 4 rwl0_14
rlabel metal1 s 7978 22536 8006 22564 4 rwl1_14
rlabel metal1 s 7978 22184 8006 22212 4 wwl0_14
rlabel metal1 s 7978 23802 8006 23830 4 rwl0_15
rlabel metal1 s 7978 23576 8006 23604 4 rwl1_15
rlabel metal1 s 7978 23928 8006 23956 4 wwl0_15
rlabel metal1 s 7978 25386 8006 25414 4 rwl0_16
rlabel metal1 s 7978 25612 8006 25640 4 rwl1_16
rlabel metal1 s 7978 25260 8006 25288 4 wwl0_16
rlabel metal1 s 7978 26878 8006 26906 4 rwl0_17
rlabel metal1 s 7978 26652 8006 26680 4 rwl1_17
rlabel metal1 s 7978 27004 8006 27032 4 wwl0_17
rlabel metal1 s 7978 28462 8006 28490 4 rwl0_18
rlabel metal1 s 7978 28688 8006 28716 4 rwl1_18
rlabel metal1 s 7978 28336 8006 28364 4 wwl0_18
rlabel metal1 s 7978 29954 8006 29982 4 rwl0_19
rlabel metal1 s 7978 29728 8006 29756 4 rwl1_19
rlabel metal1 s 7978 30080 8006 30108 4 wwl0_19
rlabel metal1 s 7978 31538 8006 31566 4 rwl0_20
rlabel metal1 s 7978 31764 8006 31792 4 rwl1_20
rlabel metal1 s 7978 31412 8006 31440 4 wwl0_20
rlabel metal1 s 7978 33030 8006 33058 4 rwl0_21
rlabel metal1 s 7978 32804 8006 32832 4 rwl1_21
rlabel metal1 s 7978 33156 8006 33184 4 wwl0_21
rlabel metal1 s 7978 34614 8006 34642 4 rwl0_22
rlabel metal1 s 7978 34840 8006 34868 4 rwl1_22
rlabel metal1 s 7978 34488 8006 34516 4 wwl0_22
rlabel metal1 s 7978 36106 8006 36134 4 rwl0_23
rlabel metal1 s 7978 35880 8006 35908 4 rwl1_23
rlabel metal1 s 7978 36232 8006 36260 4 wwl0_23
rlabel metal1 s 7978 37690 8006 37718 4 rwl0_24
rlabel metal1 s 7978 37916 8006 37944 4 rwl1_24
rlabel metal1 s 7978 37564 8006 37592 4 wwl0_24
rlabel metal1 s 7978 39182 8006 39210 4 rwl0_25
rlabel metal1 s 7978 38956 8006 38984 4 rwl1_25
rlabel metal1 s 7978 39308 8006 39336 4 wwl0_25
rlabel metal1 s 7978 40766 8006 40794 4 rwl0_26
rlabel metal1 s 7978 40992 8006 41020 4 rwl1_26
rlabel metal1 s 7978 40640 8006 40668 4 wwl0_26
rlabel metal1 s 7978 42258 8006 42286 4 rwl0_27
rlabel metal1 s 7978 42032 8006 42060 4 rwl1_27
rlabel metal1 s 7978 42384 8006 42412 4 wwl0_27
rlabel metal1 s 7978 43842 8006 43870 4 rwl0_28
rlabel metal1 s 7978 44068 8006 44096 4 rwl1_28
rlabel metal1 s 7978 43716 8006 43744 4 wwl0_28
rlabel metal1 s 7978 45334 8006 45362 4 rwl0_29
rlabel metal1 s 7978 45108 8006 45136 4 rwl1_29
rlabel metal1 s 7978 45460 8006 45488 4 wwl0_29
rlabel metal1 s 7978 46918 8006 46946 4 rwl0_30
rlabel metal1 s 7978 47144 8006 47172 4 rwl1_30
rlabel metal1 s 7978 46792 8006 46820 4 wwl0_30
rlabel metal1 s 7978 48410 8006 48438 4 rwl0_31
rlabel metal1 s 7978 48184 8006 48212 4 rwl1_31
rlabel metal1 s 7978 48536 8006 48564 4 wwl0_31
rlabel metal1 s 7978 49994 8006 50022 4 rwl0_32
rlabel metal1 s 7978 50220 8006 50248 4 rwl1_32
rlabel metal1 s 7978 49868 8006 49896 4 wwl0_32
rlabel metal1 s 7978 51486 8006 51514 4 rwl0_33
rlabel metal1 s 7978 51260 8006 51288 4 rwl1_33
rlabel metal1 s 7978 51612 8006 51640 4 wwl0_33
rlabel metal1 s 7978 53070 8006 53098 4 rwl0_34
rlabel metal1 s 7978 53296 8006 53324 4 rwl1_34
rlabel metal1 s 7978 52944 8006 52972 4 wwl0_34
rlabel metal1 s 7978 54562 8006 54590 4 rwl0_35
rlabel metal1 s 7978 54336 8006 54364 4 rwl1_35
rlabel metal1 s 7978 54688 8006 54716 4 wwl0_35
rlabel metal1 s 7978 56146 8006 56174 4 rwl0_36
rlabel metal1 s 7978 56372 8006 56400 4 rwl1_36
rlabel metal1 s 7978 56020 8006 56048 4 wwl0_36
rlabel metal1 s 7978 57638 8006 57666 4 rwl0_37
rlabel metal1 s 7978 57412 8006 57440 4 rwl1_37
rlabel metal1 s 7978 57764 8006 57792 4 wwl0_37
rlabel metal1 s 7978 59222 8006 59250 4 rwl0_38
rlabel metal1 s 7978 59448 8006 59476 4 rwl1_38
rlabel metal1 s 7978 59096 8006 59124 4 wwl0_38
rlabel metal1 s 7978 60714 8006 60742 4 rwl0_39
rlabel metal1 s 7978 60488 8006 60516 4 rwl1_39
rlabel metal1 s 7978 60840 8006 60868 4 wwl0_39
rlabel metal1 s 7978 62298 8006 62326 4 rwl0_40
rlabel metal1 s 7978 62524 8006 62552 4 rwl1_40
rlabel metal1 s 7978 62172 8006 62200 4 wwl0_40
rlabel metal1 s 7978 63790 8006 63818 4 rwl0_41
rlabel metal1 s 7978 63564 8006 63592 4 rwl1_41
rlabel metal1 s 7978 63916 8006 63944 4 wwl0_41
rlabel metal1 s 7978 65374 8006 65402 4 rwl0_42
rlabel metal1 s 7978 65600 8006 65628 4 rwl1_42
rlabel metal1 s 7978 65248 8006 65276 4 wwl0_42
rlabel metal1 s 7978 66866 8006 66894 4 rwl0_43
rlabel metal1 s 7978 66640 8006 66668 4 rwl1_43
rlabel metal1 s 7978 66992 8006 67020 4 wwl0_43
rlabel metal1 s 7978 68450 8006 68478 4 rwl0_44
rlabel metal1 s 7978 68676 8006 68704 4 rwl1_44
rlabel metal1 s 7978 68324 8006 68352 4 wwl0_44
rlabel metal1 s 7978 69942 8006 69970 4 rwl0_45
rlabel metal1 s 7978 69716 8006 69744 4 rwl1_45
rlabel metal1 s 7978 70068 8006 70096 4 wwl0_45
rlabel metal1 s 7978 71526 8006 71554 4 rwl0_46
rlabel metal1 s 7978 71752 8006 71780 4 rwl1_46
rlabel metal1 s 7978 71400 8006 71428 4 wwl0_46
rlabel metal1 s 7978 73018 8006 73046 4 rwl0_47
rlabel metal1 s 7978 72792 8006 72820 4 rwl1_47
rlabel metal1 s 7978 73144 8006 73172 4 wwl0_47
rlabel metal1 s 7978 74602 8006 74630 4 rwl0_48
rlabel metal1 s 7978 74828 8006 74856 4 rwl1_48
rlabel metal1 s 7978 74476 8006 74504 4 wwl0_48
rlabel metal1 s 7978 76094 8006 76122 4 rwl0_49
rlabel metal1 s 7978 75868 8006 75896 4 rwl1_49
rlabel metal1 s 7978 76220 8006 76248 4 wwl0_49
rlabel metal1 s 7978 77678 8006 77706 4 rwl0_50
rlabel metal1 s 7978 77904 8006 77932 4 rwl1_50
rlabel metal1 s 7978 77552 8006 77580 4 wwl0_50
rlabel metal1 s 7978 79170 8006 79198 4 rwl0_51
rlabel metal1 s 7978 78944 8006 78972 4 rwl1_51
rlabel metal1 s 7978 79296 8006 79324 4 wwl0_51
rlabel metal1 s 7978 80754 8006 80782 4 rwl0_52
rlabel metal1 s 7978 80980 8006 81008 4 rwl1_52
rlabel metal1 s 7978 80628 8006 80656 4 wwl0_52
rlabel metal1 s 7978 82246 8006 82274 4 rwl0_53
rlabel metal1 s 7978 82020 8006 82048 4 rwl1_53
rlabel metal1 s 7978 82372 8006 82400 4 wwl0_53
rlabel metal1 s 7978 83830 8006 83858 4 rwl0_54
rlabel metal1 s 7978 84056 8006 84084 4 rwl1_54
rlabel metal1 s 7978 83704 8006 83732 4 wwl0_54
rlabel metal1 s 7978 85322 8006 85350 4 rwl0_55
rlabel metal1 s 7978 85096 8006 85124 4 rwl1_55
rlabel metal1 s 7978 85448 8006 85476 4 wwl0_55
rlabel metal1 s 7978 86906 8006 86934 4 rwl0_56
rlabel metal1 s 7978 87132 8006 87160 4 rwl1_56
rlabel metal1 s 7978 86780 8006 86808 4 wwl0_56
rlabel metal1 s 7978 88398 8006 88426 4 rwl0_57
rlabel metal1 s 7978 88172 8006 88200 4 rwl1_57
rlabel metal1 s 7978 88524 8006 88552 4 wwl0_57
rlabel metal1 s 7978 89982 8006 90010 4 rwl0_58
rlabel metal1 s 7978 90208 8006 90236 4 rwl1_58
rlabel metal1 s 7978 89856 8006 89884 4 wwl0_58
rlabel metal1 s 7978 91474 8006 91502 4 rwl0_59
rlabel metal1 s 7978 91248 8006 91276 4 rwl1_59
rlabel metal1 s 7978 91600 8006 91628 4 wwl0_59
rlabel metal1 s 7978 93058 8006 93086 4 rwl0_60
rlabel metal1 s 7978 93284 8006 93312 4 rwl1_60
rlabel metal1 s 7978 92932 8006 92960 4 wwl0_60
rlabel metal1 s 7978 94550 8006 94578 4 rwl0_61
rlabel metal1 s 7978 94324 8006 94352 4 rwl1_61
rlabel metal1 s 7978 94676 8006 94704 4 wwl0_61
rlabel metal1 s 7978 96134 8006 96162 4 rwl0_62
rlabel metal1 s 7978 96360 8006 96388 4 rwl1_62
rlabel metal1 s 7978 96008 8006 96036 4 wwl0_62
rlabel metal1 s 7978 97626 8006 97654 4 rwl0_63
rlabel metal1 s 7978 97400 8006 97428 4 rwl1_63
rlabel metal1 s 7978 97752 8006 97780 4 wwl0_63
rlabel metal2 s 6802 98418 6830 98446 4 wl_en
rlabel metal3 s 7940 35337 8072 35411 4 vdd
rlabel metal3 s 1392 1503 1524 1577 4 vdd
rlabel metal3 s 7940 63021 8072 63095 4 vdd
rlabel metal3 s 7940 75325 8072 75399 4 vdd
rlabel metal3 s 6400 84553 6532 84627 4 vdd
rlabel metal3 s 6400 63021 6532 63095 4 vdd
rlabel metal3 s 6400 59945 6532 60019 4 vdd
rlabel metal3 s 1392 4583 1524 4657 4 vdd
rlabel metal3 s 6400 19957 6532 20031 4 vdd
rlabel metal3 s 2084 13819 2216 13893 4 vdd
rlabel metal3 s 7940 19957 8072 20031 4 vdd
rlabel metal3 s 7940 84553 8072 84627 4 vdd
rlabel metal3 s 6400 66097 6532 66171 4 vdd
rlabel metal3 s 1044 32295 1176 32369 4 vdd
rlabel metal3 s 6400 35337 6532 35411 4 vdd
rlabel metal3 s 7940 44565 8072 44639 4 vdd
rlabel metal3 s 7940 10729 8072 10803 4 vdd
rlabel metal3 s 6400 10729 6532 10803 4 vdd
rlabel metal3 s 7940 93781 8072 93855 4 vdd
rlabel metal3 s 1044 19979 1176 20053 4 vdd
rlabel metal3 s 2084 35375 2216 35449 4 vdd
rlabel metal3 s 7940 53793 8072 53867 4 vdd
rlabel metal3 s 2084 16899 2216 16973 4 vdd
rlabel metal3 s 6400 38413 6532 38487 4 vdd
rlabel metal3 s 7940 26109 8072 26183 4 vdd
rlabel metal3 s 7940 87629 8072 87703 4 vdd
rlabel metal3 s 7940 7653 8072 7727 4 vdd
rlabel metal3 s 7940 23033 8072 23107 4 vdd
rlabel metal3 s 6400 87629 6532 87703 4 vdd
rlabel metal3 s 6400 47641 6532 47715 4 vdd
rlabel metal3 s 6400 26109 6532 26183 4 vdd
rlabel metal3 s 7940 96857 8072 96931 4 vdd
rlabel metal3 s 6400 41489 6532 41563 4 vdd
rlabel metal3 s 7940 69173 8072 69247 4 vdd
rlabel metal3 s 6400 16881 6532 16955 4 vdd
rlabel metal3 s 7940 59945 8072 60019 4 vdd
rlabel metal3 s 1044 26135 1176 26209 4 vdd
rlabel metal3 s 6400 29185 6532 29259 4 vdd
rlabel metal3 s 6400 13805 6532 13879 4 vdd
rlabel metal3 s 6400 53793 6532 53867 4 vdd
rlabel metal3 s 6400 23033 6532 23107 4 vdd
rlabel metal3 s 7940 1501 8072 1575 4 vdd
rlabel metal3 s 7940 38413 8072 38487 4 vdd
rlabel metal3 s 7940 78401 8072 78475 4 vdd
rlabel metal3 s 1044 35375 1176 35449 4 vdd
rlabel metal3 s 6400 56869 6532 56943 4 vdd
rlabel metal3 s 7940 81477 8072 81551 4 vdd
rlabel metal3 s 7940 56869 8072 56943 4 vdd
rlabel metal3 s 1044 10739 1176 10813 4 vdd
rlabel metal3 s 6400 96857 6532 96931 4 vdd
rlabel metal3 s 7940 72249 8072 72323 4 vdd
rlabel metal3 s 2264 4583 2396 4657 4 vdd
rlabel metal3 s 1044 13819 1176 13893 4 vdd
rlabel metal3 s 2084 19979 2216 20053 4 vdd
rlabel metal3 s 7940 90705 8072 90779 4 vdd
rlabel metal3 s 7940 66097 8072 66171 4 vdd
rlabel metal3 s 7940 32261 8072 32335 4 vdd
rlabel metal3 s 7940 16881 8072 16955 4 vdd
rlabel metal3 s 6400 32261 6532 32335 4 vdd
rlabel metal3 s 6400 69173 6532 69247 4 vdd
rlabel metal3 s 2084 10739 2216 10813 4 vdd
rlabel metal3 s 6400 1501 6532 1575 4 vdd
rlabel metal3 s 6400 4577 6532 4651 4 vdd
rlabel metal3 s 6400 93781 6532 93855 4 vdd
rlabel metal3 s 6400 72249 6532 72323 4 vdd
rlabel metal3 s 2264 1503 2396 1577 4 vdd
rlabel metal3 s 6400 90705 6532 90779 4 vdd
rlabel metal3 s 2084 32295 2216 32369 4 vdd
rlabel metal3 s 7940 13805 8072 13879 4 vdd
rlabel metal3 s 6400 75325 6532 75399 4 vdd
rlabel metal3 s 7940 29185 8072 29259 4 vdd
rlabel metal3 s 1044 16899 1176 16973 4 vdd
rlabel metal3 s 6400 81477 6532 81551 4 vdd
rlabel metal3 s 7940 47641 8072 47715 4 vdd
rlabel metal3 s 6400 7653 6532 7727 4 vdd
rlabel metal3 s 7940 50717 8072 50791 4 vdd
rlabel metal3 s 6400 78401 6532 78475 4 vdd
rlabel metal3 s 2084 29215 2216 29289 4 vdd
rlabel metal3 s 6400 44565 6532 44639 4 vdd
rlabel metal3 s 6400 50717 6532 50791 4 vdd
rlabel metal3 s 7940 4577 8072 4651 4 vdd
rlabel metal3 s 7940 41489 8072 41563 4 vdd
rlabel metal3 s 2084 26135 2216 26209 4 vdd
rlabel metal3 s 1044 29215 1176 29289 4 vdd
rlabel metal3 s 7940 33799 8072 33873 4 gnd
rlabel metal3 s 6400 49179 6532 49253 4 gnd
rlabel metal3 s 7940 6115 8072 6189 4 gnd
rlabel metal3 s 7940 3039 8072 3113 4 gnd
rlabel metal3 s 6400 46103 6532 46177 4 gnd
rlabel metal3 s 6400 58407 6532 58481 4 gnd
rlabel metal3 s 2084 33835 2216 33909 4 gnd
rlabel metal3 s 7940 -37 8072 37 4 gnd
rlabel metal3 s 6400 27647 6532 27721 4 gnd
rlabel metal3 s 1044 15359 1176 15433 4 gnd
rlabel metal3 s 2084 36915 2216 36989 4 gnd
rlabel metal3 s 7940 55331 8072 55405 4 gnd
rlabel metal3 s 2264 3043 2396 3117 4 gnd
rlabel metal3 s 6400 89167 6532 89241 4 gnd
rlabel metal3 s 6400 -37 6532 37 4 gnd
rlabel metal3 s 7940 95319 8072 95393 4 gnd
rlabel metal3 s 6400 86091 6532 86165 4 gnd
rlabel metal3 s 2084 27675 2216 27749 4 gnd
rlabel metal3 s 2264 -37 2396 37 4 gnd
rlabel metal3 s 2084 12279 2216 12353 4 gnd
rlabel metal3 s 1044 33835 1176 33909 4 gnd
rlabel metal3 s 6400 73787 6532 73861 4 gnd
rlabel metal3 s 1044 27675 1176 27749 4 gnd
rlabel metal3 s 2264 6123 2396 6197 4 gnd
rlabel metal3 s 1392 -37 1524 37 4 gnd
rlabel metal3 s 6400 79939 6532 80013 4 gnd
rlabel metal3 s 1044 30755 1176 30829 4 gnd
rlabel metal3 s 1392 3043 1524 3117 4 gnd
rlabel metal3 s 7940 24571 8072 24645 4 gnd
rlabel metal3 s 6400 52255 6532 52329 4 gnd
rlabel metal3 s 7940 83015 8072 83089 4 gnd
rlabel metal3 s 2084 30755 2216 30829 4 gnd
rlabel metal3 s 1044 21519 1176 21593 4 gnd
rlabel metal3 s 7940 21495 8072 21569 4 gnd
rlabel metal3 s 7940 15343 8072 15417 4 gnd
rlabel metal3 s 7940 58407 8072 58481 4 gnd
rlabel metal3 s 7940 43027 8072 43101 4 gnd
rlabel metal3 s 6400 12267 6532 12341 4 gnd
rlabel metal3 s 6400 21495 6532 21569 4 gnd
rlabel metal3 s 2084 21519 2216 21593 4 gnd
rlabel metal3 s 6400 3039 6532 3113 4 gnd
rlabel metal3 s 2084 9199 2216 9273 4 gnd
rlabel metal3 s 2084 18439 2216 18513 4 gnd
rlabel metal3 s 6400 92243 6532 92317 4 gnd
rlabel metal3 s 7940 30723 8072 30797 4 gnd
rlabel metal3 s 6400 98395 6532 98469 4 gnd
rlabel metal3 s 1044 24595 1176 24669 4 gnd
rlabel metal3 s 7940 64559 8072 64633 4 gnd
rlabel metal3 s 6400 9191 6532 9265 4 gnd
rlabel metal3 s 7940 98395 8072 98469 4 gnd
rlabel metal3 s 7940 76863 8072 76937 4 gnd
rlabel metal3 s 7940 49179 8072 49253 4 gnd
rlabel metal3 s 1044 36915 1176 36989 4 gnd
rlabel metal3 s 6400 24571 6532 24645 4 gnd
rlabel metal3 s 1044 18439 1176 18513 4 gnd
rlabel metal3 s 7940 39951 8072 40025 4 gnd
rlabel metal3 s 7940 12267 8072 12341 4 gnd
rlabel metal3 s 7940 27647 8072 27721 4 gnd
rlabel metal3 s 6400 64559 6532 64633 4 gnd
rlabel metal3 s 7940 9191 8072 9265 4 gnd
rlabel metal3 s 7940 86091 8072 86165 4 gnd
rlabel metal3 s 6400 15343 6532 15417 4 gnd
rlabel metal3 s 7940 79939 8072 80013 4 gnd
rlabel metal3 s 6400 76863 6532 76937 4 gnd
rlabel metal3 s 7940 92243 8072 92317 4 gnd
rlabel metal3 s 1044 9199 1176 9273 4 gnd
rlabel metal3 s 6400 39951 6532 40025 4 gnd
rlabel metal3 s 7940 46103 8072 46177 4 gnd
rlabel metal3 s 6400 70711 6532 70785 4 gnd
rlabel metal3 s 6400 36875 6532 36949 4 gnd
rlabel metal3 s 6400 6115 6532 6189 4 gnd
rlabel metal3 s 6400 95319 6532 95393 4 gnd
rlabel metal3 s 7940 89167 8072 89241 4 gnd
rlabel metal3 s 2084 24595 2216 24669 4 gnd
rlabel metal3 s 6400 61483 6532 61557 4 gnd
rlabel metal3 s 7940 73787 8072 73861 4 gnd
rlabel metal3 s 6400 18419 6532 18493 4 gnd
rlabel metal3 s 7940 18419 8072 18493 4 gnd
rlabel metal3 s 6400 67635 6532 67709 4 gnd
rlabel metal3 s 1392 6123 1524 6197 4 gnd
rlabel metal3 s 6400 43027 6532 43101 4 gnd
rlabel metal3 s 7940 52255 8072 52329 4 gnd
rlabel metal3 s 6400 30723 6532 30797 4 gnd
rlabel metal3 s 7940 36875 8072 36949 4 gnd
rlabel metal3 s 6400 83015 6532 83089 4 gnd
rlabel metal3 s 7940 70711 8072 70785 4 gnd
rlabel metal3 s 1044 12279 1176 12353 4 gnd
rlabel metal3 s 6400 55331 6532 55405 4 gnd
rlabel metal3 s 6400 33799 6532 33873 4 gnd
rlabel metal3 s 7940 61483 8072 61557 4 gnd
rlabel metal3 s 2084 15359 2216 15433 4 gnd
rlabel metal3 s 7940 67635 8072 67709 4 gnd
<< properties >>
string FIXED_BBOX 0 0 8042 98460
string GDS_FILE sram_0rw2r1w_32_128_sky130A.gds
string GDS_END 2861536
string GDS_START 2728950
<< end >>
