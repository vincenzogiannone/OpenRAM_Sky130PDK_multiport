magic
tech sky130A
magscale 1 2
timestamp 1643678851
<< checkpaint >>
rect -1296 -1277 1647 2155
<< nwell >>
rect -36 402 387 895
<< locali >>
rect 0 821 351 855
rect 48 344 114 410
rect 179 360 213 394
rect 0 -17 351 17
use pinv_0  pinv_0_0
timestamp 1643678851
transform 1 0 0 0 1 0
box -36 -17 387 895
<< labels >>
rlabel locali s 196 377 196 377 4 Z
rlabel locali s 81 377 81 377 4 A
rlabel locali s 175 0 175 0 4 gnd
rlabel locali s 175 838 175 838 4 vdd
<< properties >>
string FIXED_BBOX 0 0 351 838
string GDS_FILE sram_0rw2r1w_16_128_sky130A.gds
string GDS_END 1999658
string GDS_START 1998814
<< end >>
