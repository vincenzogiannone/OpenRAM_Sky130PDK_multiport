magic
tech sky130A
magscale 1 2
timestamp 1643593061
<< checkpaint >>
rect -1260 -1260 27000 36482
<< dnwell >>
rect 1618 1524 24198 33934
<< nwell >>
rect 1534 33850 24282 34018
rect 1534 1608 1702 33850
rect 24114 1608 24282 33850
rect 1534 1440 24282 1608
<< nsubdiff >>
rect 1929 33951 1979 33975
rect 1929 33917 1937 33951
rect 1971 33917 1979 33951
rect 1929 33893 1979 33917
rect 2265 33951 2315 33975
rect 2265 33917 2273 33951
rect 2307 33917 2315 33951
rect 2265 33893 2315 33917
rect 2601 33951 2651 33975
rect 2601 33917 2609 33951
rect 2643 33917 2651 33951
rect 2601 33893 2651 33917
rect 2937 33951 2987 33975
rect 2937 33917 2945 33951
rect 2979 33917 2987 33951
rect 2937 33893 2987 33917
rect 3273 33951 3323 33975
rect 3273 33917 3281 33951
rect 3315 33917 3323 33951
rect 3273 33893 3323 33917
rect 3609 33951 3659 33975
rect 3609 33917 3617 33951
rect 3651 33917 3659 33951
rect 3609 33893 3659 33917
rect 3945 33951 3995 33975
rect 3945 33917 3953 33951
rect 3987 33917 3995 33951
rect 3945 33893 3995 33917
rect 4281 33951 4331 33975
rect 4281 33917 4289 33951
rect 4323 33917 4331 33951
rect 4281 33893 4331 33917
rect 4617 33951 4667 33975
rect 4617 33917 4625 33951
rect 4659 33917 4667 33951
rect 4617 33893 4667 33917
rect 4953 33951 5003 33975
rect 4953 33917 4961 33951
rect 4995 33917 5003 33951
rect 4953 33893 5003 33917
rect 5289 33951 5339 33975
rect 5289 33917 5297 33951
rect 5331 33917 5339 33951
rect 5289 33893 5339 33917
rect 5625 33951 5675 33975
rect 5625 33917 5633 33951
rect 5667 33917 5675 33951
rect 5625 33893 5675 33917
rect 5961 33951 6011 33975
rect 5961 33917 5969 33951
rect 6003 33917 6011 33951
rect 5961 33893 6011 33917
rect 6297 33951 6347 33975
rect 6297 33917 6305 33951
rect 6339 33917 6347 33951
rect 6297 33893 6347 33917
rect 6633 33951 6683 33975
rect 6633 33917 6641 33951
rect 6675 33917 6683 33951
rect 6633 33893 6683 33917
rect 6969 33951 7019 33975
rect 6969 33917 6977 33951
rect 7011 33917 7019 33951
rect 6969 33893 7019 33917
rect 7305 33951 7355 33975
rect 7305 33917 7313 33951
rect 7347 33917 7355 33951
rect 7305 33893 7355 33917
rect 7641 33951 7691 33975
rect 7641 33917 7649 33951
rect 7683 33917 7691 33951
rect 7641 33893 7691 33917
rect 7977 33951 8027 33975
rect 7977 33917 7985 33951
rect 8019 33917 8027 33951
rect 7977 33893 8027 33917
rect 8313 33951 8363 33975
rect 8313 33917 8321 33951
rect 8355 33917 8363 33951
rect 8313 33893 8363 33917
rect 8649 33951 8699 33975
rect 8649 33917 8657 33951
rect 8691 33917 8699 33951
rect 8649 33893 8699 33917
rect 8985 33951 9035 33975
rect 8985 33917 8993 33951
rect 9027 33917 9035 33951
rect 8985 33893 9035 33917
rect 9321 33951 9371 33975
rect 9321 33917 9329 33951
rect 9363 33917 9371 33951
rect 9321 33893 9371 33917
rect 9657 33951 9707 33975
rect 9657 33917 9665 33951
rect 9699 33917 9707 33951
rect 9657 33893 9707 33917
rect 9993 33951 10043 33975
rect 9993 33917 10001 33951
rect 10035 33917 10043 33951
rect 9993 33893 10043 33917
rect 10329 33951 10379 33975
rect 10329 33917 10337 33951
rect 10371 33917 10379 33951
rect 10329 33893 10379 33917
rect 10665 33951 10715 33975
rect 10665 33917 10673 33951
rect 10707 33917 10715 33951
rect 10665 33893 10715 33917
rect 11001 33951 11051 33975
rect 11001 33917 11009 33951
rect 11043 33917 11051 33951
rect 11001 33893 11051 33917
rect 11337 33951 11387 33975
rect 11337 33917 11345 33951
rect 11379 33917 11387 33951
rect 11337 33893 11387 33917
rect 11673 33951 11723 33975
rect 11673 33917 11681 33951
rect 11715 33917 11723 33951
rect 11673 33893 11723 33917
rect 12009 33951 12059 33975
rect 12009 33917 12017 33951
rect 12051 33917 12059 33951
rect 12009 33893 12059 33917
rect 12345 33951 12395 33975
rect 12345 33917 12353 33951
rect 12387 33917 12395 33951
rect 12345 33893 12395 33917
rect 12681 33951 12731 33975
rect 12681 33917 12689 33951
rect 12723 33917 12731 33951
rect 12681 33893 12731 33917
rect 13017 33951 13067 33975
rect 13017 33917 13025 33951
rect 13059 33917 13067 33951
rect 13017 33893 13067 33917
rect 13353 33951 13403 33975
rect 13353 33917 13361 33951
rect 13395 33917 13403 33951
rect 13353 33893 13403 33917
rect 13689 33951 13739 33975
rect 13689 33917 13697 33951
rect 13731 33917 13739 33951
rect 13689 33893 13739 33917
rect 14025 33951 14075 33975
rect 14025 33917 14033 33951
rect 14067 33917 14075 33951
rect 14025 33893 14075 33917
rect 14361 33951 14411 33975
rect 14361 33917 14369 33951
rect 14403 33917 14411 33951
rect 14361 33893 14411 33917
rect 14697 33951 14747 33975
rect 14697 33917 14705 33951
rect 14739 33917 14747 33951
rect 14697 33893 14747 33917
rect 15033 33951 15083 33975
rect 15033 33917 15041 33951
rect 15075 33917 15083 33951
rect 15033 33893 15083 33917
rect 15369 33951 15419 33975
rect 15369 33917 15377 33951
rect 15411 33917 15419 33951
rect 15369 33893 15419 33917
rect 15705 33951 15755 33975
rect 15705 33917 15713 33951
rect 15747 33917 15755 33951
rect 15705 33893 15755 33917
rect 16041 33951 16091 33975
rect 16041 33917 16049 33951
rect 16083 33917 16091 33951
rect 16041 33893 16091 33917
rect 16377 33951 16427 33975
rect 16377 33917 16385 33951
rect 16419 33917 16427 33951
rect 16377 33893 16427 33917
rect 16713 33951 16763 33975
rect 16713 33917 16721 33951
rect 16755 33917 16763 33951
rect 16713 33893 16763 33917
rect 17049 33951 17099 33975
rect 17049 33917 17057 33951
rect 17091 33917 17099 33951
rect 17049 33893 17099 33917
rect 17385 33951 17435 33975
rect 17385 33917 17393 33951
rect 17427 33917 17435 33951
rect 17385 33893 17435 33917
rect 17721 33951 17771 33975
rect 17721 33917 17729 33951
rect 17763 33917 17771 33951
rect 17721 33893 17771 33917
rect 18057 33951 18107 33975
rect 18057 33917 18065 33951
rect 18099 33917 18107 33951
rect 18057 33893 18107 33917
rect 18393 33951 18443 33975
rect 18393 33917 18401 33951
rect 18435 33917 18443 33951
rect 18393 33893 18443 33917
rect 18729 33951 18779 33975
rect 18729 33917 18737 33951
rect 18771 33917 18779 33951
rect 18729 33893 18779 33917
rect 19065 33951 19115 33975
rect 19065 33917 19073 33951
rect 19107 33917 19115 33951
rect 19065 33893 19115 33917
rect 19401 33951 19451 33975
rect 19401 33917 19409 33951
rect 19443 33917 19451 33951
rect 19401 33893 19451 33917
rect 19737 33951 19787 33975
rect 19737 33917 19745 33951
rect 19779 33917 19787 33951
rect 19737 33893 19787 33917
rect 20073 33951 20123 33975
rect 20073 33917 20081 33951
rect 20115 33917 20123 33951
rect 20073 33893 20123 33917
rect 20409 33951 20459 33975
rect 20409 33917 20417 33951
rect 20451 33917 20459 33951
rect 20409 33893 20459 33917
rect 20745 33951 20795 33975
rect 20745 33917 20753 33951
rect 20787 33917 20795 33951
rect 20745 33893 20795 33917
rect 21081 33951 21131 33975
rect 21081 33917 21089 33951
rect 21123 33917 21131 33951
rect 21081 33893 21131 33917
rect 21417 33951 21467 33975
rect 21417 33917 21425 33951
rect 21459 33917 21467 33951
rect 21417 33893 21467 33917
rect 21753 33951 21803 33975
rect 21753 33917 21761 33951
rect 21795 33917 21803 33951
rect 21753 33893 21803 33917
rect 22089 33951 22139 33975
rect 22089 33917 22097 33951
rect 22131 33917 22139 33951
rect 22089 33893 22139 33917
rect 22425 33951 22475 33975
rect 22425 33917 22433 33951
rect 22467 33917 22475 33951
rect 22425 33893 22475 33917
rect 22761 33951 22811 33975
rect 22761 33917 22769 33951
rect 22803 33917 22811 33951
rect 22761 33893 22811 33917
rect 23097 33951 23147 33975
rect 23097 33917 23105 33951
rect 23139 33917 23147 33951
rect 23097 33893 23147 33917
rect 23433 33951 23483 33975
rect 23433 33917 23441 33951
rect 23475 33917 23483 33951
rect 23433 33893 23483 33917
rect 23769 33951 23819 33975
rect 23769 33917 23777 33951
rect 23811 33917 23819 33951
rect 23769 33893 23819 33917
rect 1593 33461 1643 33485
rect 1593 33427 1601 33461
rect 1635 33427 1643 33461
rect 1593 33403 1643 33427
rect 24173 33461 24223 33485
rect 24173 33427 24181 33461
rect 24215 33427 24223 33461
rect 24173 33403 24223 33427
rect 1593 33125 1643 33149
rect 1593 33091 1601 33125
rect 1635 33091 1643 33125
rect 1593 33067 1643 33091
rect 24173 33125 24223 33149
rect 24173 33091 24181 33125
rect 24215 33091 24223 33125
rect 24173 33067 24223 33091
rect 1593 32789 1643 32813
rect 1593 32755 1601 32789
rect 1635 32755 1643 32789
rect 1593 32731 1643 32755
rect 24173 32789 24223 32813
rect 24173 32755 24181 32789
rect 24215 32755 24223 32789
rect 24173 32731 24223 32755
rect 1593 32453 1643 32477
rect 1593 32419 1601 32453
rect 1635 32419 1643 32453
rect 1593 32395 1643 32419
rect 24173 32453 24223 32477
rect 24173 32419 24181 32453
rect 24215 32419 24223 32453
rect 24173 32395 24223 32419
rect 1593 32117 1643 32141
rect 1593 32083 1601 32117
rect 1635 32083 1643 32117
rect 1593 32059 1643 32083
rect 24173 32117 24223 32141
rect 24173 32083 24181 32117
rect 24215 32083 24223 32117
rect 24173 32059 24223 32083
rect 1593 31781 1643 31805
rect 1593 31747 1601 31781
rect 1635 31747 1643 31781
rect 1593 31723 1643 31747
rect 24173 31781 24223 31805
rect 24173 31747 24181 31781
rect 24215 31747 24223 31781
rect 24173 31723 24223 31747
rect 1593 31445 1643 31469
rect 1593 31411 1601 31445
rect 1635 31411 1643 31445
rect 1593 31387 1643 31411
rect 24173 31445 24223 31469
rect 24173 31411 24181 31445
rect 24215 31411 24223 31445
rect 24173 31387 24223 31411
rect 1593 31109 1643 31133
rect 1593 31075 1601 31109
rect 1635 31075 1643 31109
rect 1593 31051 1643 31075
rect 24173 31109 24223 31133
rect 24173 31075 24181 31109
rect 24215 31075 24223 31109
rect 24173 31051 24223 31075
rect 1593 30773 1643 30797
rect 1593 30739 1601 30773
rect 1635 30739 1643 30773
rect 1593 30715 1643 30739
rect 24173 30773 24223 30797
rect 24173 30739 24181 30773
rect 24215 30739 24223 30773
rect 24173 30715 24223 30739
rect 1593 30437 1643 30461
rect 1593 30403 1601 30437
rect 1635 30403 1643 30437
rect 1593 30379 1643 30403
rect 24173 30437 24223 30461
rect 24173 30403 24181 30437
rect 24215 30403 24223 30437
rect 24173 30379 24223 30403
rect 1593 30101 1643 30125
rect 1593 30067 1601 30101
rect 1635 30067 1643 30101
rect 1593 30043 1643 30067
rect 24173 30101 24223 30125
rect 24173 30067 24181 30101
rect 24215 30067 24223 30101
rect 24173 30043 24223 30067
rect 1593 29765 1643 29789
rect 1593 29731 1601 29765
rect 1635 29731 1643 29765
rect 1593 29707 1643 29731
rect 24173 29765 24223 29789
rect 24173 29731 24181 29765
rect 24215 29731 24223 29765
rect 24173 29707 24223 29731
rect 1593 29429 1643 29453
rect 1593 29395 1601 29429
rect 1635 29395 1643 29429
rect 1593 29371 1643 29395
rect 24173 29429 24223 29453
rect 24173 29395 24181 29429
rect 24215 29395 24223 29429
rect 24173 29371 24223 29395
rect 1593 29093 1643 29117
rect 1593 29059 1601 29093
rect 1635 29059 1643 29093
rect 1593 29035 1643 29059
rect 24173 29093 24223 29117
rect 24173 29059 24181 29093
rect 24215 29059 24223 29093
rect 24173 29035 24223 29059
rect 1593 28757 1643 28781
rect 1593 28723 1601 28757
rect 1635 28723 1643 28757
rect 1593 28699 1643 28723
rect 24173 28757 24223 28781
rect 24173 28723 24181 28757
rect 24215 28723 24223 28757
rect 24173 28699 24223 28723
rect 1593 28421 1643 28445
rect 1593 28387 1601 28421
rect 1635 28387 1643 28421
rect 1593 28363 1643 28387
rect 24173 28421 24223 28445
rect 24173 28387 24181 28421
rect 24215 28387 24223 28421
rect 24173 28363 24223 28387
rect 1593 28085 1643 28109
rect 1593 28051 1601 28085
rect 1635 28051 1643 28085
rect 1593 28027 1643 28051
rect 24173 28085 24223 28109
rect 24173 28051 24181 28085
rect 24215 28051 24223 28085
rect 24173 28027 24223 28051
rect 1593 27749 1643 27773
rect 1593 27715 1601 27749
rect 1635 27715 1643 27749
rect 1593 27691 1643 27715
rect 24173 27749 24223 27773
rect 24173 27715 24181 27749
rect 24215 27715 24223 27749
rect 24173 27691 24223 27715
rect 1593 27413 1643 27437
rect 1593 27379 1601 27413
rect 1635 27379 1643 27413
rect 1593 27355 1643 27379
rect 24173 27413 24223 27437
rect 24173 27379 24181 27413
rect 24215 27379 24223 27413
rect 24173 27355 24223 27379
rect 1593 27077 1643 27101
rect 1593 27043 1601 27077
rect 1635 27043 1643 27077
rect 1593 27019 1643 27043
rect 24173 27077 24223 27101
rect 24173 27043 24181 27077
rect 24215 27043 24223 27077
rect 24173 27019 24223 27043
rect 1593 26741 1643 26765
rect 1593 26707 1601 26741
rect 1635 26707 1643 26741
rect 1593 26683 1643 26707
rect 24173 26741 24223 26765
rect 24173 26707 24181 26741
rect 24215 26707 24223 26741
rect 24173 26683 24223 26707
rect 1593 26405 1643 26429
rect 1593 26371 1601 26405
rect 1635 26371 1643 26405
rect 1593 26347 1643 26371
rect 24173 26405 24223 26429
rect 24173 26371 24181 26405
rect 24215 26371 24223 26405
rect 24173 26347 24223 26371
rect 1593 26069 1643 26093
rect 1593 26035 1601 26069
rect 1635 26035 1643 26069
rect 1593 26011 1643 26035
rect 24173 26069 24223 26093
rect 24173 26035 24181 26069
rect 24215 26035 24223 26069
rect 24173 26011 24223 26035
rect 1593 25733 1643 25757
rect 1593 25699 1601 25733
rect 1635 25699 1643 25733
rect 1593 25675 1643 25699
rect 24173 25733 24223 25757
rect 24173 25699 24181 25733
rect 24215 25699 24223 25733
rect 24173 25675 24223 25699
rect 1593 25397 1643 25421
rect 1593 25363 1601 25397
rect 1635 25363 1643 25397
rect 1593 25339 1643 25363
rect 24173 25397 24223 25421
rect 24173 25363 24181 25397
rect 24215 25363 24223 25397
rect 24173 25339 24223 25363
rect 1593 25061 1643 25085
rect 1593 25027 1601 25061
rect 1635 25027 1643 25061
rect 1593 25003 1643 25027
rect 24173 25061 24223 25085
rect 24173 25027 24181 25061
rect 24215 25027 24223 25061
rect 24173 25003 24223 25027
rect 1593 24725 1643 24749
rect 1593 24691 1601 24725
rect 1635 24691 1643 24725
rect 1593 24667 1643 24691
rect 24173 24725 24223 24749
rect 24173 24691 24181 24725
rect 24215 24691 24223 24725
rect 24173 24667 24223 24691
rect 1593 24389 1643 24413
rect 1593 24355 1601 24389
rect 1635 24355 1643 24389
rect 1593 24331 1643 24355
rect 24173 24389 24223 24413
rect 24173 24355 24181 24389
rect 24215 24355 24223 24389
rect 24173 24331 24223 24355
rect 1593 24053 1643 24077
rect 1593 24019 1601 24053
rect 1635 24019 1643 24053
rect 1593 23995 1643 24019
rect 24173 24053 24223 24077
rect 24173 24019 24181 24053
rect 24215 24019 24223 24053
rect 24173 23995 24223 24019
rect 1593 23717 1643 23741
rect 1593 23683 1601 23717
rect 1635 23683 1643 23717
rect 1593 23659 1643 23683
rect 24173 23717 24223 23741
rect 24173 23683 24181 23717
rect 24215 23683 24223 23717
rect 24173 23659 24223 23683
rect 1593 23381 1643 23405
rect 1593 23347 1601 23381
rect 1635 23347 1643 23381
rect 1593 23323 1643 23347
rect 24173 23381 24223 23405
rect 24173 23347 24181 23381
rect 24215 23347 24223 23381
rect 24173 23323 24223 23347
rect 1593 23045 1643 23069
rect 1593 23011 1601 23045
rect 1635 23011 1643 23045
rect 1593 22987 1643 23011
rect 24173 23045 24223 23069
rect 24173 23011 24181 23045
rect 24215 23011 24223 23045
rect 24173 22987 24223 23011
rect 1593 22709 1643 22733
rect 1593 22675 1601 22709
rect 1635 22675 1643 22709
rect 1593 22651 1643 22675
rect 24173 22709 24223 22733
rect 24173 22675 24181 22709
rect 24215 22675 24223 22709
rect 24173 22651 24223 22675
rect 1593 22373 1643 22397
rect 1593 22339 1601 22373
rect 1635 22339 1643 22373
rect 1593 22315 1643 22339
rect 24173 22373 24223 22397
rect 24173 22339 24181 22373
rect 24215 22339 24223 22373
rect 24173 22315 24223 22339
rect 1593 22037 1643 22061
rect 1593 22003 1601 22037
rect 1635 22003 1643 22037
rect 1593 21979 1643 22003
rect 24173 22037 24223 22061
rect 24173 22003 24181 22037
rect 24215 22003 24223 22037
rect 24173 21979 24223 22003
rect 1593 21701 1643 21725
rect 1593 21667 1601 21701
rect 1635 21667 1643 21701
rect 1593 21643 1643 21667
rect 24173 21701 24223 21725
rect 24173 21667 24181 21701
rect 24215 21667 24223 21701
rect 24173 21643 24223 21667
rect 1593 21365 1643 21389
rect 1593 21331 1601 21365
rect 1635 21331 1643 21365
rect 1593 21307 1643 21331
rect 24173 21365 24223 21389
rect 24173 21331 24181 21365
rect 24215 21331 24223 21365
rect 24173 21307 24223 21331
rect 1593 21029 1643 21053
rect 1593 20995 1601 21029
rect 1635 20995 1643 21029
rect 1593 20971 1643 20995
rect 24173 21029 24223 21053
rect 24173 20995 24181 21029
rect 24215 20995 24223 21029
rect 24173 20971 24223 20995
rect 1593 20693 1643 20717
rect 1593 20659 1601 20693
rect 1635 20659 1643 20693
rect 1593 20635 1643 20659
rect 24173 20693 24223 20717
rect 24173 20659 24181 20693
rect 24215 20659 24223 20693
rect 24173 20635 24223 20659
rect 1593 20357 1643 20381
rect 1593 20323 1601 20357
rect 1635 20323 1643 20357
rect 1593 20299 1643 20323
rect 24173 20357 24223 20381
rect 24173 20323 24181 20357
rect 24215 20323 24223 20357
rect 24173 20299 24223 20323
rect 1593 20021 1643 20045
rect 1593 19987 1601 20021
rect 1635 19987 1643 20021
rect 1593 19963 1643 19987
rect 24173 20021 24223 20045
rect 24173 19987 24181 20021
rect 24215 19987 24223 20021
rect 24173 19963 24223 19987
rect 1593 19685 1643 19709
rect 1593 19651 1601 19685
rect 1635 19651 1643 19685
rect 1593 19627 1643 19651
rect 24173 19685 24223 19709
rect 24173 19651 24181 19685
rect 24215 19651 24223 19685
rect 24173 19627 24223 19651
rect 1593 19349 1643 19373
rect 1593 19315 1601 19349
rect 1635 19315 1643 19349
rect 1593 19291 1643 19315
rect 24173 19349 24223 19373
rect 24173 19315 24181 19349
rect 24215 19315 24223 19349
rect 24173 19291 24223 19315
rect 1593 19013 1643 19037
rect 1593 18979 1601 19013
rect 1635 18979 1643 19013
rect 1593 18955 1643 18979
rect 24173 19013 24223 19037
rect 24173 18979 24181 19013
rect 24215 18979 24223 19013
rect 24173 18955 24223 18979
rect 1593 18677 1643 18701
rect 1593 18643 1601 18677
rect 1635 18643 1643 18677
rect 1593 18619 1643 18643
rect 24173 18677 24223 18701
rect 24173 18643 24181 18677
rect 24215 18643 24223 18677
rect 24173 18619 24223 18643
rect 1593 18341 1643 18365
rect 1593 18307 1601 18341
rect 1635 18307 1643 18341
rect 1593 18283 1643 18307
rect 24173 18341 24223 18365
rect 24173 18307 24181 18341
rect 24215 18307 24223 18341
rect 24173 18283 24223 18307
rect 1593 18005 1643 18029
rect 1593 17971 1601 18005
rect 1635 17971 1643 18005
rect 1593 17947 1643 17971
rect 24173 18005 24223 18029
rect 24173 17971 24181 18005
rect 24215 17971 24223 18005
rect 24173 17947 24223 17971
rect 1593 17669 1643 17693
rect 1593 17635 1601 17669
rect 1635 17635 1643 17669
rect 1593 17611 1643 17635
rect 24173 17669 24223 17693
rect 24173 17635 24181 17669
rect 24215 17635 24223 17669
rect 24173 17611 24223 17635
rect 1593 17333 1643 17357
rect 1593 17299 1601 17333
rect 1635 17299 1643 17333
rect 1593 17275 1643 17299
rect 24173 17333 24223 17357
rect 24173 17299 24181 17333
rect 24215 17299 24223 17333
rect 24173 17275 24223 17299
rect 1593 16997 1643 17021
rect 1593 16963 1601 16997
rect 1635 16963 1643 16997
rect 1593 16939 1643 16963
rect 24173 16997 24223 17021
rect 24173 16963 24181 16997
rect 24215 16963 24223 16997
rect 24173 16939 24223 16963
rect 1593 16661 1643 16685
rect 1593 16627 1601 16661
rect 1635 16627 1643 16661
rect 1593 16603 1643 16627
rect 24173 16661 24223 16685
rect 24173 16627 24181 16661
rect 24215 16627 24223 16661
rect 24173 16603 24223 16627
rect 1593 16325 1643 16349
rect 1593 16291 1601 16325
rect 1635 16291 1643 16325
rect 1593 16267 1643 16291
rect 24173 16325 24223 16349
rect 24173 16291 24181 16325
rect 24215 16291 24223 16325
rect 24173 16267 24223 16291
rect 1593 15989 1643 16013
rect 1593 15955 1601 15989
rect 1635 15955 1643 15989
rect 1593 15931 1643 15955
rect 24173 15989 24223 16013
rect 24173 15955 24181 15989
rect 24215 15955 24223 15989
rect 24173 15931 24223 15955
rect 1593 15653 1643 15677
rect 1593 15619 1601 15653
rect 1635 15619 1643 15653
rect 1593 15595 1643 15619
rect 24173 15653 24223 15677
rect 24173 15619 24181 15653
rect 24215 15619 24223 15653
rect 24173 15595 24223 15619
rect 1593 15317 1643 15341
rect 1593 15283 1601 15317
rect 1635 15283 1643 15317
rect 1593 15259 1643 15283
rect 24173 15317 24223 15341
rect 24173 15283 24181 15317
rect 24215 15283 24223 15317
rect 24173 15259 24223 15283
rect 1593 14981 1643 15005
rect 1593 14947 1601 14981
rect 1635 14947 1643 14981
rect 1593 14923 1643 14947
rect 24173 14981 24223 15005
rect 24173 14947 24181 14981
rect 24215 14947 24223 14981
rect 24173 14923 24223 14947
rect 1593 14645 1643 14669
rect 1593 14611 1601 14645
rect 1635 14611 1643 14645
rect 1593 14587 1643 14611
rect 24173 14645 24223 14669
rect 24173 14611 24181 14645
rect 24215 14611 24223 14645
rect 24173 14587 24223 14611
rect 1593 14309 1643 14333
rect 1593 14275 1601 14309
rect 1635 14275 1643 14309
rect 1593 14251 1643 14275
rect 24173 14309 24223 14333
rect 24173 14275 24181 14309
rect 24215 14275 24223 14309
rect 24173 14251 24223 14275
rect 1593 13973 1643 13997
rect 1593 13939 1601 13973
rect 1635 13939 1643 13973
rect 1593 13915 1643 13939
rect 24173 13973 24223 13997
rect 24173 13939 24181 13973
rect 24215 13939 24223 13973
rect 24173 13915 24223 13939
rect 1593 13637 1643 13661
rect 1593 13603 1601 13637
rect 1635 13603 1643 13637
rect 1593 13579 1643 13603
rect 24173 13637 24223 13661
rect 24173 13603 24181 13637
rect 24215 13603 24223 13637
rect 24173 13579 24223 13603
rect 1593 13301 1643 13325
rect 1593 13267 1601 13301
rect 1635 13267 1643 13301
rect 1593 13243 1643 13267
rect 24173 13301 24223 13325
rect 24173 13267 24181 13301
rect 24215 13267 24223 13301
rect 24173 13243 24223 13267
rect 1593 12965 1643 12989
rect 1593 12931 1601 12965
rect 1635 12931 1643 12965
rect 1593 12907 1643 12931
rect 24173 12965 24223 12989
rect 24173 12931 24181 12965
rect 24215 12931 24223 12965
rect 24173 12907 24223 12931
rect 1593 12629 1643 12653
rect 1593 12595 1601 12629
rect 1635 12595 1643 12629
rect 1593 12571 1643 12595
rect 24173 12629 24223 12653
rect 24173 12595 24181 12629
rect 24215 12595 24223 12629
rect 24173 12571 24223 12595
rect 1593 12293 1643 12317
rect 1593 12259 1601 12293
rect 1635 12259 1643 12293
rect 1593 12235 1643 12259
rect 24173 12293 24223 12317
rect 24173 12259 24181 12293
rect 24215 12259 24223 12293
rect 24173 12235 24223 12259
rect 1593 11957 1643 11981
rect 1593 11923 1601 11957
rect 1635 11923 1643 11957
rect 1593 11899 1643 11923
rect 24173 11957 24223 11981
rect 24173 11923 24181 11957
rect 24215 11923 24223 11957
rect 24173 11899 24223 11923
rect 1593 11621 1643 11645
rect 1593 11587 1601 11621
rect 1635 11587 1643 11621
rect 1593 11563 1643 11587
rect 24173 11621 24223 11645
rect 24173 11587 24181 11621
rect 24215 11587 24223 11621
rect 24173 11563 24223 11587
rect 1593 11285 1643 11309
rect 1593 11251 1601 11285
rect 1635 11251 1643 11285
rect 1593 11227 1643 11251
rect 24173 11285 24223 11309
rect 24173 11251 24181 11285
rect 24215 11251 24223 11285
rect 24173 11227 24223 11251
rect 1593 10949 1643 10973
rect 1593 10915 1601 10949
rect 1635 10915 1643 10949
rect 1593 10891 1643 10915
rect 24173 10949 24223 10973
rect 24173 10915 24181 10949
rect 24215 10915 24223 10949
rect 24173 10891 24223 10915
rect 1593 10613 1643 10637
rect 1593 10579 1601 10613
rect 1635 10579 1643 10613
rect 1593 10555 1643 10579
rect 24173 10613 24223 10637
rect 24173 10579 24181 10613
rect 24215 10579 24223 10613
rect 24173 10555 24223 10579
rect 1593 10277 1643 10301
rect 1593 10243 1601 10277
rect 1635 10243 1643 10277
rect 1593 10219 1643 10243
rect 24173 10277 24223 10301
rect 24173 10243 24181 10277
rect 24215 10243 24223 10277
rect 24173 10219 24223 10243
rect 1593 9941 1643 9965
rect 1593 9907 1601 9941
rect 1635 9907 1643 9941
rect 1593 9883 1643 9907
rect 24173 9941 24223 9965
rect 24173 9907 24181 9941
rect 24215 9907 24223 9941
rect 24173 9883 24223 9907
rect 1593 9605 1643 9629
rect 1593 9571 1601 9605
rect 1635 9571 1643 9605
rect 1593 9547 1643 9571
rect 24173 9605 24223 9629
rect 24173 9571 24181 9605
rect 24215 9571 24223 9605
rect 24173 9547 24223 9571
rect 1593 9269 1643 9293
rect 1593 9235 1601 9269
rect 1635 9235 1643 9269
rect 1593 9211 1643 9235
rect 24173 9269 24223 9293
rect 24173 9235 24181 9269
rect 24215 9235 24223 9269
rect 24173 9211 24223 9235
rect 1593 8933 1643 8957
rect 1593 8899 1601 8933
rect 1635 8899 1643 8933
rect 1593 8875 1643 8899
rect 24173 8933 24223 8957
rect 24173 8899 24181 8933
rect 24215 8899 24223 8933
rect 24173 8875 24223 8899
rect 1593 8597 1643 8621
rect 1593 8563 1601 8597
rect 1635 8563 1643 8597
rect 1593 8539 1643 8563
rect 24173 8597 24223 8621
rect 24173 8563 24181 8597
rect 24215 8563 24223 8597
rect 24173 8539 24223 8563
rect 1593 8261 1643 8285
rect 1593 8227 1601 8261
rect 1635 8227 1643 8261
rect 1593 8203 1643 8227
rect 24173 8261 24223 8285
rect 24173 8227 24181 8261
rect 24215 8227 24223 8261
rect 24173 8203 24223 8227
rect 1593 7925 1643 7949
rect 1593 7891 1601 7925
rect 1635 7891 1643 7925
rect 1593 7867 1643 7891
rect 24173 7925 24223 7949
rect 24173 7891 24181 7925
rect 24215 7891 24223 7925
rect 24173 7867 24223 7891
rect 1593 7589 1643 7613
rect 1593 7555 1601 7589
rect 1635 7555 1643 7589
rect 1593 7531 1643 7555
rect 24173 7589 24223 7613
rect 24173 7555 24181 7589
rect 24215 7555 24223 7589
rect 24173 7531 24223 7555
rect 1593 7253 1643 7277
rect 1593 7219 1601 7253
rect 1635 7219 1643 7253
rect 1593 7195 1643 7219
rect 24173 7253 24223 7277
rect 24173 7219 24181 7253
rect 24215 7219 24223 7253
rect 24173 7195 24223 7219
rect 1593 6917 1643 6941
rect 1593 6883 1601 6917
rect 1635 6883 1643 6917
rect 1593 6859 1643 6883
rect 24173 6917 24223 6941
rect 24173 6883 24181 6917
rect 24215 6883 24223 6917
rect 24173 6859 24223 6883
rect 1593 6581 1643 6605
rect 1593 6547 1601 6581
rect 1635 6547 1643 6581
rect 1593 6523 1643 6547
rect 24173 6581 24223 6605
rect 24173 6547 24181 6581
rect 24215 6547 24223 6581
rect 24173 6523 24223 6547
rect 1593 6245 1643 6269
rect 1593 6211 1601 6245
rect 1635 6211 1643 6245
rect 1593 6187 1643 6211
rect 24173 6245 24223 6269
rect 24173 6211 24181 6245
rect 24215 6211 24223 6245
rect 24173 6187 24223 6211
rect 1593 5909 1643 5933
rect 1593 5875 1601 5909
rect 1635 5875 1643 5909
rect 1593 5851 1643 5875
rect 24173 5909 24223 5933
rect 24173 5875 24181 5909
rect 24215 5875 24223 5909
rect 24173 5851 24223 5875
rect 1593 5573 1643 5597
rect 1593 5539 1601 5573
rect 1635 5539 1643 5573
rect 1593 5515 1643 5539
rect 24173 5573 24223 5597
rect 24173 5539 24181 5573
rect 24215 5539 24223 5573
rect 24173 5515 24223 5539
rect 1593 5237 1643 5261
rect 1593 5203 1601 5237
rect 1635 5203 1643 5237
rect 1593 5179 1643 5203
rect 24173 5237 24223 5261
rect 24173 5203 24181 5237
rect 24215 5203 24223 5237
rect 24173 5179 24223 5203
rect 1593 4901 1643 4925
rect 1593 4867 1601 4901
rect 1635 4867 1643 4901
rect 1593 4843 1643 4867
rect 24173 4901 24223 4925
rect 24173 4867 24181 4901
rect 24215 4867 24223 4901
rect 24173 4843 24223 4867
rect 1593 4565 1643 4589
rect 1593 4531 1601 4565
rect 1635 4531 1643 4565
rect 1593 4507 1643 4531
rect 24173 4565 24223 4589
rect 24173 4531 24181 4565
rect 24215 4531 24223 4565
rect 24173 4507 24223 4531
rect 1593 4229 1643 4253
rect 1593 4195 1601 4229
rect 1635 4195 1643 4229
rect 1593 4171 1643 4195
rect 24173 4229 24223 4253
rect 24173 4195 24181 4229
rect 24215 4195 24223 4229
rect 24173 4171 24223 4195
rect 1593 3893 1643 3917
rect 1593 3859 1601 3893
rect 1635 3859 1643 3893
rect 1593 3835 1643 3859
rect 24173 3893 24223 3917
rect 24173 3859 24181 3893
rect 24215 3859 24223 3893
rect 24173 3835 24223 3859
rect 1593 3557 1643 3581
rect 1593 3523 1601 3557
rect 1635 3523 1643 3557
rect 1593 3499 1643 3523
rect 24173 3557 24223 3581
rect 24173 3523 24181 3557
rect 24215 3523 24223 3557
rect 24173 3499 24223 3523
rect 1593 3221 1643 3245
rect 1593 3187 1601 3221
rect 1635 3187 1643 3221
rect 1593 3163 1643 3187
rect 24173 3221 24223 3245
rect 24173 3187 24181 3221
rect 24215 3187 24223 3221
rect 24173 3163 24223 3187
rect 1593 2885 1643 2909
rect 1593 2851 1601 2885
rect 1635 2851 1643 2885
rect 1593 2827 1643 2851
rect 24173 2885 24223 2909
rect 24173 2851 24181 2885
rect 24215 2851 24223 2885
rect 24173 2827 24223 2851
rect 1593 2549 1643 2573
rect 1593 2515 1601 2549
rect 1635 2515 1643 2549
rect 1593 2491 1643 2515
rect 24173 2549 24223 2573
rect 24173 2515 24181 2549
rect 24215 2515 24223 2549
rect 24173 2491 24223 2515
rect 1593 2213 1643 2237
rect 1593 2179 1601 2213
rect 1635 2179 1643 2213
rect 1593 2155 1643 2179
rect 24173 2213 24223 2237
rect 24173 2179 24181 2213
rect 24215 2179 24223 2213
rect 24173 2155 24223 2179
rect 1593 1877 1643 1901
rect 1593 1843 1601 1877
rect 1635 1843 1643 1877
rect 1593 1819 1643 1843
rect 24173 1877 24223 1901
rect 24173 1843 24181 1877
rect 24215 1843 24223 1877
rect 24173 1819 24223 1843
rect 1929 1541 1979 1565
rect 1929 1507 1937 1541
rect 1971 1507 1979 1541
rect 1929 1483 1979 1507
rect 2265 1541 2315 1565
rect 2265 1507 2273 1541
rect 2307 1507 2315 1541
rect 2265 1483 2315 1507
rect 2601 1541 2651 1565
rect 2601 1507 2609 1541
rect 2643 1507 2651 1541
rect 2601 1483 2651 1507
rect 2937 1541 2987 1565
rect 2937 1507 2945 1541
rect 2979 1507 2987 1541
rect 2937 1483 2987 1507
rect 3273 1541 3323 1565
rect 3273 1507 3281 1541
rect 3315 1507 3323 1541
rect 3273 1483 3323 1507
rect 3609 1541 3659 1565
rect 3609 1507 3617 1541
rect 3651 1507 3659 1541
rect 3609 1483 3659 1507
rect 3945 1541 3995 1565
rect 3945 1507 3953 1541
rect 3987 1507 3995 1541
rect 3945 1483 3995 1507
rect 4281 1541 4331 1565
rect 4281 1507 4289 1541
rect 4323 1507 4331 1541
rect 4281 1483 4331 1507
rect 4617 1541 4667 1565
rect 4617 1507 4625 1541
rect 4659 1507 4667 1541
rect 4617 1483 4667 1507
rect 4953 1541 5003 1565
rect 4953 1507 4961 1541
rect 4995 1507 5003 1541
rect 4953 1483 5003 1507
rect 5289 1541 5339 1565
rect 5289 1507 5297 1541
rect 5331 1507 5339 1541
rect 5289 1483 5339 1507
rect 5625 1541 5675 1565
rect 5625 1507 5633 1541
rect 5667 1507 5675 1541
rect 5625 1483 5675 1507
rect 5961 1541 6011 1565
rect 5961 1507 5969 1541
rect 6003 1507 6011 1541
rect 5961 1483 6011 1507
rect 6297 1541 6347 1565
rect 6297 1507 6305 1541
rect 6339 1507 6347 1541
rect 6297 1483 6347 1507
rect 6633 1541 6683 1565
rect 6633 1507 6641 1541
rect 6675 1507 6683 1541
rect 6633 1483 6683 1507
rect 6969 1541 7019 1565
rect 6969 1507 6977 1541
rect 7011 1507 7019 1541
rect 6969 1483 7019 1507
rect 7305 1541 7355 1565
rect 7305 1507 7313 1541
rect 7347 1507 7355 1541
rect 7305 1483 7355 1507
rect 7641 1541 7691 1565
rect 7641 1507 7649 1541
rect 7683 1507 7691 1541
rect 7641 1483 7691 1507
rect 7977 1541 8027 1565
rect 7977 1507 7985 1541
rect 8019 1507 8027 1541
rect 7977 1483 8027 1507
rect 8313 1541 8363 1565
rect 8313 1507 8321 1541
rect 8355 1507 8363 1541
rect 8313 1483 8363 1507
rect 8649 1541 8699 1565
rect 8649 1507 8657 1541
rect 8691 1507 8699 1541
rect 8649 1483 8699 1507
rect 8985 1541 9035 1565
rect 8985 1507 8993 1541
rect 9027 1507 9035 1541
rect 8985 1483 9035 1507
rect 9321 1541 9371 1565
rect 9321 1507 9329 1541
rect 9363 1507 9371 1541
rect 9321 1483 9371 1507
rect 9657 1541 9707 1565
rect 9657 1507 9665 1541
rect 9699 1507 9707 1541
rect 9657 1483 9707 1507
rect 9993 1541 10043 1565
rect 9993 1507 10001 1541
rect 10035 1507 10043 1541
rect 9993 1483 10043 1507
rect 10329 1541 10379 1565
rect 10329 1507 10337 1541
rect 10371 1507 10379 1541
rect 10329 1483 10379 1507
rect 10665 1541 10715 1565
rect 10665 1507 10673 1541
rect 10707 1507 10715 1541
rect 10665 1483 10715 1507
rect 11001 1541 11051 1565
rect 11001 1507 11009 1541
rect 11043 1507 11051 1541
rect 11001 1483 11051 1507
rect 11337 1541 11387 1565
rect 11337 1507 11345 1541
rect 11379 1507 11387 1541
rect 11337 1483 11387 1507
rect 11673 1541 11723 1565
rect 11673 1507 11681 1541
rect 11715 1507 11723 1541
rect 11673 1483 11723 1507
rect 12009 1541 12059 1565
rect 12009 1507 12017 1541
rect 12051 1507 12059 1541
rect 12009 1483 12059 1507
rect 12345 1541 12395 1565
rect 12345 1507 12353 1541
rect 12387 1507 12395 1541
rect 12345 1483 12395 1507
rect 12681 1541 12731 1565
rect 12681 1507 12689 1541
rect 12723 1507 12731 1541
rect 12681 1483 12731 1507
rect 13017 1541 13067 1565
rect 13017 1507 13025 1541
rect 13059 1507 13067 1541
rect 13017 1483 13067 1507
rect 13353 1541 13403 1565
rect 13353 1507 13361 1541
rect 13395 1507 13403 1541
rect 13353 1483 13403 1507
rect 13689 1541 13739 1565
rect 13689 1507 13697 1541
rect 13731 1507 13739 1541
rect 13689 1483 13739 1507
rect 14025 1541 14075 1565
rect 14025 1507 14033 1541
rect 14067 1507 14075 1541
rect 14025 1483 14075 1507
rect 14361 1541 14411 1565
rect 14361 1507 14369 1541
rect 14403 1507 14411 1541
rect 14361 1483 14411 1507
rect 14697 1541 14747 1565
rect 14697 1507 14705 1541
rect 14739 1507 14747 1541
rect 14697 1483 14747 1507
rect 15033 1541 15083 1565
rect 15033 1507 15041 1541
rect 15075 1507 15083 1541
rect 15033 1483 15083 1507
rect 15369 1541 15419 1565
rect 15369 1507 15377 1541
rect 15411 1507 15419 1541
rect 15369 1483 15419 1507
rect 15705 1541 15755 1565
rect 15705 1507 15713 1541
rect 15747 1507 15755 1541
rect 15705 1483 15755 1507
rect 16041 1541 16091 1565
rect 16041 1507 16049 1541
rect 16083 1507 16091 1541
rect 16041 1483 16091 1507
rect 16377 1541 16427 1565
rect 16377 1507 16385 1541
rect 16419 1507 16427 1541
rect 16377 1483 16427 1507
rect 16713 1541 16763 1565
rect 16713 1507 16721 1541
rect 16755 1507 16763 1541
rect 16713 1483 16763 1507
rect 17049 1541 17099 1565
rect 17049 1507 17057 1541
rect 17091 1507 17099 1541
rect 17049 1483 17099 1507
rect 17385 1541 17435 1565
rect 17385 1507 17393 1541
rect 17427 1507 17435 1541
rect 17385 1483 17435 1507
rect 17721 1541 17771 1565
rect 17721 1507 17729 1541
rect 17763 1507 17771 1541
rect 17721 1483 17771 1507
rect 18057 1541 18107 1565
rect 18057 1507 18065 1541
rect 18099 1507 18107 1541
rect 18057 1483 18107 1507
rect 18393 1541 18443 1565
rect 18393 1507 18401 1541
rect 18435 1507 18443 1541
rect 18393 1483 18443 1507
rect 18729 1541 18779 1565
rect 18729 1507 18737 1541
rect 18771 1507 18779 1541
rect 18729 1483 18779 1507
rect 19065 1541 19115 1565
rect 19065 1507 19073 1541
rect 19107 1507 19115 1541
rect 19065 1483 19115 1507
rect 19401 1541 19451 1565
rect 19401 1507 19409 1541
rect 19443 1507 19451 1541
rect 19401 1483 19451 1507
rect 19737 1541 19787 1565
rect 19737 1507 19745 1541
rect 19779 1507 19787 1541
rect 19737 1483 19787 1507
rect 20073 1541 20123 1565
rect 20073 1507 20081 1541
rect 20115 1507 20123 1541
rect 20073 1483 20123 1507
rect 20409 1541 20459 1565
rect 20409 1507 20417 1541
rect 20451 1507 20459 1541
rect 20409 1483 20459 1507
rect 20745 1541 20795 1565
rect 20745 1507 20753 1541
rect 20787 1507 20795 1541
rect 20745 1483 20795 1507
rect 21081 1541 21131 1565
rect 21081 1507 21089 1541
rect 21123 1507 21131 1541
rect 21081 1483 21131 1507
rect 21417 1541 21467 1565
rect 21417 1507 21425 1541
rect 21459 1507 21467 1541
rect 21417 1483 21467 1507
rect 21753 1541 21803 1565
rect 21753 1507 21761 1541
rect 21795 1507 21803 1541
rect 21753 1483 21803 1507
rect 22089 1541 22139 1565
rect 22089 1507 22097 1541
rect 22131 1507 22139 1541
rect 22089 1483 22139 1507
rect 22425 1541 22475 1565
rect 22425 1507 22433 1541
rect 22467 1507 22475 1541
rect 22425 1483 22475 1507
rect 22761 1541 22811 1565
rect 22761 1507 22769 1541
rect 22803 1507 22811 1541
rect 22761 1483 22811 1507
rect 23097 1541 23147 1565
rect 23097 1507 23105 1541
rect 23139 1507 23147 1541
rect 23097 1483 23147 1507
rect 23433 1541 23483 1565
rect 23433 1507 23441 1541
rect 23475 1507 23483 1541
rect 23433 1483 23483 1507
rect 23769 1541 23819 1565
rect 23769 1507 23777 1541
rect 23811 1507 23819 1541
rect 23769 1483 23819 1507
<< nsubdiffcont >>
rect 1937 33917 1971 33951
rect 2273 33917 2307 33951
rect 2609 33917 2643 33951
rect 2945 33917 2979 33951
rect 3281 33917 3315 33951
rect 3617 33917 3651 33951
rect 3953 33917 3987 33951
rect 4289 33917 4323 33951
rect 4625 33917 4659 33951
rect 4961 33917 4995 33951
rect 5297 33917 5331 33951
rect 5633 33917 5667 33951
rect 5969 33917 6003 33951
rect 6305 33917 6339 33951
rect 6641 33917 6675 33951
rect 6977 33917 7011 33951
rect 7313 33917 7347 33951
rect 7649 33917 7683 33951
rect 7985 33917 8019 33951
rect 8321 33917 8355 33951
rect 8657 33917 8691 33951
rect 8993 33917 9027 33951
rect 9329 33917 9363 33951
rect 9665 33917 9699 33951
rect 10001 33917 10035 33951
rect 10337 33917 10371 33951
rect 10673 33917 10707 33951
rect 11009 33917 11043 33951
rect 11345 33917 11379 33951
rect 11681 33917 11715 33951
rect 12017 33917 12051 33951
rect 12353 33917 12387 33951
rect 12689 33917 12723 33951
rect 13025 33917 13059 33951
rect 13361 33917 13395 33951
rect 13697 33917 13731 33951
rect 14033 33917 14067 33951
rect 14369 33917 14403 33951
rect 14705 33917 14739 33951
rect 15041 33917 15075 33951
rect 15377 33917 15411 33951
rect 15713 33917 15747 33951
rect 16049 33917 16083 33951
rect 16385 33917 16419 33951
rect 16721 33917 16755 33951
rect 17057 33917 17091 33951
rect 17393 33917 17427 33951
rect 17729 33917 17763 33951
rect 18065 33917 18099 33951
rect 18401 33917 18435 33951
rect 18737 33917 18771 33951
rect 19073 33917 19107 33951
rect 19409 33917 19443 33951
rect 19745 33917 19779 33951
rect 20081 33917 20115 33951
rect 20417 33917 20451 33951
rect 20753 33917 20787 33951
rect 21089 33917 21123 33951
rect 21425 33917 21459 33951
rect 21761 33917 21795 33951
rect 22097 33917 22131 33951
rect 22433 33917 22467 33951
rect 22769 33917 22803 33951
rect 23105 33917 23139 33951
rect 23441 33917 23475 33951
rect 23777 33917 23811 33951
rect 1601 33427 1635 33461
rect 24181 33427 24215 33461
rect 1601 33091 1635 33125
rect 24181 33091 24215 33125
rect 1601 32755 1635 32789
rect 24181 32755 24215 32789
rect 1601 32419 1635 32453
rect 24181 32419 24215 32453
rect 1601 32083 1635 32117
rect 24181 32083 24215 32117
rect 1601 31747 1635 31781
rect 24181 31747 24215 31781
rect 1601 31411 1635 31445
rect 24181 31411 24215 31445
rect 1601 31075 1635 31109
rect 24181 31075 24215 31109
rect 1601 30739 1635 30773
rect 24181 30739 24215 30773
rect 1601 30403 1635 30437
rect 24181 30403 24215 30437
rect 1601 30067 1635 30101
rect 24181 30067 24215 30101
rect 1601 29731 1635 29765
rect 24181 29731 24215 29765
rect 1601 29395 1635 29429
rect 24181 29395 24215 29429
rect 1601 29059 1635 29093
rect 24181 29059 24215 29093
rect 1601 28723 1635 28757
rect 24181 28723 24215 28757
rect 1601 28387 1635 28421
rect 24181 28387 24215 28421
rect 1601 28051 1635 28085
rect 24181 28051 24215 28085
rect 1601 27715 1635 27749
rect 24181 27715 24215 27749
rect 1601 27379 1635 27413
rect 24181 27379 24215 27413
rect 1601 27043 1635 27077
rect 24181 27043 24215 27077
rect 1601 26707 1635 26741
rect 24181 26707 24215 26741
rect 1601 26371 1635 26405
rect 24181 26371 24215 26405
rect 1601 26035 1635 26069
rect 24181 26035 24215 26069
rect 1601 25699 1635 25733
rect 24181 25699 24215 25733
rect 1601 25363 1635 25397
rect 24181 25363 24215 25397
rect 1601 25027 1635 25061
rect 24181 25027 24215 25061
rect 1601 24691 1635 24725
rect 24181 24691 24215 24725
rect 1601 24355 1635 24389
rect 24181 24355 24215 24389
rect 1601 24019 1635 24053
rect 24181 24019 24215 24053
rect 1601 23683 1635 23717
rect 24181 23683 24215 23717
rect 1601 23347 1635 23381
rect 24181 23347 24215 23381
rect 1601 23011 1635 23045
rect 24181 23011 24215 23045
rect 1601 22675 1635 22709
rect 24181 22675 24215 22709
rect 1601 22339 1635 22373
rect 24181 22339 24215 22373
rect 1601 22003 1635 22037
rect 24181 22003 24215 22037
rect 1601 21667 1635 21701
rect 24181 21667 24215 21701
rect 1601 21331 1635 21365
rect 24181 21331 24215 21365
rect 1601 20995 1635 21029
rect 24181 20995 24215 21029
rect 1601 20659 1635 20693
rect 24181 20659 24215 20693
rect 1601 20323 1635 20357
rect 24181 20323 24215 20357
rect 1601 19987 1635 20021
rect 24181 19987 24215 20021
rect 1601 19651 1635 19685
rect 24181 19651 24215 19685
rect 1601 19315 1635 19349
rect 24181 19315 24215 19349
rect 1601 18979 1635 19013
rect 24181 18979 24215 19013
rect 1601 18643 1635 18677
rect 24181 18643 24215 18677
rect 1601 18307 1635 18341
rect 24181 18307 24215 18341
rect 1601 17971 1635 18005
rect 24181 17971 24215 18005
rect 1601 17635 1635 17669
rect 24181 17635 24215 17669
rect 1601 17299 1635 17333
rect 24181 17299 24215 17333
rect 1601 16963 1635 16997
rect 24181 16963 24215 16997
rect 1601 16627 1635 16661
rect 24181 16627 24215 16661
rect 1601 16291 1635 16325
rect 24181 16291 24215 16325
rect 1601 15955 1635 15989
rect 24181 15955 24215 15989
rect 1601 15619 1635 15653
rect 24181 15619 24215 15653
rect 1601 15283 1635 15317
rect 24181 15283 24215 15317
rect 1601 14947 1635 14981
rect 24181 14947 24215 14981
rect 1601 14611 1635 14645
rect 24181 14611 24215 14645
rect 1601 14275 1635 14309
rect 24181 14275 24215 14309
rect 1601 13939 1635 13973
rect 24181 13939 24215 13973
rect 1601 13603 1635 13637
rect 24181 13603 24215 13637
rect 1601 13267 1635 13301
rect 24181 13267 24215 13301
rect 1601 12931 1635 12965
rect 24181 12931 24215 12965
rect 1601 12595 1635 12629
rect 24181 12595 24215 12629
rect 1601 12259 1635 12293
rect 24181 12259 24215 12293
rect 1601 11923 1635 11957
rect 24181 11923 24215 11957
rect 1601 11587 1635 11621
rect 24181 11587 24215 11621
rect 1601 11251 1635 11285
rect 24181 11251 24215 11285
rect 1601 10915 1635 10949
rect 24181 10915 24215 10949
rect 1601 10579 1635 10613
rect 24181 10579 24215 10613
rect 1601 10243 1635 10277
rect 24181 10243 24215 10277
rect 1601 9907 1635 9941
rect 24181 9907 24215 9941
rect 1601 9571 1635 9605
rect 24181 9571 24215 9605
rect 1601 9235 1635 9269
rect 24181 9235 24215 9269
rect 1601 8899 1635 8933
rect 24181 8899 24215 8933
rect 1601 8563 1635 8597
rect 24181 8563 24215 8597
rect 1601 8227 1635 8261
rect 24181 8227 24215 8261
rect 1601 7891 1635 7925
rect 24181 7891 24215 7925
rect 1601 7555 1635 7589
rect 24181 7555 24215 7589
rect 1601 7219 1635 7253
rect 24181 7219 24215 7253
rect 1601 6883 1635 6917
rect 24181 6883 24215 6917
rect 1601 6547 1635 6581
rect 24181 6547 24215 6581
rect 1601 6211 1635 6245
rect 24181 6211 24215 6245
rect 1601 5875 1635 5909
rect 24181 5875 24215 5909
rect 1601 5539 1635 5573
rect 24181 5539 24215 5573
rect 1601 5203 1635 5237
rect 24181 5203 24215 5237
rect 1601 4867 1635 4901
rect 24181 4867 24215 4901
rect 1601 4531 1635 4565
rect 24181 4531 24215 4565
rect 1601 4195 1635 4229
rect 24181 4195 24215 4229
rect 1601 3859 1635 3893
rect 24181 3859 24215 3893
rect 1601 3523 1635 3557
rect 24181 3523 24215 3557
rect 1601 3187 1635 3221
rect 24181 3187 24215 3221
rect 1601 2851 1635 2885
rect 24181 2851 24215 2885
rect 1601 2515 1635 2549
rect 24181 2515 24215 2549
rect 1601 2179 1635 2213
rect 24181 2179 24215 2213
rect 1601 1843 1635 1877
rect 24181 1843 24215 1877
rect 1937 1507 1971 1541
rect 2273 1507 2307 1541
rect 2609 1507 2643 1541
rect 2945 1507 2979 1541
rect 3281 1507 3315 1541
rect 3617 1507 3651 1541
rect 3953 1507 3987 1541
rect 4289 1507 4323 1541
rect 4625 1507 4659 1541
rect 4961 1507 4995 1541
rect 5297 1507 5331 1541
rect 5633 1507 5667 1541
rect 5969 1507 6003 1541
rect 6305 1507 6339 1541
rect 6641 1507 6675 1541
rect 6977 1507 7011 1541
rect 7313 1507 7347 1541
rect 7649 1507 7683 1541
rect 7985 1507 8019 1541
rect 8321 1507 8355 1541
rect 8657 1507 8691 1541
rect 8993 1507 9027 1541
rect 9329 1507 9363 1541
rect 9665 1507 9699 1541
rect 10001 1507 10035 1541
rect 10337 1507 10371 1541
rect 10673 1507 10707 1541
rect 11009 1507 11043 1541
rect 11345 1507 11379 1541
rect 11681 1507 11715 1541
rect 12017 1507 12051 1541
rect 12353 1507 12387 1541
rect 12689 1507 12723 1541
rect 13025 1507 13059 1541
rect 13361 1507 13395 1541
rect 13697 1507 13731 1541
rect 14033 1507 14067 1541
rect 14369 1507 14403 1541
rect 14705 1507 14739 1541
rect 15041 1507 15075 1541
rect 15377 1507 15411 1541
rect 15713 1507 15747 1541
rect 16049 1507 16083 1541
rect 16385 1507 16419 1541
rect 16721 1507 16755 1541
rect 17057 1507 17091 1541
rect 17393 1507 17427 1541
rect 17729 1507 17763 1541
rect 18065 1507 18099 1541
rect 18401 1507 18435 1541
rect 18737 1507 18771 1541
rect 19073 1507 19107 1541
rect 19409 1507 19443 1541
rect 19745 1507 19779 1541
rect 20081 1507 20115 1541
rect 20417 1507 20451 1541
rect 20753 1507 20787 1541
rect 21089 1507 21123 1541
rect 21425 1507 21459 1541
rect 21761 1507 21795 1541
rect 22097 1507 22131 1541
rect 22433 1507 22467 1541
rect 22769 1507 22803 1541
rect 23105 1507 23139 1541
rect 23441 1507 23475 1541
rect 23777 1507 23811 1541
<< locali >>
rect 1937 33951 1971 33967
rect 1937 33901 1971 33917
rect 2273 33951 2307 33967
rect 2273 33901 2307 33917
rect 2609 33951 2643 33967
rect 2609 33901 2643 33917
rect 2945 33951 2979 33967
rect 2945 33901 2979 33917
rect 3281 33951 3315 33967
rect 3281 33901 3315 33917
rect 3617 33951 3651 33967
rect 3617 33901 3651 33917
rect 3953 33951 3987 33967
rect 3953 33901 3987 33917
rect 4289 33951 4323 33967
rect 4289 33901 4323 33917
rect 4625 33951 4659 33967
rect 4625 33901 4659 33917
rect 4961 33951 4995 33967
rect 4961 33901 4995 33917
rect 5297 33951 5331 33967
rect 5297 33901 5331 33917
rect 5633 33951 5667 33967
rect 5633 33901 5667 33917
rect 5969 33951 6003 33967
rect 5969 33901 6003 33917
rect 6305 33951 6339 33967
rect 6305 33901 6339 33917
rect 6641 33951 6675 33967
rect 6641 33901 6675 33917
rect 6977 33951 7011 33967
rect 6977 33901 7011 33917
rect 7313 33951 7347 33967
rect 7313 33901 7347 33917
rect 7649 33951 7683 33967
rect 7649 33901 7683 33917
rect 7985 33951 8019 33967
rect 7985 33901 8019 33917
rect 8321 33951 8355 33967
rect 8321 33901 8355 33917
rect 8657 33951 8691 33967
rect 8657 33901 8691 33917
rect 8993 33951 9027 33967
rect 8993 33901 9027 33917
rect 9329 33951 9363 33967
rect 9329 33901 9363 33917
rect 9665 33951 9699 33967
rect 9665 33901 9699 33917
rect 10001 33951 10035 33967
rect 10001 33901 10035 33917
rect 10337 33951 10371 33967
rect 10337 33901 10371 33917
rect 10673 33951 10707 33967
rect 10673 33901 10707 33917
rect 11009 33951 11043 33967
rect 11009 33901 11043 33917
rect 11345 33951 11379 33967
rect 11345 33901 11379 33917
rect 11681 33951 11715 33967
rect 11681 33901 11715 33917
rect 12017 33951 12051 33967
rect 12017 33901 12051 33917
rect 12353 33951 12387 33967
rect 12353 33901 12387 33917
rect 12689 33951 12723 33967
rect 12689 33901 12723 33917
rect 13025 33951 13059 33967
rect 13025 33901 13059 33917
rect 13361 33951 13395 33967
rect 13361 33901 13395 33917
rect 13697 33951 13731 33967
rect 13697 33901 13731 33917
rect 14033 33951 14067 33967
rect 14033 33901 14067 33917
rect 14369 33951 14403 33967
rect 14369 33901 14403 33917
rect 14705 33951 14739 33967
rect 14705 33901 14739 33917
rect 15041 33951 15075 33967
rect 15041 33901 15075 33917
rect 15377 33951 15411 33967
rect 15377 33901 15411 33917
rect 15713 33951 15747 33967
rect 15713 33901 15747 33917
rect 16049 33951 16083 33967
rect 16049 33901 16083 33917
rect 16385 33951 16419 33967
rect 16385 33901 16419 33917
rect 16721 33951 16755 33967
rect 16721 33901 16755 33917
rect 17057 33951 17091 33967
rect 17057 33901 17091 33917
rect 17393 33951 17427 33967
rect 17393 33901 17427 33917
rect 17729 33951 17763 33967
rect 17729 33901 17763 33917
rect 18065 33951 18099 33967
rect 18065 33901 18099 33917
rect 18401 33951 18435 33967
rect 18401 33901 18435 33917
rect 18737 33951 18771 33967
rect 18737 33901 18771 33917
rect 19073 33951 19107 33967
rect 19073 33901 19107 33917
rect 19409 33951 19443 33967
rect 19409 33901 19443 33917
rect 19745 33951 19779 33967
rect 19745 33901 19779 33917
rect 20081 33951 20115 33967
rect 20081 33901 20115 33917
rect 20417 33951 20451 33967
rect 20417 33901 20451 33917
rect 20753 33951 20787 33967
rect 20753 33901 20787 33917
rect 21089 33951 21123 33967
rect 21089 33901 21123 33917
rect 21425 33951 21459 33967
rect 21425 33901 21459 33917
rect 21761 33951 21795 33967
rect 21761 33901 21795 33917
rect 22097 33951 22131 33967
rect 22097 33901 22131 33917
rect 22433 33951 22467 33967
rect 22433 33901 22467 33917
rect 22769 33951 22803 33967
rect 22769 33901 22803 33917
rect 23105 33951 23139 33967
rect 23105 33901 23139 33917
rect 23441 33951 23475 33967
rect 23441 33901 23475 33917
rect 23777 33951 23811 33967
rect 23777 33901 23811 33917
rect 1601 33461 1635 33477
rect 1601 33411 1635 33427
rect 24181 33461 24215 33477
rect 24181 33411 24215 33427
rect 1601 33125 1635 33141
rect 1601 33075 1635 33091
rect 24181 33125 24215 33141
rect 24181 33075 24215 33091
rect 1601 32789 1635 32805
rect 1601 32739 1635 32755
rect 24181 32789 24215 32805
rect 24181 32739 24215 32755
rect 1601 32453 1635 32469
rect 1601 32403 1635 32419
rect 24181 32453 24215 32469
rect 24181 32403 24215 32419
rect 1601 32117 1635 32133
rect 1601 32067 1635 32083
rect 24181 32117 24215 32133
rect 24181 32067 24215 32083
rect 1601 31781 1635 31797
rect 1601 31731 1635 31747
rect 24181 31781 24215 31797
rect 24181 31731 24215 31747
rect 1601 31445 1635 31461
rect 1601 31395 1635 31411
rect 24181 31445 24215 31461
rect 24181 31395 24215 31411
rect 1601 31109 1635 31125
rect 1601 31059 1635 31075
rect 24181 31109 24215 31125
rect 24181 31059 24215 31075
rect 1601 30773 1635 30789
rect 1601 30723 1635 30739
rect 24181 30773 24215 30789
rect 24181 30723 24215 30739
rect 1601 30437 1635 30453
rect 1601 30387 1635 30403
rect 24181 30437 24215 30453
rect 24181 30387 24215 30403
rect 1601 30101 1635 30117
rect 1601 30051 1635 30067
rect 24181 30101 24215 30117
rect 24181 30051 24215 30067
rect 1601 29765 1635 29781
rect 1601 29715 1635 29731
rect 24181 29765 24215 29781
rect 24181 29715 24215 29731
rect 1601 29429 1635 29445
rect 1601 29379 1635 29395
rect 24181 29429 24215 29445
rect 24181 29379 24215 29395
rect 1601 29093 1635 29109
rect 1601 29043 1635 29059
rect 24181 29093 24215 29109
rect 24181 29043 24215 29059
rect 1601 28757 1635 28773
rect 1601 28707 1635 28723
rect 24181 28757 24215 28773
rect 24181 28707 24215 28723
rect 1601 28421 1635 28437
rect 1601 28371 1635 28387
rect 24181 28421 24215 28437
rect 24181 28371 24215 28387
rect 1601 28085 1635 28101
rect 1601 28035 1635 28051
rect 24181 28085 24215 28101
rect 24181 28035 24215 28051
rect 1601 27749 1635 27765
rect 1601 27699 1635 27715
rect 24181 27749 24215 27765
rect 24181 27699 24215 27715
rect 1601 27413 1635 27429
rect 1601 27363 1635 27379
rect 24181 27413 24215 27429
rect 24181 27363 24215 27379
rect 1601 27077 1635 27093
rect 1601 27027 1635 27043
rect 24181 27077 24215 27093
rect 24181 27027 24215 27043
rect 1601 26741 1635 26757
rect 1601 26691 1635 26707
rect 24181 26741 24215 26757
rect 24181 26691 24215 26707
rect 1601 26405 1635 26421
rect 1601 26355 1635 26371
rect 24181 26405 24215 26421
rect 24181 26355 24215 26371
rect 1601 26069 1635 26085
rect 1601 26019 1635 26035
rect 24181 26069 24215 26085
rect 24181 26019 24215 26035
rect 1601 25733 1635 25749
rect 1601 25683 1635 25699
rect 24181 25733 24215 25749
rect 24181 25683 24215 25699
rect 1601 25397 1635 25413
rect 1601 25347 1635 25363
rect 24181 25397 24215 25413
rect 24181 25347 24215 25363
rect 1601 25061 1635 25077
rect 1601 25011 1635 25027
rect 24181 25061 24215 25077
rect 24181 25011 24215 25027
rect 1601 24725 1635 24741
rect 1601 24675 1635 24691
rect 24181 24725 24215 24741
rect 24181 24675 24215 24691
rect 1601 24389 1635 24405
rect 1601 24339 1635 24355
rect 24181 24389 24215 24405
rect 24181 24339 24215 24355
rect 1601 24053 1635 24069
rect 1601 24003 1635 24019
rect 24181 24053 24215 24069
rect 24181 24003 24215 24019
rect 1601 23717 1635 23733
rect 1601 23667 1635 23683
rect 24181 23717 24215 23733
rect 24181 23667 24215 23683
rect 1601 23381 1635 23397
rect 1601 23331 1635 23347
rect 24181 23381 24215 23397
rect 24181 23331 24215 23347
rect 1601 23045 1635 23061
rect 1601 22995 1635 23011
rect 24181 23045 24215 23061
rect 24181 22995 24215 23011
rect 1601 22709 1635 22725
rect 1601 22659 1635 22675
rect 24181 22709 24215 22725
rect 24181 22659 24215 22675
rect 1601 22373 1635 22389
rect 1601 22323 1635 22339
rect 24181 22373 24215 22389
rect 24181 22323 24215 22339
rect 1601 22037 1635 22053
rect 1601 21987 1635 22003
rect 24181 22037 24215 22053
rect 24181 21987 24215 22003
rect 1601 21701 1635 21717
rect 1601 21651 1635 21667
rect 24181 21701 24215 21717
rect 24181 21651 24215 21667
rect 1601 21365 1635 21381
rect 1601 21315 1635 21331
rect 24181 21365 24215 21381
rect 24181 21315 24215 21331
rect 1601 21029 1635 21045
rect 1601 20979 1635 20995
rect 24181 21029 24215 21045
rect 24181 20979 24215 20995
rect 1601 20693 1635 20709
rect 1601 20643 1635 20659
rect 24181 20693 24215 20709
rect 24181 20643 24215 20659
rect 1601 20357 1635 20373
rect 1601 20307 1635 20323
rect 24181 20357 24215 20373
rect 24181 20307 24215 20323
rect 1601 20021 1635 20037
rect 1601 19971 1635 19987
rect 24181 20021 24215 20037
rect 24181 19971 24215 19987
rect 1601 19685 1635 19701
rect 1601 19635 1635 19651
rect 24181 19685 24215 19701
rect 24181 19635 24215 19651
rect 1601 19349 1635 19365
rect 1601 19299 1635 19315
rect 24181 19349 24215 19365
rect 24181 19299 24215 19315
rect 1601 19013 1635 19029
rect 1601 18963 1635 18979
rect 24181 19013 24215 19029
rect 24181 18963 24215 18979
rect 1601 18677 1635 18693
rect 1601 18627 1635 18643
rect 24181 18677 24215 18693
rect 24181 18627 24215 18643
rect 1601 18341 1635 18357
rect 1601 18291 1635 18307
rect 24181 18341 24215 18357
rect 24181 18291 24215 18307
rect 1601 18005 1635 18021
rect 1601 17955 1635 17971
rect 24181 18005 24215 18021
rect 24181 17955 24215 17971
rect 1601 17669 1635 17685
rect 1601 17619 1635 17635
rect 24181 17669 24215 17685
rect 24181 17619 24215 17635
rect 1601 17333 1635 17349
rect 1601 17283 1635 17299
rect 24181 17333 24215 17349
rect 24181 17283 24215 17299
rect 1601 16997 1635 17013
rect 1601 16947 1635 16963
rect 24181 16997 24215 17013
rect 24181 16947 24215 16963
rect 1601 16661 1635 16677
rect 1601 16611 1635 16627
rect 24181 16661 24215 16677
rect 24181 16611 24215 16627
rect 1601 16325 1635 16341
rect 1601 16275 1635 16291
rect 24181 16325 24215 16341
rect 24181 16275 24215 16291
rect 1601 15989 1635 16005
rect 1601 15939 1635 15955
rect 24181 15989 24215 16005
rect 24181 15939 24215 15955
rect 1601 15653 1635 15669
rect 1601 15603 1635 15619
rect 24181 15653 24215 15669
rect 24181 15603 24215 15619
rect 1601 15317 1635 15333
rect 1601 15267 1635 15283
rect 24181 15317 24215 15333
rect 24181 15267 24215 15283
rect 1601 14981 1635 14997
rect 1601 14931 1635 14947
rect 24181 14981 24215 14997
rect 24181 14931 24215 14947
rect 1601 14645 1635 14661
rect 1601 14595 1635 14611
rect 24181 14645 24215 14661
rect 24181 14595 24215 14611
rect 1601 14309 1635 14325
rect 1601 14259 1635 14275
rect 24181 14309 24215 14325
rect 24181 14259 24215 14275
rect 1601 13973 1635 13989
rect 1601 13923 1635 13939
rect 24181 13973 24215 13989
rect 24181 13923 24215 13939
rect 1601 13637 1635 13653
rect 1601 13587 1635 13603
rect 24181 13637 24215 13653
rect 24181 13587 24215 13603
rect 1601 13301 1635 13317
rect 1601 13251 1635 13267
rect 24181 13301 24215 13317
rect 24181 13251 24215 13267
rect 1601 12965 1635 12981
rect 1601 12915 1635 12931
rect 24181 12965 24215 12981
rect 24181 12915 24215 12931
rect 1601 12629 1635 12645
rect 1601 12579 1635 12595
rect 24181 12629 24215 12645
rect 24181 12579 24215 12595
rect 1601 12293 1635 12309
rect 1601 12243 1635 12259
rect 24181 12293 24215 12309
rect 24181 12243 24215 12259
rect 1601 11957 1635 11973
rect 1601 11907 1635 11923
rect 24181 11957 24215 11973
rect 24181 11907 24215 11923
rect 1601 11621 1635 11637
rect 1601 11571 1635 11587
rect 24181 11621 24215 11637
rect 24181 11571 24215 11587
rect 1601 11285 1635 11301
rect 1601 11235 1635 11251
rect 24181 11285 24215 11301
rect 24181 11235 24215 11251
rect 1601 10949 1635 10965
rect 1601 10899 1635 10915
rect 24181 10949 24215 10965
rect 24181 10899 24215 10915
rect 1601 10613 1635 10629
rect 1601 10563 1635 10579
rect 24181 10613 24215 10629
rect 24181 10563 24215 10579
rect 1601 10277 1635 10293
rect 1601 10227 1635 10243
rect 24181 10277 24215 10293
rect 24181 10227 24215 10243
rect 1601 9941 1635 9957
rect 1601 9891 1635 9907
rect 24181 9941 24215 9957
rect 24181 9891 24215 9907
rect 1601 9605 1635 9621
rect 1601 9555 1635 9571
rect 24181 9605 24215 9621
rect 24181 9555 24215 9571
rect 1601 9269 1635 9285
rect 1601 9219 1635 9235
rect 24181 9269 24215 9285
rect 24181 9219 24215 9235
rect 1601 8933 1635 8949
rect 1601 8883 1635 8899
rect 24181 8933 24215 8949
rect 24181 8883 24215 8899
rect 1601 8597 1635 8613
rect 1601 8547 1635 8563
rect 24181 8597 24215 8613
rect 24181 8547 24215 8563
rect 1601 8261 1635 8277
rect 1601 8211 1635 8227
rect 24181 8261 24215 8277
rect 24181 8211 24215 8227
rect 1601 7925 1635 7941
rect 1601 7875 1635 7891
rect 24181 7925 24215 7941
rect 24181 7875 24215 7891
rect 1601 7589 1635 7605
rect 1601 7539 1635 7555
rect 24181 7589 24215 7605
rect 24181 7539 24215 7555
rect 1601 7253 1635 7269
rect 1601 7203 1635 7219
rect 24181 7253 24215 7269
rect 24181 7203 24215 7219
rect 1601 6917 1635 6933
rect 1601 6867 1635 6883
rect 24181 6917 24215 6933
rect 24181 6867 24215 6883
rect 1601 6581 1635 6597
rect 1601 6531 1635 6547
rect 24181 6581 24215 6597
rect 24181 6531 24215 6547
rect 1601 6245 1635 6261
rect 1601 6195 1635 6211
rect 24181 6245 24215 6261
rect 24181 6195 24215 6211
rect 1601 5909 1635 5925
rect 1601 5859 1635 5875
rect 24181 5909 24215 5925
rect 24181 5859 24215 5875
rect 1601 5573 1635 5589
rect 1601 5523 1635 5539
rect 24181 5573 24215 5589
rect 24181 5523 24215 5539
rect 1601 5237 1635 5253
rect 1601 5187 1635 5203
rect 24181 5237 24215 5253
rect 24181 5187 24215 5203
rect 1601 4901 1635 4917
rect 1601 4851 1635 4867
rect 24181 4901 24215 4917
rect 24181 4851 24215 4867
rect 1601 4565 1635 4581
rect 1601 4515 1635 4531
rect 24181 4565 24215 4581
rect 24181 4515 24215 4531
rect 1601 4229 1635 4245
rect 1601 4179 1635 4195
rect 24181 4229 24215 4245
rect 24181 4179 24215 4195
rect 1601 3893 1635 3909
rect 1601 3843 1635 3859
rect 24181 3893 24215 3909
rect 24181 3843 24215 3859
rect 1601 3557 1635 3573
rect 1601 3507 1635 3523
rect 24181 3557 24215 3573
rect 24181 3507 24215 3523
rect 1601 3221 1635 3237
rect 1601 3171 1635 3187
rect 24181 3221 24215 3237
rect 24181 3171 24215 3187
rect 1601 2885 1635 2901
rect 1601 2835 1635 2851
rect 24181 2885 24215 2901
rect 24181 2835 24215 2851
rect 1601 2549 1635 2565
rect 1601 2499 1635 2515
rect 24181 2549 24215 2565
rect 24181 2499 24215 2515
rect 1601 2213 1635 2229
rect 1601 2163 1635 2179
rect 24181 2213 24215 2229
rect 24181 2163 24215 2179
rect 1601 1877 1635 1893
rect 1601 1827 1635 1843
rect 24181 1877 24215 1893
rect 24181 1827 24215 1843
rect 1937 1541 1971 1557
rect 1937 1491 1971 1507
rect 2273 1541 2307 1557
rect 2273 1491 2307 1507
rect 2609 1541 2643 1557
rect 2609 1491 2643 1507
rect 2945 1541 2979 1557
rect 2945 1491 2979 1507
rect 3281 1541 3315 1557
rect 3281 1491 3315 1507
rect 3617 1541 3651 1557
rect 3617 1491 3651 1507
rect 3953 1541 3987 1557
rect 3953 1491 3987 1507
rect 4289 1541 4323 1557
rect 4289 1491 4323 1507
rect 4625 1541 4659 1557
rect 4625 1491 4659 1507
rect 4961 1541 4995 1557
rect 4961 1491 4995 1507
rect 5297 1541 5331 1557
rect 5297 1491 5331 1507
rect 5633 1541 5667 1557
rect 5633 1491 5667 1507
rect 5969 1541 6003 1557
rect 5969 1491 6003 1507
rect 6305 1541 6339 1557
rect 6305 1491 6339 1507
rect 6641 1541 6675 1557
rect 6641 1491 6675 1507
rect 6977 1541 7011 1557
rect 6977 1491 7011 1507
rect 7313 1541 7347 1557
rect 7313 1491 7347 1507
rect 7649 1541 7683 1557
rect 7649 1491 7683 1507
rect 7985 1541 8019 1557
rect 7985 1491 8019 1507
rect 8321 1541 8355 1557
rect 8321 1491 8355 1507
rect 8657 1541 8691 1557
rect 8657 1491 8691 1507
rect 8993 1541 9027 1557
rect 8993 1491 9027 1507
rect 9329 1541 9363 1557
rect 9329 1491 9363 1507
rect 9665 1541 9699 1557
rect 9665 1491 9699 1507
rect 10001 1541 10035 1557
rect 10001 1491 10035 1507
rect 10337 1541 10371 1557
rect 10337 1491 10371 1507
rect 10673 1541 10707 1557
rect 10673 1491 10707 1507
rect 11009 1541 11043 1557
rect 11009 1491 11043 1507
rect 11345 1541 11379 1557
rect 11345 1491 11379 1507
rect 11681 1541 11715 1557
rect 11681 1491 11715 1507
rect 12017 1541 12051 1557
rect 12017 1491 12051 1507
rect 12353 1541 12387 1557
rect 12353 1491 12387 1507
rect 12689 1541 12723 1557
rect 12689 1491 12723 1507
rect 13025 1541 13059 1557
rect 13025 1491 13059 1507
rect 13361 1541 13395 1557
rect 13361 1491 13395 1507
rect 13697 1541 13731 1557
rect 13697 1491 13731 1507
rect 14033 1541 14067 1557
rect 14033 1491 14067 1507
rect 14369 1541 14403 1557
rect 14369 1491 14403 1507
rect 14705 1541 14739 1557
rect 14705 1491 14739 1507
rect 15041 1541 15075 1557
rect 15041 1491 15075 1507
rect 15377 1541 15411 1557
rect 15377 1491 15411 1507
rect 15713 1541 15747 1557
rect 15713 1491 15747 1507
rect 16049 1541 16083 1557
rect 16049 1491 16083 1507
rect 16385 1541 16419 1557
rect 16385 1491 16419 1507
rect 16721 1541 16755 1557
rect 16721 1491 16755 1507
rect 17057 1541 17091 1557
rect 17057 1491 17091 1507
rect 17393 1541 17427 1557
rect 17393 1491 17427 1507
rect 17729 1541 17763 1557
rect 17729 1491 17763 1507
rect 18065 1541 18099 1557
rect 18065 1491 18099 1507
rect 18401 1541 18435 1557
rect 18401 1491 18435 1507
rect 18737 1541 18771 1557
rect 18737 1491 18771 1507
rect 19073 1541 19107 1557
rect 19073 1491 19107 1507
rect 19409 1541 19443 1557
rect 19409 1491 19443 1507
rect 19745 1541 19779 1557
rect 19745 1491 19779 1507
rect 20081 1541 20115 1557
rect 20081 1491 20115 1507
rect 20417 1541 20451 1557
rect 20417 1491 20451 1507
rect 20753 1541 20787 1557
rect 20753 1491 20787 1507
rect 21089 1541 21123 1557
rect 21089 1491 21123 1507
rect 21425 1541 21459 1557
rect 21425 1491 21459 1507
rect 21761 1541 21795 1557
rect 21761 1491 21795 1507
rect 22097 1541 22131 1557
rect 22097 1491 22131 1507
rect 22433 1541 22467 1557
rect 22433 1491 22467 1507
rect 22769 1541 22803 1557
rect 22769 1491 22803 1507
rect 23105 1541 23139 1557
rect 23105 1491 23139 1507
rect 23441 1541 23475 1557
rect 23441 1491 23475 1507
rect 23777 1541 23811 1557
rect 23777 1491 23811 1507
<< viali >>
rect 1937 33917 1971 33951
rect 2273 33917 2307 33951
rect 2609 33917 2643 33951
rect 2945 33917 2979 33951
rect 3281 33917 3315 33951
rect 3617 33917 3651 33951
rect 3953 33917 3987 33951
rect 4289 33917 4323 33951
rect 4625 33917 4659 33951
rect 4961 33917 4995 33951
rect 5297 33917 5331 33951
rect 5633 33917 5667 33951
rect 5969 33917 6003 33951
rect 6305 33917 6339 33951
rect 6641 33917 6675 33951
rect 6977 33917 7011 33951
rect 7313 33917 7347 33951
rect 7649 33917 7683 33951
rect 7985 33917 8019 33951
rect 8321 33917 8355 33951
rect 8657 33917 8691 33951
rect 8993 33917 9027 33951
rect 9329 33917 9363 33951
rect 9665 33917 9699 33951
rect 10001 33917 10035 33951
rect 10337 33917 10371 33951
rect 10673 33917 10707 33951
rect 11009 33917 11043 33951
rect 11345 33917 11379 33951
rect 11681 33917 11715 33951
rect 12017 33917 12051 33951
rect 12353 33917 12387 33951
rect 12689 33917 12723 33951
rect 13025 33917 13059 33951
rect 13361 33917 13395 33951
rect 13697 33917 13731 33951
rect 14033 33917 14067 33951
rect 14369 33917 14403 33951
rect 14705 33917 14739 33951
rect 15041 33917 15075 33951
rect 15377 33917 15411 33951
rect 15713 33917 15747 33951
rect 16049 33917 16083 33951
rect 16385 33917 16419 33951
rect 16721 33917 16755 33951
rect 17057 33917 17091 33951
rect 17393 33917 17427 33951
rect 17729 33917 17763 33951
rect 18065 33917 18099 33951
rect 18401 33917 18435 33951
rect 18737 33917 18771 33951
rect 19073 33917 19107 33951
rect 19409 33917 19443 33951
rect 19745 33917 19779 33951
rect 20081 33917 20115 33951
rect 20417 33917 20451 33951
rect 20753 33917 20787 33951
rect 21089 33917 21123 33951
rect 21425 33917 21459 33951
rect 21761 33917 21795 33951
rect 22097 33917 22131 33951
rect 22433 33917 22467 33951
rect 22769 33917 22803 33951
rect 23105 33917 23139 33951
rect 23441 33917 23475 33951
rect 23777 33917 23811 33951
rect 1601 33427 1635 33461
rect 24181 33427 24215 33461
rect 1601 33091 1635 33125
rect 24181 33091 24215 33125
rect 1601 32755 1635 32789
rect 24181 32755 24215 32789
rect 1601 32419 1635 32453
rect 24181 32419 24215 32453
rect 1601 32083 1635 32117
rect 24181 32083 24215 32117
rect 1601 31747 1635 31781
rect 24181 31747 24215 31781
rect 1601 31411 1635 31445
rect 24181 31411 24215 31445
rect 1601 31075 1635 31109
rect 24181 31075 24215 31109
rect 1601 30739 1635 30773
rect 24181 30739 24215 30773
rect 1601 30403 1635 30437
rect 24181 30403 24215 30437
rect 1601 30067 1635 30101
rect 24181 30067 24215 30101
rect 1601 29731 1635 29765
rect 24181 29731 24215 29765
rect 1601 29395 1635 29429
rect 24181 29395 24215 29429
rect 1601 29059 1635 29093
rect 24181 29059 24215 29093
rect 1601 28723 1635 28757
rect 24181 28723 24215 28757
rect 1601 28387 1635 28421
rect 24181 28387 24215 28421
rect 1601 28051 1635 28085
rect 24181 28051 24215 28085
rect 1601 27715 1635 27749
rect 24181 27715 24215 27749
rect 1601 27379 1635 27413
rect 24181 27379 24215 27413
rect 1601 27043 1635 27077
rect 24181 27043 24215 27077
rect 1601 26707 1635 26741
rect 24181 26707 24215 26741
rect 1601 26371 1635 26405
rect 24181 26371 24215 26405
rect 1601 26035 1635 26069
rect 24181 26035 24215 26069
rect 1601 25699 1635 25733
rect 24181 25699 24215 25733
rect 1601 25363 1635 25397
rect 24181 25363 24215 25397
rect 1601 25027 1635 25061
rect 24181 25027 24215 25061
rect 1601 24691 1635 24725
rect 24181 24691 24215 24725
rect 1601 24355 1635 24389
rect 24181 24355 24215 24389
rect 1601 24019 1635 24053
rect 24181 24019 24215 24053
rect 1601 23683 1635 23717
rect 24181 23683 24215 23717
rect 1601 23347 1635 23381
rect 24181 23347 24215 23381
rect 1601 23011 1635 23045
rect 24181 23011 24215 23045
rect 1601 22675 1635 22709
rect 24181 22675 24215 22709
rect 1601 22339 1635 22373
rect 24181 22339 24215 22373
rect 1601 22003 1635 22037
rect 24181 22003 24215 22037
rect 1601 21667 1635 21701
rect 24181 21667 24215 21701
rect 1601 21331 1635 21365
rect 24181 21331 24215 21365
rect 1601 20995 1635 21029
rect 24181 20995 24215 21029
rect 1601 20659 1635 20693
rect 24181 20659 24215 20693
rect 1601 20323 1635 20357
rect 24181 20323 24215 20357
rect 1601 19987 1635 20021
rect 24181 19987 24215 20021
rect 1601 19651 1635 19685
rect 24181 19651 24215 19685
rect 1601 19315 1635 19349
rect 24181 19315 24215 19349
rect 1601 18979 1635 19013
rect 24181 18979 24215 19013
rect 1601 18643 1635 18677
rect 24181 18643 24215 18677
rect 1601 18307 1635 18341
rect 24181 18307 24215 18341
rect 1601 17971 1635 18005
rect 24181 17971 24215 18005
rect 1601 17635 1635 17669
rect 24181 17635 24215 17669
rect 1601 17299 1635 17333
rect 24181 17299 24215 17333
rect 1601 16963 1635 16997
rect 24181 16963 24215 16997
rect 1601 16627 1635 16661
rect 24181 16627 24215 16661
rect 1601 16291 1635 16325
rect 24181 16291 24215 16325
rect 1601 15955 1635 15989
rect 24181 15955 24215 15989
rect 1601 15619 1635 15653
rect 24181 15619 24215 15653
rect 1601 15283 1635 15317
rect 24181 15283 24215 15317
rect 1601 14947 1635 14981
rect 24181 14947 24215 14981
rect 1601 14611 1635 14645
rect 24181 14611 24215 14645
rect 1601 14275 1635 14309
rect 24181 14275 24215 14309
rect 1601 13939 1635 13973
rect 24181 13939 24215 13973
rect 1601 13603 1635 13637
rect 24181 13603 24215 13637
rect 1601 13267 1635 13301
rect 24181 13267 24215 13301
rect 1601 12931 1635 12965
rect 24181 12931 24215 12965
rect 1601 12595 1635 12629
rect 24181 12595 24215 12629
rect 1601 12259 1635 12293
rect 24181 12259 24215 12293
rect 1601 11923 1635 11957
rect 24181 11923 24215 11957
rect 1601 11587 1635 11621
rect 24181 11587 24215 11621
rect 1601 11251 1635 11285
rect 24181 11251 24215 11285
rect 1601 10915 1635 10949
rect 24181 10915 24215 10949
rect 1601 10579 1635 10613
rect 24181 10579 24215 10613
rect 1601 10243 1635 10277
rect 24181 10243 24215 10277
rect 1601 9907 1635 9941
rect 24181 9907 24215 9941
rect 1601 9571 1635 9605
rect 24181 9571 24215 9605
rect 1601 9235 1635 9269
rect 24181 9235 24215 9269
rect 1601 8899 1635 8933
rect 24181 8899 24215 8933
rect 1601 8563 1635 8597
rect 24181 8563 24215 8597
rect 1601 8227 1635 8261
rect 24181 8227 24215 8261
rect 1601 7891 1635 7925
rect 24181 7891 24215 7925
rect 1601 7555 1635 7589
rect 24181 7555 24215 7589
rect 1601 7219 1635 7253
rect 24181 7219 24215 7253
rect 1601 6883 1635 6917
rect 24181 6883 24215 6917
rect 1601 6547 1635 6581
rect 24181 6547 24215 6581
rect 1601 6211 1635 6245
rect 24181 6211 24215 6245
rect 1601 5875 1635 5909
rect 24181 5875 24215 5909
rect 1601 5539 1635 5573
rect 24181 5539 24215 5573
rect 1601 5203 1635 5237
rect 24181 5203 24215 5237
rect 1601 4867 1635 4901
rect 24181 4867 24215 4901
rect 1601 4531 1635 4565
rect 24181 4531 24215 4565
rect 1601 4195 1635 4229
rect 24181 4195 24215 4229
rect 1601 3859 1635 3893
rect 24181 3859 24215 3893
rect 1601 3523 1635 3557
rect 24181 3523 24215 3557
rect 1601 3187 1635 3221
rect 24181 3187 24215 3221
rect 1601 2851 1635 2885
rect 24181 2851 24215 2885
rect 1601 2515 1635 2549
rect 24181 2515 24215 2549
rect 1601 2179 1635 2213
rect 24181 2179 24215 2213
rect 1601 1843 1635 1877
rect 24181 1843 24215 1877
rect 1937 1507 1971 1541
rect 2273 1507 2307 1541
rect 2609 1507 2643 1541
rect 2945 1507 2979 1541
rect 3281 1507 3315 1541
rect 3617 1507 3651 1541
rect 3953 1507 3987 1541
rect 4289 1507 4323 1541
rect 4625 1507 4659 1541
rect 4961 1507 4995 1541
rect 5297 1507 5331 1541
rect 5633 1507 5667 1541
rect 5969 1507 6003 1541
rect 6305 1507 6339 1541
rect 6641 1507 6675 1541
rect 6977 1507 7011 1541
rect 7313 1507 7347 1541
rect 7649 1507 7683 1541
rect 7985 1507 8019 1541
rect 8321 1507 8355 1541
rect 8657 1507 8691 1541
rect 8993 1507 9027 1541
rect 9329 1507 9363 1541
rect 9665 1507 9699 1541
rect 10001 1507 10035 1541
rect 10337 1507 10371 1541
rect 10673 1507 10707 1541
rect 11009 1507 11043 1541
rect 11345 1507 11379 1541
rect 11681 1507 11715 1541
rect 12017 1507 12051 1541
rect 12353 1507 12387 1541
rect 12689 1507 12723 1541
rect 13025 1507 13059 1541
rect 13361 1507 13395 1541
rect 13697 1507 13731 1541
rect 14033 1507 14067 1541
rect 14369 1507 14403 1541
rect 14705 1507 14739 1541
rect 15041 1507 15075 1541
rect 15377 1507 15411 1541
rect 15713 1507 15747 1541
rect 16049 1507 16083 1541
rect 16385 1507 16419 1541
rect 16721 1507 16755 1541
rect 17057 1507 17091 1541
rect 17393 1507 17427 1541
rect 17729 1507 17763 1541
rect 18065 1507 18099 1541
rect 18401 1507 18435 1541
rect 18737 1507 18771 1541
rect 19073 1507 19107 1541
rect 19409 1507 19443 1541
rect 19745 1507 19779 1541
rect 20081 1507 20115 1541
rect 20417 1507 20451 1541
rect 20753 1507 20787 1541
rect 21089 1507 21123 1541
rect 21425 1507 21459 1541
rect 21761 1507 21795 1541
rect 22097 1507 22131 1541
rect 22433 1507 22467 1541
rect 22769 1507 22803 1541
rect 23105 1507 23139 1541
rect 23441 1507 23475 1541
rect 23777 1507 23811 1541
<< metal1 >>
rect 1506 33960 24310 34046
rect 1506 33908 1928 33960
rect 1980 33951 3608 33960
rect 3660 33951 5288 33960
rect 5340 33951 6968 33960
rect 7020 33951 8648 33960
rect 8700 33951 10328 33960
rect 10380 33951 12008 33960
rect 12060 33951 13688 33960
rect 13740 33951 15368 33960
rect 15420 33951 17048 33960
rect 17100 33951 18728 33960
rect 18780 33951 20408 33960
rect 20460 33951 22088 33960
rect 22140 33951 23768 33960
rect 1980 33917 2273 33951
rect 2307 33917 2609 33951
rect 2643 33917 2945 33951
rect 2979 33917 3281 33951
rect 3315 33917 3608 33951
rect 3660 33917 3953 33951
rect 3987 33917 4289 33951
rect 4323 33917 4625 33951
rect 4659 33917 4961 33951
rect 4995 33917 5288 33951
rect 5340 33917 5633 33951
rect 5667 33917 5969 33951
rect 6003 33917 6305 33951
rect 6339 33917 6641 33951
rect 6675 33917 6968 33951
rect 7020 33917 7313 33951
rect 7347 33917 7649 33951
rect 7683 33917 7985 33951
rect 8019 33917 8321 33951
rect 8355 33917 8648 33951
rect 8700 33917 8993 33951
rect 9027 33917 9329 33951
rect 9363 33917 9665 33951
rect 9699 33917 10001 33951
rect 10035 33917 10328 33951
rect 10380 33917 10673 33951
rect 10707 33917 11009 33951
rect 11043 33917 11345 33951
rect 11379 33917 11681 33951
rect 11715 33917 12008 33951
rect 12060 33917 12353 33951
rect 12387 33917 12689 33951
rect 12723 33917 13025 33951
rect 13059 33917 13361 33951
rect 13395 33917 13688 33951
rect 13740 33917 14033 33951
rect 14067 33917 14369 33951
rect 14403 33917 14705 33951
rect 14739 33917 15041 33951
rect 15075 33917 15368 33951
rect 15420 33917 15713 33951
rect 15747 33917 16049 33951
rect 16083 33917 16385 33951
rect 16419 33917 16721 33951
rect 16755 33917 17048 33951
rect 17100 33917 17393 33951
rect 17427 33917 17729 33951
rect 17763 33917 18065 33951
rect 18099 33917 18401 33951
rect 18435 33917 18728 33951
rect 18780 33917 19073 33951
rect 19107 33917 19409 33951
rect 19443 33917 19745 33951
rect 19779 33917 20081 33951
rect 20115 33917 20408 33951
rect 20460 33917 20753 33951
rect 20787 33917 21089 33951
rect 21123 33917 21425 33951
rect 21459 33917 21761 33951
rect 21795 33917 22088 33951
rect 22140 33917 22433 33951
rect 22467 33917 22769 33951
rect 22803 33917 23105 33951
rect 23139 33917 23441 33951
rect 23475 33917 23768 33951
rect 1980 33908 3608 33917
rect 3660 33908 5288 33917
rect 5340 33908 6968 33917
rect 7020 33908 8648 33917
rect 8700 33908 10328 33917
rect 10380 33908 12008 33917
rect 12060 33908 13688 33917
rect 13740 33908 15368 33917
rect 15420 33908 17048 33917
rect 17100 33908 18728 33917
rect 18780 33908 20408 33917
rect 20460 33908 22088 33917
rect 22140 33908 23768 33917
rect 23820 33908 24310 33960
rect 1506 33822 24310 33908
rect 1586 33418 1592 33470
rect 1644 33418 1650 33470
rect 24166 33418 24172 33470
rect 24224 33418 24230 33470
rect 1586 33082 1592 33134
rect 1644 33082 1650 33134
rect 24166 33082 24172 33134
rect 24224 33082 24230 33134
rect 1586 32746 1592 32798
rect 1644 32746 1650 32798
rect 24166 32746 24172 32798
rect 24224 32746 24230 32798
rect 1586 32410 1592 32462
rect 1644 32410 1650 32462
rect 24166 32410 24172 32462
rect 24224 32410 24230 32462
rect 1586 32074 1592 32126
rect 1644 32074 1650 32126
rect 24166 32074 24172 32126
rect 24224 32074 24230 32126
rect 1586 31738 1592 31790
rect 1644 31738 1650 31790
rect 24166 31738 24172 31790
rect 24224 31738 24230 31790
rect 1586 31402 1592 31454
rect 1644 31402 1650 31454
rect 24166 31402 24172 31454
rect 24224 31402 24230 31454
rect 1586 31066 1592 31118
rect 1644 31066 1650 31118
rect 24166 31066 24172 31118
rect 24224 31066 24230 31118
rect 1586 30730 1592 30782
rect 1644 30730 1650 30782
rect 24166 30730 24172 30782
rect 24224 30730 24230 30782
rect 1586 30394 1592 30446
rect 1644 30394 1650 30446
rect 24166 30394 24172 30446
rect 24224 30394 24230 30446
rect 1586 30058 1592 30110
rect 1644 30058 1650 30110
rect 24166 30058 24172 30110
rect 24224 30058 24230 30110
rect 1586 29722 1592 29774
rect 1644 29722 1650 29774
rect 24166 29722 24172 29774
rect 24224 29722 24230 29774
rect 1586 29386 1592 29438
rect 1644 29386 1650 29438
rect 24166 29386 24172 29438
rect 24224 29386 24230 29438
rect 1586 29050 1592 29102
rect 1644 29050 1650 29102
rect 24166 29050 24172 29102
rect 24224 29050 24230 29102
rect 1586 28714 1592 28766
rect 1644 28714 1650 28766
rect 24166 28714 24172 28766
rect 24224 28714 24230 28766
rect 1586 28378 1592 28430
rect 1644 28378 1650 28430
rect 24166 28378 24172 28430
rect 24224 28378 24230 28430
rect 1586 28042 1592 28094
rect 1644 28042 1650 28094
rect 24166 28042 24172 28094
rect 24224 28042 24230 28094
rect 1586 27706 1592 27758
rect 1644 27706 1650 27758
rect 24166 27706 24172 27758
rect 24224 27706 24230 27758
rect 1586 27370 1592 27422
rect 1644 27370 1650 27422
rect 24166 27370 24172 27422
rect 24224 27370 24230 27422
rect 1586 27034 1592 27086
rect 1644 27034 1650 27086
rect 24166 27034 24172 27086
rect 24224 27034 24230 27086
rect 1586 26698 1592 26750
rect 1644 26698 1650 26750
rect 24166 26698 24172 26750
rect 24224 26698 24230 26750
rect 1586 26362 1592 26414
rect 1644 26362 1650 26414
rect 24166 26362 24172 26414
rect 24224 26362 24230 26414
rect 1586 26026 1592 26078
rect 1644 26026 1650 26078
rect 24166 26026 24172 26078
rect 24224 26026 24230 26078
rect 1586 25690 1592 25742
rect 1644 25690 1650 25742
rect 24166 25690 24172 25742
rect 24224 25690 24230 25742
rect 1586 25354 1592 25406
rect 1644 25354 1650 25406
rect 24166 25354 24172 25406
rect 24224 25354 24230 25406
rect 1586 25018 1592 25070
rect 1644 25018 1650 25070
rect 24166 25018 24172 25070
rect 24224 25018 24230 25070
rect 1586 24682 1592 24734
rect 1644 24682 1650 24734
rect 24166 24682 24172 24734
rect 24224 24682 24230 24734
rect 1586 24346 1592 24398
rect 1644 24346 1650 24398
rect 24166 24346 24172 24398
rect 24224 24346 24230 24398
rect 1586 24010 1592 24062
rect 1644 24010 1650 24062
rect 24166 24010 24172 24062
rect 24224 24010 24230 24062
rect 1586 23674 1592 23726
rect 1644 23674 1650 23726
rect 24166 23674 24172 23726
rect 24224 23674 24230 23726
rect 1586 23338 1592 23390
rect 1644 23338 1650 23390
rect 24166 23338 24172 23390
rect 24224 23338 24230 23390
rect 1586 23002 1592 23054
rect 1644 23002 1650 23054
rect 24166 23002 24172 23054
rect 24224 23002 24230 23054
rect 1586 22666 1592 22718
rect 1644 22666 1650 22718
rect 24166 22666 24172 22718
rect 24224 22666 24230 22718
rect 1586 22330 1592 22382
rect 1644 22330 1650 22382
rect 24166 22330 24172 22382
rect 24224 22330 24230 22382
rect 1586 21994 1592 22046
rect 1644 21994 1650 22046
rect 24166 21994 24172 22046
rect 24224 21994 24230 22046
rect 1586 21658 1592 21710
rect 1644 21658 1650 21710
rect 24166 21658 24172 21710
rect 24224 21658 24230 21710
rect 1586 21322 1592 21374
rect 1644 21322 1650 21374
rect 24166 21322 24172 21374
rect 24224 21322 24230 21374
rect 1586 20986 1592 21038
rect 1644 20986 1650 21038
rect 24166 20986 24172 21038
rect 24224 20986 24230 21038
rect 1586 20650 1592 20702
rect 1644 20650 1650 20702
rect 24166 20650 24172 20702
rect 24224 20650 24230 20702
rect 1586 20314 1592 20366
rect 1644 20314 1650 20366
rect 24166 20314 24172 20366
rect 24224 20314 24230 20366
rect 1586 19978 1592 20030
rect 1644 19978 1650 20030
rect 24166 19978 24172 20030
rect 24224 19978 24230 20030
rect 1586 19642 1592 19694
rect 1644 19642 1650 19694
rect 24166 19642 24172 19694
rect 24224 19642 24230 19694
rect 1586 19306 1592 19358
rect 1644 19306 1650 19358
rect 24166 19306 24172 19358
rect 24224 19306 24230 19358
rect 1586 18970 1592 19022
rect 1644 18970 1650 19022
rect 24166 18970 24172 19022
rect 24224 18970 24230 19022
rect 1586 18634 1592 18686
rect 1644 18634 1650 18686
rect 24166 18634 24172 18686
rect 24224 18634 24230 18686
rect 1586 18298 1592 18350
rect 1644 18298 1650 18350
rect 24166 18298 24172 18350
rect 24224 18298 24230 18350
rect 1586 17962 1592 18014
rect 1644 17962 1650 18014
rect 24166 17962 24172 18014
rect 24224 17962 24230 18014
rect 1586 17626 1592 17678
rect 1644 17626 1650 17678
rect 24166 17626 24172 17678
rect 24224 17626 24230 17678
rect 1586 17290 1592 17342
rect 1644 17290 1650 17342
rect 24166 17290 24172 17342
rect 24224 17290 24230 17342
rect 1586 16954 1592 17006
rect 1644 16954 1650 17006
rect 24166 16954 24172 17006
rect 24224 16954 24230 17006
rect 1586 16618 1592 16670
rect 1644 16618 1650 16670
rect 24166 16618 24172 16670
rect 24224 16618 24230 16670
rect 1586 16282 1592 16334
rect 1644 16282 1650 16334
rect 24166 16282 24172 16334
rect 24224 16282 24230 16334
rect 1586 15946 1592 15998
rect 1644 15946 1650 15998
rect 24166 15946 24172 15998
rect 24224 15946 24230 15998
rect 1586 15610 1592 15662
rect 1644 15610 1650 15662
rect 24166 15610 24172 15662
rect 24224 15610 24230 15662
rect 1586 15274 1592 15326
rect 1644 15274 1650 15326
rect 24166 15274 24172 15326
rect 24224 15274 24230 15326
rect 1586 14938 1592 14990
rect 1644 14938 1650 14990
rect 24166 14938 24172 14990
rect 24224 14938 24230 14990
rect 1586 14602 1592 14654
rect 1644 14602 1650 14654
rect 24166 14602 24172 14654
rect 24224 14602 24230 14654
rect 1586 14266 1592 14318
rect 1644 14266 1650 14318
rect 24166 14266 24172 14318
rect 24224 14266 24230 14318
rect 1586 13930 1592 13982
rect 1644 13930 1650 13982
rect 24166 13930 24172 13982
rect 24224 13930 24230 13982
rect 1586 13594 1592 13646
rect 1644 13594 1650 13646
rect 24166 13594 24172 13646
rect 24224 13594 24230 13646
rect 1586 13258 1592 13310
rect 1644 13258 1650 13310
rect 24166 13258 24172 13310
rect 24224 13258 24230 13310
rect 1586 12922 1592 12974
rect 1644 12922 1650 12974
rect 24166 12922 24172 12974
rect 24224 12922 24230 12974
rect 1586 12586 1592 12638
rect 1644 12586 1650 12638
rect 24166 12586 24172 12638
rect 24224 12586 24230 12638
rect 1586 12250 1592 12302
rect 1644 12250 1650 12302
rect 24166 12250 24172 12302
rect 24224 12250 24230 12302
rect 1586 11914 1592 11966
rect 1644 11914 1650 11966
rect 24166 11914 24172 11966
rect 24224 11914 24230 11966
rect 1586 11578 1592 11630
rect 1644 11578 1650 11630
rect 24166 11578 24172 11630
rect 24224 11578 24230 11630
rect 1586 11242 1592 11294
rect 1644 11242 1650 11294
rect 24166 11242 24172 11294
rect 24224 11242 24230 11294
rect 1586 10906 1592 10958
rect 1644 10906 1650 10958
rect 24166 10906 24172 10958
rect 24224 10906 24230 10958
rect 1586 10570 1592 10622
rect 1644 10570 1650 10622
rect 24166 10570 24172 10622
rect 24224 10570 24230 10622
rect 1586 10234 1592 10286
rect 1644 10234 1650 10286
rect 24166 10234 24172 10286
rect 24224 10234 24230 10286
rect 1586 9898 1592 9950
rect 1644 9898 1650 9950
rect 24166 9898 24172 9950
rect 24224 9898 24230 9950
rect 1586 9562 1592 9614
rect 1644 9562 1650 9614
rect 24166 9562 24172 9614
rect 24224 9562 24230 9614
rect 1586 9226 1592 9278
rect 1644 9226 1650 9278
rect 24166 9226 24172 9278
rect 24224 9226 24230 9278
rect 1586 8890 1592 8942
rect 1644 8890 1650 8942
rect 24166 8890 24172 8942
rect 24224 8890 24230 8942
rect 1586 8554 1592 8606
rect 1644 8554 1650 8606
rect 24166 8554 24172 8606
rect 24224 8554 24230 8606
rect 1586 8218 1592 8270
rect 1644 8218 1650 8270
rect 24166 8218 24172 8270
rect 24224 8218 24230 8270
rect 1586 7882 1592 7934
rect 1644 7882 1650 7934
rect 24166 7882 24172 7934
rect 24224 7882 24230 7934
rect 1586 7546 1592 7598
rect 1644 7546 1650 7598
rect 24166 7546 24172 7598
rect 24224 7546 24230 7598
rect 1586 7210 1592 7262
rect 1644 7210 1650 7262
rect 24166 7210 24172 7262
rect 24224 7210 24230 7262
rect 1586 6874 1592 6926
rect 1644 6874 1650 6926
rect 24166 6874 24172 6926
rect 24224 6874 24230 6926
rect 1586 6538 1592 6590
rect 1644 6538 1650 6590
rect 24166 6538 24172 6590
rect 24224 6538 24230 6590
rect 1586 6202 1592 6254
rect 1644 6202 1650 6254
rect 24166 6202 24172 6254
rect 24224 6202 24230 6254
rect 1586 5866 1592 5918
rect 1644 5866 1650 5918
rect 24166 5866 24172 5918
rect 24224 5866 24230 5918
rect 1586 5530 1592 5582
rect 1644 5530 1650 5582
rect 24166 5530 24172 5582
rect 24224 5530 24230 5582
rect 1586 5194 1592 5246
rect 1644 5194 1650 5246
rect 24166 5194 24172 5246
rect 24224 5194 24230 5246
rect 1586 4858 1592 4910
rect 1644 4858 1650 4910
rect 24166 4858 24172 4910
rect 24224 4858 24230 4910
rect 1586 4522 1592 4574
rect 1644 4522 1650 4574
rect 24166 4522 24172 4574
rect 24224 4522 24230 4574
rect 1586 4186 1592 4238
rect 1644 4186 1650 4238
rect 24166 4186 24172 4238
rect 24224 4186 24230 4238
rect 1586 3850 1592 3902
rect 1644 3850 1650 3902
rect 24166 3850 24172 3902
rect 24224 3850 24230 3902
rect 1586 3514 1592 3566
rect 1644 3514 1650 3566
rect 24166 3514 24172 3566
rect 24224 3514 24230 3566
rect 1586 3178 1592 3230
rect 1644 3178 1650 3230
rect 24166 3178 24172 3230
rect 24224 3178 24230 3230
rect 1586 2842 1592 2894
rect 1644 2842 1650 2894
rect 24166 2842 24172 2894
rect 24224 2842 24230 2894
rect 1586 2506 1592 2558
rect 1644 2506 1650 2558
rect 24166 2506 24172 2558
rect 24224 2506 24230 2558
rect 1586 2170 1592 2222
rect 1644 2170 1650 2222
rect 24166 2170 24172 2222
rect 24224 2170 24230 2222
rect 1586 1834 1592 1886
rect 1644 1834 1650 1886
rect 24166 1834 24172 1886
rect 24224 1834 24230 1886
rect 1506 1550 24310 1636
rect 1506 1498 1928 1550
rect 1980 1541 3608 1550
rect 3660 1541 5288 1550
rect 5340 1541 6968 1550
rect 7020 1541 8648 1550
rect 8700 1541 10328 1550
rect 10380 1541 12008 1550
rect 12060 1541 13688 1550
rect 13740 1541 15368 1550
rect 15420 1541 17048 1550
rect 17100 1541 18728 1550
rect 18780 1541 20408 1550
rect 20460 1541 22088 1550
rect 22140 1541 23768 1550
rect 1980 1507 2273 1541
rect 2307 1507 2609 1541
rect 2643 1507 2945 1541
rect 2979 1507 3281 1541
rect 3315 1507 3608 1541
rect 3660 1507 3953 1541
rect 3987 1507 4289 1541
rect 4323 1507 4625 1541
rect 4659 1507 4961 1541
rect 4995 1507 5288 1541
rect 5340 1507 5633 1541
rect 5667 1507 5969 1541
rect 6003 1507 6305 1541
rect 6339 1507 6641 1541
rect 6675 1507 6968 1541
rect 7020 1507 7313 1541
rect 7347 1507 7649 1541
rect 7683 1507 7985 1541
rect 8019 1507 8321 1541
rect 8355 1507 8648 1541
rect 8700 1507 8993 1541
rect 9027 1507 9329 1541
rect 9363 1507 9665 1541
rect 9699 1507 10001 1541
rect 10035 1507 10328 1541
rect 10380 1507 10673 1541
rect 10707 1507 11009 1541
rect 11043 1507 11345 1541
rect 11379 1507 11681 1541
rect 11715 1507 12008 1541
rect 12060 1507 12353 1541
rect 12387 1507 12689 1541
rect 12723 1507 13025 1541
rect 13059 1507 13361 1541
rect 13395 1507 13688 1541
rect 13740 1507 14033 1541
rect 14067 1507 14369 1541
rect 14403 1507 14705 1541
rect 14739 1507 15041 1541
rect 15075 1507 15368 1541
rect 15420 1507 15713 1541
rect 15747 1507 16049 1541
rect 16083 1507 16385 1541
rect 16419 1507 16721 1541
rect 16755 1507 17048 1541
rect 17100 1507 17393 1541
rect 17427 1507 17729 1541
rect 17763 1507 18065 1541
rect 18099 1507 18401 1541
rect 18435 1507 18728 1541
rect 18780 1507 19073 1541
rect 19107 1507 19409 1541
rect 19443 1507 19745 1541
rect 19779 1507 20081 1541
rect 20115 1507 20408 1541
rect 20460 1507 20753 1541
rect 20787 1507 21089 1541
rect 21123 1507 21425 1541
rect 21459 1507 21761 1541
rect 21795 1507 22088 1541
rect 22140 1507 22433 1541
rect 22467 1507 22769 1541
rect 22803 1507 23105 1541
rect 23139 1507 23441 1541
rect 23475 1507 23768 1541
rect 1980 1498 3608 1507
rect 3660 1498 5288 1507
rect 5340 1498 6968 1507
rect 7020 1498 8648 1507
rect 8700 1498 10328 1507
rect 10380 1498 12008 1507
rect 12060 1498 13688 1507
rect 13740 1498 15368 1507
rect 15420 1498 17048 1507
rect 17100 1498 18728 1507
rect 18780 1498 20408 1507
rect 20460 1498 22088 1507
rect 22140 1498 23768 1507
rect 23820 1498 24310 1550
rect 1506 1412 24310 1498
<< via1 >>
rect 1928 33951 1980 33960
rect 3608 33951 3660 33960
rect 5288 33951 5340 33960
rect 6968 33951 7020 33960
rect 8648 33951 8700 33960
rect 10328 33951 10380 33960
rect 12008 33951 12060 33960
rect 13688 33951 13740 33960
rect 15368 33951 15420 33960
rect 17048 33951 17100 33960
rect 18728 33951 18780 33960
rect 20408 33951 20460 33960
rect 22088 33951 22140 33960
rect 23768 33951 23820 33960
rect 1928 33917 1937 33951
rect 1937 33917 1971 33951
rect 1971 33917 1980 33951
rect 3608 33917 3617 33951
rect 3617 33917 3651 33951
rect 3651 33917 3660 33951
rect 5288 33917 5297 33951
rect 5297 33917 5331 33951
rect 5331 33917 5340 33951
rect 6968 33917 6977 33951
rect 6977 33917 7011 33951
rect 7011 33917 7020 33951
rect 8648 33917 8657 33951
rect 8657 33917 8691 33951
rect 8691 33917 8700 33951
rect 10328 33917 10337 33951
rect 10337 33917 10371 33951
rect 10371 33917 10380 33951
rect 12008 33917 12017 33951
rect 12017 33917 12051 33951
rect 12051 33917 12060 33951
rect 13688 33917 13697 33951
rect 13697 33917 13731 33951
rect 13731 33917 13740 33951
rect 15368 33917 15377 33951
rect 15377 33917 15411 33951
rect 15411 33917 15420 33951
rect 17048 33917 17057 33951
rect 17057 33917 17091 33951
rect 17091 33917 17100 33951
rect 18728 33917 18737 33951
rect 18737 33917 18771 33951
rect 18771 33917 18780 33951
rect 20408 33917 20417 33951
rect 20417 33917 20451 33951
rect 20451 33917 20460 33951
rect 22088 33917 22097 33951
rect 22097 33917 22131 33951
rect 22131 33917 22140 33951
rect 23768 33917 23777 33951
rect 23777 33917 23811 33951
rect 23811 33917 23820 33951
rect 1928 33908 1980 33917
rect 3608 33908 3660 33917
rect 5288 33908 5340 33917
rect 6968 33908 7020 33917
rect 8648 33908 8700 33917
rect 10328 33908 10380 33917
rect 12008 33908 12060 33917
rect 13688 33908 13740 33917
rect 15368 33908 15420 33917
rect 17048 33908 17100 33917
rect 18728 33908 18780 33917
rect 20408 33908 20460 33917
rect 22088 33908 22140 33917
rect 23768 33908 23820 33917
rect 1592 33461 1644 33470
rect 1592 33427 1601 33461
rect 1601 33427 1635 33461
rect 1635 33427 1644 33461
rect 1592 33418 1644 33427
rect 24172 33461 24224 33470
rect 24172 33427 24181 33461
rect 24181 33427 24215 33461
rect 24215 33427 24224 33461
rect 24172 33418 24224 33427
rect 1592 33125 1644 33134
rect 1592 33091 1601 33125
rect 1601 33091 1635 33125
rect 1635 33091 1644 33125
rect 1592 33082 1644 33091
rect 24172 33125 24224 33134
rect 24172 33091 24181 33125
rect 24181 33091 24215 33125
rect 24215 33091 24224 33125
rect 24172 33082 24224 33091
rect 1592 32789 1644 32798
rect 1592 32755 1601 32789
rect 1601 32755 1635 32789
rect 1635 32755 1644 32789
rect 1592 32746 1644 32755
rect 24172 32789 24224 32798
rect 24172 32755 24181 32789
rect 24181 32755 24215 32789
rect 24215 32755 24224 32789
rect 24172 32746 24224 32755
rect 1592 32453 1644 32462
rect 1592 32419 1601 32453
rect 1601 32419 1635 32453
rect 1635 32419 1644 32453
rect 1592 32410 1644 32419
rect 24172 32453 24224 32462
rect 24172 32419 24181 32453
rect 24181 32419 24215 32453
rect 24215 32419 24224 32453
rect 24172 32410 24224 32419
rect 1592 32117 1644 32126
rect 1592 32083 1601 32117
rect 1601 32083 1635 32117
rect 1635 32083 1644 32117
rect 1592 32074 1644 32083
rect 24172 32117 24224 32126
rect 24172 32083 24181 32117
rect 24181 32083 24215 32117
rect 24215 32083 24224 32117
rect 24172 32074 24224 32083
rect 1592 31781 1644 31790
rect 1592 31747 1601 31781
rect 1601 31747 1635 31781
rect 1635 31747 1644 31781
rect 1592 31738 1644 31747
rect 24172 31781 24224 31790
rect 24172 31747 24181 31781
rect 24181 31747 24215 31781
rect 24215 31747 24224 31781
rect 24172 31738 24224 31747
rect 1592 31445 1644 31454
rect 1592 31411 1601 31445
rect 1601 31411 1635 31445
rect 1635 31411 1644 31445
rect 1592 31402 1644 31411
rect 24172 31445 24224 31454
rect 24172 31411 24181 31445
rect 24181 31411 24215 31445
rect 24215 31411 24224 31445
rect 24172 31402 24224 31411
rect 1592 31109 1644 31118
rect 1592 31075 1601 31109
rect 1601 31075 1635 31109
rect 1635 31075 1644 31109
rect 1592 31066 1644 31075
rect 24172 31109 24224 31118
rect 24172 31075 24181 31109
rect 24181 31075 24215 31109
rect 24215 31075 24224 31109
rect 24172 31066 24224 31075
rect 1592 30773 1644 30782
rect 1592 30739 1601 30773
rect 1601 30739 1635 30773
rect 1635 30739 1644 30773
rect 1592 30730 1644 30739
rect 24172 30773 24224 30782
rect 24172 30739 24181 30773
rect 24181 30739 24215 30773
rect 24215 30739 24224 30773
rect 24172 30730 24224 30739
rect 1592 30437 1644 30446
rect 1592 30403 1601 30437
rect 1601 30403 1635 30437
rect 1635 30403 1644 30437
rect 1592 30394 1644 30403
rect 24172 30437 24224 30446
rect 24172 30403 24181 30437
rect 24181 30403 24215 30437
rect 24215 30403 24224 30437
rect 24172 30394 24224 30403
rect 1592 30101 1644 30110
rect 1592 30067 1601 30101
rect 1601 30067 1635 30101
rect 1635 30067 1644 30101
rect 1592 30058 1644 30067
rect 24172 30101 24224 30110
rect 24172 30067 24181 30101
rect 24181 30067 24215 30101
rect 24215 30067 24224 30101
rect 24172 30058 24224 30067
rect 1592 29765 1644 29774
rect 1592 29731 1601 29765
rect 1601 29731 1635 29765
rect 1635 29731 1644 29765
rect 1592 29722 1644 29731
rect 24172 29765 24224 29774
rect 24172 29731 24181 29765
rect 24181 29731 24215 29765
rect 24215 29731 24224 29765
rect 24172 29722 24224 29731
rect 1592 29429 1644 29438
rect 1592 29395 1601 29429
rect 1601 29395 1635 29429
rect 1635 29395 1644 29429
rect 1592 29386 1644 29395
rect 24172 29429 24224 29438
rect 24172 29395 24181 29429
rect 24181 29395 24215 29429
rect 24215 29395 24224 29429
rect 24172 29386 24224 29395
rect 1592 29093 1644 29102
rect 1592 29059 1601 29093
rect 1601 29059 1635 29093
rect 1635 29059 1644 29093
rect 1592 29050 1644 29059
rect 24172 29093 24224 29102
rect 24172 29059 24181 29093
rect 24181 29059 24215 29093
rect 24215 29059 24224 29093
rect 24172 29050 24224 29059
rect 1592 28757 1644 28766
rect 1592 28723 1601 28757
rect 1601 28723 1635 28757
rect 1635 28723 1644 28757
rect 1592 28714 1644 28723
rect 24172 28757 24224 28766
rect 24172 28723 24181 28757
rect 24181 28723 24215 28757
rect 24215 28723 24224 28757
rect 24172 28714 24224 28723
rect 1592 28421 1644 28430
rect 1592 28387 1601 28421
rect 1601 28387 1635 28421
rect 1635 28387 1644 28421
rect 1592 28378 1644 28387
rect 24172 28421 24224 28430
rect 24172 28387 24181 28421
rect 24181 28387 24215 28421
rect 24215 28387 24224 28421
rect 24172 28378 24224 28387
rect 1592 28085 1644 28094
rect 1592 28051 1601 28085
rect 1601 28051 1635 28085
rect 1635 28051 1644 28085
rect 1592 28042 1644 28051
rect 24172 28085 24224 28094
rect 24172 28051 24181 28085
rect 24181 28051 24215 28085
rect 24215 28051 24224 28085
rect 24172 28042 24224 28051
rect 1592 27749 1644 27758
rect 1592 27715 1601 27749
rect 1601 27715 1635 27749
rect 1635 27715 1644 27749
rect 1592 27706 1644 27715
rect 24172 27749 24224 27758
rect 24172 27715 24181 27749
rect 24181 27715 24215 27749
rect 24215 27715 24224 27749
rect 24172 27706 24224 27715
rect 1592 27413 1644 27422
rect 1592 27379 1601 27413
rect 1601 27379 1635 27413
rect 1635 27379 1644 27413
rect 1592 27370 1644 27379
rect 24172 27413 24224 27422
rect 24172 27379 24181 27413
rect 24181 27379 24215 27413
rect 24215 27379 24224 27413
rect 24172 27370 24224 27379
rect 1592 27077 1644 27086
rect 1592 27043 1601 27077
rect 1601 27043 1635 27077
rect 1635 27043 1644 27077
rect 1592 27034 1644 27043
rect 24172 27077 24224 27086
rect 24172 27043 24181 27077
rect 24181 27043 24215 27077
rect 24215 27043 24224 27077
rect 24172 27034 24224 27043
rect 1592 26741 1644 26750
rect 1592 26707 1601 26741
rect 1601 26707 1635 26741
rect 1635 26707 1644 26741
rect 1592 26698 1644 26707
rect 24172 26741 24224 26750
rect 24172 26707 24181 26741
rect 24181 26707 24215 26741
rect 24215 26707 24224 26741
rect 24172 26698 24224 26707
rect 1592 26405 1644 26414
rect 1592 26371 1601 26405
rect 1601 26371 1635 26405
rect 1635 26371 1644 26405
rect 1592 26362 1644 26371
rect 24172 26405 24224 26414
rect 24172 26371 24181 26405
rect 24181 26371 24215 26405
rect 24215 26371 24224 26405
rect 24172 26362 24224 26371
rect 1592 26069 1644 26078
rect 1592 26035 1601 26069
rect 1601 26035 1635 26069
rect 1635 26035 1644 26069
rect 1592 26026 1644 26035
rect 24172 26069 24224 26078
rect 24172 26035 24181 26069
rect 24181 26035 24215 26069
rect 24215 26035 24224 26069
rect 24172 26026 24224 26035
rect 1592 25733 1644 25742
rect 1592 25699 1601 25733
rect 1601 25699 1635 25733
rect 1635 25699 1644 25733
rect 1592 25690 1644 25699
rect 24172 25733 24224 25742
rect 24172 25699 24181 25733
rect 24181 25699 24215 25733
rect 24215 25699 24224 25733
rect 24172 25690 24224 25699
rect 1592 25397 1644 25406
rect 1592 25363 1601 25397
rect 1601 25363 1635 25397
rect 1635 25363 1644 25397
rect 1592 25354 1644 25363
rect 24172 25397 24224 25406
rect 24172 25363 24181 25397
rect 24181 25363 24215 25397
rect 24215 25363 24224 25397
rect 24172 25354 24224 25363
rect 1592 25061 1644 25070
rect 1592 25027 1601 25061
rect 1601 25027 1635 25061
rect 1635 25027 1644 25061
rect 1592 25018 1644 25027
rect 24172 25061 24224 25070
rect 24172 25027 24181 25061
rect 24181 25027 24215 25061
rect 24215 25027 24224 25061
rect 24172 25018 24224 25027
rect 1592 24725 1644 24734
rect 1592 24691 1601 24725
rect 1601 24691 1635 24725
rect 1635 24691 1644 24725
rect 1592 24682 1644 24691
rect 24172 24725 24224 24734
rect 24172 24691 24181 24725
rect 24181 24691 24215 24725
rect 24215 24691 24224 24725
rect 24172 24682 24224 24691
rect 1592 24389 1644 24398
rect 1592 24355 1601 24389
rect 1601 24355 1635 24389
rect 1635 24355 1644 24389
rect 1592 24346 1644 24355
rect 24172 24389 24224 24398
rect 24172 24355 24181 24389
rect 24181 24355 24215 24389
rect 24215 24355 24224 24389
rect 24172 24346 24224 24355
rect 1592 24053 1644 24062
rect 1592 24019 1601 24053
rect 1601 24019 1635 24053
rect 1635 24019 1644 24053
rect 1592 24010 1644 24019
rect 24172 24053 24224 24062
rect 24172 24019 24181 24053
rect 24181 24019 24215 24053
rect 24215 24019 24224 24053
rect 24172 24010 24224 24019
rect 1592 23717 1644 23726
rect 1592 23683 1601 23717
rect 1601 23683 1635 23717
rect 1635 23683 1644 23717
rect 1592 23674 1644 23683
rect 24172 23717 24224 23726
rect 24172 23683 24181 23717
rect 24181 23683 24215 23717
rect 24215 23683 24224 23717
rect 24172 23674 24224 23683
rect 1592 23381 1644 23390
rect 1592 23347 1601 23381
rect 1601 23347 1635 23381
rect 1635 23347 1644 23381
rect 1592 23338 1644 23347
rect 24172 23381 24224 23390
rect 24172 23347 24181 23381
rect 24181 23347 24215 23381
rect 24215 23347 24224 23381
rect 24172 23338 24224 23347
rect 1592 23045 1644 23054
rect 1592 23011 1601 23045
rect 1601 23011 1635 23045
rect 1635 23011 1644 23045
rect 1592 23002 1644 23011
rect 24172 23045 24224 23054
rect 24172 23011 24181 23045
rect 24181 23011 24215 23045
rect 24215 23011 24224 23045
rect 24172 23002 24224 23011
rect 1592 22709 1644 22718
rect 1592 22675 1601 22709
rect 1601 22675 1635 22709
rect 1635 22675 1644 22709
rect 1592 22666 1644 22675
rect 24172 22709 24224 22718
rect 24172 22675 24181 22709
rect 24181 22675 24215 22709
rect 24215 22675 24224 22709
rect 24172 22666 24224 22675
rect 1592 22373 1644 22382
rect 1592 22339 1601 22373
rect 1601 22339 1635 22373
rect 1635 22339 1644 22373
rect 1592 22330 1644 22339
rect 24172 22373 24224 22382
rect 24172 22339 24181 22373
rect 24181 22339 24215 22373
rect 24215 22339 24224 22373
rect 24172 22330 24224 22339
rect 1592 22037 1644 22046
rect 1592 22003 1601 22037
rect 1601 22003 1635 22037
rect 1635 22003 1644 22037
rect 1592 21994 1644 22003
rect 24172 22037 24224 22046
rect 24172 22003 24181 22037
rect 24181 22003 24215 22037
rect 24215 22003 24224 22037
rect 24172 21994 24224 22003
rect 1592 21701 1644 21710
rect 1592 21667 1601 21701
rect 1601 21667 1635 21701
rect 1635 21667 1644 21701
rect 1592 21658 1644 21667
rect 24172 21701 24224 21710
rect 24172 21667 24181 21701
rect 24181 21667 24215 21701
rect 24215 21667 24224 21701
rect 24172 21658 24224 21667
rect 1592 21365 1644 21374
rect 1592 21331 1601 21365
rect 1601 21331 1635 21365
rect 1635 21331 1644 21365
rect 1592 21322 1644 21331
rect 24172 21365 24224 21374
rect 24172 21331 24181 21365
rect 24181 21331 24215 21365
rect 24215 21331 24224 21365
rect 24172 21322 24224 21331
rect 1592 21029 1644 21038
rect 1592 20995 1601 21029
rect 1601 20995 1635 21029
rect 1635 20995 1644 21029
rect 1592 20986 1644 20995
rect 24172 21029 24224 21038
rect 24172 20995 24181 21029
rect 24181 20995 24215 21029
rect 24215 20995 24224 21029
rect 24172 20986 24224 20995
rect 1592 20693 1644 20702
rect 1592 20659 1601 20693
rect 1601 20659 1635 20693
rect 1635 20659 1644 20693
rect 1592 20650 1644 20659
rect 24172 20693 24224 20702
rect 24172 20659 24181 20693
rect 24181 20659 24215 20693
rect 24215 20659 24224 20693
rect 24172 20650 24224 20659
rect 1592 20357 1644 20366
rect 1592 20323 1601 20357
rect 1601 20323 1635 20357
rect 1635 20323 1644 20357
rect 1592 20314 1644 20323
rect 24172 20357 24224 20366
rect 24172 20323 24181 20357
rect 24181 20323 24215 20357
rect 24215 20323 24224 20357
rect 24172 20314 24224 20323
rect 1592 20021 1644 20030
rect 1592 19987 1601 20021
rect 1601 19987 1635 20021
rect 1635 19987 1644 20021
rect 1592 19978 1644 19987
rect 24172 20021 24224 20030
rect 24172 19987 24181 20021
rect 24181 19987 24215 20021
rect 24215 19987 24224 20021
rect 24172 19978 24224 19987
rect 1592 19685 1644 19694
rect 1592 19651 1601 19685
rect 1601 19651 1635 19685
rect 1635 19651 1644 19685
rect 1592 19642 1644 19651
rect 24172 19685 24224 19694
rect 24172 19651 24181 19685
rect 24181 19651 24215 19685
rect 24215 19651 24224 19685
rect 24172 19642 24224 19651
rect 1592 19349 1644 19358
rect 1592 19315 1601 19349
rect 1601 19315 1635 19349
rect 1635 19315 1644 19349
rect 1592 19306 1644 19315
rect 24172 19349 24224 19358
rect 24172 19315 24181 19349
rect 24181 19315 24215 19349
rect 24215 19315 24224 19349
rect 24172 19306 24224 19315
rect 1592 19013 1644 19022
rect 1592 18979 1601 19013
rect 1601 18979 1635 19013
rect 1635 18979 1644 19013
rect 1592 18970 1644 18979
rect 24172 19013 24224 19022
rect 24172 18979 24181 19013
rect 24181 18979 24215 19013
rect 24215 18979 24224 19013
rect 24172 18970 24224 18979
rect 1592 18677 1644 18686
rect 1592 18643 1601 18677
rect 1601 18643 1635 18677
rect 1635 18643 1644 18677
rect 1592 18634 1644 18643
rect 24172 18677 24224 18686
rect 24172 18643 24181 18677
rect 24181 18643 24215 18677
rect 24215 18643 24224 18677
rect 24172 18634 24224 18643
rect 1592 18341 1644 18350
rect 1592 18307 1601 18341
rect 1601 18307 1635 18341
rect 1635 18307 1644 18341
rect 1592 18298 1644 18307
rect 24172 18341 24224 18350
rect 24172 18307 24181 18341
rect 24181 18307 24215 18341
rect 24215 18307 24224 18341
rect 24172 18298 24224 18307
rect 1592 18005 1644 18014
rect 1592 17971 1601 18005
rect 1601 17971 1635 18005
rect 1635 17971 1644 18005
rect 1592 17962 1644 17971
rect 24172 18005 24224 18014
rect 24172 17971 24181 18005
rect 24181 17971 24215 18005
rect 24215 17971 24224 18005
rect 24172 17962 24224 17971
rect 1592 17669 1644 17678
rect 1592 17635 1601 17669
rect 1601 17635 1635 17669
rect 1635 17635 1644 17669
rect 1592 17626 1644 17635
rect 24172 17669 24224 17678
rect 24172 17635 24181 17669
rect 24181 17635 24215 17669
rect 24215 17635 24224 17669
rect 24172 17626 24224 17635
rect 1592 17333 1644 17342
rect 1592 17299 1601 17333
rect 1601 17299 1635 17333
rect 1635 17299 1644 17333
rect 1592 17290 1644 17299
rect 24172 17333 24224 17342
rect 24172 17299 24181 17333
rect 24181 17299 24215 17333
rect 24215 17299 24224 17333
rect 24172 17290 24224 17299
rect 1592 16997 1644 17006
rect 1592 16963 1601 16997
rect 1601 16963 1635 16997
rect 1635 16963 1644 16997
rect 1592 16954 1644 16963
rect 24172 16997 24224 17006
rect 24172 16963 24181 16997
rect 24181 16963 24215 16997
rect 24215 16963 24224 16997
rect 24172 16954 24224 16963
rect 1592 16661 1644 16670
rect 1592 16627 1601 16661
rect 1601 16627 1635 16661
rect 1635 16627 1644 16661
rect 1592 16618 1644 16627
rect 24172 16661 24224 16670
rect 24172 16627 24181 16661
rect 24181 16627 24215 16661
rect 24215 16627 24224 16661
rect 24172 16618 24224 16627
rect 1592 16325 1644 16334
rect 1592 16291 1601 16325
rect 1601 16291 1635 16325
rect 1635 16291 1644 16325
rect 1592 16282 1644 16291
rect 24172 16325 24224 16334
rect 24172 16291 24181 16325
rect 24181 16291 24215 16325
rect 24215 16291 24224 16325
rect 24172 16282 24224 16291
rect 1592 15989 1644 15998
rect 1592 15955 1601 15989
rect 1601 15955 1635 15989
rect 1635 15955 1644 15989
rect 1592 15946 1644 15955
rect 24172 15989 24224 15998
rect 24172 15955 24181 15989
rect 24181 15955 24215 15989
rect 24215 15955 24224 15989
rect 24172 15946 24224 15955
rect 1592 15653 1644 15662
rect 1592 15619 1601 15653
rect 1601 15619 1635 15653
rect 1635 15619 1644 15653
rect 1592 15610 1644 15619
rect 24172 15653 24224 15662
rect 24172 15619 24181 15653
rect 24181 15619 24215 15653
rect 24215 15619 24224 15653
rect 24172 15610 24224 15619
rect 1592 15317 1644 15326
rect 1592 15283 1601 15317
rect 1601 15283 1635 15317
rect 1635 15283 1644 15317
rect 1592 15274 1644 15283
rect 24172 15317 24224 15326
rect 24172 15283 24181 15317
rect 24181 15283 24215 15317
rect 24215 15283 24224 15317
rect 24172 15274 24224 15283
rect 1592 14981 1644 14990
rect 1592 14947 1601 14981
rect 1601 14947 1635 14981
rect 1635 14947 1644 14981
rect 1592 14938 1644 14947
rect 24172 14981 24224 14990
rect 24172 14947 24181 14981
rect 24181 14947 24215 14981
rect 24215 14947 24224 14981
rect 24172 14938 24224 14947
rect 1592 14645 1644 14654
rect 1592 14611 1601 14645
rect 1601 14611 1635 14645
rect 1635 14611 1644 14645
rect 1592 14602 1644 14611
rect 24172 14645 24224 14654
rect 24172 14611 24181 14645
rect 24181 14611 24215 14645
rect 24215 14611 24224 14645
rect 24172 14602 24224 14611
rect 1592 14309 1644 14318
rect 1592 14275 1601 14309
rect 1601 14275 1635 14309
rect 1635 14275 1644 14309
rect 1592 14266 1644 14275
rect 24172 14309 24224 14318
rect 24172 14275 24181 14309
rect 24181 14275 24215 14309
rect 24215 14275 24224 14309
rect 24172 14266 24224 14275
rect 1592 13973 1644 13982
rect 1592 13939 1601 13973
rect 1601 13939 1635 13973
rect 1635 13939 1644 13973
rect 1592 13930 1644 13939
rect 24172 13973 24224 13982
rect 24172 13939 24181 13973
rect 24181 13939 24215 13973
rect 24215 13939 24224 13973
rect 24172 13930 24224 13939
rect 1592 13637 1644 13646
rect 1592 13603 1601 13637
rect 1601 13603 1635 13637
rect 1635 13603 1644 13637
rect 1592 13594 1644 13603
rect 24172 13637 24224 13646
rect 24172 13603 24181 13637
rect 24181 13603 24215 13637
rect 24215 13603 24224 13637
rect 24172 13594 24224 13603
rect 1592 13301 1644 13310
rect 1592 13267 1601 13301
rect 1601 13267 1635 13301
rect 1635 13267 1644 13301
rect 1592 13258 1644 13267
rect 24172 13301 24224 13310
rect 24172 13267 24181 13301
rect 24181 13267 24215 13301
rect 24215 13267 24224 13301
rect 24172 13258 24224 13267
rect 1592 12965 1644 12974
rect 1592 12931 1601 12965
rect 1601 12931 1635 12965
rect 1635 12931 1644 12965
rect 1592 12922 1644 12931
rect 24172 12965 24224 12974
rect 24172 12931 24181 12965
rect 24181 12931 24215 12965
rect 24215 12931 24224 12965
rect 24172 12922 24224 12931
rect 1592 12629 1644 12638
rect 1592 12595 1601 12629
rect 1601 12595 1635 12629
rect 1635 12595 1644 12629
rect 1592 12586 1644 12595
rect 24172 12629 24224 12638
rect 24172 12595 24181 12629
rect 24181 12595 24215 12629
rect 24215 12595 24224 12629
rect 24172 12586 24224 12595
rect 1592 12293 1644 12302
rect 1592 12259 1601 12293
rect 1601 12259 1635 12293
rect 1635 12259 1644 12293
rect 1592 12250 1644 12259
rect 24172 12293 24224 12302
rect 24172 12259 24181 12293
rect 24181 12259 24215 12293
rect 24215 12259 24224 12293
rect 24172 12250 24224 12259
rect 1592 11957 1644 11966
rect 1592 11923 1601 11957
rect 1601 11923 1635 11957
rect 1635 11923 1644 11957
rect 1592 11914 1644 11923
rect 24172 11957 24224 11966
rect 24172 11923 24181 11957
rect 24181 11923 24215 11957
rect 24215 11923 24224 11957
rect 24172 11914 24224 11923
rect 1592 11621 1644 11630
rect 1592 11587 1601 11621
rect 1601 11587 1635 11621
rect 1635 11587 1644 11621
rect 1592 11578 1644 11587
rect 24172 11621 24224 11630
rect 24172 11587 24181 11621
rect 24181 11587 24215 11621
rect 24215 11587 24224 11621
rect 24172 11578 24224 11587
rect 1592 11285 1644 11294
rect 1592 11251 1601 11285
rect 1601 11251 1635 11285
rect 1635 11251 1644 11285
rect 1592 11242 1644 11251
rect 24172 11285 24224 11294
rect 24172 11251 24181 11285
rect 24181 11251 24215 11285
rect 24215 11251 24224 11285
rect 24172 11242 24224 11251
rect 1592 10949 1644 10958
rect 1592 10915 1601 10949
rect 1601 10915 1635 10949
rect 1635 10915 1644 10949
rect 1592 10906 1644 10915
rect 24172 10949 24224 10958
rect 24172 10915 24181 10949
rect 24181 10915 24215 10949
rect 24215 10915 24224 10949
rect 24172 10906 24224 10915
rect 1592 10613 1644 10622
rect 1592 10579 1601 10613
rect 1601 10579 1635 10613
rect 1635 10579 1644 10613
rect 1592 10570 1644 10579
rect 24172 10613 24224 10622
rect 24172 10579 24181 10613
rect 24181 10579 24215 10613
rect 24215 10579 24224 10613
rect 24172 10570 24224 10579
rect 1592 10277 1644 10286
rect 1592 10243 1601 10277
rect 1601 10243 1635 10277
rect 1635 10243 1644 10277
rect 1592 10234 1644 10243
rect 24172 10277 24224 10286
rect 24172 10243 24181 10277
rect 24181 10243 24215 10277
rect 24215 10243 24224 10277
rect 24172 10234 24224 10243
rect 1592 9941 1644 9950
rect 1592 9907 1601 9941
rect 1601 9907 1635 9941
rect 1635 9907 1644 9941
rect 1592 9898 1644 9907
rect 24172 9941 24224 9950
rect 24172 9907 24181 9941
rect 24181 9907 24215 9941
rect 24215 9907 24224 9941
rect 24172 9898 24224 9907
rect 1592 9605 1644 9614
rect 1592 9571 1601 9605
rect 1601 9571 1635 9605
rect 1635 9571 1644 9605
rect 1592 9562 1644 9571
rect 24172 9605 24224 9614
rect 24172 9571 24181 9605
rect 24181 9571 24215 9605
rect 24215 9571 24224 9605
rect 24172 9562 24224 9571
rect 1592 9269 1644 9278
rect 1592 9235 1601 9269
rect 1601 9235 1635 9269
rect 1635 9235 1644 9269
rect 1592 9226 1644 9235
rect 24172 9269 24224 9278
rect 24172 9235 24181 9269
rect 24181 9235 24215 9269
rect 24215 9235 24224 9269
rect 24172 9226 24224 9235
rect 1592 8933 1644 8942
rect 1592 8899 1601 8933
rect 1601 8899 1635 8933
rect 1635 8899 1644 8933
rect 1592 8890 1644 8899
rect 24172 8933 24224 8942
rect 24172 8899 24181 8933
rect 24181 8899 24215 8933
rect 24215 8899 24224 8933
rect 24172 8890 24224 8899
rect 1592 8597 1644 8606
rect 1592 8563 1601 8597
rect 1601 8563 1635 8597
rect 1635 8563 1644 8597
rect 1592 8554 1644 8563
rect 24172 8597 24224 8606
rect 24172 8563 24181 8597
rect 24181 8563 24215 8597
rect 24215 8563 24224 8597
rect 24172 8554 24224 8563
rect 1592 8261 1644 8270
rect 1592 8227 1601 8261
rect 1601 8227 1635 8261
rect 1635 8227 1644 8261
rect 1592 8218 1644 8227
rect 24172 8261 24224 8270
rect 24172 8227 24181 8261
rect 24181 8227 24215 8261
rect 24215 8227 24224 8261
rect 24172 8218 24224 8227
rect 1592 7925 1644 7934
rect 1592 7891 1601 7925
rect 1601 7891 1635 7925
rect 1635 7891 1644 7925
rect 1592 7882 1644 7891
rect 24172 7925 24224 7934
rect 24172 7891 24181 7925
rect 24181 7891 24215 7925
rect 24215 7891 24224 7925
rect 24172 7882 24224 7891
rect 1592 7589 1644 7598
rect 1592 7555 1601 7589
rect 1601 7555 1635 7589
rect 1635 7555 1644 7589
rect 1592 7546 1644 7555
rect 24172 7589 24224 7598
rect 24172 7555 24181 7589
rect 24181 7555 24215 7589
rect 24215 7555 24224 7589
rect 24172 7546 24224 7555
rect 1592 7253 1644 7262
rect 1592 7219 1601 7253
rect 1601 7219 1635 7253
rect 1635 7219 1644 7253
rect 1592 7210 1644 7219
rect 24172 7253 24224 7262
rect 24172 7219 24181 7253
rect 24181 7219 24215 7253
rect 24215 7219 24224 7253
rect 24172 7210 24224 7219
rect 1592 6917 1644 6926
rect 1592 6883 1601 6917
rect 1601 6883 1635 6917
rect 1635 6883 1644 6917
rect 1592 6874 1644 6883
rect 24172 6917 24224 6926
rect 24172 6883 24181 6917
rect 24181 6883 24215 6917
rect 24215 6883 24224 6917
rect 24172 6874 24224 6883
rect 1592 6581 1644 6590
rect 1592 6547 1601 6581
rect 1601 6547 1635 6581
rect 1635 6547 1644 6581
rect 1592 6538 1644 6547
rect 24172 6581 24224 6590
rect 24172 6547 24181 6581
rect 24181 6547 24215 6581
rect 24215 6547 24224 6581
rect 24172 6538 24224 6547
rect 1592 6245 1644 6254
rect 1592 6211 1601 6245
rect 1601 6211 1635 6245
rect 1635 6211 1644 6245
rect 1592 6202 1644 6211
rect 24172 6245 24224 6254
rect 24172 6211 24181 6245
rect 24181 6211 24215 6245
rect 24215 6211 24224 6245
rect 24172 6202 24224 6211
rect 1592 5909 1644 5918
rect 1592 5875 1601 5909
rect 1601 5875 1635 5909
rect 1635 5875 1644 5909
rect 1592 5866 1644 5875
rect 24172 5909 24224 5918
rect 24172 5875 24181 5909
rect 24181 5875 24215 5909
rect 24215 5875 24224 5909
rect 24172 5866 24224 5875
rect 1592 5573 1644 5582
rect 1592 5539 1601 5573
rect 1601 5539 1635 5573
rect 1635 5539 1644 5573
rect 1592 5530 1644 5539
rect 24172 5573 24224 5582
rect 24172 5539 24181 5573
rect 24181 5539 24215 5573
rect 24215 5539 24224 5573
rect 24172 5530 24224 5539
rect 1592 5237 1644 5246
rect 1592 5203 1601 5237
rect 1601 5203 1635 5237
rect 1635 5203 1644 5237
rect 1592 5194 1644 5203
rect 24172 5237 24224 5246
rect 24172 5203 24181 5237
rect 24181 5203 24215 5237
rect 24215 5203 24224 5237
rect 24172 5194 24224 5203
rect 1592 4901 1644 4910
rect 1592 4867 1601 4901
rect 1601 4867 1635 4901
rect 1635 4867 1644 4901
rect 1592 4858 1644 4867
rect 24172 4901 24224 4910
rect 24172 4867 24181 4901
rect 24181 4867 24215 4901
rect 24215 4867 24224 4901
rect 24172 4858 24224 4867
rect 1592 4565 1644 4574
rect 1592 4531 1601 4565
rect 1601 4531 1635 4565
rect 1635 4531 1644 4565
rect 1592 4522 1644 4531
rect 24172 4565 24224 4574
rect 24172 4531 24181 4565
rect 24181 4531 24215 4565
rect 24215 4531 24224 4565
rect 24172 4522 24224 4531
rect 1592 4229 1644 4238
rect 1592 4195 1601 4229
rect 1601 4195 1635 4229
rect 1635 4195 1644 4229
rect 1592 4186 1644 4195
rect 24172 4229 24224 4238
rect 24172 4195 24181 4229
rect 24181 4195 24215 4229
rect 24215 4195 24224 4229
rect 24172 4186 24224 4195
rect 1592 3893 1644 3902
rect 1592 3859 1601 3893
rect 1601 3859 1635 3893
rect 1635 3859 1644 3893
rect 1592 3850 1644 3859
rect 24172 3893 24224 3902
rect 24172 3859 24181 3893
rect 24181 3859 24215 3893
rect 24215 3859 24224 3893
rect 24172 3850 24224 3859
rect 1592 3557 1644 3566
rect 1592 3523 1601 3557
rect 1601 3523 1635 3557
rect 1635 3523 1644 3557
rect 1592 3514 1644 3523
rect 24172 3557 24224 3566
rect 24172 3523 24181 3557
rect 24181 3523 24215 3557
rect 24215 3523 24224 3557
rect 24172 3514 24224 3523
rect 1592 3221 1644 3230
rect 1592 3187 1601 3221
rect 1601 3187 1635 3221
rect 1635 3187 1644 3221
rect 1592 3178 1644 3187
rect 24172 3221 24224 3230
rect 24172 3187 24181 3221
rect 24181 3187 24215 3221
rect 24215 3187 24224 3221
rect 24172 3178 24224 3187
rect 1592 2885 1644 2894
rect 1592 2851 1601 2885
rect 1601 2851 1635 2885
rect 1635 2851 1644 2885
rect 1592 2842 1644 2851
rect 24172 2885 24224 2894
rect 24172 2851 24181 2885
rect 24181 2851 24215 2885
rect 24215 2851 24224 2885
rect 24172 2842 24224 2851
rect 1592 2549 1644 2558
rect 1592 2515 1601 2549
rect 1601 2515 1635 2549
rect 1635 2515 1644 2549
rect 1592 2506 1644 2515
rect 24172 2549 24224 2558
rect 24172 2515 24181 2549
rect 24181 2515 24215 2549
rect 24215 2515 24224 2549
rect 24172 2506 24224 2515
rect 1592 2213 1644 2222
rect 1592 2179 1601 2213
rect 1601 2179 1635 2213
rect 1635 2179 1644 2213
rect 1592 2170 1644 2179
rect 24172 2213 24224 2222
rect 24172 2179 24181 2213
rect 24181 2179 24215 2213
rect 24215 2179 24224 2213
rect 24172 2170 24224 2179
rect 1592 1877 1644 1886
rect 1592 1843 1601 1877
rect 1601 1843 1635 1877
rect 1635 1843 1644 1877
rect 1592 1834 1644 1843
rect 24172 1877 24224 1886
rect 24172 1843 24181 1877
rect 24181 1843 24215 1877
rect 24215 1843 24224 1877
rect 24172 1834 24224 1843
rect 1928 1541 1980 1550
rect 3608 1541 3660 1550
rect 5288 1541 5340 1550
rect 6968 1541 7020 1550
rect 8648 1541 8700 1550
rect 10328 1541 10380 1550
rect 12008 1541 12060 1550
rect 13688 1541 13740 1550
rect 15368 1541 15420 1550
rect 17048 1541 17100 1550
rect 18728 1541 18780 1550
rect 20408 1541 20460 1550
rect 22088 1541 22140 1550
rect 23768 1541 23820 1550
rect 1928 1507 1937 1541
rect 1937 1507 1971 1541
rect 1971 1507 1980 1541
rect 3608 1507 3617 1541
rect 3617 1507 3651 1541
rect 3651 1507 3660 1541
rect 5288 1507 5297 1541
rect 5297 1507 5331 1541
rect 5331 1507 5340 1541
rect 6968 1507 6977 1541
rect 6977 1507 7011 1541
rect 7011 1507 7020 1541
rect 8648 1507 8657 1541
rect 8657 1507 8691 1541
rect 8691 1507 8700 1541
rect 10328 1507 10337 1541
rect 10337 1507 10371 1541
rect 10371 1507 10380 1541
rect 12008 1507 12017 1541
rect 12017 1507 12051 1541
rect 12051 1507 12060 1541
rect 13688 1507 13697 1541
rect 13697 1507 13731 1541
rect 13731 1507 13740 1541
rect 15368 1507 15377 1541
rect 15377 1507 15411 1541
rect 15411 1507 15420 1541
rect 17048 1507 17057 1541
rect 17057 1507 17091 1541
rect 17091 1507 17100 1541
rect 18728 1507 18737 1541
rect 18737 1507 18771 1541
rect 18771 1507 18780 1541
rect 20408 1507 20417 1541
rect 20417 1507 20451 1541
rect 20451 1507 20460 1541
rect 22088 1507 22097 1541
rect 22097 1507 22131 1541
rect 22131 1507 22140 1541
rect 23768 1507 23777 1541
rect 23777 1507 23811 1541
rect 23811 1507 23820 1541
rect 1928 1498 1980 1507
rect 3608 1498 3660 1507
rect 5288 1498 5340 1507
rect 6968 1498 7020 1507
rect 8648 1498 8700 1507
rect 10328 1498 10380 1507
rect 12008 1498 12060 1507
rect 13688 1498 13740 1507
rect 15368 1498 15420 1507
rect 17048 1498 17100 1507
rect 18728 1498 18780 1507
rect 20408 1498 20460 1507
rect 22088 1498 22140 1507
rect 23768 1498 23820 1507
<< metal2 >>
rect 1506 33470 1730 34046
rect 1506 33418 1592 33470
rect 1644 33418 1730 33470
rect 1506 33134 1730 33418
rect 1506 33082 1592 33134
rect 1644 33082 1730 33134
rect 1506 32798 1730 33082
rect 24086 33470 24310 34046
rect 24086 33418 24172 33470
rect 24224 33418 24310 33470
rect 24086 33134 24310 33418
rect 24086 33082 24172 33134
rect 24224 33082 24310 33134
rect 1506 32746 1592 32798
rect 1644 32746 1730 32798
rect 1506 32462 1730 32746
rect 1506 32410 1592 32462
rect 1644 32410 1730 32462
rect 1506 32128 1730 32410
rect 1506 32072 1590 32128
rect 1646 32072 1730 32128
rect 1506 31790 1730 32072
rect 1506 31738 1592 31790
rect 1644 31738 1730 31790
rect 1506 31454 1730 31738
rect 1506 31402 1592 31454
rect 1644 31402 1730 31454
rect 1506 31118 1730 31402
rect 1506 31066 1592 31118
rect 1644 31066 1730 31118
rect 1506 30782 1730 31066
rect 1506 30730 1592 30782
rect 1644 30730 1730 30782
rect 1506 30448 1730 30730
rect 1506 30392 1590 30448
rect 1646 30392 1730 30448
rect 1506 30110 1730 30392
rect 1506 30058 1592 30110
rect 1644 30058 1730 30110
rect 1506 29774 1730 30058
rect 1506 29722 1592 29774
rect 1644 29722 1730 29774
rect 1506 29438 1730 29722
rect 1506 29386 1592 29438
rect 1644 29386 1730 29438
rect 1506 29102 1730 29386
rect 1506 29050 1592 29102
rect 1644 29050 1730 29102
rect 1506 28768 1730 29050
rect 1506 28712 1590 28768
rect 1646 28712 1730 28768
rect 1506 28430 1730 28712
rect 1506 28378 1592 28430
rect 1644 28378 1730 28430
rect 1506 28094 1730 28378
rect 1506 28042 1592 28094
rect 1644 28042 1730 28094
rect 1506 27758 1730 28042
rect 1506 27706 1592 27758
rect 1644 27706 1730 27758
rect 1506 27422 1730 27706
rect 1506 27370 1592 27422
rect 1644 27370 1730 27422
rect 1506 27088 1730 27370
rect 1506 27032 1590 27088
rect 1646 27032 1730 27088
rect 1506 26750 1730 27032
rect 1506 26698 1592 26750
rect 1644 26698 1730 26750
rect 1506 26414 1730 26698
rect 1506 26362 1592 26414
rect 1644 26362 1730 26414
rect 1506 26078 1730 26362
rect 1506 26026 1592 26078
rect 1644 26026 1730 26078
rect 1506 25742 1730 26026
rect 1506 25690 1592 25742
rect 1644 25690 1730 25742
rect 1506 25408 1730 25690
rect 1506 25352 1590 25408
rect 1646 25352 1730 25408
rect 1506 25070 1730 25352
rect 1506 25018 1592 25070
rect 1644 25018 1730 25070
rect 1506 24734 1730 25018
rect 1506 24682 1592 24734
rect 1644 24682 1730 24734
rect 1506 24398 1730 24682
rect 1506 24346 1592 24398
rect 1644 24346 1730 24398
rect 1506 24062 1730 24346
rect 1506 24010 1592 24062
rect 1644 24010 1730 24062
rect 1506 23728 1730 24010
rect 1506 23672 1590 23728
rect 1646 23672 1730 23728
rect 1506 23390 1730 23672
rect 1506 23338 1592 23390
rect 1644 23338 1730 23390
rect 1506 23054 1730 23338
rect 1506 23002 1592 23054
rect 1644 23002 1730 23054
rect 1506 22718 1730 23002
rect 1506 22666 1592 22718
rect 1644 22666 1730 22718
rect 1506 22382 1730 22666
rect 1506 22330 1592 22382
rect 1644 22330 1730 22382
rect 1506 22048 1730 22330
rect 1506 21992 1590 22048
rect 1646 21992 1730 22048
rect 1506 21710 1730 21992
rect 1506 21658 1592 21710
rect 1644 21658 1730 21710
rect 1506 21374 1730 21658
rect 1506 21322 1592 21374
rect 1644 21322 1730 21374
rect 1506 21038 1730 21322
rect 1506 20986 1592 21038
rect 1644 20986 1730 21038
rect 1506 20702 1730 20986
rect 1506 20650 1592 20702
rect 1644 20650 1730 20702
rect 1506 20368 1730 20650
rect 1506 20312 1590 20368
rect 1646 20312 1730 20368
rect 1506 20030 1730 20312
rect 1506 19978 1592 20030
rect 1644 19978 1730 20030
rect 1506 19694 1730 19978
rect 1506 19642 1592 19694
rect 1644 19642 1730 19694
rect 1506 19358 1730 19642
rect 1506 19306 1592 19358
rect 1644 19306 1730 19358
rect 1506 19022 1730 19306
rect 1506 18970 1592 19022
rect 1644 18970 1730 19022
rect 1506 18688 1730 18970
rect 1506 18632 1590 18688
rect 1646 18632 1730 18688
rect 1506 18350 1730 18632
rect 1506 18298 1592 18350
rect 1644 18298 1730 18350
rect 1506 18014 1730 18298
rect 1506 17962 1592 18014
rect 1644 17962 1730 18014
rect 1506 17678 1730 17962
rect 1506 17626 1592 17678
rect 1644 17626 1730 17678
rect 1506 17342 1730 17626
rect 1506 17290 1592 17342
rect 1644 17290 1730 17342
rect 1506 17008 1730 17290
rect 1506 16952 1590 17008
rect 1646 16952 1730 17008
rect 1506 16670 1730 16952
rect 1506 16618 1592 16670
rect 1644 16618 1730 16670
rect 1506 16334 1730 16618
rect 1506 16282 1592 16334
rect 1644 16282 1730 16334
rect 1506 15998 1730 16282
rect 1506 15946 1592 15998
rect 1644 15946 1730 15998
rect 1506 15662 1730 15946
rect 1506 15610 1592 15662
rect 1644 15610 1730 15662
rect 1506 15328 1730 15610
rect 1506 15272 1590 15328
rect 1646 15272 1730 15328
rect 1506 14990 1730 15272
rect 1506 14938 1592 14990
rect 1644 14938 1730 14990
rect 1506 14654 1730 14938
rect 1506 14602 1592 14654
rect 1644 14602 1730 14654
rect 1506 14318 1730 14602
rect 1506 14266 1592 14318
rect 1644 14266 1730 14318
rect 1506 13982 1730 14266
rect 1506 13930 1592 13982
rect 1644 13930 1730 13982
rect 1506 13648 1730 13930
rect 1506 13592 1590 13648
rect 1646 13592 1730 13648
rect 1506 13310 1730 13592
rect 1506 13258 1592 13310
rect 1644 13258 1730 13310
rect 1506 12974 1730 13258
rect 1506 12922 1592 12974
rect 1644 12922 1730 12974
rect 1506 12638 1730 12922
rect 1506 12586 1592 12638
rect 1644 12586 1730 12638
rect 1506 12302 1730 12586
rect 1506 12250 1592 12302
rect 1644 12250 1730 12302
rect 1506 11968 1730 12250
rect 1506 11912 1590 11968
rect 1646 11912 1730 11968
rect 1506 11630 1730 11912
rect 1506 11578 1592 11630
rect 1644 11578 1730 11630
rect 1506 11294 1730 11578
rect 1506 11242 1592 11294
rect 1644 11242 1730 11294
rect 1506 10958 1730 11242
rect 1506 10906 1592 10958
rect 1644 10906 1730 10958
rect 1506 10622 1730 10906
rect 1506 10570 1592 10622
rect 1644 10570 1730 10622
rect 1506 10288 1730 10570
rect 1506 10232 1590 10288
rect 1646 10232 1730 10288
rect 1506 9950 1730 10232
rect 1506 9898 1592 9950
rect 1644 9898 1730 9950
rect 1506 9614 1730 9898
rect 1506 9562 1592 9614
rect 1644 9562 1730 9614
rect 1506 9278 1730 9562
rect 1506 9226 1592 9278
rect 1644 9226 1730 9278
rect 1506 8942 1730 9226
rect 1506 8890 1592 8942
rect 1644 8890 1730 8942
rect 1506 8608 1730 8890
rect 1506 8552 1590 8608
rect 1646 8552 1730 8608
rect 1506 8270 1730 8552
rect 1506 8218 1592 8270
rect 1644 8218 1730 8270
rect 1506 7934 1730 8218
rect 1506 7882 1592 7934
rect 1644 7882 1730 7934
rect 1506 7598 1730 7882
rect 1506 7546 1592 7598
rect 1644 7546 1730 7598
rect 1506 7262 1730 7546
rect 1506 7210 1592 7262
rect 1644 7210 1730 7262
rect 1506 6928 1730 7210
rect 1506 6872 1590 6928
rect 1646 6872 1730 6928
rect 1506 6590 1730 6872
rect 1506 6538 1592 6590
rect 1644 6538 1730 6590
rect 1506 6254 1730 6538
rect 1506 6202 1592 6254
rect 1644 6202 1730 6254
rect 1506 5918 1730 6202
rect 1506 5866 1592 5918
rect 1644 5866 1730 5918
rect 1506 5582 1730 5866
rect 1506 5530 1592 5582
rect 1644 5530 1730 5582
rect 1506 5248 1730 5530
rect 1506 5192 1590 5248
rect 1646 5192 1730 5248
rect 1506 4910 1730 5192
rect 1506 4858 1592 4910
rect 1644 4858 1730 4910
rect 1506 4574 1730 4858
rect 1506 4522 1592 4574
rect 1644 4522 1730 4574
rect 1506 4238 1730 4522
rect 1506 4186 1592 4238
rect 1644 4186 1730 4238
rect 1506 3902 1730 4186
rect 1506 3850 1592 3902
rect 1644 3850 1730 3902
rect 1506 3568 1730 3850
rect 1506 3512 1590 3568
rect 1646 3512 1730 3568
rect 8002 3587 8030 8790
rect 9768 8788 9796 20666
rect 9852 9980 9880 20666
rect 9936 10464 9964 20666
rect 10020 11656 10048 20666
rect 10104 12140 10132 20666
rect 10188 13332 10216 20666
rect 14944 7881 14972 32958
rect 24086 32798 24310 33082
rect 24086 32746 24172 32798
rect 24224 32746 24310 32798
rect 24086 32462 24310 32746
rect 24086 32410 24172 32462
rect 24224 32410 24310 32462
rect 24086 32128 24310 32410
rect 24086 32072 24170 32128
rect 24226 32072 24310 32128
rect 24086 31790 24310 32072
rect 24086 31738 24172 31790
rect 24224 31738 24310 31790
rect 24086 31454 24310 31738
rect 24086 31402 24172 31454
rect 24224 31402 24310 31454
rect 24086 31118 24310 31402
rect 24086 31066 24172 31118
rect 24224 31066 24310 31118
rect 24086 30782 24310 31066
rect 24086 30730 24172 30782
rect 24224 30730 24310 30782
rect 24086 30448 24310 30730
rect 24086 30392 24170 30448
rect 24226 30392 24310 30448
rect 24086 30110 24310 30392
rect 24086 30058 24172 30110
rect 24224 30058 24310 30110
rect 24086 29774 24310 30058
rect 24086 29722 24172 29774
rect 24224 29722 24310 29774
rect 24086 29438 24310 29722
rect 24086 29386 24172 29438
rect 24224 29386 24310 29438
rect 24086 29102 24310 29386
rect 24086 29050 24172 29102
rect 24224 29050 24310 29102
rect 24086 28768 24310 29050
rect 24086 28712 24170 28768
rect 24226 28712 24310 28768
rect 24086 28430 24310 28712
rect 24086 28378 24172 28430
rect 24224 28378 24310 28430
rect 24086 28094 24310 28378
rect 24086 28042 24172 28094
rect 24224 28042 24310 28094
rect 24086 27758 24310 28042
rect 24086 27706 24172 27758
rect 24224 27706 24310 27758
rect 24086 27422 24310 27706
rect 24086 27370 24172 27422
rect 24224 27370 24310 27422
rect 24086 27088 24310 27370
rect 24086 27032 24170 27088
rect 24226 27032 24310 27088
rect 24086 26750 24310 27032
rect 24086 26698 24172 26750
rect 24224 26698 24310 26750
rect 24086 26414 24310 26698
rect 24086 26362 24172 26414
rect 24224 26362 24310 26414
rect 24086 26078 24310 26362
rect 24086 26026 24172 26078
rect 24224 26026 24310 26078
rect 24086 25742 24310 26026
rect 24086 25690 24172 25742
rect 24224 25690 24310 25742
rect 24086 25408 24310 25690
rect 24086 25352 24170 25408
rect 24226 25352 24310 25408
rect 24086 25070 24310 25352
rect 24086 25018 24172 25070
rect 24224 25018 24310 25070
rect 24086 24734 24310 25018
rect 24086 24682 24172 24734
rect 24224 24682 24310 24734
rect 24086 24398 24310 24682
rect 24086 24346 24172 24398
rect 24224 24346 24310 24398
rect 24086 24062 24310 24346
rect 24086 24010 24172 24062
rect 24224 24010 24310 24062
rect 24086 23728 24310 24010
rect 24086 23672 24170 23728
rect 24226 23672 24310 23728
rect 24086 23390 24310 23672
rect 24086 23338 24172 23390
rect 24224 23338 24310 23390
rect 24086 23054 24310 23338
rect 24086 23002 24172 23054
rect 24224 23002 24310 23054
rect 24086 22718 24310 23002
rect 24086 22666 24172 22718
rect 24224 22666 24310 22718
rect 24086 22382 24310 22666
rect 24086 22330 24172 22382
rect 24224 22330 24310 22382
rect 24086 22048 24310 22330
rect 24086 21992 24170 22048
rect 24226 21992 24310 22048
rect 24086 21710 24310 21992
rect 24086 21658 24172 21710
rect 24224 21658 24310 21710
rect 24086 21374 24310 21658
rect 24086 21322 24172 21374
rect 24224 21322 24310 21374
rect 24086 21038 24310 21322
rect 24086 20986 24172 21038
rect 24224 20986 24310 21038
rect 24086 20702 24310 20986
rect 24086 20650 24172 20702
rect 24224 20650 24310 20702
rect 24086 20368 24310 20650
rect 24086 20312 24170 20368
rect 24226 20312 24310 20368
rect 24086 20030 24310 20312
rect 24086 19978 24172 20030
rect 24224 19978 24310 20030
rect 24086 19694 24310 19978
rect 24086 19642 24172 19694
rect 24224 19642 24310 19694
rect 24086 19358 24310 19642
rect 24086 19306 24172 19358
rect 24224 19306 24310 19358
rect 24086 19022 24310 19306
rect 24086 18970 24172 19022
rect 24224 18970 24310 19022
rect 24086 18688 24310 18970
rect 24086 18632 24170 18688
rect 24226 18632 24310 18688
rect 24086 18350 24310 18632
rect 24086 18298 24172 18350
rect 24224 18298 24310 18350
rect 24086 18014 24310 18298
rect 24086 17962 24172 18014
rect 24224 17962 24310 18014
rect 24086 17678 24310 17962
rect 24086 17626 24172 17678
rect 24224 17626 24310 17678
rect 24086 17342 24310 17626
rect 24086 17290 24172 17342
rect 24224 17290 24310 17342
rect 24086 17008 24310 17290
rect 24086 16952 24170 17008
rect 24226 16952 24310 17008
rect 24086 16670 24310 16952
rect 24086 16618 24172 16670
rect 24224 16618 24310 16670
rect 24086 16334 24310 16618
rect 24086 16282 24172 16334
rect 24224 16282 24310 16334
rect 24086 15998 24310 16282
rect 24086 15946 24172 15998
rect 24224 15946 24310 15998
rect 24086 15662 24310 15946
rect 24086 15610 24172 15662
rect 24224 15610 24310 15662
rect 24086 15328 24310 15610
rect 24086 15272 24170 15328
rect 24226 15272 24310 15328
rect 24086 14990 24310 15272
rect 24086 14938 24172 14990
rect 24224 14938 24310 14990
rect 24086 14654 24310 14938
rect 24086 14602 24172 14654
rect 24224 14602 24310 14654
rect 24086 14318 24310 14602
rect 24086 14266 24172 14318
rect 24224 14266 24310 14318
rect 24086 13982 24310 14266
rect 24086 13930 24172 13982
rect 24224 13930 24310 13982
rect 24086 13648 24310 13930
rect 24086 13592 24170 13648
rect 24226 13592 24310 13648
rect 24086 13310 24310 13592
rect 24086 13258 24172 13310
rect 24224 13258 24310 13310
rect 24086 12974 24310 13258
rect 24086 12922 24172 12974
rect 24224 12922 24310 12974
rect 24086 12638 24310 12922
rect 24086 12586 24172 12638
rect 24224 12586 24310 12638
rect 24086 12302 24310 12586
rect 24086 12250 24172 12302
rect 24224 12250 24310 12302
rect 24086 11968 24310 12250
rect 24086 11912 24170 11968
rect 24226 11912 24310 11968
rect 24086 11630 24310 11912
rect 24086 11578 24172 11630
rect 24224 11578 24310 11630
rect 24086 11294 24310 11578
rect 24086 11242 24172 11294
rect 24224 11242 24310 11294
rect 24086 10958 24310 11242
rect 24086 10906 24172 10958
rect 24224 10906 24310 10958
rect 24086 10622 24310 10906
rect 24086 10570 24172 10622
rect 24224 10570 24310 10622
rect 24086 10288 24310 10570
rect 24086 10232 24170 10288
rect 24226 10232 24310 10288
rect 24086 9950 24310 10232
rect 24086 9898 24172 9950
rect 24224 9898 24310 9950
rect 24086 9614 24310 9898
rect 24086 9562 24172 9614
rect 24224 9562 24310 9614
rect 24086 9278 24310 9562
rect 24086 9226 24172 9278
rect 24224 9226 24310 9278
rect 24086 8942 24310 9226
rect 24086 8890 24172 8942
rect 24224 8890 24310 8942
rect 24086 8608 24310 8890
rect 24086 8552 24170 8608
rect 24226 8552 24310 8608
rect 24086 8270 24310 8552
rect 24086 8218 24172 8270
rect 24224 8218 24310 8270
rect 24086 7934 24310 8218
rect 24086 7882 24172 7934
rect 24224 7882 24310 7934
rect 24086 7598 24310 7882
rect 24086 7546 24172 7598
rect 24224 7546 24310 7598
rect 24086 7262 24310 7546
rect 24086 7210 24172 7262
rect 24224 7210 24310 7262
rect 24086 6928 24310 7210
rect 16078 4456 16106 6153
rect 18294 4456 18322 6903
rect 24086 6872 24170 6928
rect 24226 6872 24310 6928
rect 24086 6590 24310 6872
rect 24086 6538 24172 6590
rect 24224 6538 24310 6590
rect 24086 6254 24310 6538
rect 24086 6202 24172 6254
rect 24224 6202 24310 6254
rect 24086 5918 24310 6202
rect 24086 5866 24172 5918
rect 24224 5866 24310 5918
rect 24086 5582 24310 5866
rect 24086 5530 24172 5582
rect 24224 5530 24310 5582
rect 24086 5248 24310 5530
rect 24086 5192 24170 5248
rect 24226 5192 24310 5248
rect 24086 4910 24310 5192
rect 24086 4858 24172 4910
rect 24224 4858 24310 4910
rect 24086 4574 24310 4858
rect 24086 4522 24172 4574
rect 24224 4522 24310 4574
rect 24086 4238 24310 4522
rect 24086 4186 24172 4238
rect 24224 4186 24310 4238
rect 24086 3902 24310 4186
rect 24086 3850 24172 3902
rect 24224 3850 24310 3902
rect 8002 3573 8596 3587
rect 7986 3559 8596 3573
rect 24086 3568 24310 3850
rect 1506 3230 1730 3512
rect 1506 3178 1592 3230
rect 1644 3178 1730 3230
rect 1506 2894 1730 3178
rect 1506 2842 1592 2894
rect 1644 2842 1730 2894
rect 1506 2558 1730 2842
rect 7986 2692 8046 3559
rect 7986 2664 7988 2692
rect 8044 2664 8046 2692
rect 24086 3512 24170 3568
rect 24226 3512 24310 3568
rect 24086 3230 24310 3512
rect 24086 3178 24172 3230
rect 24224 3178 24310 3230
rect 24086 2894 24310 3178
rect 24086 2842 24172 2894
rect 24224 2842 24310 2894
rect 1506 2506 1592 2558
rect 1644 2506 1730 2558
rect 1506 2222 1730 2506
rect 1506 2170 1592 2222
rect 1644 2170 1730 2222
rect 1506 1888 1730 2170
rect 1506 1832 1590 1888
rect 1646 1832 1730 1888
rect 1506 1412 1730 1832
rect 24086 2558 24310 2842
rect 24086 2506 24172 2558
rect 24224 2506 24310 2558
rect 24086 2222 24310 2506
rect 24086 2170 24172 2222
rect 24224 2170 24310 2222
rect 24086 1888 24310 2170
rect 24086 1832 24170 1888
rect 24226 1832 24310 1888
rect 24086 1412 24310 1832
<< via2 >>
rect 1926 33960 1982 33962
rect 1926 33908 1928 33960
rect 1928 33908 1980 33960
rect 1980 33908 1982 33960
rect 1926 33906 1982 33908
rect 3606 33960 3662 33962
rect 3606 33908 3608 33960
rect 3608 33908 3660 33960
rect 3660 33908 3662 33960
rect 3606 33906 3662 33908
rect 5286 33960 5342 33962
rect 5286 33908 5288 33960
rect 5288 33908 5340 33960
rect 5340 33908 5342 33960
rect 5286 33906 5342 33908
rect 6966 33960 7022 33962
rect 6966 33908 6968 33960
rect 6968 33908 7020 33960
rect 7020 33908 7022 33960
rect 6966 33906 7022 33908
rect 8646 33960 8702 33962
rect 8646 33908 8648 33960
rect 8648 33908 8700 33960
rect 8700 33908 8702 33960
rect 8646 33906 8702 33908
rect 10326 33960 10382 33962
rect 10326 33908 10328 33960
rect 10328 33908 10380 33960
rect 10380 33908 10382 33960
rect 10326 33906 10382 33908
rect 12006 33960 12062 33962
rect 12006 33908 12008 33960
rect 12008 33908 12060 33960
rect 12060 33908 12062 33960
rect 12006 33906 12062 33908
rect 13686 33960 13742 33962
rect 13686 33908 13688 33960
rect 13688 33908 13740 33960
rect 13740 33908 13742 33960
rect 13686 33906 13742 33908
rect 15366 33960 15422 33962
rect 15366 33908 15368 33960
rect 15368 33908 15420 33960
rect 15420 33908 15422 33960
rect 15366 33906 15422 33908
rect 17046 33960 17102 33962
rect 17046 33908 17048 33960
rect 17048 33908 17100 33960
rect 17100 33908 17102 33960
rect 17046 33906 17102 33908
rect 18726 33960 18782 33962
rect 18726 33908 18728 33960
rect 18728 33908 18780 33960
rect 18780 33908 18782 33960
rect 18726 33906 18782 33908
rect 20406 33960 20462 33962
rect 20406 33908 20408 33960
rect 20408 33908 20460 33960
rect 20460 33908 20462 33960
rect 20406 33906 20462 33908
rect 22086 33960 22142 33962
rect 22086 33908 22088 33960
rect 22088 33908 22140 33960
rect 22140 33908 22142 33960
rect 22086 33906 22142 33908
rect 23766 33960 23822 33962
rect 23766 33908 23768 33960
rect 23768 33908 23820 33960
rect 23820 33908 23822 33960
rect 23766 33906 23822 33908
rect 1590 32126 1646 32128
rect 1590 32074 1592 32126
rect 1592 32074 1644 32126
rect 1644 32074 1646 32126
rect 1590 32072 1646 32074
rect 1590 30446 1646 30448
rect 1590 30394 1592 30446
rect 1592 30394 1644 30446
rect 1644 30394 1646 30446
rect 1590 30392 1646 30394
rect 1590 28766 1646 28768
rect 1590 28714 1592 28766
rect 1592 28714 1644 28766
rect 1644 28714 1646 28766
rect 1590 28712 1646 28714
rect 1590 27086 1646 27088
rect 1590 27034 1592 27086
rect 1592 27034 1644 27086
rect 1644 27034 1646 27086
rect 1590 27032 1646 27034
rect 1590 25406 1646 25408
rect 1590 25354 1592 25406
rect 1592 25354 1644 25406
rect 1644 25354 1646 25406
rect 1590 25352 1646 25354
rect 1590 23726 1646 23728
rect 1590 23674 1592 23726
rect 1592 23674 1644 23726
rect 1644 23674 1646 23726
rect 1590 23672 1646 23674
rect 1590 22046 1646 22048
rect 1590 21994 1592 22046
rect 1592 21994 1644 22046
rect 1644 21994 1646 22046
rect 1590 21992 1646 21994
rect 1590 20366 1646 20368
rect 1590 20314 1592 20366
rect 1592 20314 1644 20366
rect 1644 20314 1646 20366
rect 1590 20312 1646 20314
rect 1590 18686 1646 18688
rect 1590 18634 1592 18686
rect 1592 18634 1644 18686
rect 1644 18634 1646 18686
rect 1590 18632 1646 18634
rect 1590 17006 1646 17008
rect 1590 16954 1592 17006
rect 1592 16954 1644 17006
rect 1644 16954 1646 17006
rect 1590 16952 1646 16954
rect 1590 15326 1646 15328
rect 1590 15274 1592 15326
rect 1592 15274 1644 15326
rect 1644 15274 1646 15326
rect 1590 15272 1646 15274
rect 1590 13646 1646 13648
rect 1590 13594 1592 13646
rect 1592 13594 1644 13646
rect 1644 13594 1646 13646
rect 1590 13592 1646 13594
rect 8279 13272 8335 13328
rect 9359 13276 9415 13332
rect 8279 12088 8335 12144
rect 9359 12084 9415 12140
rect 1590 11966 1646 11968
rect 1590 11914 1592 11966
rect 1592 11914 1644 11966
rect 1644 11914 1646 11966
rect 1590 11912 1646 11914
rect 8279 11596 8335 11652
rect 9359 11600 9415 11656
rect 8279 10412 8335 10468
rect 9359 10408 9415 10464
rect 1590 10286 1646 10288
rect 1590 10234 1592 10286
rect 1592 10234 1644 10286
rect 1644 10234 1646 10286
rect 1590 10232 1646 10234
rect 8279 9920 8335 9976
rect 9359 9924 9415 9980
rect 7988 8790 8044 8846
rect 1590 8606 1646 8608
rect 1590 8554 1592 8606
rect 1592 8554 1644 8606
rect 1644 8554 1646 8606
rect 1590 8552 1646 8554
rect 1590 6926 1646 6928
rect 1590 6874 1592 6926
rect 1592 6874 1644 6926
rect 1644 6874 1646 6926
rect 1590 6872 1646 6874
rect 1590 5246 1646 5248
rect 1590 5194 1592 5246
rect 1592 5194 1644 5246
rect 1644 5194 1646 5246
rect 1590 5192 1646 5194
rect 2637 3766 2693 3822
rect 1590 3566 1646 3568
rect 1590 3514 1592 3566
rect 1592 3514 1644 3566
rect 1644 3514 1646 3566
rect 1590 3512 1646 3514
rect 6159 3551 6215 3607
rect 8279 8736 8335 8792
rect 10174 13276 10230 13332
rect 10090 12084 10146 12140
rect 10006 11600 10062 11656
rect 9922 10408 9978 10464
rect 9838 9924 9894 9980
rect 9359 8732 9415 8788
rect 9754 8732 9810 8788
rect 24170 32126 24226 32128
rect 24170 32074 24172 32126
rect 24172 32074 24224 32126
rect 24224 32074 24226 32126
rect 24170 32072 24226 32074
rect 24170 30446 24226 30448
rect 24170 30394 24172 30446
rect 24172 30394 24224 30446
rect 24224 30394 24226 30446
rect 24170 30392 24226 30394
rect 24170 28766 24226 28768
rect 24170 28714 24172 28766
rect 24172 28714 24224 28766
rect 24224 28714 24226 28766
rect 24170 28712 24226 28714
rect 24170 27086 24226 27088
rect 24170 27034 24172 27086
rect 24172 27034 24224 27086
rect 24224 27034 24226 27086
rect 24170 27032 24226 27034
rect 24170 25406 24226 25408
rect 24170 25354 24172 25406
rect 24172 25354 24224 25406
rect 24224 25354 24226 25406
rect 24170 25352 24226 25354
rect 24170 23726 24226 23728
rect 24170 23674 24172 23726
rect 24172 23674 24224 23726
rect 24224 23674 24226 23726
rect 24170 23672 24226 23674
rect 24170 22046 24226 22048
rect 24170 21994 24172 22046
rect 24172 21994 24224 22046
rect 24224 21994 24226 22046
rect 24170 21992 24226 21994
rect 24170 20366 24226 20368
rect 24170 20314 24172 20366
rect 24172 20314 24224 20366
rect 24224 20314 24226 20366
rect 24170 20312 24226 20314
rect 24170 18686 24226 18688
rect 24170 18634 24172 18686
rect 24172 18634 24224 18686
rect 24224 18634 24226 18686
rect 24170 18632 24226 18634
rect 24170 17006 24226 17008
rect 24170 16954 24172 17006
rect 24172 16954 24224 17006
rect 24224 16954 24226 17006
rect 24170 16952 24226 16954
rect 24170 15326 24226 15328
rect 24170 15274 24172 15326
rect 24172 15274 24224 15326
rect 24224 15274 24226 15326
rect 24170 15272 24226 15274
rect 24170 13646 24226 13648
rect 24170 13594 24172 13646
rect 24172 13594 24224 13646
rect 24224 13594 24226 13646
rect 24170 13592 24226 13594
rect 24170 11966 24226 11968
rect 24170 11914 24172 11966
rect 24172 11914 24224 11966
rect 24224 11914 24226 11966
rect 24170 11912 24226 11914
rect 24170 10286 24226 10288
rect 24170 10234 24172 10286
rect 24172 10234 24224 10286
rect 24224 10234 24226 10286
rect 24170 10232 24226 10234
rect 24170 8606 24226 8608
rect 24170 8554 24172 8606
rect 24172 8554 24224 8606
rect 24224 8554 24226 8606
rect 24170 8552 24226 8554
rect 9554 7825 9610 7881
rect 14930 7825 14986 7881
rect 9554 6903 9610 6959
rect 18280 6903 18336 6959
rect 21174 6914 21230 6970
rect 21634 6914 21690 6970
rect 9554 6153 9610 6209
rect 16064 6153 16120 6209
rect 24170 6926 24226 6928
rect 24170 6874 24172 6926
rect 24172 6874 24224 6926
rect 24224 6874 24226 6926
rect 24170 6872 24226 6874
rect 24170 5246 24226 5248
rect 24170 5194 24172 5246
rect 24172 5194 24224 5246
rect 24224 5194 24226 5246
rect 24170 5192 24226 5194
rect 2637 2582 2693 2638
rect 7988 2636 8044 2692
rect 24170 3566 24226 3568
rect 24170 3514 24172 3566
rect 24172 3514 24224 3566
rect 24224 3514 24226 3566
rect 24170 3512 24226 3514
rect 11243 2582 11299 2638
rect 12725 2582 12781 2638
rect 1590 1886 1646 1888
rect 1590 1834 1592 1886
rect 1592 1834 1644 1886
rect 1644 1834 1646 1886
rect 1590 1832 1646 1834
rect 24170 1886 24226 1888
rect 24170 1834 24172 1886
rect 24172 1834 24224 1886
rect 24224 1834 24226 1886
rect 24170 1832 24226 1834
rect 1926 1550 1982 1552
rect 1926 1498 1928 1550
rect 1928 1498 1980 1550
rect 1980 1498 1982 1550
rect 1926 1496 1982 1498
rect 3606 1550 3662 1552
rect 3606 1498 3608 1550
rect 3608 1498 3660 1550
rect 3660 1498 3662 1550
rect 3606 1496 3662 1498
rect 5286 1550 5342 1552
rect 5286 1498 5288 1550
rect 5288 1498 5340 1550
rect 5340 1498 5342 1550
rect 5286 1496 5342 1498
rect 6966 1550 7022 1552
rect 6966 1498 6968 1550
rect 6968 1498 7020 1550
rect 7020 1498 7022 1550
rect 6966 1496 7022 1498
rect 8646 1550 8702 1552
rect 8646 1498 8648 1550
rect 8648 1498 8700 1550
rect 8700 1498 8702 1550
rect 8646 1496 8702 1498
rect 10326 1550 10382 1552
rect 10326 1498 10328 1550
rect 10328 1498 10380 1550
rect 10380 1498 10382 1550
rect 10326 1496 10382 1498
rect 12006 1550 12062 1552
rect 12006 1498 12008 1550
rect 12008 1498 12060 1550
rect 12060 1498 12062 1550
rect 12006 1496 12062 1498
rect 13686 1550 13742 1552
rect 13686 1498 13688 1550
rect 13688 1498 13740 1550
rect 13740 1498 13742 1550
rect 13686 1496 13742 1498
rect 15366 1550 15422 1552
rect 15366 1498 15368 1550
rect 15368 1498 15420 1550
rect 15420 1498 15422 1550
rect 15366 1496 15422 1498
rect 17046 1550 17102 1552
rect 17046 1498 17048 1550
rect 17048 1498 17100 1550
rect 17100 1498 17102 1550
rect 17046 1496 17102 1498
rect 18726 1550 18782 1552
rect 18726 1498 18728 1550
rect 18728 1498 18780 1550
rect 18780 1498 18782 1550
rect 18726 1496 18782 1498
rect 20406 1550 20462 1552
rect 20406 1498 20408 1550
rect 20408 1498 20460 1550
rect 20460 1498 20462 1550
rect 20406 1496 20462 1498
rect 22086 1550 22142 1552
rect 22086 1498 22088 1550
rect 22088 1498 22140 1550
rect 22140 1498 22142 1550
rect 22086 1496 22142 1498
rect 23766 1550 23822 1552
rect 23766 1498 23768 1550
rect 23768 1498 23820 1550
rect 23820 1498 23822 1550
rect 23766 1496 23822 1498
<< metal3 >>
rect 302 35158 358 35220
rect 422 35158 478 35220
rect 542 35158 25198 35220
rect 25262 35158 25318 35220
rect 25382 35158 25438 35220
rect 240 35102 25500 35158
rect 302 35038 358 35102
rect 422 35038 478 35102
rect 542 35038 25198 35102
rect 25262 35038 25318 35102
rect 25382 35038 25438 35102
rect 240 34982 25500 35038
rect 302 34920 358 34982
rect 422 34920 478 34982
rect 542 34920 10558 34982
rect 10622 34920 16198 34982
rect 16262 34920 25198 34982
rect 25262 34920 25318 34982
rect 25382 34920 25438 34982
rect 902 34558 958 34620
rect 1022 34558 1078 34620
rect 1142 34558 24598 34620
rect 24662 34558 24718 34620
rect 24782 34558 24838 34620
rect 840 34502 24900 34558
rect 902 34438 958 34502
rect 1022 34438 1078 34502
rect 1142 34438 24598 34502
rect 24662 34438 24718 34502
rect 24782 34438 24838 34502
rect 840 34382 24900 34438
rect 902 34320 958 34382
rect 1022 34320 1078 34382
rect 1142 34320 1918 34382
rect 1982 34320 3718 34382
rect 3782 34320 5278 34382
rect 5342 34320 7078 34382
rect 7142 34320 8758 34382
rect 8822 34320 10318 34382
rect 10382 34320 11998 34382
rect 12062 34320 13678 34382
rect 13742 34320 15358 34382
rect 15422 34320 17038 34382
rect 17102 34320 18838 34382
rect 18902 34320 20398 34382
rect 20462 34320 22198 34382
rect 22262 34320 23758 34382
rect 23822 34320 24598 34382
rect 24662 34320 24718 34382
rect 24782 34320 24838 34382
rect 1920 33906 1926 33958
rect 1982 33906 2100 34020
rect 1920 33840 2100 33906
rect 3600 33962 3718 34020
rect 3600 33906 3606 33962
rect 3662 33958 3718 33962
rect 3662 33906 3780 33958
rect 3600 33840 3780 33906
rect 5280 33906 5286 33958
rect 5342 33906 5460 34020
rect 5280 33840 5460 33906
rect 6960 33962 7078 34020
rect 6960 33906 6966 33962
rect 7022 33958 7078 33962
rect 8640 33962 8758 34020
rect 7022 33906 7140 33958
rect 6960 33840 7140 33906
rect 8640 33906 8646 33962
rect 8702 33958 8758 33962
rect 8702 33906 8820 33958
rect 8640 33840 8820 33906
rect 10320 33906 10326 33958
rect 10382 33906 10500 34020
rect 10320 33840 10500 33906
rect 12000 33906 12006 33958
rect 12062 33906 12180 34020
rect 12000 33902 12180 33906
rect 12062 33840 12180 33902
rect 13680 33906 13686 33958
rect 13742 33906 13860 34020
rect 13680 33840 13860 33906
rect 15360 33906 15366 33958
rect 15422 33906 15540 34020
rect 15360 33900 15540 33906
rect 17040 33906 17046 33958
rect 17102 33906 17220 34020
rect 15360 33840 16078 33900
rect 17040 33840 17220 33906
rect 18720 33962 18838 34020
rect 18720 33906 18726 33962
rect 18782 33958 18838 33962
rect 18782 33906 18900 33958
rect 18720 33840 18900 33906
rect 20400 33906 20406 33958
rect 20462 33906 20580 34020
rect 20400 33840 20580 33906
rect 22080 33962 22198 34020
rect 22080 33906 22086 33962
rect 22142 33958 22198 33962
rect 22142 33906 22260 33958
rect 22080 33840 22260 33906
rect 23760 33906 23766 33958
rect 23822 33906 23940 34020
rect 23760 33840 23940 33906
rect 10622 33000 11580 33060
rect 10622 32998 10740 33000
rect 10560 32880 10740 32998
rect 11400 32940 11580 33000
rect 11342 32880 11580 32940
rect 16080 32998 16198 33060
rect 16080 32880 16260 32998
rect 16080 32700 16140 32880
rect 14880 32640 16140 32700
rect 14880 32580 15060 32640
rect 14880 32520 16198 32580
rect 1142 32160 1740 32220
rect 1560 32128 1740 32160
rect 1560 32072 1590 32128
rect 1646 32072 1740 32128
rect 1560 32040 1740 32072
rect 24120 32160 24598 32220
rect 24120 32128 24300 32160
rect 24120 32072 24170 32128
rect 24226 32072 24300 32128
rect 24120 32040 24300 32072
rect 10560 31382 10740 31500
rect 10622 31380 10740 31382
rect 11400 31440 11998 31500
rect 11400 31380 11580 31440
rect 16142 31438 16260 31500
rect 16080 31382 16260 31438
rect 10622 31320 11580 31380
rect 16142 31320 16260 31382
rect 14880 31080 16078 31140
rect 14880 31020 15060 31080
rect 14880 30960 16078 31020
rect 1142 30480 1740 30540
rect 1560 30448 1740 30480
rect 1560 30392 1590 30448
rect 1646 30392 1740 30448
rect 1560 30360 1740 30392
rect 24120 30448 24300 30540
rect 24120 30392 24170 30448
rect 24226 30420 24300 30448
rect 24226 30392 24598 30420
rect 24120 30360 24598 30392
rect 10560 29880 11278 29940
rect 10560 29820 10740 29880
rect 11400 29822 11580 29940
rect 16080 29878 16198 29940
rect 11400 29820 11518 29822
rect 10560 29760 11518 29820
rect 16080 29760 16260 29878
rect 16080 29580 16140 29760
rect 14880 29520 16140 29580
rect 14880 29460 15060 29520
rect 14880 29400 16198 29460
rect 1560 28768 1740 28860
rect 1560 28740 1590 28768
rect 1142 28712 1590 28740
rect 1646 28712 1740 28768
rect 1142 28680 1740 28712
rect 24120 28800 24598 28860
rect 24120 28768 24300 28800
rect 24120 28712 24170 28768
rect 24226 28712 24300 28768
rect 24120 28680 24300 28712
rect 10622 28440 11580 28500
rect 10622 28438 10740 28440
rect 10560 28320 10740 28438
rect 11400 28320 11580 28440
rect 16142 28318 16260 28380
rect 16080 28200 16260 28318
rect 16080 28140 16140 28200
rect 14880 28080 16140 28140
rect 14880 28020 15060 28080
rect 14880 27960 16078 28020
rect 1560 27088 1740 27180
rect 1560 27060 1590 27088
rect 1142 27032 1590 27060
rect 1646 27032 1740 27088
rect 1142 27000 1740 27032
rect 24120 27088 24300 27180
rect 24120 27032 24170 27088
rect 24226 27060 24300 27088
rect 24226 27032 24598 27060
rect 24120 27000 24598 27032
rect 10560 26822 10740 26940
rect 10622 26820 10740 26822
rect 11400 26878 11518 26940
rect 16080 26878 16198 26940
rect 11400 26820 11580 26878
rect 10622 26760 11580 26820
rect 16080 26760 16260 26878
rect 16080 26580 16140 26760
rect 14880 26520 16140 26580
rect 14880 26460 15060 26520
rect 14880 26400 16198 26460
rect 1560 25408 1740 25500
rect 1560 25380 1590 25408
rect 1142 25352 1590 25380
rect 1646 25352 1740 25408
rect 24120 25440 24598 25500
rect 24120 25408 24300 25440
rect 1142 25320 1740 25352
rect 16142 25318 16260 25380
rect 24120 25352 24170 25408
rect 24226 25352 24300 25408
rect 24120 25320 24300 25352
rect 16080 25200 16260 25318
rect 16080 25140 16140 25200
rect 14880 25080 16140 25140
rect 14880 25020 15060 25080
rect 14880 24960 16078 25020
rect 1142 23760 1740 23820
rect 1560 23728 1740 23760
rect 10622 23760 11580 23820
rect 10622 23758 10740 23760
rect 1560 23672 1590 23728
rect 1646 23672 1740 23728
rect 1560 23640 1740 23672
rect 10560 23640 10740 23758
rect 11400 23702 11580 23760
rect 16080 23758 16198 23820
rect 24120 23760 24598 23820
rect 11400 23640 11518 23702
rect 16080 23640 16260 23758
rect 24120 23728 24300 23760
rect 24120 23672 24170 23728
rect 24226 23672 24300 23728
rect 24120 23640 24300 23672
rect 16080 23580 16140 23640
rect 14880 23520 16140 23580
rect 14880 23462 15060 23520
rect 14942 23400 15060 23462
rect 10560 22142 10740 22260
rect 1142 22080 1740 22140
rect 10560 22080 10678 22142
rect 1560 22048 1740 22080
rect 11400 22140 11580 22260
rect 16142 22198 16260 22260
rect 10742 22080 11580 22140
rect 16080 22080 16260 22198
rect 24120 22080 24598 22140
rect 1560 21992 1590 22048
rect 1646 21992 1740 22048
rect 16080 22020 16140 22080
rect 1560 21960 1740 21992
rect 14880 21960 16140 22020
rect 24120 22048 24300 22080
rect 24120 21992 24170 22048
rect 24226 21992 24300 22048
rect 24120 21960 24300 21992
rect 14880 21900 15060 21960
rect 14880 21840 16078 21900
rect 10560 20640 11518 20700
rect 10560 20580 10740 20640
rect 11400 20638 11518 20640
rect 10560 20520 11278 20580
rect 11400 20520 11580 20638
rect 16080 20580 16260 20700
rect 14942 20520 16260 20580
rect 14942 20518 15060 20520
rect 14880 20462 15060 20518
rect 1142 20400 1740 20460
rect 14880 20400 14998 20462
rect 1560 20368 1740 20400
rect 1560 20312 1590 20368
rect 1646 20312 1740 20368
rect 1560 20280 1740 20312
rect 24120 20368 24300 20460
rect 24120 20312 24170 20368
rect 24226 20340 24300 20368
rect 24226 20312 24598 20340
rect 24120 20280 24598 20312
rect 10560 19198 10678 19260
rect 10742 19200 11580 19260
rect 10560 19080 10740 19198
rect 11400 19140 11580 19200
rect 16142 19198 16260 19260
rect 11400 19080 12060 19140
rect 12000 19020 12060 19080
rect 16080 19080 16260 19198
rect 16080 19020 16140 19080
rect 12000 18960 16140 19020
rect 14880 18902 15060 18960
rect 14942 18840 15060 18902
rect 1560 18688 1740 18780
rect 1560 18660 1590 18688
rect 1142 18632 1590 18660
rect 1646 18632 1740 18688
rect 1142 18600 1740 18632
rect 24120 18688 24300 18780
rect 24120 18632 24170 18688
rect 24226 18660 24300 18688
rect 24226 18632 24598 18660
rect 24120 18600 24598 18632
rect 10560 17582 10740 17700
rect 11342 17640 11580 17700
rect 10622 17580 10740 17582
rect 11400 17580 11580 17640
rect 10622 17520 11580 17580
rect 14880 17518 14998 17580
rect 16080 17580 16260 17700
rect 15062 17520 16260 17580
rect 14880 17462 15060 17518
rect 14880 17400 14998 17462
rect 1560 17008 1740 17100
rect 1560 16980 1590 17008
rect 1142 16952 1590 16980
rect 1646 16952 1740 17008
rect 1142 16920 1740 16952
rect 24120 17008 24300 17100
rect 24120 16952 24170 17008
rect 24226 16980 24300 17008
rect 24226 16952 24598 16980
rect 24120 16920 24598 16952
rect 16080 16020 16260 16140
rect 14942 15960 16260 16020
rect 14942 15958 15060 15960
rect 14880 15902 15060 15958
rect 14942 15840 15060 15902
rect 1560 15328 1740 15420
rect 1560 15300 1590 15328
rect 1142 15272 1590 15300
rect 1646 15272 1740 15328
rect 24120 15360 24598 15420
rect 24120 15328 24300 15360
rect 1142 15240 1740 15272
rect 8760 15240 10558 15300
rect 8760 15182 8940 15240
rect 24120 15272 24170 15328
rect 24226 15272 24300 15328
rect 24120 15240 24300 15272
rect 8760 15120 8878 15182
rect 8942 15120 10558 15180
rect 10622 14518 10740 14580
rect 10560 14460 10740 14518
rect 11400 14460 11580 14580
rect 8760 14342 8940 14460
rect 10560 14400 11580 14460
rect 8822 14280 8940 14342
rect 14880 14398 14998 14460
rect 16080 14460 16260 14580
rect 15062 14400 16260 14460
rect 14880 14342 15060 14398
rect 14880 14280 14998 14342
rect 1142 13680 1740 13740
rect 1560 13648 1740 13680
rect 1560 13592 1590 13648
rect 1646 13592 1740 13648
rect 24120 13680 24598 13740
rect 24120 13648 24300 13680
rect 1560 13560 1740 13592
rect 8760 13558 8878 13620
rect 24120 13592 24170 13648
rect 24226 13592 24300 13648
rect 24120 13560 24300 13592
rect 8760 13500 8940 13558
rect 8702 13440 8940 13500
rect 8160 13328 8340 13380
rect 8160 13272 8279 13328
rect 8335 13272 8340 13328
rect 9357 13332 10232 13334
rect 9357 13276 9359 13332
rect 9415 13276 10174 13332
rect 10230 13276 10232 13332
rect 9357 13274 10232 13276
rect 8160 13260 8340 13272
rect 0 13200 8340 13260
rect 10560 12960 11580 13020
rect 10560 12840 10740 12960
rect 11400 12840 11580 12960
rect 14942 12958 15060 13020
rect 14880 12900 15060 12958
rect 16080 12902 16260 13020
rect 16080 12900 16198 12902
rect 14880 12840 16198 12900
rect 10560 12780 10620 12840
rect 8822 12720 10620 12780
rect 8822 12718 8940 12720
rect 8760 12662 8940 12718
rect 8760 12600 8878 12662
rect 0 12144 8340 12180
rect 0 12120 8279 12144
rect 8160 12088 8279 12120
rect 8335 12088 8340 12144
rect 1142 12000 1740 12060
rect 8160 12000 8340 12088
rect 9357 12140 10148 12142
rect 9357 12084 9359 12140
rect 9415 12084 10090 12140
rect 10146 12084 10148 12140
rect 9357 12082 10148 12084
rect 24120 12000 24598 12060
rect 1560 11968 1740 12000
rect 1560 11912 1590 11968
rect 1646 11912 1740 11968
rect 24120 11968 24300 12000
rect 1560 11880 1740 11912
rect 8702 11880 8940 11940
rect 24120 11912 24170 11968
rect 24226 11912 24300 11968
rect 24120 11880 24300 11912
rect 8760 11822 8940 11880
rect 8822 11820 8940 11822
rect 8822 11760 10558 11820
rect 0 11652 8340 11700
rect 0 11640 8279 11652
rect 8160 11596 8279 11640
rect 8335 11596 8340 11652
rect 9357 11656 10064 11658
rect 9357 11600 9359 11656
rect 9415 11600 10006 11656
rect 10062 11600 10064 11656
rect 9357 11598 10064 11600
rect 8160 11520 8340 11596
rect 10622 11520 10740 11580
rect 10622 11518 10638 11520
rect 10560 11340 10638 11518
rect 11400 11340 11580 11580
rect 14880 11398 14998 11460
rect 14880 11342 15060 11398
rect 10560 11280 11580 11340
rect 14942 11340 15060 11342
rect 16080 11340 16260 11460
rect 14942 11280 16260 11340
rect 8760 11038 8878 11100
rect 8760 10982 8940 11038
rect 8760 10920 8878 10982
rect 0 10468 8340 10500
rect 0 10440 8279 10468
rect 8160 10412 8279 10440
rect 8335 10412 8340 10468
rect 1142 10320 1740 10380
rect 8160 10320 8340 10412
rect 9357 10464 9980 10466
rect 9357 10408 9359 10464
rect 9415 10408 9922 10464
rect 9978 10408 9980 10464
rect 9357 10406 9980 10408
rect 1560 10288 1740 10320
rect 1560 10232 1590 10288
rect 1646 10232 1740 10288
rect 24120 10288 24300 10380
rect 1560 10200 1740 10232
rect 8822 10198 8940 10260
rect 24120 10232 24170 10288
rect 24226 10260 24300 10288
rect 24226 10232 24598 10260
rect 24120 10200 24598 10232
rect 8760 10142 8940 10198
rect 8822 10080 8940 10142
rect 8160 9976 8340 10020
rect 8160 9920 8279 9976
rect 8335 9920 8340 9976
rect 9357 9980 9896 9982
rect 9357 9924 9359 9980
rect 9415 9924 9838 9980
rect 9894 9924 9896 9980
rect 9357 9922 9896 9924
rect 8160 9900 8340 9920
rect 10560 9902 10740 10020
rect 0 9840 8340 9900
rect 10622 9900 10740 9902
rect 11400 9900 11580 10020
rect 16080 9958 16198 10020
rect 16080 9900 16260 9958
rect 10622 9840 12060 9900
rect 12000 9780 12060 9840
rect 14880 9840 16678 9900
rect 14880 9780 15060 9840
rect 12000 9720 15060 9780
rect 8760 9358 8878 9420
rect 8942 9360 10558 9420
rect 8760 9240 8940 9358
rect 7986 8846 8100 8848
rect 0 8760 1860 8820
rect 7986 8790 7988 8846
rect 8044 8790 8100 8846
rect 7986 8788 8100 8790
rect 8277 8792 8337 8794
rect 1800 8700 1860 8760
rect 8277 8736 8279 8792
rect 8335 8736 8337 8792
rect 8277 8700 8337 8736
rect 9357 8788 9812 8790
rect 9357 8732 9359 8788
rect 9415 8732 9754 8788
rect 9810 8732 9812 8788
rect 9357 8730 9812 8732
rect 1560 8608 1740 8700
rect 1800 8640 8340 8700
rect 1560 8580 1590 8608
rect 1142 8552 1590 8580
rect 1646 8552 1740 8608
rect 24120 8608 24300 8700
rect 1142 8520 1740 8552
rect 8822 8518 8940 8580
rect 24120 8552 24170 8608
rect 24226 8580 24300 8608
rect 24226 8552 24598 8580
rect 24120 8520 24598 8552
rect 8760 8460 8940 8518
rect 8760 8400 10740 8460
rect 10560 8340 10740 8400
rect 11400 8340 11580 8460
rect 14942 8398 15060 8460
rect 10560 8280 11580 8340
rect 14880 8340 15060 8398
rect 16080 8340 16260 8460
rect 14880 8280 16860 8340
rect 16680 8220 16860 8280
rect 17520 8220 17700 8340
rect 16680 8160 17700 8220
rect 9552 7881 14988 7883
rect 9552 7825 9554 7881
rect 9610 7825 14930 7881
rect 14986 7825 14988 7881
rect 9552 7823 14988 7825
rect 16742 7440 17700 7500
rect 16742 7438 16860 7440
rect 16680 7380 16860 7438
rect 16680 7320 17278 7380
rect 17520 7320 17700 7440
rect 21120 7200 21540 7260
rect 21120 7140 21180 7200
rect 21000 7080 21180 7140
rect 21480 7140 21540 7200
rect 21600 7200 22620 7260
rect 21600 7140 21660 7200
rect 21480 7080 21660 7140
rect 22560 7140 22620 7200
rect 22560 7080 25198 7140
rect 1560 6928 1740 7020
rect 21000 6998 21152 7080
rect 1560 6900 1590 6928
rect 1142 6872 1590 6900
rect 1646 6872 1740 6928
rect 9552 6959 18338 6961
rect 21000 6960 21060 6998
rect 21240 6972 21300 7020
rect 21552 6998 21612 7080
rect 21720 6972 21780 7020
rect 22648 6998 22708 7080
rect 23108 6998 23168 7080
rect 24240 6990 24598 7020
rect 21172 6970 21300 6972
rect 9552 6903 9554 6959
rect 9610 6903 18280 6959
rect 18336 6903 18338 6959
rect 9552 6901 18338 6903
rect 21172 6914 21174 6970
rect 21230 6914 21300 6970
rect 21172 6900 21300 6914
rect 21632 6970 21780 6972
rect 21632 6914 21634 6970
rect 21690 6914 21780 6970
rect 24198 6960 24598 6990
rect 24198 6930 24270 6960
rect 1142 6840 1740 6872
rect 21120 6840 21478 6900
rect 21632 6900 21780 6914
rect 24168 6928 24270 6930
rect 21600 6840 24060 6900
rect 24168 6872 24170 6928
rect 24226 6900 24270 6928
rect 24226 6872 24228 6900
rect 24168 6870 24228 6872
rect 24000 6780 24060 6840
rect 24000 6720 25740 6780
rect 21542 6600 25740 6660
rect 9552 6209 16122 6211
rect 9552 6153 9554 6209
rect 9610 6153 16064 6209
rect 16120 6153 16122 6209
rect 9552 6151 16122 6153
rect 21000 6060 21180 6180
rect 21480 6120 22740 6180
rect 21480 6060 21660 6120
rect 21000 6000 21660 6060
rect 22560 6060 22740 6120
rect 23040 6060 23220 6180
rect 22560 6000 24118 6060
rect 1560 5248 1740 5340
rect 24182 5280 24598 5340
rect 24182 5278 24300 5280
rect 1560 5220 1590 5248
rect 1142 5192 1590 5220
rect 1646 5192 1740 5248
rect 1142 5160 1740 5192
rect 24120 5248 24300 5278
rect 24120 5192 24170 5248
rect 24226 5192 24300 5248
rect 24120 5160 24300 5192
rect 16560 4860 16740 4980
rect 17342 4920 18300 4980
rect 17342 4918 17460 4920
rect 17280 4860 17460 4918
rect 16560 4800 17460 4860
rect 18120 4800 18300 4920
rect 542 4080 2580 4140
rect 2400 4022 2580 4080
rect 2400 3960 2518 4022
rect 2635 3822 2695 3824
rect 2635 3766 2637 3822
rect 2693 3766 2695 3822
rect 2635 3764 2695 3766
rect 1560 3568 1740 3660
rect 1560 3540 1590 3568
rect 1142 3512 1590 3540
rect 1646 3540 1740 3568
rect 6120 3607 6300 3660
rect 6120 3551 6159 3607
rect 6215 3551 6300 3607
rect 6120 3542 6300 3551
rect 24120 3600 24598 3660
rect 24120 3568 24300 3600
rect 1646 3512 2398 3540
rect 1142 3480 2398 3512
rect 6120 3480 6238 3542
rect 24120 3512 24170 3568
rect 24226 3512 24300 3568
rect 24120 3480 24300 3512
rect 2462 3238 2580 3300
rect 2400 3120 2580 3238
rect 11760 3240 13380 3300
rect 11760 3180 11940 3240
rect 11760 3120 11998 3180
rect 13200 3120 13380 3240
rect 11280 2694 11340 2700
rect 7986 2692 12546 2694
rect 2635 2638 2695 2640
rect 2635 2582 2637 2638
rect 2693 2582 2695 2638
rect 7986 2636 7988 2692
rect 8044 2638 12546 2692
rect 12720 2640 12780 2700
rect 8044 2636 11243 2638
rect 7986 2634 11243 2636
rect 2635 2580 2695 2582
rect 11241 2582 11243 2634
rect 11299 2634 12546 2638
rect 12723 2638 12783 2640
rect 11299 2582 11301 2634
rect 12723 2582 12725 2638
rect 12781 2582 12783 2638
rect 11241 2580 11278 2582
rect 12782 2580 12783 2582
rect 2400 2398 2518 2460
rect 11760 2400 13380 2460
rect 2400 2280 2580 2398
rect 11760 2280 11940 2400
rect 13200 2342 13380 2400
rect 13200 2280 13318 2342
rect 1560 1888 1740 1980
rect 1560 1832 1590 1888
rect 1646 1860 1740 1888
rect 24120 1920 24598 1980
rect 24120 1888 24300 1920
rect 24120 1862 24170 1888
rect 1646 1832 1918 1860
rect 1560 1800 1918 1832
rect 24226 1832 24300 1888
rect 24182 1800 24300 1832
rect 1982 1558 2100 1620
rect 1920 1552 2100 1558
rect 1920 1502 1926 1552
rect 1982 1440 2100 1552
rect 3600 1552 3780 1620
rect 3600 1496 3606 1552
rect 3662 1502 3780 1552
rect 5280 1552 5460 1620
rect 3662 1496 3718 1502
rect 3600 1440 3718 1496
rect 5280 1496 5286 1552
rect 5342 1502 5460 1552
rect 6960 1552 7140 1620
rect 5342 1496 5398 1502
rect 5280 1440 5398 1496
rect 6960 1496 6966 1552
rect 7022 1502 7140 1552
rect 8640 1552 8820 1620
rect 7022 1496 7078 1502
rect 6960 1440 7078 1496
rect 8640 1496 8646 1552
rect 8702 1502 8820 1552
rect 10320 1552 10500 1620
rect 12062 1558 12180 1620
rect 10320 1502 10326 1552
rect 8702 1496 8758 1502
rect 8640 1440 8758 1496
rect 10382 1440 10500 1552
rect 12000 1552 12180 1558
rect 12000 1502 12006 1552
rect 12062 1440 12180 1552
rect 13680 1552 13860 1620
rect 13680 1502 13686 1552
rect 13742 1440 13860 1552
rect 15360 1552 15540 1620
rect 15360 1502 15366 1552
rect 15422 1440 15540 1552
rect 17040 1552 17220 1620
rect 17040 1502 17046 1552
rect 17102 1440 17220 1552
rect 18720 1552 18900 1620
rect 18720 1496 18726 1552
rect 18782 1502 18900 1552
rect 20400 1552 20580 1620
rect 20400 1502 20406 1552
rect 18782 1496 18838 1502
rect 18720 1440 18838 1496
rect 20462 1440 20580 1552
rect 22080 1552 22260 1620
rect 22080 1502 22086 1552
rect 22142 1440 22260 1552
rect 23760 1560 24118 1620
rect 23760 1552 23940 1560
rect 23760 1496 23766 1552
rect 23822 1496 23940 1552
rect 23760 1440 23940 1496
rect 902 1078 958 1140
rect 1022 1078 1078 1140
rect 1142 1078 1918 1140
rect 1982 1078 3718 1140
rect 3782 1078 5398 1140
rect 5462 1078 7078 1140
rect 7142 1078 8758 1140
rect 8822 1078 10318 1140
rect 10382 1078 11998 1140
rect 12062 1078 13678 1140
rect 13742 1078 15358 1140
rect 15422 1078 17038 1140
rect 17102 1078 18838 1140
rect 18902 1078 20398 1140
rect 20462 1078 22078 1140
rect 22142 1078 24598 1140
rect 24662 1078 24718 1140
rect 24782 1078 24838 1140
rect 840 1022 24900 1078
rect 902 958 958 1022
rect 1022 958 1078 1022
rect 1142 958 24598 1022
rect 24662 958 24718 1022
rect 24782 958 24838 1022
rect 840 902 24900 958
rect 902 840 958 902
rect 1022 840 1078 902
rect 1142 840 24598 902
rect 24662 840 24718 902
rect 24782 840 24838 902
rect 302 478 358 540
rect 422 478 478 540
rect 542 478 13318 540
rect 13382 478 25198 540
rect 25262 478 25318 540
rect 25382 478 25438 540
rect 240 422 25500 478
rect 302 358 358 422
rect 422 358 478 422
rect 542 358 25198 422
rect 25262 358 25318 422
rect 25382 358 25438 422
rect 240 302 25500 358
rect 302 240 358 302
rect 422 240 478 302
rect 542 240 25198 302
rect 25262 240 25318 302
rect 25382 240 25438 302
<< via3 >>
rect 238 35158 302 35222
rect 358 35158 422 35222
rect 478 35158 542 35222
rect 25198 35158 25262 35222
rect 25318 35158 25382 35222
rect 25438 35158 25502 35222
rect 238 35038 302 35102
rect 358 35038 422 35102
rect 478 35038 542 35102
rect 25198 35038 25262 35102
rect 25318 35038 25382 35102
rect 25438 35038 25502 35102
rect 238 34918 302 34982
rect 358 34918 422 34982
rect 478 34918 542 34982
rect 10558 34918 10622 34982
rect 16198 34918 16262 34982
rect 25198 34918 25262 34982
rect 25318 34918 25382 34982
rect 25438 34918 25502 34982
rect 838 34558 902 34622
rect 958 34558 1022 34622
rect 1078 34558 1142 34622
rect 24598 34558 24662 34622
rect 24718 34558 24782 34622
rect 24838 34558 24902 34622
rect 838 34438 902 34502
rect 958 34438 1022 34502
rect 1078 34438 1142 34502
rect 24598 34438 24662 34502
rect 24718 34438 24782 34502
rect 24838 34438 24902 34502
rect 838 34318 902 34382
rect 958 34318 1022 34382
rect 1078 34318 1142 34382
rect 1918 34318 1982 34382
rect 3718 34318 3782 34382
rect 5278 34318 5342 34382
rect 7078 34318 7142 34382
rect 8758 34318 8822 34382
rect 10318 34318 10382 34382
rect 11998 34318 12062 34382
rect 13678 34318 13742 34382
rect 15358 34318 15422 34382
rect 17038 34318 17102 34382
rect 18838 34318 18902 34382
rect 20398 34318 20462 34382
rect 22198 34318 22262 34382
rect 23758 34318 23822 34382
rect 24598 34318 24662 34382
rect 24718 34318 24782 34382
rect 24838 34318 24902 34382
rect 1918 33962 1982 34022
rect 1918 33958 1926 33962
rect 1926 33958 1982 33962
rect 3718 33958 3782 34022
rect 5278 33962 5342 34022
rect 5278 33958 5286 33962
rect 5286 33958 5342 33962
rect 7078 33958 7142 34022
rect 8758 33958 8822 34022
rect 10318 33962 10382 34022
rect 10318 33958 10326 33962
rect 10326 33958 10382 33962
rect 11998 33962 12062 34022
rect 11998 33958 12006 33962
rect 12006 33958 12062 33962
rect 13678 33962 13742 34022
rect 13678 33958 13686 33962
rect 13686 33958 13742 33962
rect 11998 33838 12062 33902
rect 15358 33962 15422 34022
rect 15358 33958 15366 33962
rect 15366 33958 15422 33962
rect 17038 33962 17102 34022
rect 17038 33958 17046 33962
rect 17046 33958 17102 33962
rect 16078 33838 16142 33902
rect 18838 33958 18902 34022
rect 20398 33962 20462 34022
rect 20398 33958 20406 33962
rect 20406 33958 20462 33962
rect 22198 33958 22262 34022
rect 23758 33962 23822 34022
rect 23758 33958 23766 33962
rect 23766 33958 23822 33962
rect 10558 32998 10622 33062
rect 11278 32878 11342 32942
rect 16198 32998 16262 33062
rect 16198 32518 16262 32582
rect 1078 32158 1142 32222
rect 24598 32158 24662 32222
rect 10558 31318 10622 31382
rect 11998 31438 12062 31502
rect 16078 31438 16142 31502
rect 16078 31318 16142 31382
rect 16078 31078 16142 31142
rect 16078 30958 16142 31022
rect 1078 30478 1142 30542
rect 24598 30358 24662 30422
rect 11278 29878 11342 29942
rect 16198 29878 16262 29942
rect 11518 29758 11582 29822
rect 16198 29398 16262 29462
rect 1078 28678 1142 28742
rect 24598 28798 24662 28862
rect 10558 28438 10622 28502
rect 16078 28318 16142 28382
rect 16078 27958 16142 28022
rect 1078 26998 1142 27062
rect 24598 26998 24662 27062
rect 10558 26758 10622 26822
rect 11518 26878 11582 26942
rect 16198 26878 16262 26942
rect 16198 26398 16262 26462
rect 1078 25318 1142 25382
rect 24598 25438 24662 25502
rect 16078 25318 16142 25382
rect 16078 24958 16142 25022
rect 1078 23758 1142 23822
rect 10558 23758 10622 23822
rect 16198 23758 16262 23822
rect 11518 23638 11582 23702
rect 24598 23758 24662 23822
rect 14878 23398 14942 23462
rect 1078 22078 1142 22142
rect 10678 22078 10742 22142
rect 16078 22198 16142 22262
rect 24598 22078 24662 22142
rect 16078 21838 16142 21902
rect 11518 20638 11582 20702
rect 11278 20518 11342 20582
rect 14878 20518 14942 20582
rect 1078 20398 1142 20462
rect 14998 20398 15062 20462
rect 24598 20278 24662 20342
rect 10678 19198 10742 19262
rect 16078 19198 16142 19262
rect 14878 18838 14942 18902
rect 1078 18598 1142 18662
rect 24598 18598 24662 18662
rect 11278 17638 11342 17702
rect 10558 17518 10622 17582
rect 14998 17518 15062 17582
rect 14998 17398 15062 17462
rect 1078 16918 1142 16982
rect 24598 16918 24662 16982
rect 14878 15958 14942 16022
rect 14878 15838 14942 15902
rect 1078 15238 1142 15302
rect 24598 15358 24662 15422
rect 10558 15238 10622 15302
rect 8878 15118 8942 15182
rect 10558 15118 10622 15182
rect 10558 14518 10622 14582
rect 8758 14278 8822 14342
rect 14998 14398 15062 14462
rect 14998 14278 15062 14342
rect 1078 13678 1142 13742
rect 24598 13678 24662 13742
rect 8878 13558 8942 13622
rect 8638 13438 8702 13502
rect 14878 12958 14942 13022
rect 8758 12718 8822 12782
rect 16198 12838 16262 12902
rect 8878 12598 8942 12662
rect 1078 11998 1142 12062
rect 24598 11998 24662 12062
rect 8638 11878 8702 11942
rect 8758 11758 8822 11822
rect 10558 11758 10622 11822
rect 10558 11518 10622 11582
rect 14998 11398 15062 11462
rect 14878 11278 14942 11342
rect 8878 11038 8942 11102
rect 8878 10918 8942 10982
rect 1078 10318 1142 10382
rect 8758 10198 8822 10262
rect 24598 10198 24662 10262
rect 8758 10078 8822 10142
rect 10558 9838 10622 9902
rect 16198 9958 16262 10022
rect 16678 9838 16742 9902
rect 8878 9358 8942 9422
rect 10558 9358 10622 9422
rect 1078 8518 1142 8582
rect 8758 8518 8822 8582
rect 24598 8518 24662 8582
rect 14878 8398 14942 8462
rect 16678 7438 16742 7502
rect 17278 7318 17342 7382
rect 1078 6838 1142 6902
rect 25198 7078 25262 7142
rect 24598 6958 24662 7022
rect 21478 6838 21542 6902
rect 21478 6598 21542 6662
rect 24118 5998 24182 6062
rect 24118 5278 24182 5342
rect 24598 5278 24662 5342
rect 1078 5158 1142 5222
rect 17278 4918 17342 4982
rect 478 4078 542 4142
rect 2518 3958 2582 4022
rect 1078 3478 1142 3542
rect 24598 3598 24662 3662
rect 2398 3478 2462 3542
rect 6238 3478 6302 3542
rect 2398 3238 2462 3302
rect 11998 3118 12062 3182
rect 11278 2518 11342 2582
rect 12718 2518 12782 2582
rect 2518 2398 2582 2462
rect 13318 2278 13382 2342
rect 24598 1918 24662 1982
rect 1918 1798 1982 1862
rect 24118 1832 24170 1862
rect 24170 1832 24182 1862
rect 24118 1798 24182 1832
rect 1918 1558 1982 1622
rect 1918 1496 1926 1502
rect 1926 1496 1982 1502
rect 1918 1438 1982 1496
rect 3718 1438 3782 1502
rect 5398 1438 5462 1502
rect 7078 1438 7142 1502
rect 11998 1558 12062 1622
rect 8758 1438 8822 1502
rect 10318 1496 10326 1502
rect 10326 1496 10382 1502
rect 10318 1438 10382 1496
rect 11998 1496 12006 1502
rect 12006 1496 12062 1502
rect 11998 1438 12062 1496
rect 13678 1496 13686 1502
rect 13686 1496 13742 1502
rect 13678 1438 13742 1496
rect 15358 1496 15366 1502
rect 15366 1496 15422 1502
rect 15358 1438 15422 1496
rect 17038 1496 17046 1502
rect 17046 1496 17102 1502
rect 17038 1438 17102 1496
rect 18838 1438 18902 1502
rect 20398 1496 20406 1502
rect 20406 1496 20462 1502
rect 20398 1438 20462 1496
rect 22078 1496 22086 1502
rect 22086 1496 22142 1502
rect 22078 1438 22142 1496
rect 24118 1558 24182 1622
rect 838 1078 902 1142
rect 958 1078 1022 1142
rect 1078 1078 1142 1142
rect 1918 1078 1982 1142
rect 3718 1078 3782 1142
rect 5398 1078 5462 1142
rect 7078 1078 7142 1142
rect 8758 1078 8822 1142
rect 10318 1078 10382 1142
rect 11998 1078 12062 1142
rect 13678 1078 13742 1142
rect 15358 1078 15422 1142
rect 17038 1078 17102 1142
rect 18838 1078 18902 1142
rect 20398 1078 20462 1142
rect 22078 1078 22142 1142
rect 24598 1078 24662 1142
rect 24718 1078 24782 1142
rect 24838 1078 24902 1142
rect 838 958 902 1022
rect 958 958 1022 1022
rect 1078 958 1142 1022
rect 24598 958 24662 1022
rect 24718 958 24782 1022
rect 24838 958 24902 1022
rect 838 838 902 902
rect 958 838 1022 902
rect 1078 838 1142 902
rect 24598 838 24662 902
rect 24718 838 24782 902
rect 24838 838 24902 902
rect 238 478 302 542
rect 358 478 422 542
rect 478 478 542 542
rect 13318 478 13382 542
rect 25198 478 25262 542
rect 25318 478 25382 542
rect 25438 478 25502 542
rect 238 358 302 422
rect 358 358 422 422
rect 478 358 542 422
rect 25198 358 25262 422
rect 25318 358 25382 422
rect 25438 358 25502 422
rect 238 238 302 302
rect 358 238 422 302
rect 478 238 542 302
rect 25198 238 25262 302
rect 25318 238 25382 302
rect 25438 238 25502 302
<< metal4 >>
rect 302 35158 358 35220
rect 422 35158 478 35220
rect 25262 35158 25318 35220
rect 25382 35158 25438 35220
rect 240 35102 540 35158
rect 25200 35102 25500 35158
rect 302 35038 358 35102
rect 422 35038 478 35102
rect 25262 35038 25318 35102
rect 25382 35038 25438 35102
rect 240 34982 540 35038
rect 25200 34982 25500 35038
rect 302 34918 358 34982
rect 422 34918 478 34982
rect 25262 34918 25318 34982
rect 25382 34918 25438 34982
rect 240 4142 540 34918
rect 902 34558 958 34620
rect 1022 34558 1078 34620
rect 840 34502 1140 34558
rect 902 34438 958 34502
rect 1022 34438 1078 34502
rect 840 34382 1140 34438
rect 902 34318 958 34382
rect 1022 34318 1078 34382
rect 840 32222 1140 34318
rect 1920 34022 1980 34318
rect 3720 34022 3780 34318
rect 5280 34022 5340 34318
rect 7080 34022 7140 34318
rect 8760 34022 8820 34318
rect 10320 34022 10380 34318
rect 10560 33062 10620 34918
rect 12000 34022 12060 34318
rect 13680 34022 13740 34318
rect 15360 34022 15420 34318
rect 840 32158 1078 32222
rect 840 30542 1140 32158
rect 840 30478 1078 30542
rect 840 28742 1140 30478
rect 840 28678 1078 28742
rect 840 27062 1140 28678
rect 10560 28502 10620 31318
rect 11280 29942 11340 32878
rect 12000 31502 12060 33838
rect 16080 31502 16140 33838
rect 16200 33062 16260 34918
rect 24662 34558 24718 34620
rect 24782 34558 24838 34620
rect 24600 34502 24900 34558
rect 24662 34438 24718 34502
rect 24782 34438 24838 34502
rect 24600 34382 24900 34438
rect 24662 34318 24718 34382
rect 24782 34318 24838 34382
rect 17040 34022 17100 34318
rect 18840 34022 18900 34318
rect 20400 34022 20460 34318
rect 22200 34022 22260 34318
rect 23760 34022 23820 34318
rect 16080 31142 16140 31318
rect 840 26998 1078 27062
rect 840 25382 1140 26998
rect 11520 26942 11580 29758
rect 16080 28382 16140 30958
rect 16200 29942 16260 32518
rect 24600 32222 24900 34318
rect 24662 32158 24900 32222
rect 24600 30422 24900 32158
rect 24662 30358 24900 30422
rect 840 25318 1078 25382
rect 840 23822 1140 25318
rect 10560 23822 10620 26758
rect 16080 25382 16140 27958
rect 16200 26942 16260 29398
rect 24600 28862 24900 30358
rect 24662 28798 24900 28862
rect 24600 27062 24900 28798
rect 24662 26998 24900 27062
rect 840 23758 1078 23822
rect 840 22142 1140 23758
rect 840 22078 1078 22142
rect 840 20462 1140 22078
rect 840 20398 1078 20462
rect 840 18662 1140 20398
rect 10680 19262 10740 22078
rect 11520 20702 11580 23638
rect 14880 20582 14940 23398
rect 16080 22262 16140 24958
rect 16200 23822 16260 26398
rect 24600 25502 24900 26998
rect 24662 25438 24900 25502
rect 24600 23822 24900 25438
rect 24662 23758 24900 23822
rect 24600 22142 24900 23758
rect 24662 22078 24900 22142
rect 840 18598 1078 18662
rect 840 16982 1140 18598
rect 11280 17702 11340 20518
rect 840 16918 1078 16982
rect 840 15302 1140 16918
rect 10560 15302 10620 17518
rect 14880 16022 14940 18838
rect 15000 17582 15060 20398
rect 16080 19262 16140 21838
rect 24600 20342 24900 22078
rect 24662 20278 24900 20342
rect 24600 18662 24900 20278
rect 24662 18598 24900 18662
rect 840 15238 1078 15302
rect 840 13742 1140 15238
rect 840 13678 1078 13742
rect 840 12062 1140 13678
rect 840 11998 1078 12062
rect 840 10382 1140 11998
rect 8640 11942 8700 13438
rect 8760 12782 8820 14278
rect 8880 13622 8940 15118
rect 10560 14582 10620 15118
rect 14880 13022 14940 15838
rect 15000 14462 15060 17398
rect 24600 16982 24900 18598
rect 24662 16918 24900 16982
rect 24600 15422 24900 16918
rect 24662 15358 24900 15422
rect 840 10318 1078 10382
rect 840 8582 1140 10318
rect 8760 10262 8820 11758
rect 8880 11102 8940 12598
rect 10560 11582 10620 11758
rect 15000 11462 15060 14278
rect 24600 13742 24900 15358
rect 24662 13678 24900 13742
rect 8760 8582 8820 10078
rect 8880 9422 8940 10918
rect 10560 9422 10620 9838
rect 840 8518 1078 8582
rect 840 6902 1140 8518
rect 14880 8462 14940 11278
rect 16200 10022 16260 12838
rect 24600 12062 24900 13678
rect 24662 11998 24900 12062
rect 24600 10262 24900 11998
rect 24662 10198 24900 10262
rect 16680 7502 16740 9838
rect 24600 8582 24900 10198
rect 24662 8518 24900 8582
rect 840 6838 1078 6902
rect 840 5222 1140 6838
rect 840 5158 1078 5222
rect 240 4078 478 4142
rect 240 542 540 4078
rect 840 3542 1140 5158
rect 17280 4982 17340 7318
rect 24600 7022 24900 8518
rect 25200 7142 25500 34918
rect 25262 7078 25500 7142
rect 24662 6958 24900 7022
rect 21480 6662 21540 6838
rect 24120 5342 24180 5998
rect 24600 5342 24900 6958
rect 24662 5278 24900 5342
rect 840 3478 1078 3542
rect 840 1142 1140 3478
rect 2400 3302 2460 3478
rect 2520 2462 2580 3958
rect 24600 3662 24900 5278
rect 24662 3598 24900 3662
rect 1920 1622 1980 1798
rect 1920 1142 1980 1438
rect 3720 1142 3780 1438
rect 5400 1142 5460 1438
rect 902 1078 958 1142
rect 1022 1078 1078 1142
rect 840 1022 1140 1078
rect 902 958 958 1022
rect 1022 958 1078 1022
rect 840 902 1140 958
rect 902 840 958 902
rect 1022 840 1078 902
rect 302 478 358 542
rect 422 478 478 542
rect 240 422 540 478
rect 302 358 358 422
rect 422 358 478 422
rect 240 302 540 358
rect 302 240 358 302
rect 422 240 478 302
rect 6240 0 6300 3478
rect 7080 1142 7140 1438
rect 8760 1142 8820 1438
rect 10320 1142 10380 1438
rect 11280 0 11340 2518
rect 12000 1622 12060 3118
rect 12000 1142 12060 1438
rect 12720 0 12780 2518
rect 13320 542 13380 2278
rect 24600 1982 24900 3598
rect 24662 1918 24900 1982
rect 24120 1622 24180 1798
rect 13680 1142 13740 1438
rect 15360 1142 15420 1438
rect 17040 1142 17100 1438
rect 18840 1142 18900 1438
rect 20400 1142 20460 1438
rect 22080 1142 22140 1438
rect 24600 1142 24900 1918
rect 24662 1078 24718 1142
rect 24782 1078 24838 1142
rect 24600 1022 24900 1078
rect 24662 958 24718 1022
rect 24782 958 24838 1022
rect 24600 902 24900 958
rect 24662 840 24718 902
rect 24782 840 24838 902
rect 25200 542 25500 7078
rect 25262 478 25318 542
rect 25382 478 25438 542
rect 25200 422 25500 478
rect 25262 358 25318 422
rect 25382 358 25438 422
rect 25200 302 25500 358
rect 25262 240 25318 302
rect 25382 240 25438 302
use contact_28  contact_28_0
timestamp 1643593061
transform 1 0 25200 0 1 7080
box 0 0 1 1
use contact_28  contact_28_1
timestamp 1643593061
transform 1 0 16200 0 1 34920
box 0 0 1 1
use contact_28  contact_28_2
timestamp 1643593061
transform 1 0 16200 0 1 33000
box 0 0 1 1
use contact_28  contact_28_3
timestamp 1643593061
transform 1 0 16200 0 1 26880
box 0 0 1 1
use contact_28  contact_28_4
timestamp 1643593061
transform 1 0 16200 0 1 29400
box 0 0 1 1
use contact_28  contact_28_5
timestamp 1643593061
transform 1 0 16200 0 1 23760
box 0 0 1 1
use contact_28  contact_28_6
timestamp 1643593061
transform 1 0 16200 0 1 26400
box 0 0 1 1
use contact_28  contact_28_7
timestamp 1643593061
transform 1 0 15000 0 1 20400
box 0 0 1 1
use contact_28  contact_28_8
timestamp 1643593061
transform 1 0 15000 0 1 17520
box 0 0 1 1
use contact_28  contact_28_9
timestamp 1643593061
transform 1 0 15000 0 1 11400
box 0 0 1 1
use contact_28  contact_28_10
timestamp 1643593061
transform 1 0 15000 0 1 14280
box 0 0 1 1
use contact_28  contact_28_11
timestamp 1643593061
transform 1 0 15000 0 1 17400
box 0 0 1 1
use contact_28  contact_28_12
timestamp 1643593061
transform 1 0 15000 0 1 14400
box 0 0 1 1
use contact_28  contact_28_13
timestamp 1643593061
transform 1 0 16200 0 1 29880
box 0 0 1 1
use contact_28  contact_28_14
timestamp 1643593061
transform 1 0 16200 0 1 32520
box 0 0 1 1
use contact_28  contact_28_15
timestamp 1643593061
transform 1 0 14880 0 1 11280
box 0 0 1 1
use contact_28  contact_28_16
timestamp 1643593061
transform 1 0 14880 0 1 8400
box 0 0 1 1
use contact_28  contact_28_17
timestamp 1643593061
transform 1 0 14880 0 1 20520
box 0 0 1 1
use contact_28  contact_28_18
timestamp 1643593061
transform 1 0 14880 0 1 23400
box 0 0 1 1
use contact_28  contact_28_19
timestamp 1643593061
transform 1 0 13320 0 1 480
box 0 0 1 1
use contact_28  contact_28_20
timestamp 1643593061
transform 1 0 13320 0 1 2280
box 0 0 1 1
use contact_28  contact_28_21
timestamp 1643593061
transform 1 0 11520 0 1 29760
box 0 0 1 1
use contact_28  contact_28_22
timestamp 1643593061
transform 1 0 11520 0 1 26880
box 0 0 1 1
use contact_28  contact_28_23
timestamp 1643593061
transform 1 0 11520 0 1 20640
box 0 0 1 1
use contact_28  contact_28_24
timestamp 1643593061
transform 1 0 11520 0 1 23640
box 0 0 1 1
use contact_28  contact_28_25
timestamp 1643593061
transform 1 0 10560 0 1 34920
box 0 0 1 1
use contact_28  contact_28_26
timestamp 1643593061
transform 1 0 10560 0 1 33000
box 0 0 1 1
use contact_28  contact_28_27
timestamp 1643593061
transform 1 0 11280 0 1 17640
box 0 0 1 1
use contact_28  contact_28_28
timestamp 1643593061
transform 1 0 11280 0 1 20520
box 0 0 1 1
use contact_28  contact_28_29
timestamp 1643593061
transform 1 0 10560 0 1 23760
box 0 0 1 1
use contact_28  contact_28_30
timestamp 1643593061
transform 1 0 10560 0 1 26760
box 0 0 1 1
use contact_28  contact_28_31
timestamp 1643593061
transform 1 0 11280 0 1 32880
box 0 0 1 1
use contact_28  contact_28_32
timestamp 1643593061
transform 1 0 11280 0 1 29880
box 0 0 1 1
use contact_28  contact_28_33
timestamp 1643593061
transform 1 0 10560 0 1 11520
box 0 0 1 1
use contact_28  contact_28_34
timestamp 1643593061
transform 1 0 10560 0 1 11760
box 0 0 1 1
use contact_28  contact_28_35
timestamp 1643593061
transform 1 0 8640 0 1 11880
box 0 0 1 1
use contact_28  contact_28_36
timestamp 1643593061
transform 1 0 8640 0 1 13440
box 0 0 1 1
use contact_28  contact_28_37
timestamp 1643593061
transform 1 0 8760 0 1 11760
box 0 0 1 1
use contact_28  contact_28_38
timestamp 1643593061
transform 1 0 8760 0 1 10200
box 0 0 1 1
use contact_28  contact_28_39
timestamp 1643593061
transform 1 0 8760 0 1 8520
box 0 0 1 1
use contact_28  contact_28_40
timestamp 1643593061
transform 1 0 8760 0 1 10080
box 0 0 1 1
use contact_28  contact_28_41
timestamp 1643593061
transform 1 0 10560 0 1 17520
box 0 0 1 1
use contact_28  contact_28_42
timestamp 1643593061
transform 1 0 10560 0 1 15240
box 0 0 1 1
use contact_28  contact_28_43
timestamp 1643593061
transform 1 0 10560 0 1 14520
box 0 0 1 1
use contact_28  contact_28_44
timestamp 1643593061
transform 1 0 10560 0 1 15120
box 0 0 1 1
use contact_28  contact_28_45
timestamp 1643593061
transform 1 0 8880 0 1 13560
box 0 0 1 1
use contact_28  contact_28_46
timestamp 1643593061
transform 1 0 8880 0 1 15120
box 0 0 1 1
use contact_28  contact_28_47
timestamp 1643593061
transform 1 0 480 0 1 4080
box 0 0 1 1
use contact_28  contact_28_48
timestamp 1643593061
transform 1 0 2520 0 1 3960
box 0 0 1 1
use contact_28  contact_28_49
timestamp 1643593061
transform 1 0 2520 0 1 2400
box 0 0 1 1
use contact_28  contact_28_50
timestamp 1643593061
transform 1 0 24600 0 1 6960
box 0 0 1 1
use contact_28  contact_28_51
timestamp 1643593061
transform 1 0 24600 0 1 23760
box 0 0 1 1
use contact_28  contact_28_52
timestamp 1643593061
transform 1 0 24600 0 1 18600
box 0 0 1 1
use contact_28  contact_28_53
timestamp 1643593061
transform 1 0 24600 0 1 15360
box 0 0 1 1
use contact_28  contact_28_54
timestamp 1643593061
transform 1 0 24600 0 1 27000
box 0 0 1 1
use contact_28  contact_28_55
timestamp 1643593061
transform 1 0 24600 0 1 3600
box 0 0 1 1
use contact_28  contact_28_56
timestamp 1643593061
transform 1 0 24600 0 1 25440
box 0 0 1 1
use contact_28  contact_28_57
timestamp 1643593061
transform 1 0 24600 0 1 10200
box 0 0 1 1
use contact_28  contact_28_58
timestamp 1643593061
transform 1 0 24600 0 1 20280
box 0 0 1 1
use contact_28  contact_28_59
timestamp 1643593061
transform 1 0 24600 0 1 28800
box 0 0 1 1
use contact_28  contact_28_60
timestamp 1643593061
transform 1 0 24600 0 1 8520
box 0 0 1 1
use contact_28  contact_28_61
timestamp 1643593061
transform 1 0 24600 0 1 22080
box 0 0 1 1
use contact_28  contact_28_62
timestamp 1643593061
transform 1 0 24600 0 1 13680
box 0 0 1 1
use contact_28  contact_28_63
timestamp 1643593061
transform 1 0 24600 0 1 1920
box 0 0 1 1
use contact_28  contact_28_64
timestamp 1643593061
transform 1 0 24600 0 1 16920
box 0 0 1 1
use contact_28  contact_28_65
timestamp 1643593061
transform 1 0 24600 0 1 30360
box 0 0 1 1
use contact_28  contact_28_66
timestamp 1643593061
transform 1 0 24600 0 1 12000
box 0 0 1 1
use contact_28  contact_28_67
timestamp 1643593061
transform 1 0 24600 0 1 5280
box 0 0 1 1
use contact_28  contact_28_68
timestamp 1643593061
transform 1 0 24600 0 1 32160
box 0 0 1 1
use contact_28  contact_28_69
timestamp 1643593061
transform 1 0 23760 0 1 34320
box 0 0 1 1
use contact_28  contact_28_70
timestamp 1643593061
transform 1 0 23760 0 1 33960
box 0 0 1 1
use contact_28  contact_28_71
timestamp 1643593061
transform 1 0 24120 0 1 1800
box 0 0 1 1
use contact_28  contact_28_72
timestamp 1643593061
transform 1 0 24120 0 1 1560
box 0 0 1 1
use contact_28  contact_28_73
timestamp 1643593061
transform 1 0 24120 0 1 5280
box 0 0 1 1
use contact_28  contact_28_74
timestamp 1643593061
transform 1 0 24120 0 1 6000
box 0 0 1 1
use contact_28  contact_28_75
timestamp 1643593061
transform 1 0 22080 0 1 1080
box 0 0 1 1
use contact_28  contact_28_76
timestamp 1643593061
transform 1 0 22080 0 1 1440
box 0 0 1 1
use contact_28  contact_28_77
timestamp 1643593061
transform 1 0 22200 0 1 34320
box 0 0 1 1
use contact_28  contact_28_78
timestamp 1643593061
transform 1 0 22200 0 1 33960
box 0 0 1 1
use contact_28  contact_28_79
timestamp 1643593061
transform 1 0 20400 0 1 34320
box 0 0 1 1
use contact_28  contact_28_80
timestamp 1643593061
transform 1 0 20400 0 1 33960
box 0 0 1 1
use contact_28  contact_28_81
timestamp 1643593061
transform 1 0 20400 0 1 1080
box 0 0 1 1
use contact_28  contact_28_82
timestamp 1643593061
transform 1 0 20400 0 1 1440
box 0 0 1 1
use contact_28  contact_28_83
timestamp 1643593061
transform 1 0 18840 0 1 1080
box 0 0 1 1
use contact_28  contact_28_84
timestamp 1643593061
transform 1 0 18840 0 1 1440
box 0 0 1 1
use contact_28  contact_28_85
timestamp 1643593061
transform 1 0 18840 0 1 34320
box 0 0 1 1
use contact_28  contact_28_86
timestamp 1643593061
transform 1 0 18840 0 1 33960
box 0 0 1 1
use contact_28  contact_28_87
timestamp 1643593061
transform 1 0 17040 0 1 1080
box 0 0 1 1
use contact_28  contact_28_88
timestamp 1643593061
transform 1 0 17040 0 1 1440
box 0 0 1 1
use contact_28  contact_28_89
timestamp 1643593061
transform 1 0 17040 0 1 34320
box 0 0 1 1
use contact_28  contact_28_90
timestamp 1643593061
transform 1 0 17040 0 1 33960
box 0 0 1 1
use contact_28  contact_28_91
timestamp 1643593061
transform 1 0 17280 0 1 4920
box 0 0 1 1
use contact_28  contact_28_92
timestamp 1643593061
transform 1 0 17280 0 1 7320
box 0 0 1 1
use contact_28  contact_28_93
timestamp 1643593061
transform 1 0 16680 0 1 7440
box 0 0 1 1
use contact_28  contact_28_94
timestamp 1643593061
transform 1 0 16680 0 1 9840
box 0 0 1 1
use contact_28  contact_28_95
timestamp 1643593061
transform 1 0 16200 0 1 9960
box 0 0 1 1
use contact_28  contact_28_96
timestamp 1643593061
transform 1 0 16200 0 1 12840
box 0 0 1 1
use contact_28  contact_28_97
timestamp 1643593061
transform 1 0 15360 0 1 1080
box 0 0 1 1
use contact_28  contact_28_98
timestamp 1643593061
transform 1 0 15360 0 1 1440
box 0 0 1 1
use contact_28  contact_28_99
timestamp 1643593061
transform 1 0 15360 0 1 34320
box 0 0 1 1
use contact_28  contact_28_100
timestamp 1643593061
transform 1 0 15360 0 1 33960
box 0 0 1 1
use contact_28  contact_28_101
timestamp 1643593061
transform 1 0 16080 0 1 31440
box 0 0 1 1
use contact_28  contact_28_102
timestamp 1643593061
transform 1 0 16080 0 1 33840
box 0 0 1 1
use contact_28  contact_28_103
timestamp 1643593061
transform 1 0 16080 0 1 19200
box 0 0 1 1
use contact_28  contact_28_104
timestamp 1643593061
transform 1 0 16080 0 1 21840
box 0 0 1 1
use contact_28  contact_28_105
timestamp 1643593061
transform 1 0 16080 0 1 25320
box 0 0 1 1
use contact_28  contact_28_106
timestamp 1643593061
transform 1 0 16080 0 1 27960
box 0 0 1 1
use contact_28  contact_28_107
timestamp 1643593061
transform 1 0 14880 0 1 12960
box 0 0 1 1
use contact_28  contact_28_108
timestamp 1643593061
transform 1 0 14880 0 1 15840
box 0 0 1 1
use contact_28  contact_28_109
timestamp 1643593061
transform 1 0 16080 0 1 31320
box 0 0 1 1
use contact_28  contact_28_110
timestamp 1643593061
transform 1 0 16080 0 1 31080
box 0 0 1 1
use contact_28  contact_28_111
timestamp 1643593061
transform 1 0 16080 0 1 28320
box 0 0 1 1
use contact_28  contact_28_112
timestamp 1643593061
transform 1 0 16080 0 1 30960
box 0 0 1 1
use contact_28  contact_28_113
timestamp 1643593061
transform 1 0 14880 0 1 15960
box 0 0 1 1
use contact_28  contact_28_114
timestamp 1643593061
transform 1 0 14880 0 1 18840
box 0 0 1 1
use contact_28  contact_28_115
timestamp 1643593061
transform 1 0 16080 0 1 22200
box 0 0 1 1
use contact_28  contact_28_116
timestamp 1643593061
transform 1 0 16080 0 1 24960
box 0 0 1 1
use contact_28  contact_28_117
timestamp 1643593061
transform 1 0 13680 0 1 34320
box 0 0 1 1
use contact_28  contact_28_118
timestamp 1643593061
transform 1 0 13680 0 1 33960
box 0 0 1 1
use contact_28  contact_28_119
timestamp 1643593061
transform 1 0 13680 0 1 1080
box 0 0 1 1
use contact_28  contact_28_120
timestamp 1643593061
transform 1 0 13680 0 1 1440
box 0 0 1 1
use contact_28  contact_28_121
timestamp 1643593061
transform 1 0 12000 0 1 1080
box 0 0 1 1
use contact_28  contact_28_122
timestamp 1643593061
transform 1 0 12000 0 1 1440
box 0 0 1 1
use contact_28  contact_28_123
timestamp 1643593061
transform 1 0 12000 0 1 34320
box 0 0 1 1
use contact_28  contact_28_124
timestamp 1643593061
transform 1 0 12000 0 1 33960
box 0 0 1 1
use contact_28  contact_28_125
timestamp 1643593061
transform 1 0 12000 0 1 1560
box 0 0 1 1
use contact_28  contact_28_126
timestamp 1643593061
transform 1 0 12000 0 1 3120
box 0 0 1 1
use contact_28  contact_28_127
timestamp 1643593061
transform 1 0 12000 0 1 33840
box 0 0 1 1
use contact_28  contact_28_128
timestamp 1643593061
transform 1 0 12000 0 1 31440
box 0 0 1 1
use contact_28  contact_28_129
timestamp 1643593061
transform 1 0 10560 0 1 31320
box 0 0 1 1
use contact_28  contact_28_130
timestamp 1643593061
transform 1 0 10560 0 1 28440
box 0 0 1 1
use contact_28  contact_28_131
timestamp 1643593061
transform 1 0 10680 0 1 19200
box 0 0 1 1
use contact_28  contact_28_132
timestamp 1643593061
transform 1 0 10680 0 1 22080
box 0 0 1 1
use contact_28  contact_28_133
timestamp 1643593061
transform 1 0 10320 0 1 34320
box 0 0 1 1
use contact_28  contact_28_134
timestamp 1643593061
transform 1 0 10320 0 1 33960
box 0 0 1 1
use contact_28  contact_28_135
timestamp 1643593061
transform 1 0 10320 0 1 1080
box 0 0 1 1
use contact_28  contact_28_136
timestamp 1643593061
transform 1 0 10320 0 1 1440
box 0 0 1 1
use contact_28  contact_28_137
timestamp 1643593061
transform 1 0 10560 0 1 9840
box 0 0 1 1
use contact_28  contact_28_138
timestamp 1643593061
transform 1 0 10560 0 1 9360
box 0 0 1 1
use contact_28  contact_28_139
timestamp 1643593061
transform 1 0 8880 0 1 9360
box 0 0 1 1
use contact_28  contact_28_140
timestamp 1643593061
transform 1 0 8880 0 1 10920
box 0 0 1 1
use contact_28  contact_28_141
timestamp 1643593061
transform 1 0 8760 0 1 14280
box 0 0 1 1
use contact_28  contact_28_142
timestamp 1643593061
transform 1 0 8760 0 1 12720
box 0 0 1 1
use contact_28  contact_28_143
timestamp 1643593061
transform 1 0 8880 0 1 11040
box 0 0 1 1
use contact_28  contact_28_144
timestamp 1643593061
transform 1 0 8880 0 1 12600
box 0 0 1 1
use contact_28  contact_28_145
timestamp 1643593061
transform 1 0 8760 0 1 34320
box 0 0 1 1
use contact_28  contact_28_146
timestamp 1643593061
transform 1 0 8760 0 1 33960
box 0 0 1 1
use contact_28  contact_28_147
timestamp 1643593061
transform 1 0 8760 0 1 1080
box 0 0 1 1
use contact_28  contact_28_148
timestamp 1643593061
transform 1 0 8760 0 1 1440
box 0 0 1 1
use contact_28  contact_28_149
timestamp 1643593061
transform 1 0 7080 0 1 34320
box 0 0 1 1
use contact_28  contact_28_150
timestamp 1643593061
transform 1 0 7080 0 1 33960
box 0 0 1 1
use contact_28  contact_28_151
timestamp 1643593061
transform 1 0 7080 0 1 1080
box 0 0 1 1
use contact_28  contact_28_152
timestamp 1643593061
transform 1 0 7080 0 1 1440
box 0 0 1 1
use contact_28  contact_28_153
timestamp 1643593061
transform 1 0 5280 0 1 34320
box 0 0 1 1
use contact_28  contact_28_154
timestamp 1643593061
transform 1 0 5280 0 1 33960
box 0 0 1 1
use contact_28  contact_28_155
timestamp 1643593061
transform 1 0 5400 0 1 1080
box 0 0 1 1
use contact_28  contact_28_156
timestamp 1643593061
transform 1 0 5400 0 1 1440
box 0 0 1 1
use contact_28  contact_28_157
timestamp 1643593061
transform 1 0 3720 0 1 34320
box 0 0 1 1
use contact_28  contact_28_158
timestamp 1643593061
transform 1 0 3720 0 1 33960
box 0 0 1 1
use contact_28  contact_28_159
timestamp 1643593061
transform 1 0 3720 0 1 1080
box 0 0 1 1
use contact_28  contact_28_160
timestamp 1643593061
transform 1 0 3720 0 1 1440
box 0 0 1 1
use contact_28  contact_28_161
timestamp 1643593061
transform 1 0 1920 0 1 1080
box 0 0 1 1
use contact_28  contact_28_162
timestamp 1643593061
transform 1 0 1920 0 1 1440
box 0 0 1 1
use contact_28  contact_28_163
timestamp 1643593061
transform 1 0 1920 0 1 34320
box 0 0 1 1
use contact_28  contact_28_164
timestamp 1643593061
transform 1 0 1920 0 1 33960
box 0 0 1 1
use contact_28  contact_28_165
timestamp 1643593061
transform 1 0 1080 0 1 25320
box 0 0 1 1
use contact_28  contact_28_166
timestamp 1643593061
transform 1 0 1080 0 1 22080
box 0 0 1 1
use contact_28  contact_28_167
timestamp 1643593061
transform 1 0 1080 0 1 5160
box 0 0 1 1
use contact_28  contact_28_168
timestamp 1643593061
transform 1 0 1080 0 1 27000
box 0 0 1 1
use contact_28  contact_28_169
timestamp 1643593061
transform 1 0 1080 0 1 12000
box 0 0 1 1
use contact_28  contact_28_170
timestamp 1643593061
transform 1 0 1920 0 1 1560
box 0 0 1 1
use contact_28  contact_28_171
timestamp 1643593061
transform 1 0 1920 0 1 1800
box 0 0 1 1
use contact_28  contact_28_172
timestamp 1643593061
transform 1 0 1080 0 1 30480
box 0 0 1 1
use contact_28  contact_28_173
timestamp 1643593061
transform 1 0 1080 0 1 28680
box 0 0 1 1
use contact_28  contact_28_174
timestamp 1643593061
transform 1 0 1080 0 1 3480
box 0 0 1 1
use contact_28  contact_28_175
timestamp 1643593061
transform 1 0 2400 0 1 3240
box 0 0 1 1
use contact_28  contact_28_176
timestamp 1643593061
transform 1 0 2400 0 1 3480
box 0 0 1 1
use contact_28  contact_28_177
timestamp 1643593061
transform 1 0 1080 0 1 8520
box 0 0 1 1
use contact_28  contact_28_178
timestamp 1643593061
transform 1 0 1080 0 1 23760
box 0 0 1 1
use contact_28  contact_28_179
timestamp 1643593061
transform 1 0 1080 0 1 15240
box 0 0 1 1
use contact_28  contact_28_180
timestamp 1643593061
transform 1 0 1080 0 1 13680
box 0 0 1 1
use contact_28  contact_28_181
timestamp 1643593061
transform 1 0 1080 0 1 32160
box 0 0 1 1
use contact_28  contact_28_182
timestamp 1643593061
transform 1 0 1080 0 1 18600
box 0 0 1 1
use contact_28  contact_28_183
timestamp 1643593061
transform 1 0 1080 0 1 16920
box 0 0 1 1
use contact_28  contact_28_184
timestamp 1643593061
transform 1 0 1080 0 1 6840
box 0 0 1 1
use contact_28  contact_28_185
timestamp 1643593061
transform 1 0 1080 0 1 20400
box 0 0 1 1
use contact_28  contact_28_186
timestamp 1643593061
transform 1 0 1080 0 1 10320
box 0 0 1 1
use contact_34  contact_34_0
timestamp 1643593061
transform 1 0 480 0 1 360
box 0 0 1 1
use contact_34  contact_34_1
timestamp 1643593061
transform 1 0 25200 0 1 35040
box 0 0 1 1
use contact_34  contact_34_2
timestamp 1643593061
transform 1 0 360 0 1 35040
box 0 0 1 1
use contact_34  contact_34_3
timestamp 1643593061
transform 1 0 25440 0 1 35040
box 0 0 1 1
use contact_34  contact_34_4
timestamp 1643593061
transform 1 0 240 0 1 35040
box 0 0 1 1
use contact_34  contact_34_5
timestamp 1643593061
transform 1 0 360 0 1 480
box 0 0 1 1
use contact_34  contact_34_6
timestamp 1643593061
transform 1 0 25320 0 1 35040
box 0 0 1 1
use contact_34  contact_34_7
timestamp 1643593061
transform 1 0 25440 0 1 480
box 0 0 1 1
use contact_34  contact_34_8
timestamp 1643593061
transform 1 0 25440 0 1 240
box 0 0 1 1
use contact_34  contact_34_9
timestamp 1643593061
transform 1 0 25200 0 1 480
box 0 0 1 1
use contact_34  contact_34_10
timestamp 1643593061
transform 1 0 240 0 1 480
box 0 0 1 1
use contact_34  contact_34_11
timestamp 1643593061
transform 1 0 25200 0 1 240
box 0 0 1 1
use contact_34  contact_34_12
timestamp 1643593061
transform 1 0 360 0 1 240
box 0 0 1 1
use contact_34  contact_34_13
timestamp 1643593061
transform 1 0 25320 0 1 480
box 0 0 1 1
use contact_34  contact_34_14
timestamp 1643593061
transform 1 0 240 0 1 240
box 0 0 1 1
use contact_34  contact_34_15
timestamp 1643593061
transform 1 0 360 0 1 35160
box 0 0 1 1
use contact_34  contact_34_16
timestamp 1643593061
transform 1 0 25320 0 1 240
box 0 0 1 1
use contact_34  contact_34_17
timestamp 1643593061
transform 1 0 480 0 1 35040
box 0 0 1 1
use contact_34  contact_34_18
timestamp 1643593061
transform 1 0 25440 0 1 35160
box 0 0 1 1
use contact_34  contact_34_19
timestamp 1643593061
transform 1 0 240 0 1 35160
box 0 0 1 1
use contact_34  contact_34_20
timestamp 1643593061
transform 1 0 25440 0 1 34920
box 0 0 1 1
use contact_34  contact_34_21
timestamp 1643593061
transform 1 0 480 0 1 480
box 0 0 1 1
use contact_34  contact_34_22
timestamp 1643593061
transform 1 0 480 0 1 240
box 0 0 1 1
use contact_34  contact_34_23
timestamp 1643593061
transform 1 0 25200 0 1 34920
box 0 0 1 1
use contact_34  contact_34_24
timestamp 1643593061
transform 1 0 360 0 1 34920
box 0 0 1 1
use contact_34  contact_34_25
timestamp 1643593061
transform 1 0 25320 0 1 35160
box 0 0 1 1
use contact_34  contact_34_26
timestamp 1643593061
transform 1 0 240 0 1 34920
box 0 0 1 1
use contact_34  contact_34_27
timestamp 1643593061
transform 1 0 25320 0 1 34920
box 0 0 1 1
use contact_34  contact_34_28
timestamp 1643593061
transform 1 0 25440 0 1 360
box 0 0 1 1
use contact_34  contact_34_29
timestamp 1643593061
transform 1 0 25200 0 1 35160
box 0 0 1 1
use contact_34  contact_34_30
timestamp 1643593061
transform 1 0 480 0 1 35160
box 0 0 1 1
use contact_34  contact_34_31
timestamp 1643593061
transform 1 0 25200 0 1 360
box 0 0 1 1
use contact_34  contact_34_32
timestamp 1643593061
transform 1 0 360 0 1 360
box 0 0 1 1
use contact_34  contact_34_33
timestamp 1643593061
transform 1 0 480 0 1 34920
box 0 0 1 1
use contact_34  contact_34_34
timestamp 1643593061
transform 1 0 240 0 1 360
box 0 0 1 1
use contact_34  contact_34_35
timestamp 1643593061
transform 1 0 25320 0 1 360
box 0 0 1 1
use contact_34  contact_34_36
timestamp 1643593061
transform 1 0 24600 0 1 1080
box 0 0 1 1
use contact_34  contact_34_37
timestamp 1643593061
transform 1 0 960 0 1 840
box 0 0 1 1
use contact_34  contact_34_38
timestamp 1643593061
transform 1 0 840 0 1 34440
box 0 0 1 1
use contact_34  contact_34_39
timestamp 1643593061
transform 1 0 24600 0 1 840
box 0 0 1 1
use contact_34  contact_34_40
timestamp 1643593061
transform 1 0 24720 0 1 1080
box 0 0 1 1
use contact_34  contact_34_41
timestamp 1643593061
transform 1 0 24840 0 1 840
box 0 0 1 1
use contact_34  contact_34_42
timestamp 1643593061
transform 1 0 1080 0 1 840
box 0 0 1 1
use contact_34  contact_34_43
timestamp 1643593061
transform 1 0 24720 0 1 840
box 0 0 1 1
use contact_34  contact_34_44
timestamp 1643593061
transform 1 0 840 0 1 960
box 0 0 1 1
use contact_34  contact_34_45
timestamp 1643593061
transform 1 0 24720 0 1 34320
box 0 0 1 1
use contact_34  contact_34_46
timestamp 1643593061
transform 1 0 24840 0 1 34440
box 0 0 1 1
use contact_34  contact_34_47
timestamp 1643593061
transform 1 0 1080 0 1 34440
box 0 0 1 1
use contact_34  contact_34_48
timestamp 1643593061
transform 1 0 840 0 1 34560
box 0 0 1 1
use contact_34  contact_34_49
timestamp 1643593061
transform 1 0 24720 0 1 34440
box 0 0 1 1
use contact_34  contact_34_50
timestamp 1643593061
transform 1 0 960 0 1 34440
box 0 0 1 1
use contact_34  contact_34_51
timestamp 1643593061
transform 1 0 24600 0 1 34440
box 0 0 1 1
use contact_34  contact_34_52
timestamp 1643593061
transform 1 0 960 0 1 1080
box 0 0 1 1
use contact_34  contact_34_53
timestamp 1643593061
transform 1 0 840 0 1 34320
box 0 0 1 1
use contact_34  contact_34_54
timestamp 1643593061
transform 1 0 24840 0 1 960
box 0 0 1 1
use contact_34  contact_34_55
timestamp 1643593061
transform 1 0 1080 0 1 960
box 0 0 1 1
use contact_34  contact_34_56
timestamp 1643593061
transform 1 0 24720 0 1 960
box 0 0 1 1
use contact_34  contact_34_57
timestamp 1643593061
transform 1 0 840 0 1 1080
box 0 0 1 1
use contact_34  contact_34_58
timestamp 1643593061
transform 1 0 960 0 1 960
box 0 0 1 1
use contact_34  contact_34_59
timestamp 1643593061
transform 1 0 24840 0 1 34320
box 0 0 1 1
use contact_34  contact_34_60
timestamp 1643593061
transform 1 0 24600 0 1 960
box 0 0 1 1
use contact_34  contact_34_61
timestamp 1643593061
transform 1 0 960 0 1 34560
box 0 0 1 1
use contact_34  contact_34_62
timestamp 1643593061
transform 1 0 960 0 1 34320
box 0 0 1 1
use contact_34  contact_34_63
timestamp 1643593061
transform 1 0 840 0 1 840
box 0 0 1 1
use contact_34  contact_34_64
timestamp 1643593061
transform 1 0 24840 0 1 34560
box 0 0 1 1
use contact_34  contact_34_65
timestamp 1643593061
transform 1 0 24600 0 1 34320
box 0 0 1 1
use contact_34  contact_34_66
timestamp 1643593061
transform 1 0 1080 0 1 34560
box 0 0 1 1
use contact_34  contact_34_67
timestamp 1643593061
transform 1 0 24720 0 1 34560
box 0 0 1 1
use contact_34  contact_34_68
timestamp 1643593061
transform 1 0 1080 0 1 34320
box 0 0 1 1
use contact_34  contact_34_69
timestamp 1643593061
transform 1 0 24840 0 1 1080
box 0 0 1 1
use contact_34  contact_34_70
timestamp 1643593061
transform 1 0 1080 0 1 1080
box 0 0 1 1
use contact_34  contact_34_71
timestamp 1643593061
transform 1 0 24600 0 1 34560
box 0 0 1 1
use contact_28  contact_28_187
timestamp 1643593061
transform 1 0 21480 0 1 6600
box 0 0 1 1
use contact_28  contact_28_188
timestamp 1643593061
transform 1 0 21480 0 1 6840
box 0 0 1 1
use contact_28  contact_28_189
timestamp 1643593061
transform 1 0 6240 0 1 3480
box 0 0 1 1
use contact_28  contact_28_190
timestamp 1643593061
transform 1 0 12720 0 1 2520
box 0 0 1 1
use contact_28  contact_28_191
timestamp 1643593061
transform 1 0 11280 0 1 2520
box 0 0 1 1
use contact_32  contact_32_0
timestamp 1643593061
transform 1 0 1522 0 1 33844
box 0 0 192 180
use contact_32  contact_32_1
timestamp 1643593061
transform 1 0 24102 0 1 33844
box 0 0 192 180
use contact_32  contact_32_2
timestamp 1643593061
transform 1 0 24102 0 1 1434
box 0 0 192 180
use contact_32  contact_32_3
timestamp 1643593061
transform 1 0 1522 0 1 1434
box 0 0 192 180
use contact_17  contact_17_0
timestamp 1643593061
transform 1 0 24166 0 1 33418
box 0 0 1 1
use contact_13  contact_13_0
timestamp 1643593061
transform 1 0 24169 0 1 33421
box 0 0 1 1
use contact_21  contact_21_0
timestamp 1643593061
transform 1 0 24173 0 1 33403
box 0 0 1 1
use contact_17  contact_17_1
timestamp 1643593061
transform 1 0 24166 0 1 33082
box 0 0 1 1
use contact_13  contact_13_1
timestamp 1643593061
transform 1 0 24169 0 1 33085
box 0 0 1 1
use contact_21  contact_21_1
timestamp 1643593061
transform 1 0 24173 0 1 33067
box 0 0 1 1
use contact_17  contact_17_2
timestamp 1643593061
transform 1 0 24166 0 1 32746
box 0 0 1 1
use contact_13  contact_13_2
timestamp 1643593061
transform 1 0 24169 0 1 32749
box 0 0 1 1
use contact_21  contact_21_2
timestamp 1643593061
transform 1 0 24173 0 1 32731
box 0 0 1 1
use contact_17  contact_17_3
timestamp 1643593061
transform 1 0 24166 0 1 32410
box 0 0 1 1
use contact_13  contact_13_3
timestamp 1643593061
transform 1 0 24169 0 1 32413
box 0 0 1 1
use contact_21  contact_21_3
timestamp 1643593061
transform 1 0 24173 0 1 32395
box 0 0 1 1
use contact_18  contact_18_0
timestamp 1643593061
transform 1 0 24168 0 1 32070
box 0 0 1 1
use contact_17  contact_17_4
timestamp 1643593061
transform 1 0 24166 0 1 32074
box 0 0 1 1
use contact_13  contact_13_4
timestamp 1643593061
transform 1 0 24169 0 1 32077
box 0 0 1 1
use contact_21  contact_21_4
timestamp 1643593061
transform 1 0 24173 0 1 32059
box 0 0 1 1
use contact_17  contact_17_5
timestamp 1643593061
transform 1 0 24166 0 1 31738
box 0 0 1 1
use contact_13  contact_13_5
timestamp 1643593061
transform 1 0 24169 0 1 31741
box 0 0 1 1
use contact_21  contact_21_5
timestamp 1643593061
transform 1 0 24173 0 1 31723
box 0 0 1 1
use contact_17  contact_17_6
timestamp 1643593061
transform 1 0 24166 0 1 31402
box 0 0 1 1
use contact_13  contact_13_6
timestamp 1643593061
transform 1 0 24169 0 1 31405
box 0 0 1 1
use contact_21  contact_21_6
timestamp 1643593061
transform 1 0 24173 0 1 31387
box 0 0 1 1
use contact_17  contact_17_7
timestamp 1643593061
transform 1 0 24166 0 1 31066
box 0 0 1 1
use contact_13  contact_13_7
timestamp 1643593061
transform 1 0 24169 0 1 31069
box 0 0 1 1
use contact_21  contact_21_7
timestamp 1643593061
transform 1 0 24173 0 1 31051
box 0 0 1 1
use contact_17  contact_17_8
timestamp 1643593061
transform 1 0 24166 0 1 30730
box 0 0 1 1
use contact_13  contact_13_8
timestamp 1643593061
transform 1 0 24169 0 1 30733
box 0 0 1 1
use contact_21  contact_21_8
timestamp 1643593061
transform 1 0 24173 0 1 30715
box 0 0 1 1
use contact_18  contact_18_1
timestamp 1643593061
transform 1 0 24168 0 1 30390
box 0 0 1 1
use contact_17  contact_17_9
timestamp 1643593061
transform 1 0 24166 0 1 30394
box 0 0 1 1
use contact_13  contact_13_9
timestamp 1643593061
transform 1 0 24169 0 1 30397
box 0 0 1 1
use contact_21  contact_21_9
timestamp 1643593061
transform 1 0 24173 0 1 30379
box 0 0 1 1
use contact_17  contact_17_10
timestamp 1643593061
transform 1 0 24166 0 1 30058
box 0 0 1 1
use contact_13  contact_13_10
timestamp 1643593061
transform 1 0 24169 0 1 30061
box 0 0 1 1
use contact_21  contact_21_10
timestamp 1643593061
transform 1 0 24173 0 1 30043
box 0 0 1 1
use contact_17  contact_17_11
timestamp 1643593061
transform 1 0 24166 0 1 29722
box 0 0 1 1
use contact_13  contact_13_11
timestamp 1643593061
transform 1 0 24169 0 1 29725
box 0 0 1 1
use contact_21  contact_21_11
timestamp 1643593061
transform 1 0 24173 0 1 29707
box 0 0 1 1
use contact_17  contact_17_12
timestamp 1643593061
transform 1 0 24166 0 1 29386
box 0 0 1 1
use contact_13  contact_13_12
timestamp 1643593061
transform 1 0 24169 0 1 29389
box 0 0 1 1
use contact_21  contact_21_12
timestamp 1643593061
transform 1 0 24173 0 1 29371
box 0 0 1 1
use contact_17  contact_17_13
timestamp 1643593061
transform 1 0 24166 0 1 29050
box 0 0 1 1
use contact_13  contact_13_13
timestamp 1643593061
transform 1 0 24169 0 1 29053
box 0 0 1 1
use contact_21  contact_21_13
timestamp 1643593061
transform 1 0 24173 0 1 29035
box 0 0 1 1
use contact_18  contact_18_2
timestamp 1643593061
transform 1 0 24168 0 1 28710
box 0 0 1 1
use contact_17  contact_17_14
timestamp 1643593061
transform 1 0 24166 0 1 28714
box 0 0 1 1
use contact_13  contact_13_14
timestamp 1643593061
transform 1 0 24169 0 1 28717
box 0 0 1 1
use contact_21  contact_21_14
timestamp 1643593061
transform 1 0 24173 0 1 28699
box 0 0 1 1
use contact_17  contact_17_15
timestamp 1643593061
transform 1 0 24166 0 1 28378
box 0 0 1 1
use contact_13  contact_13_15
timestamp 1643593061
transform 1 0 24169 0 1 28381
box 0 0 1 1
use contact_21  contact_21_15
timestamp 1643593061
transform 1 0 24173 0 1 28363
box 0 0 1 1
use contact_17  contact_17_16
timestamp 1643593061
transform 1 0 24166 0 1 28042
box 0 0 1 1
use contact_13  contact_13_16
timestamp 1643593061
transform 1 0 24169 0 1 28045
box 0 0 1 1
use contact_21  contact_21_16
timestamp 1643593061
transform 1 0 24173 0 1 28027
box 0 0 1 1
use contact_17  contact_17_17
timestamp 1643593061
transform 1 0 24166 0 1 27706
box 0 0 1 1
use contact_13  contact_13_17
timestamp 1643593061
transform 1 0 24169 0 1 27709
box 0 0 1 1
use contact_21  contact_21_17
timestamp 1643593061
transform 1 0 24173 0 1 27691
box 0 0 1 1
use contact_17  contact_17_18
timestamp 1643593061
transform 1 0 24166 0 1 27370
box 0 0 1 1
use contact_13  contact_13_18
timestamp 1643593061
transform 1 0 24169 0 1 27373
box 0 0 1 1
use contact_21  contact_21_18
timestamp 1643593061
transform 1 0 24173 0 1 27355
box 0 0 1 1
use contact_18  contact_18_3
timestamp 1643593061
transform 1 0 24168 0 1 27030
box 0 0 1 1
use contact_17  contact_17_19
timestamp 1643593061
transform 1 0 24166 0 1 27034
box 0 0 1 1
use contact_13  contact_13_19
timestamp 1643593061
transform 1 0 24169 0 1 27037
box 0 0 1 1
use contact_21  contact_21_19
timestamp 1643593061
transform 1 0 24173 0 1 27019
box 0 0 1 1
use contact_17  contact_17_20
timestamp 1643593061
transform 1 0 24166 0 1 26698
box 0 0 1 1
use contact_13  contact_13_20
timestamp 1643593061
transform 1 0 24169 0 1 26701
box 0 0 1 1
use contact_21  contact_21_20
timestamp 1643593061
transform 1 0 24173 0 1 26683
box 0 0 1 1
use contact_17  contact_17_21
timestamp 1643593061
transform 1 0 24166 0 1 26362
box 0 0 1 1
use contact_13  contact_13_21
timestamp 1643593061
transform 1 0 24169 0 1 26365
box 0 0 1 1
use contact_21  contact_21_21
timestamp 1643593061
transform 1 0 24173 0 1 26347
box 0 0 1 1
use contact_17  contact_17_22
timestamp 1643593061
transform 1 0 24166 0 1 26026
box 0 0 1 1
use contact_13  contact_13_22
timestamp 1643593061
transform 1 0 24169 0 1 26029
box 0 0 1 1
use contact_21  contact_21_22
timestamp 1643593061
transform 1 0 24173 0 1 26011
box 0 0 1 1
use contact_17  contact_17_23
timestamp 1643593061
transform 1 0 24166 0 1 25690
box 0 0 1 1
use contact_13  contact_13_23
timestamp 1643593061
transform 1 0 24169 0 1 25693
box 0 0 1 1
use contact_21  contact_21_23
timestamp 1643593061
transform 1 0 24173 0 1 25675
box 0 0 1 1
use contact_18  contact_18_4
timestamp 1643593061
transform 1 0 24168 0 1 25350
box 0 0 1 1
use contact_17  contact_17_24
timestamp 1643593061
transform 1 0 24166 0 1 25354
box 0 0 1 1
use contact_13  contact_13_24
timestamp 1643593061
transform 1 0 24169 0 1 25357
box 0 0 1 1
use contact_21  contact_21_24
timestamp 1643593061
transform 1 0 24173 0 1 25339
box 0 0 1 1
use contact_17  contact_17_25
timestamp 1643593061
transform 1 0 24166 0 1 25018
box 0 0 1 1
use contact_13  contact_13_25
timestamp 1643593061
transform 1 0 24169 0 1 25021
box 0 0 1 1
use contact_21  contact_21_25
timestamp 1643593061
transform 1 0 24173 0 1 25003
box 0 0 1 1
use contact_17  contact_17_26
timestamp 1643593061
transform 1 0 24166 0 1 24682
box 0 0 1 1
use contact_13  contact_13_26
timestamp 1643593061
transform 1 0 24169 0 1 24685
box 0 0 1 1
use contact_21  contact_21_26
timestamp 1643593061
transform 1 0 24173 0 1 24667
box 0 0 1 1
use contact_17  contact_17_27
timestamp 1643593061
transform 1 0 24166 0 1 24346
box 0 0 1 1
use contact_13  contact_13_27
timestamp 1643593061
transform 1 0 24169 0 1 24349
box 0 0 1 1
use contact_21  contact_21_27
timestamp 1643593061
transform 1 0 24173 0 1 24331
box 0 0 1 1
use contact_17  contact_17_28
timestamp 1643593061
transform 1 0 24166 0 1 24010
box 0 0 1 1
use contact_13  contact_13_28
timestamp 1643593061
transform 1 0 24169 0 1 24013
box 0 0 1 1
use contact_21  contact_21_28
timestamp 1643593061
transform 1 0 24173 0 1 23995
box 0 0 1 1
use contact_18  contact_18_5
timestamp 1643593061
transform 1 0 24168 0 1 23670
box 0 0 1 1
use contact_17  contact_17_29
timestamp 1643593061
transform 1 0 24166 0 1 23674
box 0 0 1 1
use contact_13  contact_13_29
timestamp 1643593061
transform 1 0 24169 0 1 23677
box 0 0 1 1
use contact_21  contact_21_29
timestamp 1643593061
transform 1 0 24173 0 1 23659
box 0 0 1 1
use contact_17  contact_17_30
timestamp 1643593061
transform 1 0 24166 0 1 23338
box 0 0 1 1
use contact_13  contact_13_30
timestamp 1643593061
transform 1 0 24169 0 1 23341
box 0 0 1 1
use contact_21  contact_21_30
timestamp 1643593061
transform 1 0 24173 0 1 23323
box 0 0 1 1
use contact_17  contact_17_31
timestamp 1643593061
transform 1 0 24166 0 1 23002
box 0 0 1 1
use contact_13  contact_13_31
timestamp 1643593061
transform 1 0 24169 0 1 23005
box 0 0 1 1
use contact_21  contact_21_31
timestamp 1643593061
transform 1 0 24173 0 1 22987
box 0 0 1 1
use contact_17  contact_17_32
timestamp 1643593061
transform 1 0 24166 0 1 22666
box 0 0 1 1
use contact_13  contact_13_32
timestamp 1643593061
transform 1 0 24169 0 1 22669
box 0 0 1 1
use contact_21  contact_21_32
timestamp 1643593061
transform 1 0 24173 0 1 22651
box 0 0 1 1
use contact_17  contact_17_33
timestamp 1643593061
transform 1 0 24166 0 1 22330
box 0 0 1 1
use contact_13  contact_13_33
timestamp 1643593061
transform 1 0 24169 0 1 22333
box 0 0 1 1
use contact_21  contact_21_33
timestamp 1643593061
transform 1 0 24173 0 1 22315
box 0 0 1 1
use contact_18  contact_18_6
timestamp 1643593061
transform 1 0 24168 0 1 21990
box 0 0 1 1
use contact_17  contact_17_34
timestamp 1643593061
transform 1 0 24166 0 1 21994
box 0 0 1 1
use contact_13  contact_13_34
timestamp 1643593061
transform 1 0 24169 0 1 21997
box 0 0 1 1
use contact_21  contact_21_34
timestamp 1643593061
transform 1 0 24173 0 1 21979
box 0 0 1 1
use contact_17  contact_17_35
timestamp 1643593061
transform 1 0 24166 0 1 21658
box 0 0 1 1
use contact_13  contact_13_35
timestamp 1643593061
transform 1 0 24169 0 1 21661
box 0 0 1 1
use contact_21  contact_21_35
timestamp 1643593061
transform 1 0 24173 0 1 21643
box 0 0 1 1
use contact_17  contact_17_36
timestamp 1643593061
transform 1 0 24166 0 1 21322
box 0 0 1 1
use contact_13  contact_13_36
timestamp 1643593061
transform 1 0 24169 0 1 21325
box 0 0 1 1
use contact_21  contact_21_36
timestamp 1643593061
transform 1 0 24173 0 1 21307
box 0 0 1 1
use contact_17  contact_17_37
timestamp 1643593061
transform 1 0 24166 0 1 20986
box 0 0 1 1
use contact_13  contact_13_37
timestamp 1643593061
transform 1 0 24169 0 1 20989
box 0 0 1 1
use contact_21  contact_21_37
timestamp 1643593061
transform 1 0 24173 0 1 20971
box 0 0 1 1
use contact_17  contact_17_38
timestamp 1643593061
transform 1 0 24166 0 1 20650
box 0 0 1 1
use contact_13  contact_13_38
timestamp 1643593061
transform 1 0 24169 0 1 20653
box 0 0 1 1
use contact_21  contact_21_38
timestamp 1643593061
transform 1 0 24173 0 1 20635
box 0 0 1 1
use contact_18  contact_18_7
timestamp 1643593061
transform 1 0 24168 0 1 20310
box 0 0 1 1
use contact_17  contact_17_39
timestamp 1643593061
transform 1 0 24166 0 1 20314
box 0 0 1 1
use contact_13  contact_13_39
timestamp 1643593061
transform 1 0 24169 0 1 20317
box 0 0 1 1
use contact_21  contact_21_39
timestamp 1643593061
transform 1 0 24173 0 1 20299
box 0 0 1 1
use contact_17  contact_17_40
timestamp 1643593061
transform 1 0 24166 0 1 19978
box 0 0 1 1
use contact_13  contact_13_40
timestamp 1643593061
transform 1 0 24169 0 1 19981
box 0 0 1 1
use contact_21  contact_21_40
timestamp 1643593061
transform 1 0 24173 0 1 19963
box 0 0 1 1
use contact_17  contact_17_41
timestamp 1643593061
transform 1 0 24166 0 1 19642
box 0 0 1 1
use contact_13  contact_13_41
timestamp 1643593061
transform 1 0 24169 0 1 19645
box 0 0 1 1
use contact_21  contact_21_41
timestamp 1643593061
transform 1 0 24173 0 1 19627
box 0 0 1 1
use contact_17  contact_17_42
timestamp 1643593061
transform 1 0 24166 0 1 19306
box 0 0 1 1
use contact_13  contact_13_42
timestamp 1643593061
transform 1 0 24169 0 1 19309
box 0 0 1 1
use contact_21  contact_21_42
timestamp 1643593061
transform 1 0 24173 0 1 19291
box 0 0 1 1
use contact_17  contact_17_43
timestamp 1643593061
transform 1 0 24166 0 1 18970
box 0 0 1 1
use contact_13  contact_13_43
timestamp 1643593061
transform 1 0 24169 0 1 18973
box 0 0 1 1
use contact_21  contact_21_43
timestamp 1643593061
transform 1 0 24173 0 1 18955
box 0 0 1 1
use contact_18  contact_18_8
timestamp 1643593061
transform 1 0 24168 0 1 18630
box 0 0 1 1
use contact_17  contact_17_44
timestamp 1643593061
transform 1 0 24166 0 1 18634
box 0 0 1 1
use contact_13  contact_13_44
timestamp 1643593061
transform 1 0 24169 0 1 18637
box 0 0 1 1
use contact_21  contact_21_44
timestamp 1643593061
transform 1 0 24173 0 1 18619
box 0 0 1 1
use contact_17  contact_17_45
timestamp 1643593061
transform 1 0 24166 0 1 18298
box 0 0 1 1
use contact_13  contact_13_45
timestamp 1643593061
transform 1 0 24169 0 1 18301
box 0 0 1 1
use contact_21  contact_21_45
timestamp 1643593061
transform 1 0 24173 0 1 18283
box 0 0 1 1
use contact_17  contact_17_46
timestamp 1643593061
transform 1 0 24166 0 1 17962
box 0 0 1 1
use contact_13  contact_13_46
timestamp 1643593061
transform 1 0 24169 0 1 17965
box 0 0 1 1
use contact_21  contact_21_46
timestamp 1643593061
transform 1 0 24173 0 1 17947
box 0 0 1 1
use contact_17  contact_17_47
timestamp 1643593061
transform 1 0 24166 0 1 17626
box 0 0 1 1
use contact_13  contact_13_47
timestamp 1643593061
transform 1 0 24169 0 1 17629
box 0 0 1 1
use contact_21  contact_21_47
timestamp 1643593061
transform 1 0 24173 0 1 17611
box 0 0 1 1
use contact_17  contact_17_48
timestamp 1643593061
transform 1 0 24166 0 1 17290
box 0 0 1 1
use contact_13  contact_13_48
timestamp 1643593061
transform 1 0 24169 0 1 17293
box 0 0 1 1
use contact_21  contact_21_48
timestamp 1643593061
transform 1 0 24173 0 1 17275
box 0 0 1 1
use contact_18  contact_18_9
timestamp 1643593061
transform 1 0 24168 0 1 16950
box 0 0 1 1
use contact_17  contact_17_49
timestamp 1643593061
transform 1 0 24166 0 1 16954
box 0 0 1 1
use contact_13  contact_13_49
timestamp 1643593061
transform 1 0 24169 0 1 16957
box 0 0 1 1
use contact_21  contact_21_49
timestamp 1643593061
transform 1 0 24173 0 1 16939
box 0 0 1 1
use contact_17  contact_17_50
timestamp 1643593061
transform 1 0 24166 0 1 16618
box 0 0 1 1
use contact_13  contact_13_50
timestamp 1643593061
transform 1 0 24169 0 1 16621
box 0 0 1 1
use contact_21  contact_21_50
timestamp 1643593061
transform 1 0 24173 0 1 16603
box 0 0 1 1
use contact_17  contact_17_51
timestamp 1643593061
transform 1 0 24166 0 1 16282
box 0 0 1 1
use contact_13  contact_13_51
timestamp 1643593061
transform 1 0 24169 0 1 16285
box 0 0 1 1
use contact_21  contact_21_51
timestamp 1643593061
transform 1 0 24173 0 1 16267
box 0 0 1 1
use contact_17  contact_17_52
timestamp 1643593061
transform 1 0 24166 0 1 15946
box 0 0 1 1
use contact_13  contact_13_52
timestamp 1643593061
transform 1 0 24169 0 1 15949
box 0 0 1 1
use contact_21  contact_21_52
timestamp 1643593061
transform 1 0 24173 0 1 15931
box 0 0 1 1
use contact_17  contact_17_53
timestamp 1643593061
transform 1 0 24166 0 1 15610
box 0 0 1 1
use contact_13  contact_13_53
timestamp 1643593061
transform 1 0 24169 0 1 15613
box 0 0 1 1
use contact_21  contact_21_53
timestamp 1643593061
transform 1 0 24173 0 1 15595
box 0 0 1 1
use contact_18  contact_18_10
timestamp 1643593061
transform 1 0 24168 0 1 15270
box 0 0 1 1
use contact_17  contact_17_54
timestamp 1643593061
transform 1 0 24166 0 1 15274
box 0 0 1 1
use contact_13  contact_13_54
timestamp 1643593061
transform 1 0 24169 0 1 15277
box 0 0 1 1
use contact_21  contact_21_54
timestamp 1643593061
transform 1 0 24173 0 1 15259
box 0 0 1 1
use contact_17  contact_17_55
timestamp 1643593061
transform 1 0 24166 0 1 14938
box 0 0 1 1
use contact_13  contact_13_55
timestamp 1643593061
transform 1 0 24169 0 1 14941
box 0 0 1 1
use contact_21  contact_21_55
timestamp 1643593061
transform 1 0 24173 0 1 14923
box 0 0 1 1
use contact_17  contact_17_56
timestamp 1643593061
transform 1 0 24166 0 1 14602
box 0 0 1 1
use contact_13  contact_13_56
timestamp 1643593061
transform 1 0 24169 0 1 14605
box 0 0 1 1
use contact_21  contact_21_56
timestamp 1643593061
transform 1 0 24173 0 1 14587
box 0 0 1 1
use contact_17  contact_17_57
timestamp 1643593061
transform 1 0 24166 0 1 14266
box 0 0 1 1
use contact_13  contact_13_57
timestamp 1643593061
transform 1 0 24169 0 1 14269
box 0 0 1 1
use contact_21  contact_21_57
timestamp 1643593061
transform 1 0 24173 0 1 14251
box 0 0 1 1
use contact_17  contact_17_58
timestamp 1643593061
transform 1 0 24166 0 1 13930
box 0 0 1 1
use contact_13  contact_13_58
timestamp 1643593061
transform 1 0 24169 0 1 13933
box 0 0 1 1
use contact_21  contact_21_58
timestamp 1643593061
transform 1 0 24173 0 1 13915
box 0 0 1 1
use contact_18  contact_18_11
timestamp 1643593061
transform 1 0 24168 0 1 13590
box 0 0 1 1
use contact_17  contact_17_59
timestamp 1643593061
transform 1 0 24166 0 1 13594
box 0 0 1 1
use contact_13  contact_13_59
timestamp 1643593061
transform 1 0 24169 0 1 13597
box 0 0 1 1
use contact_21  contact_21_59
timestamp 1643593061
transform 1 0 24173 0 1 13579
box 0 0 1 1
use contact_17  contact_17_60
timestamp 1643593061
transform 1 0 24166 0 1 13258
box 0 0 1 1
use contact_13  contact_13_60
timestamp 1643593061
transform 1 0 24169 0 1 13261
box 0 0 1 1
use contact_21  contact_21_60
timestamp 1643593061
transform 1 0 24173 0 1 13243
box 0 0 1 1
use contact_17  contact_17_61
timestamp 1643593061
transform 1 0 24166 0 1 12922
box 0 0 1 1
use contact_13  contact_13_61
timestamp 1643593061
transform 1 0 24169 0 1 12925
box 0 0 1 1
use contact_21  contact_21_61
timestamp 1643593061
transform 1 0 24173 0 1 12907
box 0 0 1 1
use contact_17  contact_17_62
timestamp 1643593061
transform 1 0 24166 0 1 12586
box 0 0 1 1
use contact_13  contact_13_62
timestamp 1643593061
transform 1 0 24169 0 1 12589
box 0 0 1 1
use contact_21  contact_21_62
timestamp 1643593061
transform 1 0 24173 0 1 12571
box 0 0 1 1
use contact_17  contact_17_63
timestamp 1643593061
transform 1 0 24166 0 1 12250
box 0 0 1 1
use contact_13  contact_13_63
timestamp 1643593061
transform 1 0 24169 0 1 12253
box 0 0 1 1
use contact_21  contact_21_63
timestamp 1643593061
transform 1 0 24173 0 1 12235
box 0 0 1 1
use contact_18  contact_18_12
timestamp 1643593061
transform 1 0 24168 0 1 11910
box 0 0 1 1
use contact_17  contact_17_64
timestamp 1643593061
transform 1 0 24166 0 1 11914
box 0 0 1 1
use contact_13  contact_13_64
timestamp 1643593061
transform 1 0 24169 0 1 11917
box 0 0 1 1
use contact_21  contact_21_64
timestamp 1643593061
transform 1 0 24173 0 1 11899
box 0 0 1 1
use contact_17  contact_17_65
timestamp 1643593061
transform 1 0 24166 0 1 11578
box 0 0 1 1
use contact_13  contact_13_65
timestamp 1643593061
transform 1 0 24169 0 1 11581
box 0 0 1 1
use contact_21  contact_21_65
timestamp 1643593061
transform 1 0 24173 0 1 11563
box 0 0 1 1
use contact_17  contact_17_66
timestamp 1643593061
transform 1 0 24166 0 1 11242
box 0 0 1 1
use contact_13  contact_13_66
timestamp 1643593061
transform 1 0 24169 0 1 11245
box 0 0 1 1
use contact_21  contact_21_66
timestamp 1643593061
transform 1 0 24173 0 1 11227
box 0 0 1 1
use contact_17  contact_17_67
timestamp 1643593061
transform 1 0 24166 0 1 10906
box 0 0 1 1
use contact_13  contact_13_67
timestamp 1643593061
transform 1 0 24169 0 1 10909
box 0 0 1 1
use contact_21  contact_21_67
timestamp 1643593061
transform 1 0 24173 0 1 10891
box 0 0 1 1
use contact_17  contact_17_68
timestamp 1643593061
transform 1 0 24166 0 1 10570
box 0 0 1 1
use contact_13  contact_13_68
timestamp 1643593061
transform 1 0 24169 0 1 10573
box 0 0 1 1
use contact_21  contact_21_68
timestamp 1643593061
transform 1 0 24173 0 1 10555
box 0 0 1 1
use contact_18  contact_18_13
timestamp 1643593061
transform 1 0 24168 0 1 10230
box 0 0 1 1
use contact_17  contact_17_69
timestamp 1643593061
transform 1 0 24166 0 1 10234
box 0 0 1 1
use contact_13  contact_13_69
timestamp 1643593061
transform 1 0 24169 0 1 10237
box 0 0 1 1
use contact_21  contact_21_69
timestamp 1643593061
transform 1 0 24173 0 1 10219
box 0 0 1 1
use contact_17  contact_17_70
timestamp 1643593061
transform 1 0 24166 0 1 9898
box 0 0 1 1
use contact_13  contact_13_70
timestamp 1643593061
transform 1 0 24169 0 1 9901
box 0 0 1 1
use contact_21  contact_21_70
timestamp 1643593061
transform 1 0 24173 0 1 9883
box 0 0 1 1
use contact_17  contact_17_71
timestamp 1643593061
transform 1 0 24166 0 1 9562
box 0 0 1 1
use contact_13  contact_13_71
timestamp 1643593061
transform 1 0 24169 0 1 9565
box 0 0 1 1
use contact_21  contact_21_71
timestamp 1643593061
transform 1 0 24173 0 1 9547
box 0 0 1 1
use contact_17  contact_17_72
timestamp 1643593061
transform 1 0 24166 0 1 9226
box 0 0 1 1
use contact_13  contact_13_72
timestamp 1643593061
transform 1 0 24169 0 1 9229
box 0 0 1 1
use contact_21  contact_21_72
timestamp 1643593061
transform 1 0 24173 0 1 9211
box 0 0 1 1
use contact_17  contact_17_73
timestamp 1643593061
transform 1 0 24166 0 1 8890
box 0 0 1 1
use contact_13  contact_13_73
timestamp 1643593061
transform 1 0 24169 0 1 8893
box 0 0 1 1
use contact_21  contact_21_73
timestamp 1643593061
transform 1 0 24173 0 1 8875
box 0 0 1 1
use contact_18  contact_18_14
timestamp 1643593061
transform 1 0 24168 0 1 8550
box 0 0 1 1
use contact_17  contact_17_74
timestamp 1643593061
transform 1 0 24166 0 1 8554
box 0 0 1 1
use contact_13  contact_13_74
timestamp 1643593061
transform 1 0 24169 0 1 8557
box 0 0 1 1
use contact_21  contact_21_74
timestamp 1643593061
transform 1 0 24173 0 1 8539
box 0 0 1 1
use contact_17  contact_17_75
timestamp 1643593061
transform 1 0 24166 0 1 8218
box 0 0 1 1
use contact_13  contact_13_75
timestamp 1643593061
transform 1 0 24169 0 1 8221
box 0 0 1 1
use contact_21  contact_21_75
timestamp 1643593061
transform 1 0 24173 0 1 8203
box 0 0 1 1
use contact_17  contact_17_76
timestamp 1643593061
transform 1 0 24166 0 1 7882
box 0 0 1 1
use contact_13  contact_13_76
timestamp 1643593061
transform 1 0 24169 0 1 7885
box 0 0 1 1
use contact_21  contact_21_76
timestamp 1643593061
transform 1 0 24173 0 1 7867
box 0 0 1 1
use contact_17  contact_17_77
timestamp 1643593061
transform 1 0 24166 0 1 7546
box 0 0 1 1
use contact_13  contact_13_77
timestamp 1643593061
transform 1 0 24169 0 1 7549
box 0 0 1 1
use contact_21  contact_21_77
timestamp 1643593061
transform 1 0 24173 0 1 7531
box 0 0 1 1
use contact_17  contact_17_78
timestamp 1643593061
transform 1 0 24166 0 1 7210
box 0 0 1 1
use contact_13  contact_13_78
timestamp 1643593061
transform 1 0 24169 0 1 7213
box 0 0 1 1
use contact_21  contact_21_78
timestamp 1643593061
transform 1 0 24173 0 1 7195
box 0 0 1 1
use contact_18  contact_18_15
timestamp 1643593061
transform 1 0 24168 0 1 6870
box 0 0 1 1
use contact_17  contact_17_79
timestamp 1643593061
transform 1 0 24166 0 1 6874
box 0 0 1 1
use contact_13  contact_13_79
timestamp 1643593061
transform 1 0 24169 0 1 6877
box 0 0 1 1
use contact_21  contact_21_79
timestamp 1643593061
transform 1 0 24173 0 1 6859
box 0 0 1 1
use contact_17  contact_17_80
timestamp 1643593061
transform 1 0 24166 0 1 6538
box 0 0 1 1
use contact_13  contact_13_80
timestamp 1643593061
transform 1 0 24169 0 1 6541
box 0 0 1 1
use contact_21  contact_21_80
timestamp 1643593061
transform 1 0 24173 0 1 6523
box 0 0 1 1
use contact_17  contact_17_81
timestamp 1643593061
transform 1 0 24166 0 1 6202
box 0 0 1 1
use contact_13  contact_13_81
timestamp 1643593061
transform 1 0 24169 0 1 6205
box 0 0 1 1
use contact_21  contact_21_81
timestamp 1643593061
transform 1 0 24173 0 1 6187
box 0 0 1 1
use contact_17  contact_17_82
timestamp 1643593061
transform 1 0 24166 0 1 5866
box 0 0 1 1
use contact_13  contact_13_82
timestamp 1643593061
transform 1 0 24169 0 1 5869
box 0 0 1 1
use contact_21  contact_21_82
timestamp 1643593061
transform 1 0 24173 0 1 5851
box 0 0 1 1
use contact_17  contact_17_83
timestamp 1643593061
transform 1 0 24166 0 1 5530
box 0 0 1 1
use contact_13  contact_13_83
timestamp 1643593061
transform 1 0 24169 0 1 5533
box 0 0 1 1
use contact_21  contact_21_83
timestamp 1643593061
transform 1 0 24173 0 1 5515
box 0 0 1 1
use contact_18  contact_18_16
timestamp 1643593061
transform 1 0 24168 0 1 5190
box 0 0 1 1
use contact_17  contact_17_84
timestamp 1643593061
transform 1 0 24166 0 1 5194
box 0 0 1 1
use contact_13  contact_13_84
timestamp 1643593061
transform 1 0 24169 0 1 5197
box 0 0 1 1
use contact_21  contact_21_84
timestamp 1643593061
transform 1 0 24173 0 1 5179
box 0 0 1 1
use contact_17  contact_17_85
timestamp 1643593061
transform 1 0 24166 0 1 4858
box 0 0 1 1
use contact_13  contact_13_85
timestamp 1643593061
transform 1 0 24169 0 1 4861
box 0 0 1 1
use contact_21  contact_21_85
timestamp 1643593061
transform 1 0 24173 0 1 4843
box 0 0 1 1
use contact_17  contact_17_86
timestamp 1643593061
transform 1 0 24166 0 1 4522
box 0 0 1 1
use contact_13  contact_13_86
timestamp 1643593061
transform 1 0 24169 0 1 4525
box 0 0 1 1
use contact_21  contact_21_86
timestamp 1643593061
transform 1 0 24173 0 1 4507
box 0 0 1 1
use contact_17  contact_17_87
timestamp 1643593061
transform 1 0 24166 0 1 4186
box 0 0 1 1
use contact_13  contact_13_87
timestamp 1643593061
transform 1 0 24169 0 1 4189
box 0 0 1 1
use contact_21  contact_21_87
timestamp 1643593061
transform 1 0 24173 0 1 4171
box 0 0 1 1
use contact_17  contact_17_88
timestamp 1643593061
transform 1 0 24166 0 1 3850
box 0 0 1 1
use contact_13  contact_13_88
timestamp 1643593061
transform 1 0 24169 0 1 3853
box 0 0 1 1
use contact_21  contact_21_88
timestamp 1643593061
transform 1 0 24173 0 1 3835
box 0 0 1 1
use contact_18  contact_18_17
timestamp 1643593061
transform 1 0 24168 0 1 3510
box 0 0 1 1
use contact_17  contact_17_89
timestamp 1643593061
transform 1 0 24166 0 1 3514
box 0 0 1 1
use contact_13  contact_13_89
timestamp 1643593061
transform 1 0 24169 0 1 3517
box 0 0 1 1
use contact_21  contact_21_89
timestamp 1643593061
transform 1 0 24173 0 1 3499
box 0 0 1 1
use contact_17  contact_17_90
timestamp 1643593061
transform 1 0 24166 0 1 3178
box 0 0 1 1
use contact_13  contact_13_90
timestamp 1643593061
transform 1 0 24169 0 1 3181
box 0 0 1 1
use contact_21  contact_21_90
timestamp 1643593061
transform 1 0 24173 0 1 3163
box 0 0 1 1
use contact_17  contact_17_91
timestamp 1643593061
transform 1 0 24166 0 1 2842
box 0 0 1 1
use contact_13  contact_13_91
timestamp 1643593061
transform 1 0 24169 0 1 2845
box 0 0 1 1
use contact_21  contact_21_91
timestamp 1643593061
transform 1 0 24173 0 1 2827
box 0 0 1 1
use contact_17  contact_17_92
timestamp 1643593061
transform 1 0 24166 0 1 2506
box 0 0 1 1
use contact_13  contact_13_92
timestamp 1643593061
transform 1 0 24169 0 1 2509
box 0 0 1 1
use contact_21  contact_21_92
timestamp 1643593061
transform 1 0 24173 0 1 2491
box 0 0 1 1
use contact_17  contact_17_93
timestamp 1643593061
transform 1 0 24166 0 1 2170
box 0 0 1 1
use contact_13  contact_13_93
timestamp 1643593061
transform 1 0 24169 0 1 2173
box 0 0 1 1
use contact_21  contact_21_93
timestamp 1643593061
transform 1 0 24173 0 1 2155
box 0 0 1 1
use contact_18  contact_18_18
timestamp 1643593061
transform 1 0 24168 0 1 1830
box 0 0 1 1
use contact_17  contact_17_94
timestamp 1643593061
transform 1 0 24166 0 1 1834
box 0 0 1 1
use contact_13  contact_13_94
timestamp 1643593061
transform 1 0 24169 0 1 1837
box 0 0 1 1
use contact_21  contact_21_94
timestamp 1643593061
transform 1 0 24173 0 1 1819
box 0 0 1 1
use contact_17  contact_17_95
timestamp 1643593061
transform 1 0 1586 0 1 33418
box 0 0 1 1
use contact_13  contact_13_95
timestamp 1643593061
transform 1 0 1589 0 1 33421
box 0 0 1 1
use contact_21  contact_21_95
timestamp 1643593061
transform 1 0 1593 0 1 33403
box 0 0 1 1
use contact_17  contact_17_96
timestamp 1643593061
transform 1 0 1586 0 1 33082
box 0 0 1 1
use contact_13  contact_13_96
timestamp 1643593061
transform 1 0 1589 0 1 33085
box 0 0 1 1
use contact_21  contact_21_96
timestamp 1643593061
transform 1 0 1593 0 1 33067
box 0 0 1 1
use contact_17  contact_17_97
timestamp 1643593061
transform 1 0 1586 0 1 32746
box 0 0 1 1
use contact_13  contact_13_97
timestamp 1643593061
transform 1 0 1589 0 1 32749
box 0 0 1 1
use contact_21  contact_21_97
timestamp 1643593061
transform 1 0 1593 0 1 32731
box 0 0 1 1
use contact_17  contact_17_98
timestamp 1643593061
transform 1 0 1586 0 1 32410
box 0 0 1 1
use contact_13  contact_13_98
timestamp 1643593061
transform 1 0 1589 0 1 32413
box 0 0 1 1
use contact_21  contact_21_98
timestamp 1643593061
transform 1 0 1593 0 1 32395
box 0 0 1 1
use contact_18  contact_18_19
timestamp 1643593061
transform 1 0 1588 0 1 32070
box 0 0 1 1
use contact_17  contact_17_99
timestamp 1643593061
transform 1 0 1586 0 1 32074
box 0 0 1 1
use contact_13  contact_13_99
timestamp 1643593061
transform 1 0 1589 0 1 32077
box 0 0 1 1
use contact_21  contact_21_99
timestamp 1643593061
transform 1 0 1593 0 1 32059
box 0 0 1 1
use contact_17  contact_17_100
timestamp 1643593061
transform 1 0 1586 0 1 31738
box 0 0 1 1
use contact_13  contact_13_100
timestamp 1643593061
transform 1 0 1589 0 1 31741
box 0 0 1 1
use contact_21  contact_21_100
timestamp 1643593061
transform 1 0 1593 0 1 31723
box 0 0 1 1
use contact_17  contact_17_101
timestamp 1643593061
transform 1 0 1586 0 1 31402
box 0 0 1 1
use contact_13  contact_13_101
timestamp 1643593061
transform 1 0 1589 0 1 31405
box 0 0 1 1
use contact_21  contact_21_101
timestamp 1643593061
transform 1 0 1593 0 1 31387
box 0 0 1 1
use contact_17  contact_17_102
timestamp 1643593061
transform 1 0 1586 0 1 31066
box 0 0 1 1
use contact_13  contact_13_102
timestamp 1643593061
transform 1 0 1589 0 1 31069
box 0 0 1 1
use contact_21  contact_21_102
timestamp 1643593061
transform 1 0 1593 0 1 31051
box 0 0 1 1
use contact_17  contact_17_103
timestamp 1643593061
transform 1 0 1586 0 1 30730
box 0 0 1 1
use contact_13  contact_13_103
timestamp 1643593061
transform 1 0 1589 0 1 30733
box 0 0 1 1
use contact_21  contact_21_103
timestamp 1643593061
transform 1 0 1593 0 1 30715
box 0 0 1 1
use contact_18  contact_18_20
timestamp 1643593061
transform 1 0 1588 0 1 30390
box 0 0 1 1
use contact_17  contact_17_104
timestamp 1643593061
transform 1 0 1586 0 1 30394
box 0 0 1 1
use contact_13  contact_13_104
timestamp 1643593061
transform 1 0 1589 0 1 30397
box 0 0 1 1
use contact_21  contact_21_104
timestamp 1643593061
transform 1 0 1593 0 1 30379
box 0 0 1 1
use contact_17  contact_17_105
timestamp 1643593061
transform 1 0 1586 0 1 30058
box 0 0 1 1
use contact_13  contact_13_105
timestamp 1643593061
transform 1 0 1589 0 1 30061
box 0 0 1 1
use contact_21  contact_21_105
timestamp 1643593061
transform 1 0 1593 0 1 30043
box 0 0 1 1
use contact_17  contact_17_106
timestamp 1643593061
transform 1 0 1586 0 1 29722
box 0 0 1 1
use contact_13  contact_13_106
timestamp 1643593061
transform 1 0 1589 0 1 29725
box 0 0 1 1
use contact_21  contact_21_106
timestamp 1643593061
transform 1 0 1593 0 1 29707
box 0 0 1 1
use contact_17  contact_17_107
timestamp 1643593061
transform 1 0 1586 0 1 29386
box 0 0 1 1
use contact_13  contact_13_107
timestamp 1643593061
transform 1 0 1589 0 1 29389
box 0 0 1 1
use contact_21  contact_21_107
timestamp 1643593061
transform 1 0 1593 0 1 29371
box 0 0 1 1
use contact_17  contact_17_108
timestamp 1643593061
transform 1 0 1586 0 1 29050
box 0 0 1 1
use contact_13  contact_13_108
timestamp 1643593061
transform 1 0 1589 0 1 29053
box 0 0 1 1
use contact_21  contact_21_108
timestamp 1643593061
transform 1 0 1593 0 1 29035
box 0 0 1 1
use contact_18  contact_18_21
timestamp 1643593061
transform 1 0 1588 0 1 28710
box 0 0 1 1
use contact_17  contact_17_109
timestamp 1643593061
transform 1 0 1586 0 1 28714
box 0 0 1 1
use contact_13  contact_13_109
timestamp 1643593061
transform 1 0 1589 0 1 28717
box 0 0 1 1
use contact_21  contact_21_109
timestamp 1643593061
transform 1 0 1593 0 1 28699
box 0 0 1 1
use contact_17  contact_17_110
timestamp 1643593061
transform 1 0 1586 0 1 28378
box 0 0 1 1
use contact_13  contact_13_110
timestamp 1643593061
transform 1 0 1589 0 1 28381
box 0 0 1 1
use contact_21  contact_21_110
timestamp 1643593061
transform 1 0 1593 0 1 28363
box 0 0 1 1
use contact_17  contact_17_111
timestamp 1643593061
transform 1 0 1586 0 1 28042
box 0 0 1 1
use contact_13  contact_13_111
timestamp 1643593061
transform 1 0 1589 0 1 28045
box 0 0 1 1
use contact_21  contact_21_111
timestamp 1643593061
transform 1 0 1593 0 1 28027
box 0 0 1 1
use contact_17  contact_17_112
timestamp 1643593061
transform 1 0 1586 0 1 27706
box 0 0 1 1
use contact_13  contact_13_112
timestamp 1643593061
transform 1 0 1589 0 1 27709
box 0 0 1 1
use contact_21  contact_21_112
timestamp 1643593061
transform 1 0 1593 0 1 27691
box 0 0 1 1
use contact_17  contact_17_113
timestamp 1643593061
transform 1 0 1586 0 1 27370
box 0 0 1 1
use contact_13  contact_13_113
timestamp 1643593061
transform 1 0 1589 0 1 27373
box 0 0 1 1
use contact_21  contact_21_113
timestamp 1643593061
transform 1 0 1593 0 1 27355
box 0 0 1 1
use contact_18  contact_18_22
timestamp 1643593061
transform 1 0 1588 0 1 27030
box 0 0 1 1
use contact_17  contact_17_114
timestamp 1643593061
transform 1 0 1586 0 1 27034
box 0 0 1 1
use contact_13  contact_13_114
timestamp 1643593061
transform 1 0 1589 0 1 27037
box 0 0 1 1
use contact_21  contact_21_114
timestamp 1643593061
transform 1 0 1593 0 1 27019
box 0 0 1 1
use contact_17  contact_17_115
timestamp 1643593061
transform 1 0 1586 0 1 26698
box 0 0 1 1
use contact_13  contact_13_115
timestamp 1643593061
transform 1 0 1589 0 1 26701
box 0 0 1 1
use contact_21  contact_21_115
timestamp 1643593061
transform 1 0 1593 0 1 26683
box 0 0 1 1
use contact_17  contact_17_116
timestamp 1643593061
transform 1 0 1586 0 1 26362
box 0 0 1 1
use contact_13  contact_13_116
timestamp 1643593061
transform 1 0 1589 0 1 26365
box 0 0 1 1
use contact_21  contact_21_116
timestamp 1643593061
transform 1 0 1593 0 1 26347
box 0 0 1 1
use contact_17  contact_17_117
timestamp 1643593061
transform 1 0 1586 0 1 26026
box 0 0 1 1
use contact_13  contact_13_117
timestamp 1643593061
transform 1 0 1589 0 1 26029
box 0 0 1 1
use contact_21  contact_21_117
timestamp 1643593061
transform 1 0 1593 0 1 26011
box 0 0 1 1
use contact_17  contact_17_118
timestamp 1643593061
transform 1 0 1586 0 1 25690
box 0 0 1 1
use contact_13  contact_13_118
timestamp 1643593061
transform 1 0 1589 0 1 25693
box 0 0 1 1
use contact_21  contact_21_118
timestamp 1643593061
transform 1 0 1593 0 1 25675
box 0 0 1 1
use contact_18  contact_18_23
timestamp 1643593061
transform 1 0 1588 0 1 25350
box 0 0 1 1
use contact_17  contact_17_119
timestamp 1643593061
transform 1 0 1586 0 1 25354
box 0 0 1 1
use contact_13  contact_13_119
timestamp 1643593061
transform 1 0 1589 0 1 25357
box 0 0 1 1
use contact_21  contact_21_119
timestamp 1643593061
transform 1 0 1593 0 1 25339
box 0 0 1 1
use contact_17  contact_17_120
timestamp 1643593061
transform 1 0 1586 0 1 25018
box 0 0 1 1
use contact_13  contact_13_120
timestamp 1643593061
transform 1 0 1589 0 1 25021
box 0 0 1 1
use contact_21  contact_21_120
timestamp 1643593061
transform 1 0 1593 0 1 25003
box 0 0 1 1
use contact_17  contact_17_121
timestamp 1643593061
transform 1 0 1586 0 1 24682
box 0 0 1 1
use contact_13  contact_13_121
timestamp 1643593061
transform 1 0 1589 0 1 24685
box 0 0 1 1
use contact_21  contact_21_121
timestamp 1643593061
transform 1 0 1593 0 1 24667
box 0 0 1 1
use contact_17  contact_17_122
timestamp 1643593061
transform 1 0 1586 0 1 24346
box 0 0 1 1
use contact_13  contact_13_122
timestamp 1643593061
transform 1 0 1589 0 1 24349
box 0 0 1 1
use contact_21  contact_21_122
timestamp 1643593061
transform 1 0 1593 0 1 24331
box 0 0 1 1
use contact_17  contact_17_123
timestamp 1643593061
transform 1 0 1586 0 1 24010
box 0 0 1 1
use contact_13  contact_13_123
timestamp 1643593061
transform 1 0 1589 0 1 24013
box 0 0 1 1
use contact_21  contact_21_123
timestamp 1643593061
transform 1 0 1593 0 1 23995
box 0 0 1 1
use contact_18  contact_18_24
timestamp 1643593061
transform 1 0 1588 0 1 23670
box 0 0 1 1
use contact_17  contact_17_124
timestamp 1643593061
transform 1 0 1586 0 1 23674
box 0 0 1 1
use contact_13  contact_13_124
timestamp 1643593061
transform 1 0 1589 0 1 23677
box 0 0 1 1
use contact_21  contact_21_124
timestamp 1643593061
transform 1 0 1593 0 1 23659
box 0 0 1 1
use contact_17  contact_17_125
timestamp 1643593061
transform 1 0 1586 0 1 23338
box 0 0 1 1
use contact_13  contact_13_125
timestamp 1643593061
transform 1 0 1589 0 1 23341
box 0 0 1 1
use contact_21  contact_21_125
timestamp 1643593061
transform 1 0 1593 0 1 23323
box 0 0 1 1
use contact_17  contact_17_126
timestamp 1643593061
transform 1 0 1586 0 1 23002
box 0 0 1 1
use contact_13  contact_13_126
timestamp 1643593061
transform 1 0 1589 0 1 23005
box 0 0 1 1
use contact_21  contact_21_126
timestamp 1643593061
transform 1 0 1593 0 1 22987
box 0 0 1 1
use contact_17  contact_17_127
timestamp 1643593061
transform 1 0 1586 0 1 22666
box 0 0 1 1
use contact_13  contact_13_127
timestamp 1643593061
transform 1 0 1589 0 1 22669
box 0 0 1 1
use contact_21  contact_21_127
timestamp 1643593061
transform 1 0 1593 0 1 22651
box 0 0 1 1
use contact_17  contact_17_128
timestamp 1643593061
transform 1 0 1586 0 1 22330
box 0 0 1 1
use contact_13  contact_13_128
timestamp 1643593061
transform 1 0 1589 0 1 22333
box 0 0 1 1
use contact_21  contact_21_128
timestamp 1643593061
transform 1 0 1593 0 1 22315
box 0 0 1 1
use contact_18  contact_18_25
timestamp 1643593061
transform 1 0 1588 0 1 21990
box 0 0 1 1
use contact_17  contact_17_129
timestamp 1643593061
transform 1 0 1586 0 1 21994
box 0 0 1 1
use contact_13  contact_13_129
timestamp 1643593061
transform 1 0 1589 0 1 21997
box 0 0 1 1
use contact_21  contact_21_129
timestamp 1643593061
transform 1 0 1593 0 1 21979
box 0 0 1 1
use contact_17  contact_17_130
timestamp 1643593061
transform 1 0 1586 0 1 21658
box 0 0 1 1
use contact_13  contact_13_130
timestamp 1643593061
transform 1 0 1589 0 1 21661
box 0 0 1 1
use contact_21  contact_21_130
timestamp 1643593061
transform 1 0 1593 0 1 21643
box 0 0 1 1
use contact_17  contact_17_131
timestamp 1643593061
transform 1 0 1586 0 1 21322
box 0 0 1 1
use contact_13  contact_13_131
timestamp 1643593061
transform 1 0 1589 0 1 21325
box 0 0 1 1
use contact_21  contact_21_131
timestamp 1643593061
transform 1 0 1593 0 1 21307
box 0 0 1 1
use contact_17  contact_17_132
timestamp 1643593061
transform 1 0 1586 0 1 20986
box 0 0 1 1
use contact_13  contact_13_132
timestamp 1643593061
transform 1 0 1589 0 1 20989
box 0 0 1 1
use contact_21  contact_21_132
timestamp 1643593061
transform 1 0 1593 0 1 20971
box 0 0 1 1
use contact_17  contact_17_133
timestamp 1643593061
transform 1 0 1586 0 1 20650
box 0 0 1 1
use contact_13  contact_13_133
timestamp 1643593061
transform 1 0 1589 0 1 20653
box 0 0 1 1
use contact_21  contact_21_133
timestamp 1643593061
transform 1 0 1593 0 1 20635
box 0 0 1 1
use contact_18  contact_18_26
timestamp 1643593061
transform 1 0 1588 0 1 20310
box 0 0 1 1
use contact_17  contact_17_134
timestamp 1643593061
transform 1 0 1586 0 1 20314
box 0 0 1 1
use contact_13  contact_13_134
timestamp 1643593061
transform 1 0 1589 0 1 20317
box 0 0 1 1
use contact_21  contact_21_134
timestamp 1643593061
transform 1 0 1593 0 1 20299
box 0 0 1 1
use contact_17  contact_17_135
timestamp 1643593061
transform 1 0 1586 0 1 19978
box 0 0 1 1
use contact_13  contact_13_135
timestamp 1643593061
transform 1 0 1589 0 1 19981
box 0 0 1 1
use contact_21  contact_21_135
timestamp 1643593061
transform 1 0 1593 0 1 19963
box 0 0 1 1
use contact_17  contact_17_136
timestamp 1643593061
transform 1 0 1586 0 1 19642
box 0 0 1 1
use contact_13  contact_13_136
timestamp 1643593061
transform 1 0 1589 0 1 19645
box 0 0 1 1
use contact_21  contact_21_136
timestamp 1643593061
transform 1 0 1593 0 1 19627
box 0 0 1 1
use contact_17  contact_17_137
timestamp 1643593061
transform 1 0 1586 0 1 19306
box 0 0 1 1
use contact_13  contact_13_137
timestamp 1643593061
transform 1 0 1589 0 1 19309
box 0 0 1 1
use contact_21  contact_21_137
timestamp 1643593061
transform 1 0 1593 0 1 19291
box 0 0 1 1
use contact_17  contact_17_138
timestamp 1643593061
transform 1 0 1586 0 1 18970
box 0 0 1 1
use contact_13  contact_13_138
timestamp 1643593061
transform 1 0 1589 0 1 18973
box 0 0 1 1
use contact_21  contact_21_138
timestamp 1643593061
transform 1 0 1593 0 1 18955
box 0 0 1 1
use contact_18  contact_18_27
timestamp 1643593061
transform 1 0 1588 0 1 18630
box 0 0 1 1
use contact_17  contact_17_139
timestamp 1643593061
transform 1 0 1586 0 1 18634
box 0 0 1 1
use contact_13  contact_13_139
timestamp 1643593061
transform 1 0 1589 0 1 18637
box 0 0 1 1
use contact_21  contact_21_139
timestamp 1643593061
transform 1 0 1593 0 1 18619
box 0 0 1 1
use contact_17  contact_17_140
timestamp 1643593061
transform 1 0 1586 0 1 18298
box 0 0 1 1
use contact_13  contact_13_140
timestamp 1643593061
transform 1 0 1589 0 1 18301
box 0 0 1 1
use contact_21  contact_21_140
timestamp 1643593061
transform 1 0 1593 0 1 18283
box 0 0 1 1
use contact_17  contact_17_141
timestamp 1643593061
transform 1 0 1586 0 1 17962
box 0 0 1 1
use contact_13  contact_13_141
timestamp 1643593061
transform 1 0 1589 0 1 17965
box 0 0 1 1
use contact_21  contact_21_141
timestamp 1643593061
transform 1 0 1593 0 1 17947
box 0 0 1 1
use contact_17  contact_17_142
timestamp 1643593061
transform 1 0 1586 0 1 17626
box 0 0 1 1
use contact_13  contact_13_142
timestamp 1643593061
transform 1 0 1589 0 1 17629
box 0 0 1 1
use contact_21  contact_21_142
timestamp 1643593061
transform 1 0 1593 0 1 17611
box 0 0 1 1
use contact_17  contact_17_143
timestamp 1643593061
transform 1 0 1586 0 1 17290
box 0 0 1 1
use contact_13  contact_13_143
timestamp 1643593061
transform 1 0 1589 0 1 17293
box 0 0 1 1
use contact_21  contact_21_143
timestamp 1643593061
transform 1 0 1593 0 1 17275
box 0 0 1 1
use contact_18  contact_18_28
timestamp 1643593061
transform 1 0 1588 0 1 16950
box 0 0 1 1
use contact_17  contact_17_144
timestamp 1643593061
transform 1 0 1586 0 1 16954
box 0 0 1 1
use contact_13  contact_13_144
timestamp 1643593061
transform 1 0 1589 0 1 16957
box 0 0 1 1
use contact_21  contact_21_144
timestamp 1643593061
transform 1 0 1593 0 1 16939
box 0 0 1 1
use contact_17  contact_17_145
timestamp 1643593061
transform 1 0 1586 0 1 16618
box 0 0 1 1
use contact_13  contact_13_145
timestamp 1643593061
transform 1 0 1589 0 1 16621
box 0 0 1 1
use contact_21  contact_21_145
timestamp 1643593061
transform 1 0 1593 0 1 16603
box 0 0 1 1
use contact_17  contact_17_146
timestamp 1643593061
transform 1 0 1586 0 1 16282
box 0 0 1 1
use contact_13  contact_13_146
timestamp 1643593061
transform 1 0 1589 0 1 16285
box 0 0 1 1
use contact_21  contact_21_146
timestamp 1643593061
transform 1 0 1593 0 1 16267
box 0 0 1 1
use contact_17  contact_17_147
timestamp 1643593061
transform 1 0 1586 0 1 15946
box 0 0 1 1
use contact_13  contact_13_147
timestamp 1643593061
transform 1 0 1589 0 1 15949
box 0 0 1 1
use contact_21  contact_21_147
timestamp 1643593061
transform 1 0 1593 0 1 15931
box 0 0 1 1
use contact_17  contact_17_148
timestamp 1643593061
transform 1 0 1586 0 1 15610
box 0 0 1 1
use contact_13  contact_13_148
timestamp 1643593061
transform 1 0 1589 0 1 15613
box 0 0 1 1
use contact_21  contact_21_148
timestamp 1643593061
transform 1 0 1593 0 1 15595
box 0 0 1 1
use contact_18  contact_18_29
timestamp 1643593061
transform 1 0 1588 0 1 15270
box 0 0 1 1
use contact_17  contact_17_149
timestamp 1643593061
transform 1 0 1586 0 1 15274
box 0 0 1 1
use contact_13  contact_13_149
timestamp 1643593061
transform 1 0 1589 0 1 15277
box 0 0 1 1
use contact_21  contact_21_149
timestamp 1643593061
transform 1 0 1593 0 1 15259
box 0 0 1 1
use contact_17  contact_17_150
timestamp 1643593061
transform 1 0 1586 0 1 14938
box 0 0 1 1
use contact_13  contact_13_150
timestamp 1643593061
transform 1 0 1589 0 1 14941
box 0 0 1 1
use contact_21  contact_21_150
timestamp 1643593061
transform 1 0 1593 0 1 14923
box 0 0 1 1
use contact_17  contact_17_151
timestamp 1643593061
transform 1 0 1586 0 1 14602
box 0 0 1 1
use contact_13  contact_13_151
timestamp 1643593061
transform 1 0 1589 0 1 14605
box 0 0 1 1
use contact_21  contact_21_151
timestamp 1643593061
transform 1 0 1593 0 1 14587
box 0 0 1 1
use contact_17  contact_17_152
timestamp 1643593061
transform 1 0 1586 0 1 14266
box 0 0 1 1
use contact_13  contact_13_152
timestamp 1643593061
transform 1 0 1589 0 1 14269
box 0 0 1 1
use contact_21  contact_21_152
timestamp 1643593061
transform 1 0 1593 0 1 14251
box 0 0 1 1
use contact_17  contact_17_153
timestamp 1643593061
transform 1 0 1586 0 1 13930
box 0 0 1 1
use contact_13  contact_13_153
timestamp 1643593061
transform 1 0 1589 0 1 13933
box 0 0 1 1
use contact_21  contact_21_153
timestamp 1643593061
transform 1 0 1593 0 1 13915
box 0 0 1 1
use contact_18  contact_18_30
timestamp 1643593061
transform 1 0 1588 0 1 13590
box 0 0 1 1
use contact_17  contact_17_154
timestamp 1643593061
transform 1 0 1586 0 1 13594
box 0 0 1 1
use contact_13  contact_13_154
timestamp 1643593061
transform 1 0 1589 0 1 13597
box 0 0 1 1
use contact_21  contact_21_154
timestamp 1643593061
transform 1 0 1593 0 1 13579
box 0 0 1 1
use contact_17  contact_17_155
timestamp 1643593061
transform 1 0 1586 0 1 13258
box 0 0 1 1
use contact_13  contact_13_155
timestamp 1643593061
transform 1 0 1589 0 1 13261
box 0 0 1 1
use contact_21  contact_21_155
timestamp 1643593061
transform 1 0 1593 0 1 13243
box 0 0 1 1
use contact_17  contact_17_156
timestamp 1643593061
transform 1 0 1586 0 1 12922
box 0 0 1 1
use contact_13  contact_13_156
timestamp 1643593061
transform 1 0 1589 0 1 12925
box 0 0 1 1
use contact_21  contact_21_156
timestamp 1643593061
transform 1 0 1593 0 1 12907
box 0 0 1 1
use contact_17  contact_17_157
timestamp 1643593061
transform 1 0 1586 0 1 12586
box 0 0 1 1
use contact_13  contact_13_157
timestamp 1643593061
transform 1 0 1589 0 1 12589
box 0 0 1 1
use contact_21  contact_21_157
timestamp 1643593061
transform 1 0 1593 0 1 12571
box 0 0 1 1
use contact_17  contact_17_158
timestamp 1643593061
transform 1 0 1586 0 1 12250
box 0 0 1 1
use contact_13  contact_13_158
timestamp 1643593061
transform 1 0 1589 0 1 12253
box 0 0 1 1
use contact_21  contact_21_158
timestamp 1643593061
transform 1 0 1593 0 1 12235
box 0 0 1 1
use contact_18  contact_18_31
timestamp 1643593061
transform 1 0 1588 0 1 11910
box 0 0 1 1
use contact_17  contact_17_159
timestamp 1643593061
transform 1 0 1586 0 1 11914
box 0 0 1 1
use contact_13  contact_13_159
timestamp 1643593061
transform 1 0 1589 0 1 11917
box 0 0 1 1
use contact_21  contact_21_159
timestamp 1643593061
transform 1 0 1593 0 1 11899
box 0 0 1 1
use contact_17  contact_17_160
timestamp 1643593061
transform 1 0 1586 0 1 11578
box 0 0 1 1
use contact_13  contact_13_160
timestamp 1643593061
transform 1 0 1589 0 1 11581
box 0 0 1 1
use contact_21  contact_21_160
timestamp 1643593061
transform 1 0 1593 0 1 11563
box 0 0 1 1
use contact_17  contact_17_161
timestamp 1643593061
transform 1 0 1586 0 1 11242
box 0 0 1 1
use contact_13  contact_13_161
timestamp 1643593061
transform 1 0 1589 0 1 11245
box 0 0 1 1
use contact_21  contact_21_161
timestamp 1643593061
transform 1 0 1593 0 1 11227
box 0 0 1 1
use contact_17  contact_17_162
timestamp 1643593061
transform 1 0 1586 0 1 10906
box 0 0 1 1
use contact_13  contact_13_162
timestamp 1643593061
transform 1 0 1589 0 1 10909
box 0 0 1 1
use contact_21  contact_21_162
timestamp 1643593061
transform 1 0 1593 0 1 10891
box 0 0 1 1
use contact_17  contact_17_163
timestamp 1643593061
transform 1 0 1586 0 1 10570
box 0 0 1 1
use contact_13  contact_13_163
timestamp 1643593061
transform 1 0 1589 0 1 10573
box 0 0 1 1
use contact_21  contact_21_163
timestamp 1643593061
transform 1 0 1593 0 1 10555
box 0 0 1 1
use contact_18  contact_18_32
timestamp 1643593061
transform 1 0 1588 0 1 10230
box 0 0 1 1
use contact_17  contact_17_164
timestamp 1643593061
transform 1 0 1586 0 1 10234
box 0 0 1 1
use contact_13  contact_13_164
timestamp 1643593061
transform 1 0 1589 0 1 10237
box 0 0 1 1
use contact_21  contact_21_164
timestamp 1643593061
transform 1 0 1593 0 1 10219
box 0 0 1 1
use contact_17  contact_17_165
timestamp 1643593061
transform 1 0 1586 0 1 9898
box 0 0 1 1
use contact_13  contact_13_165
timestamp 1643593061
transform 1 0 1589 0 1 9901
box 0 0 1 1
use contact_21  contact_21_165
timestamp 1643593061
transform 1 0 1593 0 1 9883
box 0 0 1 1
use contact_17  contact_17_166
timestamp 1643593061
transform 1 0 1586 0 1 9562
box 0 0 1 1
use contact_13  contact_13_166
timestamp 1643593061
transform 1 0 1589 0 1 9565
box 0 0 1 1
use contact_21  contact_21_166
timestamp 1643593061
transform 1 0 1593 0 1 9547
box 0 0 1 1
use contact_17  contact_17_167
timestamp 1643593061
transform 1 0 1586 0 1 9226
box 0 0 1 1
use contact_13  contact_13_167
timestamp 1643593061
transform 1 0 1589 0 1 9229
box 0 0 1 1
use contact_21  contact_21_167
timestamp 1643593061
transform 1 0 1593 0 1 9211
box 0 0 1 1
use contact_17  contact_17_168
timestamp 1643593061
transform 1 0 1586 0 1 8890
box 0 0 1 1
use contact_13  contact_13_168
timestamp 1643593061
transform 1 0 1589 0 1 8893
box 0 0 1 1
use contact_21  contact_21_168
timestamp 1643593061
transform 1 0 1593 0 1 8875
box 0 0 1 1
use contact_18  contact_18_33
timestamp 1643593061
transform 1 0 1588 0 1 8550
box 0 0 1 1
use contact_17  contact_17_169
timestamp 1643593061
transform 1 0 1586 0 1 8554
box 0 0 1 1
use contact_13  contact_13_169
timestamp 1643593061
transform 1 0 1589 0 1 8557
box 0 0 1 1
use contact_21  contact_21_169
timestamp 1643593061
transform 1 0 1593 0 1 8539
box 0 0 1 1
use contact_17  contact_17_170
timestamp 1643593061
transform 1 0 1586 0 1 8218
box 0 0 1 1
use contact_13  contact_13_170
timestamp 1643593061
transform 1 0 1589 0 1 8221
box 0 0 1 1
use contact_21  contact_21_170
timestamp 1643593061
transform 1 0 1593 0 1 8203
box 0 0 1 1
use contact_17  contact_17_171
timestamp 1643593061
transform 1 0 1586 0 1 7882
box 0 0 1 1
use contact_13  contact_13_171
timestamp 1643593061
transform 1 0 1589 0 1 7885
box 0 0 1 1
use contact_21  contact_21_171
timestamp 1643593061
transform 1 0 1593 0 1 7867
box 0 0 1 1
use contact_17  contact_17_172
timestamp 1643593061
transform 1 0 1586 0 1 7546
box 0 0 1 1
use contact_13  contact_13_172
timestamp 1643593061
transform 1 0 1589 0 1 7549
box 0 0 1 1
use contact_21  contact_21_172
timestamp 1643593061
transform 1 0 1593 0 1 7531
box 0 0 1 1
use contact_17  contact_17_173
timestamp 1643593061
transform 1 0 1586 0 1 7210
box 0 0 1 1
use contact_13  contact_13_173
timestamp 1643593061
transform 1 0 1589 0 1 7213
box 0 0 1 1
use contact_21  contact_21_173
timestamp 1643593061
transform 1 0 1593 0 1 7195
box 0 0 1 1
use contact_18  contact_18_34
timestamp 1643593061
transform 1 0 1588 0 1 6870
box 0 0 1 1
use contact_17  contact_17_174
timestamp 1643593061
transform 1 0 1586 0 1 6874
box 0 0 1 1
use contact_13  contact_13_174
timestamp 1643593061
transform 1 0 1589 0 1 6877
box 0 0 1 1
use contact_21  contact_21_174
timestamp 1643593061
transform 1 0 1593 0 1 6859
box 0 0 1 1
use contact_17  contact_17_175
timestamp 1643593061
transform 1 0 1586 0 1 6538
box 0 0 1 1
use contact_13  contact_13_175
timestamp 1643593061
transform 1 0 1589 0 1 6541
box 0 0 1 1
use contact_21  contact_21_175
timestamp 1643593061
transform 1 0 1593 0 1 6523
box 0 0 1 1
use contact_17  contact_17_176
timestamp 1643593061
transform 1 0 1586 0 1 6202
box 0 0 1 1
use contact_13  contact_13_176
timestamp 1643593061
transform 1 0 1589 0 1 6205
box 0 0 1 1
use contact_21  contact_21_176
timestamp 1643593061
transform 1 0 1593 0 1 6187
box 0 0 1 1
use contact_17  contact_17_177
timestamp 1643593061
transform 1 0 1586 0 1 5866
box 0 0 1 1
use contact_13  contact_13_177
timestamp 1643593061
transform 1 0 1589 0 1 5869
box 0 0 1 1
use contact_21  contact_21_177
timestamp 1643593061
transform 1 0 1593 0 1 5851
box 0 0 1 1
use contact_17  contact_17_178
timestamp 1643593061
transform 1 0 1586 0 1 5530
box 0 0 1 1
use contact_13  contact_13_178
timestamp 1643593061
transform 1 0 1589 0 1 5533
box 0 0 1 1
use contact_21  contact_21_178
timestamp 1643593061
transform 1 0 1593 0 1 5515
box 0 0 1 1
use contact_18  contact_18_35
timestamp 1643593061
transform 1 0 1588 0 1 5190
box 0 0 1 1
use contact_17  contact_17_179
timestamp 1643593061
transform 1 0 1586 0 1 5194
box 0 0 1 1
use contact_13  contact_13_179
timestamp 1643593061
transform 1 0 1589 0 1 5197
box 0 0 1 1
use contact_21  contact_21_179
timestamp 1643593061
transform 1 0 1593 0 1 5179
box 0 0 1 1
use contact_17  contact_17_180
timestamp 1643593061
transform 1 0 1586 0 1 4858
box 0 0 1 1
use contact_13  contact_13_180
timestamp 1643593061
transform 1 0 1589 0 1 4861
box 0 0 1 1
use contact_21  contact_21_180
timestamp 1643593061
transform 1 0 1593 0 1 4843
box 0 0 1 1
use contact_17  contact_17_181
timestamp 1643593061
transform 1 0 1586 0 1 4522
box 0 0 1 1
use contact_13  contact_13_181
timestamp 1643593061
transform 1 0 1589 0 1 4525
box 0 0 1 1
use contact_21  contact_21_181
timestamp 1643593061
transform 1 0 1593 0 1 4507
box 0 0 1 1
use contact_17  contact_17_182
timestamp 1643593061
transform 1 0 1586 0 1 4186
box 0 0 1 1
use contact_13  contact_13_182
timestamp 1643593061
transform 1 0 1589 0 1 4189
box 0 0 1 1
use contact_21  contact_21_182
timestamp 1643593061
transform 1 0 1593 0 1 4171
box 0 0 1 1
use contact_17  contact_17_183
timestamp 1643593061
transform 1 0 1586 0 1 3850
box 0 0 1 1
use contact_13  contact_13_183
timestamp 1643593061
transform 1 0 1589 0 1 3853
box 0 0 1 1
use contact_21  contact_21_183
timestamp 1643593061
transform 1 0 1593 0 1 3835
box 0 0 1 1
use contact_18  contact_18_36
timestamp 1643593061
transform 1 0 1588 0 1 3510
box 0 0 1 1
use contact_17  contact_17_184
timestamp 1643593061
transform 1 0 1586 0 1 3514
box 0 0 1 1
use contact_13  contact_13_184
timestamp 1643593061
transform 1 0 1589 0 1 3517
box 0 0 1 1
use contact_21  contact_21_184
timestamp 1643593061
transform 1 0 1593 0 1 3499
box 0 0 1 1
use contact_17  contact_17_185
timestamp 1643593061
transform 1 0 1586 0 1 3178
box 0 0 1 1
use contact_13  contact_13_185
timestamp 1643593061
transform 1 0 1589 0 1 3181
box 0 0 1 1
use contact_21  contact_21_185
timestamp 1643593061
transform 1 0 1593 0 1 3163
box 0 0 1 1
use contact_17  contact_17_186
timestamp 1643593061
transform 1 0 1586 0 1 2842
box 0 0 1 1
use contact_13  contact_13_186
timestamp 1643593061
transform 1 0 1589 0 1 2845
box 0 0 1 1
use contact_21  contact_21_186
timestamp 1643593061
transform 1 0 1593 0 1 2827
box 0 0 1 1
use contact_17  contact_17_187
timestamp 1643593061
transform 1 0 1586 0 1 2506
box 0 0 1 1
use contact_13  contact_13_187
timestamp 1643593061
transform 1 0 1589 0 1 2509
box 0 0 1 1
use contact_21  contact_21_187
timestamp 1643593061
transform 1 0 1593 0 1 2491
box 0 0 1 1
use contact_17  contact_17_188
timestamp 1643593061
transform 1 0 1586 0 1 2170
box 0 0 1 1
use contact_13  contact_13_188
timestamp 1643593061
transform 1 0 1589 0 1 2173
box 0 0 1 1
use contact_21  contact_21_188
timestamp 1643593061
transform 1 0 1593 0 1 2155
box 0 0 1 1
use contact_18  contact_18_37
timestamp 1643593061
transform 1 0 1588 0 1 1830
box 0 0 1 1
use contact_17  contact_17_189
timestamp 1643593061
transform 1 0 1586 0 1 1834
box 0 0 1 1
use contact_13  contact_13_189
timestamp 1643593061
transform 1 0 1589 0 1 1837
box 0 0 1 1
use contact_21  contact_21_189
timestamp 1643593061
transform 1 0 1593 0 1 1819
box 0 0 1 1
use contact_18  contact_18_38
timestamp 1643593061
transform 1 0 23764 0 1 33904
box 0 0 1 1
use contact_17  contact_17_190
timestamp 1643593061
transform 1 0 23762 0 1 33908
box 0 0 1 1
use contact_13  contact_13_190
timestamp 1643593061
transform 1 0 23765 0 1 33911
box 0 0 1 1
use contact_21  contact_21_190
timestamp 1643593061
transform 1 0 23769 0 1 33893
box 0 0 1 1
use contact_13  contact_13_191
timestamp 1643593061
transform 1 0 23429 0 1 33911
box 0 0 1 1
use contact_21  contact_21_191
timestamp 1643593061
transform 1 0 23433 0 1 33893
box 0 0 1 1
use contact_13  contact_13_192
timestamp 1643593061
transform 1 0 23093 0 1 33911
box 0 0 1 1
use contact_21  contact_21_192
timestamp 1643593061
transform 1 0 23097 0 1 33893
box 0 0 1 1
use contact_13  contact_13_193
timestamp 1643593061
transform 1 0 22757 0 1 33911
box 0 0 1 1
use contact_21  contact_21_193
timestamp 1643593061
transform 1 0 22761 0 1 33893
box 0 0 1 1
use contact_13  contact_13_194
timestamp 1643593061
transform 1 0 22421 0 1 33911
box 0 0 1 1
use contact_21  contact_21_194
timestamp 1643593061
transform 1 0 22425 0 1 33893
box 0 0 1 1
use contact_18  contact_18_39
timestamp 1643593061
transform 1 0 22084 0 1 33904
box 0 0 1 1
use contact_17  contact_17_191
timestamp 1643593061
transform 1 0 22082 0 1 33908
box 0 0 1 1
use contact_13  contact_13_195
timestamp 1643593061
transform 1 0 22085 0 1 33911
box 0 0 1 1
use contact_21  contact_21_195
timestamp 1643593061
transform 1 0 22089 0 1 33893
box 0 0 1 1
use contact_13  contact_13_196
timestamp 1643593061
transform 1 0 21749 0 1 33911
box 0 0 1 1
use contact_21  contact_21_196
timestamp 1643593061
transform 1 0 21753 0 1 33893
box 0 0 1 1
use contact_13  contact_13_197
timestamp 1643593061
transform 1 0 21413 0 1 33911
box 0 0 1 1
use contact_21  contact_21_197
timestamp 1643593061
transform 1 0 21417 0 1 33893
box 0 0 1 1
use contact_13  contact_13_198
timestamp 1643593061
transform 1 0 21077 0 1 33911
box 0 0 1 1
use contact_21  contact_21_198
timestamp 1643593061
transform 1 0 21081 0 1 33893
box 0 0 1 1
use contact_13  contact_13_199
timestamp 1643593061
transform 1 0 20741 0 1 33911
box 0 0 1 1
use contact_21  contact_21_199
timestamp 1643593061
transform 1 0 20745 0 1 33893
box 0 0 1 1
use contact_18  contact_18_40
timestamp 1643593061
transform 1 0 20404 0 1 33904
box 0 0 1 1
use contact_17  contact_17_192
timestamp 1643593061
transform 1 0 20402 0 1 33908
box 0 0 1 1
use contact_13  contact_13_200
timestamp 1643593061
transform 1 0 20405 0 1 33911
box 0 0 1 1
use contact_21  contact_21_200
timestamp 1643593061
transform 1 0 20409 0 1 33893
box 0 0 1 1
use contact_13  contact_13_201
timestamp 1643593061
transform 1 0 20069 0 1 33911
box 0 0 1 1
use contact_21  contact_21_201
timestamp 1643593061
transform 1 0 20073 0 1 33893
box 0 0 1 1
use contact_13  contact_13_202
timestamp 1643593061
transform 1 0 19733 0 1 33911
box 0 0 1 1
use contact_21  contact_21_202
timestamp 1643593061
transform 1 0 19737 0 1 33893
box 0 0 1 1
use contact_13  contact_13_203
timestamp 1643593061
transform 1 0 19397 0 1 33911
box 0 0 1 1
use contact_21  contact_21_203
timestamp 1643593061
transform 1 0 19401 0 1 33893
box 0 0 1 1
use contact_13  contact_13_204
timestamp 1643593061
transform 1 0 19061 0 1 33911
box 0 0 1 1
use contact_21  contact_21_204
timestamp 1643593061
transform 1 0 19065 0 1 33893
box 0 0 1 1
use contact_18  contact_18_41
timestamp 1643593061
transform 1 0 18724 0 1 33904
box 0 0 1 1
use contact_17  contact_17_193
timestamp 1643593061
transform 1 0 18722 0 1 33908
box 0 0 1 1
use contact_13  contact_13_205
timestamp 1643593061
transform 1 0 18725 0 1 33911
box 0 0 1 1
use contact_21  contact_21_205
timestamp 1643593061
transform 1 0 18729 0 1 33893
box 0 0 1 1
use contact_13  contact_13_206
timestamp 1643593061
transform 1 0 18389 0 1 33911
box 0 0 1 1
use contact_21  contact_21_206
timestamp 1643593061
transform 1 0 18393 0 1 33893
box 0 0 1 1
use contact_13  contact_13_207
timestamp 1643593061
transform 1 0 18053 0 1 33911
box 0 0 1 1
use contact_21  contact_21_207
timestamp 1643593061
transform 1 0 18057 0 1 33893
box 0 0 1 1
use contact_13  contact_13_208
timestamp 1643593061
transform 1 0 17717 0 1 33911
box 0 0 1 1
use contact_21  contact_21_208
timestamp 1643593061
transform 1 0 17721 0 1 33893
box 0 0 1 1
use contact_13  contact_13_209
timestamp 1643593061
transform 1 0 17381 0 1 33911
box 0 0 1 1
use contact_21  contact_21_209
timestamp 1643593061
transform 1 0 17385 0 1 33893
box 0 0 1 1
use contact_18  contact_18_42
timestamp 1643593061
transform 1 0 17044 0 1 33904
box 0 0 1 1
use contact_17  contact_17_194
timestamp 1643593061
transform 1 0 17042 0 1 33908
box 0 0 1 1
use contact_13  contact_13_210
timestamp 1643593061
transform 1 0 17045 0 1 33911
box 0 0 1 1
use contact_21  contact_21_210
timestamp 1643593061
transform 1 0 17049 0 1 33893
box 0 0 1 1
use contact_13  contact_13_211
timestamp 1643593061
transform 1 0 16709 0 1 33911
box 0 0 1 1
use contact_21  contact_21_211
timestamp 1643593061
transform 1 0 16713 0 1 33893
box 0 0 1 1
use contact_13  contact_13_212
timestamp 1643593061
transform 1 0 16373 0 1 33911
box 0 0 1 1
use contact_21  contact_21_212
timestamp 1643593061
transform 1 0 16377 0 1 33893
box 0 0 1 1
use contact_13  contact_13_213
timestamp 1643593061
transform 1 0 16037 0 1 33911
box 0 0 1 1
use contact_21  contact_21_213
timestamp 1643593061
transform 1 0 16041 0 1 33893
box 0 0 1 1
use contact_13  contact_13_214
timestamp 1643593061
transform 1 0 15701 0 1 33911
box 0 0 1 1
use contact_21  contact_21_214
timestamp 1643593061
transform 1 0 15705 0 1 33893
box 0 0 1 1
use contact_18  contact_18_43
timestamp 1643593061
transform 1 0 15364 0 1 33904
box 0 0 1 1
use contact_17  contact_17_195
timestamp 1643593061
transform 1 0 15362 0 1 33908
box 0 0 1 1
use contact_13  contact_13_215
timestamp 1643593061
transform 1 0 15365 0 1 33911
box 0 0 1 1
use contact_21  contact_21_215
timestamp 1643593061
transform 1 0 15369 0 1 33893
box 0 0 1 1
use contact_13  contact_13_216
timestamp 1643593061
transform 1 0 15029 0 1 33911
box 0 0 1 1
use contact_21  contact_21_216
timestamp 1643593061
transform 1 0 15033 0 1 33893
box 0 0 1 1
use contact_13  contact_13_217
timestamp 1643593061
transform 1 0 14693 0 1 33911
box 0 0 1 1
use contact_21  contact_21_217
timestamp 1643593061
transform 1 0 14697 0 1 33893
box 0 0 1 1
use contact_13  contact_13_218
timestamp 1643593061
transform 1 0 14357 0 1 33911
box 0 0 1 1
use contact_21  contact_21_218
timestamp 1643593061
transform 1 0 14361 0 1 33893
box 0 0 1 1
use contact_13  contact_13_219
timestamp 1643593061
transform 1 0 14021 0 1 33911
box 0 0 1 1
use contact_21  contact_21_219
timestamp 1643593061
transform 1 0 14025 0 1 33893
box 0 0 1 1
use contact_18  contact_18_44
timestamp 1643593061
transform 1 0 13684 0 1 33904
box 0 0 1 1
use contact_17  contact_17_196
timestamp 1643593061
transform 1 0 13682 0 1 33908
box 0 0 1 1
use contact_13  contact_13_220
timestamp 1643593061
transform 1 0 13685 0 1 33911
box 0 0 1 1
use contact_21  contact_21_220
timestamp 1643593061
transform 1 0 13689 0 1 33893
box 0 0 1 1
use contact_13  contact_13_221
timestamp 1643593061
transform 1 0 13349 0 1 33911
box 0 0 1 1
use contact_21  contact_21_221
timestamp 1643593061
transform 1 0 13353 0 1 33893
box 0 0 1 1
use contact_13  contact_13_222
timestamp 1643593061
transform 1 0 13013 0 1 33911
box 0 0 1 1
use contact_21  contact_21_222
timestamp 1643593061
transform 1 0 13017 0 1 33893
box 0 0 1 1
use contact_13  contact_13_223
timestamp 1643593061
transform 1 0 12677 0 1 33911
box 0 0 1 1
use contact_21  contact_21_223
timestamp 1643593061
transform 1 0 12681 0 1 33893
box 0 0 1 1
use contact_13  contact_13_224
timestamp 1643593061
transform 1 0 12341 0 1 33911
box 0 0 1 1
use contact_21  contact_21_224
timestamp 1643593061
transform 1 0 12345 0 1 33893
box 0 0 1 1
use contact_18  contact_18_45
timestamp 1643593061
transform 1 0 12004 0 1 33904
box 0 0 1 1
use contact_17  contact_17_197
timestamp 1643593061
transform 1 0 12002 0 1 33908
box 0 0 1 1
use contact_13  contact_13_225
timestamp 1643593061
transform 1 0 12005 0 1 33911
box 0 0 1 1
use contact_21  contact_21_225
timestamp 1643593061
transform 1 0 12009 0 1 33893
box 0 0 1 1
use contact_13  contact_13_226
timestamp 1643593061
transform 1 0 11669 0 1 33911
box 0 0 1 1
use contact_21  contact_21_226
timestamp 1643593061
transform 1 0 11673 0 1 33893
box 0 0 1 1
use contact_13  contact_13_227
timestamp 1643593061
transform 1 0 11333 0 1 33911
box 0 0 1 1
use contact_21  contact_21_227
timestamp 1643593061
transform 1 0 11337 0 1 33893
box 0 0 1 1
use contact_13  contact_13_228
timestamp 1643593061
transform 1 0 10997 0 1 33911
box 0 0 1 1
use contact_21  contact_21_228
timestamp 1643593061
transform 1 0 11001 0 1 33893
box 0 0 1 1
use contact_13  contact_13_229
timestamp 1643593061
transform 1 0 10661 0 1 33911
box 0 0 1 1
use contact_21  contact_21_229
timestamp 1643593061
transform 1 0 10665 0 1 33893
box 0 0 1 1
use contact_18  contact_18_46
timestamp 1643593061
transform 1 0 10324 0 1 33904
box 0 0 1 1
use contact_17  contact_17_198
timestamp 1643593061
transform 1 0 10322 0 1 33908
box 0 0 1 1
use contact_13  contact_13_230
timestamp 1643593061
transform 1 0 10325 0 1 33911
box 0 0 1 1
use contact_21  contact_21_230
timestamp 1643593061
transform 1 0 10329 0 1 33893
box 0 0 1 1
use contact_13  contact_13_231
timestamp 1643593061
transform 1 0 9989 0 1 33911
box 0 0 1 1
use contact_21  contact_21_231
timestamp 1643593061
transform 1 0 9993 0 1 33893
box 0 0 1 1
use contact_13  contact_13_232
timestamp 1643593061
transform 1 0 9653 0 1 33911
box 0 0 1 1
use contact_21  contact_21_232
timestamp 1643593061
transform 1 0 9657 0 1 33893
box 0 0 1 1
use contact_13  contact_13_233
timestamp 1643593061
transform 1 0 9317 0 1 33911
box 0 0 1 1
use contact_21  contact_21_233
timestamp 1643593061
transform 1 0 9321 0 1 33893
box 0 0 1 1
use contact_13  contact_13_234
timestamp 1643593061
transform 1 0 8981 0 1 33911
box 0 0 1 1
use contact_21  contact_21_234
timestamp 1643593061
transform 1 0 8985 0 1 33893
box 0 0 1 1
use contact_18  contact_18_47
timestamp 1643593061
transform 1 0 8644 0 1 33904
box 0 0 1 1
use contact_17  contact_17_199
timestamp 1643593061
transform 1 0 8642 0 1 33908
box 0 0 1 1
use contact_13  contact_13_235
timestamp 1643593061
transform 1 0 8645 0 1 33911
box 0 0 1 1
use contact_21  contact_21_235
timestamp 1643593061
transform 1 0 8649 0 1 33893
box 0 0 1 1
use contact_13  contact_13_236
timestamp 1643593061
transform 1 0 8309 0 1 33911
box 0 0 1 1
use contact_21  contact_21_236
timestamp 1643593061
transform 1 0 8313 0 1 33893
box 0 0 1 1
use contact_13  contact_13_237
timestamp 1643593061
transform 1 0 7973 0 1 33911
box 0 0 1 1
use contact_21  contact_21_237
timestamp 1643593061
transform 1 0 7977 0 1 33893
box 0 0 1 1
use contact_13  contact_13_238
timestamp 1643593061
transform 1 0 7637 0 1 33911
box 0 0 1 1
use contact_21  contact_21_238
timestamp 1643593061
transform 1 0 7641 0 1 33893
box 0 0 1 1
use contact_13  contact_13_239
timestamp 1643593061
transform 1 0 7301 0 1 33911
box 0 0 1 1
use contact_21  contact_21_239
timestamp 1643593061
transform 1 0 7305 0 1 33893
box 0 0 1 1
use contact_18  contact_18_48
timestamp 1643593061
transform 1 0 6964 0 1 33904
box 0 0 1 1
use contact_17  contact_17_200
timestamp 1643593061
transform 1 0 6962 0 1 33908
box 0 0 1 1
use contact_13  contact_13_240
timestamp 1643593061
transform 1 0 6965 0 1 33911
box 0 0 1 1
use contact_21  contact_21_240
timestamp 1643593061
transform 1 0 6969 0 1 33893
box 0 0 1 1
use contact_13  contact_13_241
timestamp 1643593061
transform 1 0 6629 0 1 33911
box 0 0 1 1
use contact_21  contact_21_241
timestamp 1643593061
transform 1 0 6633 0 1 33893
box 0 0 1 1
use contact_13  contact_13_242
timestamp 1643593061
transform 1 0 6293 0 1 33911
box 0 0 1 1
use contact_21  contact_21_242
timestamp 1643593061
transform 1 0 6297 0 1 33893
box 0 0 1 1
use contact_13  contact_13_243
timestamp 1643593061
transform 1 0 5957 0 1 33911
box 0 0 1 1
use contact_21  contact_21_243
timestamp 1643593061
transform 1 0 5961 0 1 33893
box 0 0 1 1
use contact_13  contact_13_244
timestamp 1643593061
transform 1 0 5621 0 1 33911
box 0 0 1 1
use contact_21  contact_21_244
timestamp 1643593061
transform 1 0 5625 0 1 33893
box 0 0 1 1
use contact_18  contact_18_49
timestamp 1643593061
transform 1 0 5284 0 1 33904
box 0 0 1 1
use contact_17  contact_17_201
timestamp 1643593061
transform 1 0 5282 0 1 33908
box 0 0 1 1
use contact_13  contact_13_245
timestamp 1643593061
transform 1 0 5285 0 1 33911
box 0 0 1 1
use contact_21  contact_21_245
timestamp 1643593061
transform 1 0 5289 0 1 33893
box 0 0 1 1
use contact_13  contact_13_246
timestamp 1643593061
transform 1 0 4949 0 1 33911
box 0 0 1 1
use contact_21  contact_21_246
timestamp 1643593061
transform 1 0 4953 0 1 33893
box 0 0 1 1
use contact_13  contact_13_247
timestamp 1643593061
transform 1 0 4613 0 1 33911
box 0 0 1 1
use contact_21  contact_21_247
timestamp 1643593061
transform 1 0 4617 0 1 33893
box 0 0 1 1
use contact_13  contact_13_248
timestamp 1643593061
transform 1 0 4277 0 1 33911
box 0 0 1 1
use contact_21  contact_21_248
timestamp 1643593061
transform 1 0 4281 0 1 33893
box 0 0 1 1
use contact_13  contact_13_249
timestamp 1643593061
transform 1 0 3941 0 1 33911
box 0 0 1 1
use contact_21  contact_21_249
timestamp 1643593061
transform 1 0 3945 0 1 33893
box 0 0 1 1
use contact_18  contact_18_50
timestamp 1643593061
transform 1 0 3604 0 1 33904
box 0 0 1 1
use contact_17  contact_17_202
timestamp 1643593061
transform 1 0 3602 0 1 33908
box 0 0 1 1
use contact_13  contact_13_250
timestamp 1643593061
transform 1 0 3605 0 1 33911
box 0 0 1 1
use contact_21  contact_21_250
timestamp 1643593061
transform 1 0 3609 0 1 33893
box 0 0 1 1
use contact_13  contact_13_251
timestamp 1643593061
transform 1 0 3269 0 1 33911
box 0 0 1 1
use contact_21  contact_21_251
timestamp 1643593061
transform 1 0 3273 0 1 33893
box 0 0 1 1
use contact_13  contact_13_252
timestamp 1643593061
transform 1 0 2933 0 1 33911
box 0 0 1 1
use contact_21  contact_21_252
timestamp 1643593061
transform 1 0 2937 0 1 33893
box 0 0 1 1
use contact_13  contact_13_253
timestamp 1643593061
transform 1 0 2597 0 1 33911
box 0 0 1 1
use contact_21  contact_21_253
timestamp 1643593061
transform 1 0 2601 0 1 33893
box 0 0 1 1
use contact_13  contact_13_254
timestamp 1643593061
transform 1 0 2261 0 1 33911
box 0 0 1 1
use contact_21  contact_21_254
timestamp 1643593061
transform 1 0 2265 0 1 33893
box 0 0 1 1
use contact_18  contact_18_51
timestamp 1643593061
transform 1 0 1924 0 1 33904
box 0 0 1 1
use contact_17  contact_17_203
timestamp 1643593061
transform 1 0 1922 0 1 33908
box 0 0 1 1
use contact_13  contact_13_255
timestamp 1643593061
transform 1 0 1925 0 1 33911
box 0 0 1 1
use contact_21  contact_21_255
timestamp 1643593061
transform 1 0 1929 0 1 33893
box 0 0 1 1
use contact_18  contact_18_52
timestamp 1643593061
transform 1 0 23764 0 1 1494
box 0 0 1 1
use contact_17  contact_17_204
timestamp 1643593061
transform 1 0 23762 0 1 1498
box 0 0 1 1
use contact_13  contact_13_256
timestamp 1643593061
transform 1 0 23765 0 1 1501
box 0 0 1 1
use contact_21  contact_21_256
timestamp 1643593061
transform 1 0 23769 0 1 1483
box 0 0 1 1
use contact_13  contact_13_257
timestamp 1643593061
transform 1 0 23429 0 1 1501
box 0 0 1 1
use contact_21  contact_21_257
timestamp 1643593061
transform 1 0 23433 0 1 1483
box 0 0 1 1
use contact_13  contact_13_258
timestamp 1643593061
transform 1 0 23093 0 1 1501
box 0 0 1 1
use contact_21  contact_21_258
timestamp 1643593061
transform 1 0 23097 0 1 1483
box 0 0 1 1
use contact_13  contact_13_259
timestamp 1643593061
transform 1 0 22757 0 1 1501
box 0 0 1 1
use contact_21  contact_21_259
timestamp 1643593061
transform 1 0 22761 0 1 1483
box 0 0 1 1
use contact_13  contact_13_260
timestamp 1643593061
transform 1 0 22421 0 1 1501
box 0 0 1 1
use contact_21  contact_21_260
timestamp 1643593061
transform 1 0 22425 0 1 1483
box 0 0 1 1
use contact_18  contact_18_53
timestamp 1643593061
transform 1 0 22084 0 1 1494
box 0 0 1 1
use contact_17  contact_17_205
timestamp 1643593061
transform 1 0 22082 0 1 1498
box 0 0 1 1
use contact_13  contact_13_261
timestamp 1643593061
transform 1 0 22085 0 1 1501
box 0 0 1 1
use contact_21  contact_21_261
timestamp 1643593061
transform 1 0 22089 0 1 1483
box 0 0 1 1
use contact_13  contact_13_262
timestamp 1643593061
transform 1 0 21749 0 1 1501
box 0 0 1 1
use contact_21  contact_21_262
timestamp 1643593061
transform 1 0 21753 0 1 1483
box 0 0 1 1
use contact_13  contact_13_263
timestamp 1643593061
transform 1 0 21413 0 1 1501
box 0 0 1 1
use contact_21  contact_21_263
timestamp 1643593061
transform 1 0 21417 0 1 1483
box 0 0 1 1
use contact_13  contact_13_264
timestamp 1643593061
transform 1 0 21077 0 1 1501
box 0 0 1 1
use contact_21  contact_21_264
timestamp 1643593061
transform 1 0 21081 0 1 1483
box 0 0 1 1
use contact_13  contact_13_265
timestamp 1643593061
transform 1 0 20741 0 1 1501
box 0 0 1 1
use contact_21  contact_21_265
timestamp 1643593061
transform 1 0 20745 0 1 1483
box 0 0 1 1
use contact_18  contact_18_54
timestamp 1643593061
transform 1 0 20404 0 1 1494
box 0 0 1 1
use contact_17  contact_17_206
timestamp 1643593061
transform 1 0 20402 0 1 1498
box 0 0 1 1
use contact_13  contact_13_266
timestamp 1643593061
transform 1 0 20405 0 1 1501
box 0 0 1 1
use contact_21  contact_21_266
timestamp 1643593061
transform 1 0 20409 0 1 1483
box 0 0 1 1
use contact_13  contact_13_267
timestamp 1643593061
transform 1 0 20069 0 1 1501
box 0 0 1 1
use contact_21  contact_21_267
timestamp 1643593061
transform 1 0 20073 0 1 1483
box 0 0 1 1
use contact_13  contact_13_268
timestamp 1643593061
transform 1 0 19733 0 1 1501
box 0 0 1 1
use contact_21  contact_21_268
timestamp 1643593061
transform 1 0 19737 0 1 1483
box 0 0 1 1
use contact_13  contact_13_269
timestamp 1643593061
transform 1 0 19397 0 1 1501
box 0 0 1 1
use contact_21  contact_21_269
timestamp 1643593061
transform 1 0 19401 0 1 1483
box 0 0 1 1
use contact_13  contact_13_270
timestamp 1643593061
transform 1 0 19061 0 1 1501
box 0 0 1 1
use contact_21  contact_21_270
timestamp 1643593061
transform 1 0 19065 0 1 1483
box 0 0 1 1
use contact_18  contact_18_55
timestamp 1643593061
transform 1 0 18724 0 1 1494
box 0 0 1 1
use contact_17  contact_17_207
timestamp 1643593061
transform 1 0 18722 0 1 1498
box 0 0 1 1
use contact_13  contact_13_271
timestamp 1643593061
transform 1 0 18725 0 1 1501
box 0 0 1 1
use contact_21  contact_21_271
timestamp 1643593061
transform 1 0 18729 0 1 1483
box 0 0 1 1
use contact_13  contact_13_272
timestamp 1643593061
transform 1 0 18389 0 1 1501
box 0 0 1 1
use contact_21  contact_21_272
timestamp 1643593061
transform 1 0 18393 0 1 1483
box 0 0 1 1
use contact_13  contact_13_273
timestamp 1643593061
transform 1 0 18053 0 1 1501
box 0 0 1 1
use contact_21  contact_21_273
timestamp 1643593061
transform 1 0 18057 0 1 1483
box 0 0 1 1
use contact_13  contact_13_274
timestamp 1643593061
transform 1 0 17717 0 1 1501
box 0 0 1 1
use contact_21  contact_21_274
timestamp 1643593061
transform 1 0 17721 0 1 1483
box 0 0 1 1
use contact_13  contact_13_275
timestamp 1643593061
transform 1 0 17381 0 1 1501
box 0 0 1 1
use contact_21  contact_21_275
timestamp 1643593061
transform 1 0 17385 0 1 1483
box 0 0 1 1
use contact_18  contact_18_56
timestamp 1643593061
transform 1 0 17044 0 1 1494
box 0 0 1 1
use contact_17  contact_17_208
timestamp 1643593061
transform 1 0 17042 0 1 1498
box 0 0 1 1
use contact_13  contact_13_276
timestamp 1643593061
transform 1 0 17045 0 1 1501
box 0 0 1 1
use contact_21  contact_21_276
timestamp 1643593061
transform 1 0 17049 0 1 1483
box 0 0 1 1
use contact_13  contact_13_277
timestamp 1643593061
transform 1 0 16709 0 1 1501
box 0 0 1 1
use contact_21  contact_21_277
timestamp 1643593061
transform 1 0 16713 0 1 1483
box 0 0 1 1
use contact_13  contact_13_278
timestamp 1643593061
transform 1 0 16373 0 1 1501
box 0 0 1 1
use contact_21  contact_21_278
timestamp 1643593061
transform 1 0 16377 0 1 1483
box 0 0 1 1
use contact_13  contact_13_279
timestamp 1643593061
transform 1 0 16037 0 1 1501
box 0 0 1 1
use contact_21  contact_21_279
timestamp 1643593061
transform 1 0 16041 0 1 1483
box 0 0 1 1
use contact_13  contact_13_280
timestamp 1643593061
transform 1 0 15701 0 1 1501
box 0 0 1 1
use contact_21  contact_21_280
timestamp 1643593061
transform 1 0 15705 0 1 1483
box 0 0 1 1
use contact_18  contact_18_57
timestamp 1643593061
transform 1 0 15364 0 1 1494
box 0 0 1 1
use contact_17  contact_17_209
timestamp 1643593061
transform 1 0 15362 0 1 1498
box 0 0 1 1
use contact_13  contact_13_281
timestamp 1643593061
transform 1 0 15365 0 1 1501
box 0 0 1 1
use contact_21  contact_21_281
timestamp 1643593061
transform 1 0 15369 0 1 1483
box 0 0 1 1
use contact_13  contact_13_282
timestamp 1643593061
transform 1 0 15029 0 1 1501
box 0 0 1 1
use contact_21  contact_21_282
timestamp 1643593061
transform 1 0 15033 0 1 1483
box 0 0 1 1
use contact_13  contact_13_283
timestamp 1643593061
transform 1 0 14693 0 1 1501
box 0 0 1 1
use contact_21  contact_21_283
timestamp 1643593061
transform 1 0 14697 0 1 1483
box 0 0 1 1
use contact_13  contact_13_284
timestamp 1643593061
transform 1 0 14357 0 1 1501
box 0 0 1 1
use contact_21  contact_21_284
timestamp 1643593061
transform 1 0 14361 0 1 1483
box 0 0 1 1
use contact_13  contact_13_285
timestamp 1643593061
transform 1 0 14021 0 1 1501
box 0 0 1 1
use contact_21  contact_21_285
timestamp 1643593061
transform 1 0 14025 0 1 1483
box 0 0 1 1
use contact_18  contact_18_58
timestamp 1643593061
transform 1 0 13684 0 1 1494
box 0 0 1 1
use contact_17  contact_17_210
timestamp 1643593061
transform 1 0 13682 0 1 1498
box 0 0 1 1
use contact_13  contact_13_286
timestamp 1643593061
transform 1 0 13685 0 1 1501
box 0 0 1 1
use contact_21  contact_21_286
timestamp 1643593061
transform 1 0 13689 0 1 1483
box 0 0 1 1
use contact_13  contact_13_287
timestamp 1643593061
transform 1 0 13349 0 1 1501
box 0 0 1 1
use contact_21  contact_21_287
timestamp 1643593061
transform 1 0 13353 0 1 1483
box 0 0 1 1
use contact_13  contact_13_288
timestamp 1643593061
transform 1 0 13013 0 1 1501
box 0 0 1 1
use contact_21  contact_21_288
timestamp 1643593061
transform 1 0 13017 0 1 1483
box 0 0 1 1
use contact_13  contact_13_289
timestamp 1643593061
transform 1 0 12677 0 1 1501
box 0 0 1 1
use contact_21  contact_21_289
timestamp 1643593061
transform 1 0 12681 0 1 1483
box 0 0 1 1
use contact_13  contact_13_290
timestamp 1643593061
transform 1 0 12341 0 1 1501
box 0 0 1 1
use contact_21  contact_21_290
timestamp 1643593061
transform 1 0 12345 0 1 1483
box 0 0 1 1
use contact_18  contact_18_59
timestamp 1643593061
transform 1 0 12004 0 1 1494
box 0 0 1 1
use contact_17  contact_17_211
timestamp 1643593061
transform 1 0 12002 0 1 1498
box 0 0 1 1
use contact_13  contact_13_291
timestamp 1643593061
transform 1 0 12005 0 1 1501
box 0 0 1 1
use contact_21  contact_21_291
timestamp 1643593061
transform 1 0 12009 0 1 1483
box 0 0 1 1
use contact_13  contact_13_292
timestamp 1643593061
transform 1 0 11669 0 1 1501
box 0 0 1 1
use contact_21  contact_21_292
timestamp 1643593061
transform 1 0 11673 0 1 1483
box 0 0 1 1
use contact_13  contact_13_293
timestamp 1643593061
transform 1 0 11333 0 1 1501
box 0 0 1 1
use contact_21  contact_21_293
timestamp 1643593061
transform 1 0 11337 0 1 1483
box 0 0 1 1
use contact_13  contact_13_294
timestamp 1643593061
transform 1 0 10997 0 1 1501
box 0 0 1 1
use contact_21  contact_21_294
timestamp 1643593061
transform 1 0 11001 0 1 1483
box 0 0 1 1
use contact_13  contact_13_295
timestamp 1643593061
transform 1 0 10661 0 1 1501
box 0 0 1 1
use contact_21  contact_21_295
timestamp 1643593061
transform 1 0 10665 0 1 1483
box 0 0 1 1
use contact_18  contact_18_60
timestamp 1643593061
transform 1 0 10324 0 1 1494
box 0 0 1 1
use contact_17  contact_17_212
timestamp 1643593061
transform 1 0 10322 0 1 1498
box 0 0 1 1
use contact_13  contact_13_296
timestamp 1643593061
transform 1 0 10325 0 1 1501
box 0 0 1 1
use contact_21  contact_21_296
timestamp 1643593061
transform 1 0 10329 0 1 1483
box 0 0 1 1
use contact_13  contact_13_297
timestamp 1643593061
transform 1 0 9989 0 1 1501
box 0 0 1 1
use contact_21  contact_21_297
timestamp 1643593061
transform 1 0 9993 0 1 1483
box 0 0 1 1
use contact_13  contact_13_298
timestamp 1643593061
transform 1 0 9653 0 1 1501
box 0 0 1 1
use contact_21  contact_21_298
timestamp 1643593061
transform 1 0 9657 0 1 1483
box 0 0 1 1
use contact_13  contact_13_299
timestamp 1643593061
transform 1 0 9317 0 1 1501
box 0 0 1 1
use contact_21  contact_21_299
timestamp 1643593061
transform 1 0 9321 0 1 1483
box 0 0 1 1
use contact_13  contact_13_300
timestamp 1643593061
transform 1 0 8981 0 1 1501
box 0 0 1 1
use contact_21  contact_21_300
timestamp 1643593061
transform 1 0 8985 0 1 1483
box 0 0 1 1
use contact_18  contact_18_61
timestamp 1643593061
transform 1 0 8644 0 1 1494
box 0 0 1 1
use contact_17  contact_17_213
timestamp 1643593061
transform 1 0 8642 0 1 1498
box 0 0 1 1
use contact_13  contact_13_301
timestamp 1643593061
transform 1 0 8645 0 1 1501
box 0 0 1 1
use contact_21  contact_21_301
timestamp 1643593061
transform 1 0 8649 0 1 1483
box 0 0 1 1
use contact_13  contact_13_302
timestamp 1643593061
transform 1 0 8309 0 1 1501
box 0 0 1 1
use contact_21  contact_21_302
timestamp 1643593061
transform 1 0 8313 0 1 1483
box 0 0 1 1
use contact_13  contact_13_303
timestamp 1643593061
transform 1 0 7973 0 1 1501
box 0 0 1 1
use contact_21  contact_21_303
timestamp 1643593061
transform 1 0 7977 0 1 1483
box 0 0 1 1
use contact_13  contact_13_304
timestamp 1643593061
transform 1 0 7637 0 1 1501
box 0 0 1 1
use contact_21  contact_21_304
timestamp 1643593061
transform 1 0 7641 0 1 1483
box 0 0 1 1
use contact_13  contact_13_305
timestamp 1643593061
transform 1 0 7301 0 1 1501
box 0 0 1 1
use contact_21  contact_21_305
timestamp 1643593061
transform 1 0 7305 0 1 1483
box 0 0 1 1
use contact_18  contact_18_62
timestamp 1643593061
transform 1 0 6964 0 1 1494
box 0 0 1 1
use contact_17  contact_17_214
timestamp 1643593061
transform 1 0 6962 0 1 1498
box 0 0 1 1
use contact_13  contact_13_306
timestamp 1643593061
transform 1 0 6965 0 1 1501
box 0 0 1 1
use contact_21  contact_21_306
timestamp 1643593061
transform 1 0 6969 0 1 1483
box 0 0 1 1
use contact_13  contact_13_307
timestamp 1643593061
transform 1 0 6629 0 1 1501
box 0 0 1 1
use contact_21  contact_21_307
timestamp 1643593061
transform 1 0 6633 0 1 1483
box 0 0 1 1
use contact_13  contact_13_308
timestamp 1643593061
transform 1 0 6293 0 1 1501
box 0 0 1 1
use contact_21  contact_21_308
timestamp 1643593061
transform 1 0 6297 0 1 1483
box 0 0 1 1
use contact_13  contact_13_309
timestamp 1643593061
transform 1 0 5957 0 1 1501
box 0 0 1 1
use contact_21  contact_21_309
timestamp 1643593061
transform 1 0 5961 0 1 1483
box 0 0 1 1
use contact_13  contact_13_310
timestamp 1643593061
transform 1 0 5621 0 1 1501
box 0 0 1 1
use contact_21  contact_21_310
timestamp 1643593061
transform 1 0 5625 0 1 1483
box 0 0 1 1
use contact_18  contact_18_63
timestamp 1643593061
transform 1 0 5284 0 1 1494
box 0 0 1 1
use contact_17  contact_17_215
timestamp 1643593061
transform 1 0 5282 0 1 1498
box 0 0 1 1
use contact_13  contact_13_311
timestamp 1643593061
transform 1 0 5285 0 1 1501
box 0 0 1 1
use contact_21  contact_21_311
timestamp 1643593061
transform 1 0 5289 0 1 1483
box 0 0 1 1
use contact_13  contact_13_312
timestamp 1643593061
transform 1 0 4949 0 1 1501
box 0 0 1 1
use contact_21  contact_21_312
timestamp 1643593061
transform 1 0 4953 0 1 1483
box 0 0 1 1
use contact_13  contact_13_313
timestamp 1643593061
transform 1 0 4613 0 1 1501
box 0 0 1 1
use contact_21  contact_21_313
timestamp 1643593061
transform 1 0 4617 0 1 1483
box 0 0 1 1
use contact_13  contact_13_314
timestamp 1643593061
transform 1 0 4277 0 1 1501
box 0 0 1 1
use contact_21  contact_21_314
timestamp 1643593061
transform 1 0 4281 0 1 1483
box 0 0 1 1
use contact_13  contact_13_315
timestamp 1643593061
transform 1 0 3941 0 1 1501
box 0 0 1 1
use contact_21  contact_21_315
timestamp 1643593061
transform 1 0 3945 0 1 1483
box 0 0 1 1
use contact_18  contact_18_64
timestamp 1643593061
transform 1 0 3604 0 1 1494
box 0 0 1 1
use contact_17  contact_17_216
timestamp 1643593061
transform 1 0 3602 0 1 1498
box 0 0 1 1
use contact_13  contact_13_316
timestamp 1643593061
transform 1 0 3605 0 1 1501
box 0 0 1 1
use contact_21  contact_21_316
timestamp 1643593061
transform 1 0 3609 0 1 1483
box 0 0 1 1
use contact_13  contact_13_317
timestamp 1643593061
transform 1 0 3269 0 1 1501
box 0 0 1 1
use contact_21  contact_21_317
timestamp 1643593061
transform 1 0 3273 0 1 1483
box 0 0 1 1
use contact_13  contact_13_318
timestamp 1643593061
transform 1 0 2933 0 1 1501
box 0 0 1 1
use contact_21  contact_21_318
timestamp 1643593061
transform 1 0 2937 0 1 1483
box 0 0 1 1
use contact_13  contact_13_319
timestamp 1643593061
transform 1 0 2597 0 1 1501
box 0 0 1 1
use contact_21  contact_21_319
timestamp 1643593061
transform 1 0 2601 0 1 1483
box 0 0 1 1
use contact_13  contact_13_320
timestamp 1643593061
transform 1 0 2261 0 1 1501
box 0 0 1 1
use contact_21  contact_21_320
timestamp 1643593061
transform 1 0 2265 0 1 1483
box 0 0 1 1
use contact_18  contact_18_65
timestamp 1643593061
transform 1 0 1924 0 1 1494
box 0 0 1 1
use contact_17  contact_17_217
timestamp 1643593061
transform 1 0 1922 0 1 1498
box 0 0 1 1
use contact_13  contact_13_321
timestamp 1643593061
transform 1 0 1925 0 1 1501
box 0 0 1 1
use contact_21  contact_21_321
timestamp 1643593061
transform 1 0 1929 0 1 1483
box 0 0 1 1
use contact_18  contact_18_66
timestamp 1643593061
transform 1 0 8277 0 1 13270
box 0 0 1 1
use contact_18  contact_18_67
timestamp 1643593061
transform 1 0 8277 0 1 12086
box 0 0 1 1
use contact_18  contact_18_68
timestamp 1643593061
transform 1 0 8277 0 1 11594
box 0 0 1 1
use contact_18  contact_18_69
timestamp 1643593061
transform 1 0 8277 0 1 10410
box 0 0 1 1
use contact_18  contact_18_70
timestamp 1643593061
transform 1 0 8277 0 1 9918
box 0 0 1 1
use contact_18  contact_18_71
timestamp 1643593061
transform 1 0 8277 0 1 8734
box 0 0 1 1
use contact_18  contact_18_72
timestamp 1643593061
transform 1 0 21632 0 1 6912
box 0 0 1 1
use contact_18  contact_18_73
timestamp 1643593061
transform 1 0 21632 0 1 6912
box 0 0 1 1
use contact_18  contact_18_74
timestamp 1643593061
transform 1 0 21172 0 1 6912
box 0 0 1 1
use contact_18  contact_18_75
timestamp 1643593061
transform 1 0 21172 0 1 6912
box 0 0 1 1
use contact_18  contact_18_76
timestamp 1643593061
transform 1 0 12723 0 1 2580
box 0 0 1 1
use contact_18  contact_18_77
timestamp 1643593061
transform 1 0 11241 0 1 2580
box 0 0 1 1
use contact_18  contact_18_78
timestamp 1643593061
transform 1 0 6157 0 1 3549
box 0 0 1 1
use contact_18  contact_18_79
timestamp 1643593061
transform 1 0 2635 0 1 3764
box 0 0 1 1
use contact_18  contact_18_80
timestamp 1643593061
transform 1 0 2635 0 1 2580
box 0 0 1 1
use contact_18  contact_18_81
timestamp 1643593061
transform 1 0 10172 0 1 13274
box 0 0 1 1
use contact_18  contact_18_82
timestamp 1643593061
transform 1 0 9357 0 1 13274
box 0 0 1 1
use contact_18  contact_18_83
timestamp 1643593061
transform 1 0 10088 0 1 12082
box 0 0 1 1
use contact_18  contact_18_84
timestamp 1643593061
transform 1 0 9357 0 1 12082
box 0 0 1 1
use contact_18  contact_18_85
timestamp 1643593061
transform 1 0 10004 0 1 11598
box 0 0 1 1
use contact_18  contact_18_86
timestamp 1643593061
transform 1 0 9357 0 1 11598
box 0 0 1 1
use contact_18  contact_18_87
timestamp 1643593061
transform 1 0 9920 0 1 10406
box 0 0 1 1
use contact_18  contact_18_88
timestamp 1643593061
transform 1 0 9357 0 1 10406
box 0 0 1 1
use contact_18  contact_18_89
timestamp 1643593061
transform 1 0 9836 0 1 9922
box 0 0 1 1
use contact_18  contact_18_90
timestamp 1643593061
transform 1 0 9357 0 1 9922
box 0 0 1 1
use contact_18  contact_18_91
timestamp 1643593061
transform 1 0 9752 0 1 8730
box 0 0 1 1
use contact_18  contact_18_92
timestamp 1643593061
transform 1 0 9357 0 1 8730
box 0 0 1 1
use contact_18  contact_18_93
timestamp 1643593061
transform 1 0 14928 0 1 7823
box 0 0 1 1
use contact_18  contact_18_94
timestamp 1643593061
transform 1 0 9552 0 1 7823
box 0 0 1 1
use contact_18  contact_18_95
timestamp 1643593061
transform 1 0 18278 0 1 6901
box 0 0 1 1
use contact_18  contact_18_96
timestamp 1643593061
transform 1 0 9552 0 1 6901
box 0 0 1 1
use contact_18  contact_18_97
timestamp 1643593061
transform 1 0 16062 0 1 6151
box 0 0 1 1
use contact_18  contact_18_98
timestamp 1643593061
transform 1 0 9552 0 1 6151
box 0 0 1 1
use contact_26  contact_26_0
timestamp 1643593061
transform 1 0 7986 0 1 2634
box 0 0 1 1
use contact_26  contact_26_1
timestamp 1643593061
transform 1 0 7986 0 1 8788
box 0 0 1 1
use data_dff  data_dff_0
timestamp 1643593061
transform 1 0 11064 0 1 2364
box -3 -42 2964 916
use row_addr_dff  row_addr_dff_0
timestamp 1643593061
transform 1 0 8100 0 1 8518
box -3 -42 1482 6746
use control_logic_multiport  control_logic_multiport_0
timestamp 1643593061
transform 1 0 2458 0 1 2364
box -32 -42 7124 5902
use bank  bank_0
timestamp 1643593061
transform 1 0 9750 0 1 4470
box 0 0 13524 28624
<< labels >>
rlabel metal3 s 2634 2580 2694 2640 4 web
rlabel metal3 s 2634 3764 2694 3824 4 csb
rlabel metal4 s 6240 0 6300 180 4 clk
rlabel metal4 s 11280 0 11340 180 4 din0[0]
rlabel metal4 s 12720 0 12780 180 4 din0[1]
rlabel metal3 s 25560 6600 25740 6660 4 dout0[0]
rlabel metal3 s 21172 6912 21232 6972 4 dout1[0]
rlabel metal3 s 25560 6720 25740 6780 4 dout0[1]
rlabel metal3 s 21632 6912 21692 6972 4 dout1[1]
rlabel metal3 s 0 8760 180 8820 4 addr1[0]
rlabel metal3 s 0 9840 180 9900 4 addr1[1]
rlabel metal3 s 0 10440 180 10500 4 addr1[2]
rlabel metal3 s 0 11640 180 11700 4 addr1[3]
rlabel metal3 s 0 12120 180 12180 4 addr1[4]
rlabel metal3 s 0 13200 180 13260 4 addr1[5]
rlabel metal4 s 24600 840 24900 34620 4 vdd
rlabel metal4 s 840 840 1140 34620 4 vdd
rlabel metal3 s 840 840 24900 1140 4 vdd
rlabel metal3 s 840 34320 24900 34620 4 vdd
rlabel metal4 s 25200 240 25500 35220 4 gnd
rlabel metal4 s 240 240 540 35220 4 gnd
rlabel metal3 s 240 34920 25500 35220 4 gnd
rlabel metal3 s 240 240 25500 540 4 gnd
<< properties >>
string FIXED_BBOX 0 0 25740 35220
string GDS_FILE sram_0rw2r1w_2_16_sky130A.gds
string GDS_END 148712
string GDS_START 126
<< end >>
