VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO sram_0rw2r1w_16_128_sky130A
   CLASS BLOCK ;
   SIZE 606.02 BY 317.7 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  96.46 0.0 97.22 1.82 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  102.82 0.0 103.58 1.82 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  110.24 0.0 111.0 1.82 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  118.72 0.0 119.48 1.82 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  126.14 0.0 126.9 1.82 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  133.56 0.0 134.32 1.82 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  140.98 0.0 141.74 1.82 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  147.34 0.0 148.1 1.82 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  154.76 0.0 155.52 1.82 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  162.18 0.0 162.94 1.82 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  169.6 0.0 170.36 1.82 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  178.08 0.0 178.84 1.82 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  184.44 0.0 185.2 1.82 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  192.92 0.0 193.68 1.82 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  199.28 0.0 200.04 1.82 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  207.76 0.0 208.52 1.82 ;
      END
   END din0[15]
   PIN addr[0]
      DIRECTION INPUT ;
      PORT
      END
   END addr[0]
   PIN addr[1]
      DIRECTION INPUT ;
      PORT
      END
   END addr[1]
   PIN addr[2]
      DIRECTION INPUT ;
      PORT
      END
   END addr[2]
   PIN addr[3]
      DIRECTION INPUT ;
      PORT
      END
   END addr[3]
   PIN addr[4]
      DIRECTION INPUT ;
      PORT
      END
   END addr[4]
   PIN addr[5]
      DIRECTION INPUT ;
      PORT
      END
   END addr[5]
   PIN addr[6]
      DIRECTION INPUT ;
      PORT
      END
   END addr[6]
   PIN addr[7]
      DIRECTION INPUT ;
      PORT
      END
   END addr[7]
   PIN addr[8]
      DIRECTION INPUT ;
      PORT
      END
   END addr[8]
   PIN csb
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  14.125 37.105 14.785 37.435 ;
      END
   END csb
   PIN web
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  14.125 31.185 14.785 31.515 ;
      END
   END web
   PIN clk
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  30.74 0.0 31.5 1.82 ;
      END
   END clk
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  111.3 0.0 112.06 1.82 ;
      END
   END dout0[0]
   PIN dout1[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  111.3 53.185 111.96 53.515 ;
      END
   END dout1[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  127.2 0.0 127.96 1.82 ;
      END
   END dout0[1]
   PIN dout1[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  126.86 53.185 127.52 53.515 ;
      END
   END dout1[1]
   PIN dout0[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  143.1 0.0 143.86 1.82 ;
      END
   END dout0[2]
   PIN dout1[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  142.42 53.185 143.08 53.515 ;
      END
   END dout1[2]
   PIN dout0[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  157.94 0.0 158.7 1.82 ;
      END
   END dout0[3]
   PIN dout1[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  157.98 53.185 158.64 53.515 ;
      END
   END dout1[3]
   PIN dout0[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  172.78 0.0 173.54 1.82 ;
      END
   END dout0[4]
   PIN dout1[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  173.54 53.185 174.2 53.515 ;
      END
   END dout1[4]
   PIN dout0[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  189.74 0.0 190.5 1.82 ;
      END
   END dout0[5]
   PIN dout1[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  189.1 53.185 189.76 53.515 ;
      END
   END dout1[5]
   PIN dout0[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  204.58 0.0 205.34 1.82 ;
      END
   END dout0[6]
   PIN dout1[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  204.66 53.185 205.32 53.515 ;
      END
   END dout1[6]
   PIN dout0[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  219.42 0.0 220.18 1.82 ;
      END
   END dout0[7]
   PIN dout1[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  220.22 53.185 220.88 53.515 ;
      END
   END dout1[7]
   PIN dout0[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  235.32 0.0 236.08 1.82 ;
      END
   END dout0[8]
   PIN dout1[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  235.78 53.185 236.44 53.515 ;
      END
   END dout1[8]
   PIN dout0[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  252.28 0.0 253.04 1.82 ;
      END
   END dout0[9]
   PIN dout1[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  251.34 53.185 252.0 53.515 ;
      END
   END dout1[9]
   PIN dout0[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  266.06 0.0 266.82 1.82 ;
      END
   END dout0[10]
   PIN dout1[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  266.9 53.185 267.56 53.515 ;
      END
   END dout1[10]
   PIN dout0[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  281.96 0.0 282.72 1.82 ;
      END
   END dout0[11]
   PIN dout1[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  282.46 53.185 283.12 53.515 ;
      END
   END dout1[11]
   PIN dout0[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  298.92 0.0 299.68 1.82 ;
      END
   END dout0[12]
   PIN dout1[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  298.02 53.185 298.68 53.515 ;
      END
   END dout1[12]
   PIN dout0[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  312.7 0.0 313.46 1.82 ;
      END
   END dout0[13]
   PIN dout1[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  313.58 53.185 314.24 53.515 ;
      END
   END dout1[13]
   PIN dout0[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  328.6 0.0 329.36 1.82 ;
      END
   END dout0[14]
   PIN dout1[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  329.14 53.185 329.8 53.515 ;
      END
   END dout1[14]
   PIN dout0[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  344.5 0.0 345.26 1.82 ;
      END
   END dout0[15]
   PIN dout1[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  344.7 53.185 345.36 53.515 ;
      END
   END dout1[15]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met3 ;
         RECT  7.42 7.42 600.72 10.3 ;
         LAYER met3 ;
         RECT  7.42 309.52 600.72 312.4 ;
         LAYER met4 ;
         RECT  7.42 7.42 10.3 312.4 ;
         LAYER met4 ;
         RECT  597.84 7.42 600.72 312.4 ;
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met4 ;
         RECT  603.14 2.12 606.02 317.7 ;
         LAYER met4 ;
         RECT  2.12 2.12 5.0 317.7 ;
         LAYER met3 ;
         RECT  2.12 314.82 606.02 317.7 ;
         LAYER met3 ;
         RECT  2.12 2.12 606.02 5.0 ;
      END
   END gnd
   OBS
   LAYER  met1 ;
      RECT  0.62 0.62 605.4 317.08 ;
   LAYER  met2 ;
      RECT  0.62 0.62 605.4 317.08 ;
   LAYER  met3 ;
      RECT  0.62 36.505 13.525 38.035 ;
      RECT  15.385 36.505 605.4 38.035 ;
      RECT  13.525 32.115 15.385 36.505 ;
      RECT  15.385 38.035 110.7 52.585 ;
      RECT  15.385 52.585 110.7 54.115 ;
      RECT  110.7 38.035 112.56 52.585 ;
      RECT  112.56 38.035 605.4 52.585 ;
      RECT  112.56 52.585 126.26 54.115 ;
      RECT  128.12 52.585 141.82 54.115 ;
      RECT  143.68 52.585 157.38 54.115 ;
      RECT  159.24 52.585 172.94 54.115 ;
      RECT  174.8 52.585 188.5 54.115 ;
      RECT  190.36 52.585 204.06 54.115 ;
      RECT  205.92 52.585 219.62 54.115 ;
      RECT  221.48 52.585 235.18 54.115 ;
      RECT  237.04 52.585 250.74 54.115 ;
      RECT  252.6 52.585 266.3 54.115 ;
      RECT  268.16 52.585 281.86 54.115 ;
      RECT  283.72 52.585 297.42 54.115 ;
      RECT  299.28 52.585 312.98 54.115 ;
      RECT  314.84 52.585 328.54 54.115 ;
      RECT  330.4 52.585 344.1 54.115 ;
      RECT  345.96 52.585 605.4 54.115 ;
      RECT  0.62 6.82 6.82 10.9 ;
      RECT  0.62 10.9 6.82 36.505 ;
      RECT  6.82 10.9 13.525 36.505 ;
      RECT  15.385 10.9 601.32 36.505 ;
      RECT  601.32 6.82 605.4 10.9 ;
      RECT  601.32 10.9 605.4 36.505 ;
      RECT  13.525 10.9 15.385 30.585 ;
      RECT  0.62 38.035 6.82 308.92 ;
      RECT  0.62 308.92 6.82 313.0 ;
      RECT  6.82 38.035 13.525 308.92 ;
      RECT  13.525 38.035 15.385 308.92 ;
      RECT  15.385 54.115 110.7 308.92 ;
      RECT  110.7 54.115 112.56 308.92 ;
      RECT  112.56 54.115 601.32 308.92 ;
      RECT  601.32 54.115 605.4 308.92 ;
      RECT  601.32 308.92 605.4 313.0 ;
      RECT  0.62 313.0 1.52 314.22 ;
      RECT  0.62 314.22 1.52 317.08 ;
      RECT  1.52 313.0 6.82 314.22 ;
      RECT  6.82 313.0 13.525 314.22 ;
      RECT  13.525 313.0 15.385 314.22 ;
      RECT  15.385 313.0 110.7 314.22 ;
      RECT  110.7 313.0 112.56 314.22 ;
      RECT  112.56 313.0 601.32 314.22 ;
      RECT  601.32 313.0 605.4 314.22 ;
      RECT  0.62 0.62 1.52 1.52 ;
      RECT  0.62 1.52 1.52 5.6 ;
      RECT  0.62 5.6 1.52 6.82 ;
      RECT  1.52 0.62 6.82 1.52 ;
      RECT  1.52 5.6 6.82 6.82 ;
      RECT  6.82 0.62 13.525 1.52 ;
      RECT  6.82 5.6 13.525 6.82 ;
      RECT  15.385 0.62 601.32 1.52 ;
      RECT  15.385 5.6 601.32 6.82 ;
      RECT  601.32 0.62 605.4 1.52 ;
      RECT  601.32 5.6 605.4 6.82 ;
      RECT  13.525 0.62 15.385 1.52 ;
      RECT  13.525 5.6 15.385 6.82 ;
   LAYER  met4 ;
      RECT  95.86 2.42 97.82 317.08 ;
      RECT  97.82 0.62 102.22 2.42 ;
      RECT  104.18 0.62 109.64 2.42 ;
      RECT  120.08 0.62 125.54 2.42 ;
      RECT  134.92 0.62 140.38 2.42 ;
      RECT  148.7 0.62 154.16 2.42 ;
      RECT  163.54 0.62 169.0 2.42 ;
      RECT  179.44 0.62 183.84 2.42 ;
      RECT  194.28 0.62 198.68 2.42 ;
      RECT  32.1 0.62 95.86 2.42 ;
      RECT  112.66 0.62 118.12 2.42 ;
      RECT  128.56 0.62 132.96 2.42 ;
      RECT  142.34 0.62 142.5 2.42 ;
      RECT  144.46 0.62 146.74 2.42 ;
      RECT  156.12 0.62 157.34 2.42 ;
      RECT  159.3 0.62 161.58 2.42 ;
      RECT  170.96 0.62 172.18 2.42 ;
      RECT  174.14 0.62 177.48 2.42 ;
      RECT  185.8 0.62 189.14 2.42 ;
      RECT  191.1 0.62 192.32 2.42 ;
      RECT  200.64 0.62 203.98 2.42 ;
      RECT  205.94 0.62 207.16 2.42 ;
      RECT  209.12 0.62 218.82 2.42 ;
      RECT  220.78 0.62 234.72 2.42 ;
      RECT  236.68 0.62 251.68 2.42 ;
      RECT  253.64 0.62 265.46 2.42 ;
      RECT  267.42 0.62 281.36 2.42 ;
      RECT  283.32 0.62 298.32 2.42 ;
      RECT  300.28 0.62 312.1 2.42 ;
      RECT  314.06 0.62 328.0 2.42 ;
      RECT  329.96 0.62 343.9 2.42 ;
      RECT  6.82 2.42 10.9 6.82 ;
      RECT  6.82 313.0 10.9 317.08 ;
      RECT  10.9 2.42 95.86 6.82 ;
      RECT  10.9 6.82 95.86 313.0 ;
      RECT  10.9 313.0 95.86 317.08 ;
      RECT  97.82 2.42 597.24 6.82 ;
      RECT  97.82 6.82 597.24 313.0 ;
      RECT  97.82 313.0 597.24 317.08 ;
      RECT  597.24 2.42 601.32 6.82 ;
      RECT  597.24 313.0 601.32 317.08 ;
      RECT  345.86 0.62 602.54 1.52 ;
      RECT  345.86 1.52 602.54 2.42 ;
      RECT  602.54 0.62 605.4 1.52 ;
      RECT  601.32 2.42 602.54 6.82 ;
      RECT  601.32 6.82 602.54 313.0 ;
      RECT  601.32 313.0 602.54 317.08 ;
      RECT  0.62 0.62 1.52 1.52 ;
      RECT  0.62 1.52 1.52 2.42 ;
      RECT  1.52 0.62 5.6 1.52 ;
      RECT  5.6 0.62 30.14 1.52 ;
      RECT  5.6 1.52 30.14 2.42 ;
      RECT  0.62 2.42 1.52 6.82 ;
      RECT  5.6 2.42 6.82 6.82 ;
      RECT  0.62 6.82 1.52 313.0 ;
      RECT  5.6 6.82 6.82 313.0 ;
      RECT  0.62 313.0 1.52 317.08 ;
      RECT  5.6 313.0 6.82 317.08 ;
   END
END    sram_0rw2r1w_16_128_sky130A
END    LIBRARY
