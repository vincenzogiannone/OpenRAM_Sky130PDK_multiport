magic
tech sky130A
magscale 1 2
timestamp 1643593061
<< checkpaint >>
rect -1292 -1302 4272 2978
<< metal1 >>
rect 0 1702 2976 1706
rect -32 1650 -26 1702
rect 26 1650 2976 1702
rect 0 1646 2976 1650
rect 0 864 2976 868
rect -32 812 -26 864
rect 26 812 2976 864
rect 0 808 2976 812
rect 0 26 2976 30
rect -32 -26 -26 26
rect 26 -26 2976 26
rect 0 -30 2976 -26
<< via1 >>
rect -26 1650 26 1702
rect -26 812 26 864
rect -26 -26 26 26
<< metal2 >>
rect 0 866 28 1648
rect 2662 1453 2690 1481
rect 180 1416 234 1444
rect 2172 1117 2200 1145
rect 0 28 28 810
rect 2172 531 2200 559
rect 180 232 234 260
rect 2662 195 2690 223
<< via2 >>
rect -28 1702 28 1704
rect -28 1650 -26 1702
rect -26 1650 26 1702
rect 26 1650 28 1702
rect -28 1648 28 1650
rect -28 864 28 866
rect -28 812 -26 864
rect -26 812 26 864
rect 26 812 28 864
rect -28 810 28 812
rect -28 26 28 28
rect -28 -26 -26 26
rect -26 -26 26 26
rect 26 -26 28 26
rect -28 -28 28 -26
<< metal3 >>
rect -30 1704 30 1706
rect -30 1648 -28 1704
rect 28 1648 30 1704
rect -30 1646 30 1648
rect -30 866 30 868
rect -30 810 -28 866
rect 28 810 30 866
rect -30 808 30 810
rect -30 28 30 30
rect -30 -28 -28 28
rect 28 -28 30 28
rect -30 -30 30 -28
use contact_18  contact_18_0
timestamp 1643593061
transform 1 0 -30 0 1 1646
box 0 0 1 1
use contact_17  contact_17_0
timestamp 1643593061
transform 1 0 -32 0 1 1650
box 0 0 1 1
use contact_18  contact_18_1
timestamp 1643593061
transform 1 0 -30 0 1 808
box 0 0 1 1
use contact_17  contact_17_1
timestamp 1643593061
transform 1 0 -32 0 1 812
box 0 0 1 1
use contact_18  contact_18_2
timestamp 1643593061
transform 1 0 -30 0 1 -30
box 0 0 1 1
use contact_17  contact_17_2
timestamp 1643593061
transform 1 0 -32 0 1 -26
box 0 0 1 1
use contact_18  contact_18_3
timestamp 1643593061
transform 1 0 -30 0 1 808
box 0 0 1 1
use contact_17  contact_17_3
timestamp 1643593061
transform 1 0 -32 0 1 812
box 0 0 1 1
use dff_buf_0  dff_buf_0_0
timestamp 1643593061
transform 1 0 0 0 -1 1676
box 0 -42 3012 916
use dff_buf_0  dff_buf_0_1
timestamp 1643593061
transform 1 0 0 0 1 0
box 0 -42 3012 916
<< labels >>
rlabel metal3 s -30 808 30 868 4 vdd
rlabel metal3 s 0 838 0 838 4 vdd
rlabel metal3 s -30 -30 30 30 4 gnd
rlabel metal3 s -30 1646 30 1706 4 gnd
rlabel metal2 s 180 232 234 260 4 din_0
rlabel metal2 s 2662 195 2690 223 4 dout_0
rlabel metal2 s 2172 531 2200 559 4 dout_bar_0
rlabel metal2 s 180 1416 234 1444 4 din_1
rlabel metal2 s 2662 1453 2690 1481 4 dout_1
rlabel metal2 s 2172 1117 2200 1145 4 dout_bar_1
rlabel metal2 s 0 0 28 1676 4 clk
<< properties >>
string FIXED_BBOX -30 -30 30 -26
string GDS_FILE sram_0rw2r1w_2_16_sky130A.gds
string GDS_END 492072
string GDS_START 488962
<< end >>
