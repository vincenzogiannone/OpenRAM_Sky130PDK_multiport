magic
tech sky130A
magscale 1 2
timestamp 1644969367
<< checkpaint >>
rect -1319 -1316 2117 1602
<< nwell >>
rect -54 228 852 342
rect -59 60 857 228
rect -54 -54 852 60
<< scpmos >>
rect 60 0 90 288
rect 168 0 198 288
rect 276 0 306 288
rect 384 0 414 288
rect 492 0 522 288
rect 600 0 630 288
rect 708 0 738 288
<< pdiff >>
rect 0 161 60 288
rect 0 127 8 161
rect 42 127 60 161
rect 0 0 60 127
rect 90 161 168 288
rect 90 127 112 161
rect 146 127 168 161
rect 90 0 168 127
rect 198 161 276 288
rect 198 127 220 161
rect 254 127 276 161
rect 198 0 276 127
rect 306 161 384 288
rect 306 127 328 161
rect 362 127 384 161
rect 306 0 384 127
rect 414 161 492 288
rect 414 127 436 161
rect 470 127 492 161
rect 414 0 492 127
rect 522 161 600 288
rect 522 127 544 161
rect 578 127 600 161
rect 522 0 600 127
rect 630 161 708 288
rect 630 127 652 161
rect 686 127 708 161
rect 630 0 708 127
rect 738 161 798 288
rect 738 127 756 161
rect 790 127 798 161
rect 738 0 798 127
<< pdiffc >>
rect 8 127 42 161
rect 112 127 146 161
rect 220 127 254 161
rect 328 127 362 161
rect 436 127 470 161
rect 544 127 578 161
rect 652 127 686 161
rect 756 127 790 161
<< poly >>
rect 60 288 90 314
rect 168 288 198 314
rect 276 288 306 314
rect 384 288 414 314
rect 492 288 522 314
rect 600 288 630 314
rect 708 288 738 314
rect 60 -26 90 0
rect 168 -26 198 0
rect 276 -26 306 0
rect 384 -26 414 0
rect 492 -26 522 0
rect 600 -26 630 0
rect 708 -26 738 0
rect 60 -56 738 -26
<< locali >>
rect 8 161 42 177
rect 8 111 42 127
rect 112 161 146 177
rect 112 77 146 127
rect 220 161 254 177
rect 220 111 254 127
rect 328 161 362 177
rect 328 77 362 127
rect 436 161 470 177
rect 436 111 470 127
rect 544 161 578 177
rect 544 77 578 127
rect 652 161 686 177
rect 652 111 686 127
rect 756 161 790 177
rect 756 77 790 127
rect 112 43 790 77
use contact_9  contact_9_0
timestamp 1644969367
transform 1 0 748 0 1 103
box 0 0 2 2
use contact_9  contact_9_1
timestamp 1644969367
transform 1 0 644 0 1 103
box 0 0 2 2
use contact_9  contact_9_2
timestamp 1644969367
transform 1 0 536 0 1 103
box 0 0 2 2
use contact_9  contact_9_3
timestamp 1644969367
transform 1 0 428 0 1 103
box 0 0 2 2
use contact_9  contact_9_4
timestamp 1644969367
transform 1 0 320 0 1 103
box 0 0 2 2
use contact_9  contact_9_5
timestamp 1644969367
transform 1 0 212 0 1 103
box 0 0 2 2
use contact_9  contact_9_6
timestamp 1644969367
transform 1 0 104 0 1 103
box 0 0 2 2
use contact_9  contact_9_7
timestamp 1644969367
transform 1 0 0 0 1 103
box 0 0 2 2
<< labels >>
rlabel mvvaractor s 399 -41 399 -41 4 G
rlabel locali s 237 144 237 144 4 S
rlabel locali s 25 144 25 144 4 S
rlabel locali s 453 144 453 144 4 S
rlabel locali s 669 144 669 144 4 S
rlabel locali s 451 60 451 60 4 D
<< properties >>
string FIXED_BBOX -54 -56 852 60
string GDS_FILE sram_0rw2r1w_32_128_sky130A.gds
string GDS_END 3315094
string GDS_START 3313026
<< end >>
