magic
tech sky130A
magscale 1 2
timestamp 1643593061
<< checkpaint >>
rect -1296 -1277 2906 2155
<< locali >>
rect 0 821 1610 855
rect 196 497 262 563
rect 330 390 364 561
rect 330 356 459 390
rect 991 356 1025 390
rect 96 257 162 323
rect 0 -17 1610 17
use pdriver_2  pdriver_2_0
timestamp 1643593061
transform 1 0 378 0 1 0
box -36 -17 1268 895
use pnand2_0  pnand2_0_0
timestamp 1643593061
transform 1 0 0 0 1 0
box -36 -17 414 895
<< labels >>
rlabel locali s 1008 373 1008 373 4 Z
rlabel locali s 129 290 129 290 4 A
rlabel locali s 229 530 229 530 4 B
rlabel locali s 805 0 805 0 4 gnd
rlabel locali s 805 838 805 838 4 vdd
<< properties >>
string FIXED_BBOX 0 0 1610 838
string GDS_FILE sram_0rw2r1w_2_16_sky130A.gds
string GDS_END 559198
string GDS_START 558064
<< end >>
