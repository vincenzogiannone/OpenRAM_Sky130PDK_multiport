magic
tech sky130A
timestamp 1642430334
<< nwell >>
rect 0 236 349 476
<< nmos >>
rect 54 69 69 111
rect 110 69 125 111
rect 224 69 239 111
rect 280 69 295 111
<< pmos >>
rect 54 254 69 389
rect 110 254 125 389
rect 224 254 239 389
rect 280 254 295 389
<< ndiff >>
rect 18 98 54 111
rect 18 81 25 98
rect 42 81 54 98
rect 18 69 54 81
rect 69 98 110 111
rect 69 81 81 98
rect 98 81 110 98
rect 69 69 110 81
rect 125 98 161 111
rect 125 81 137 98
rect 154 81 161 98
rect 125 69 161 81
rect 188 98 224 111
rect 188 81 195 98
rect 212 81 224 98
rect 188 69 224 81
rect 239 69 280 111
rect 295 98 331 111
rect 295 81 307 98
rect 324 81 331 98
rect 295 69 331 81
<< pdiff >>
rect 18 368 54 389
rect 18 351 25 368
rect 42 351 54 368
rect 18 330 54 351
rect 18 313 25 330
rect 42 313 54 330
rect 18 292 54 313
rect 18 275 25 292
rect 42 275 54 292
rect 18 254 54 275
rect 69 368 110 389
rect 69 351 81 368
rect 98 351 110 368
rect 69 330 110 351
rect 69 313 81 330
rect 98 313 110 330
rect 69 292 110 313
rect 69 275 81 292
rect 98 275 110 292
rect 69 254 110 275
rect 125 368 161 389
rect 125 351 137 368
rect 154 351 161 368
rect 125 330 161 351
rect 125 313 137 330
rect 154 313 161 330
rect 125 292 161 313
rect 125 275 137 292
rect 154 275 161 292
rect 125 254 161 275
rect 188 368 224 389
rect 188 351 195 368
rect 212 351 224 368
rect 188 330 224 351
rect 188 313 195 330
rect 212 313 224 330
rect 188 292 224 313
rect 188 275 195 292
rect 212 275 224 292
rect 188 254 224 275
rect 239 254 280 389
rect 295 368 331 389
rect 295 351 307 368
rect 324 351 331 368
rect 295 330 331 351
rect 295 313 307 330
rect 324 313 331 330
rect 295 292 331 313
rect 295 275 307 292
rect 324 275 331 292
rect 295 254 331 275
<< ndiffc >>
rect 25 81 42 98
rect 81 81 98 98
rect 137 81 154 98
rect 195 81 212 98
rect 307 81 324 98
<< pdiffc >>
rect 25 351 42 368
rect 25 313 42 330
rect 25 275 42 292
rect 81 351 98 368
rect 81 313 98 330
rect 81 275 98 292
rect 137 351 154 368
rect 137 313 154 330
rect 137 275 154 292
rect 195 351 212 368
rect 195 313 212 330
rect 195 275 212 292
rect 307 351 324 368
rect 307 313 324 330
rect 307 275 324 292
<< psubdiff >>
rect 61 30 97 42
rect 61 12 70 30
rect 88 12 97 30
rect 61 0 97 12
rect 157 30 193 42
rect 157 12 166 30
rect 184 12 193 30
rect 157 0 193 12
rect 253 30 289 42
rect 253 12 262 30
rect 280 12 289 30
rect 253 0 289 12
<< nsubdiff >>
rect 61 446 97 458
rect 61 428 70 446
rect 88 428 97 446
rect 61 416 97 428
rect 157 446 193 458
rect 157 428 166 446
rect 184 428 193 446
rect 157 416 193 428
rect 253 446 289 458
rect 253 428 262 446
rect 280 428 289 446
rect 253 416 289 428
<< psubdiffcont >>
rect 70 12 88 30
rect 166 12 184 30
rect 262 12 280 30
<< nsubdiffcont >>
rect 70 428 88 446
rect 166 428 184 446
rect 262 428 280 446
<< poly >>
rect 54 389 69 402
rect 110 389 125 402
rect 224 389 239 402
rect 280 389 295 402
rect 54 203 69 254
rect 4 195 69 203
rect 4 178 9 195
rect 26 188 69 195
rect 26 178 31 188
rect 4 170 31 178
rect 54 111 69 188
rect 110 161 125 254
rect 224 237 239 254
rect 280 237 295 254
rect 212 229 239 237
rect 212 212 217 229
rect 234 212 239 229
rect 212 204 239 212
rect 268 229 295 237
rect 268 212 273 229
rect 290 212 295 229
rect 268 204 295 212
rect 98 153 125 161
rect 98 136 103 153
rect 120 136 125 153
rect 98 128 125 136
rect 110 111 125 128
rect 224 111 239 204
rect 268 153 295 161
rect 268 136 273 153
rect 290 136 295 153
rect 268 128 295 136
rect 280 111 295 128
rect 54 56 69 69
rect 110 56 125 69
rect 224 56 239 69
rect 280 56 295 69
<< polycont >>
rect 9 178 26 195
rect 217 212 234 229
rect 273 212 290 229
rect 103 136 120 153
rect 273 136 290 153
<< locali >>
rect 70 446 91 454
rect 88 428 91 446
rect 70 420 91 428
rect 166 446 184 454
rect 262 446 280 454
rect 184 428 205 437
rect 166 420 205 428
rect 262 420 280 428
rect 74 389 91 420
rect 188 389 205 420
rect 18 368 49 389
rect 18 351 25 368
rect 42 351 49 368
rect 18 330 49 351
rect 18 313 25 330
rect 42 313 49 330
rect 18 292 49 313
rect 18 275 25 292
rect 42 275 49 292
rect 18 254 49 275
rect 74 368 105 389
rect 74 351 81 368
rect 98 351 105 368
rect 74 330 105 351
rect 74 313 81 330
rect 98 313 105 330
rect 74 292 105 313
rect 74 275 81 292
rect 98 275 105 292
rect 74 254 105 275
rect 130 368 161 389
rect 130 351 137 368
rect 154 351 161 368
rect 130 330 161 351
rect 130 313 137 330
rect 154 313 161 330
rect 130 292 161 313
rect 130 275 137 292
rect 154 275 161 292
rect 130 254 161 275
rect 188 368 219 389
rect 188 351 195 368
rect 212 351 219 368
rect 188 330 219 351
rect 188 313 195 330
rect 212 313 219 330
rect 188 292 219 313
rect 188 275 195 292
rect 212 275 219 292
rect 188 254 219 275
rect 300 368 331 389
rect 300 351 307 368
rect 324 351 331 368
rect 300 330 331 351
rect 300 313 307 330
rect 324 313 331 330
rect 300 292 331 313
rect 300 275 307 292
rect 324 275 331 292
rect 300 254 331 275
rect 32 237 49 254
rect 32 220 69 237
rect 9 195 26 203
rect 9 170 26 178
rect 52 147 69 220
rect 144 230 161 254
rect 217 230 234 237
rect 144 229 234 230
rect 144 212 217 229
rect 32 129 69 147
rect 103 153 120 161
rect 32 111 49 129
rect 103 128 120 136
rect 144 111 161 212
rect 217 204 234 212
rect 273 229 290 237
rect 273 204 290 212
rect 273 153 290 161
rect 273 128 290 136
rect 314 153 331 254
rect 314 111 331 136
rect 18 98 49 111
rect 18 81 25 98
rect 42 81 49 98
rect 18 69 49 81
rect 74 98 105 111
rect 74 81 81 98
rect 98 81 105 98
rect 74 69 105 81
rect 130 98 161 111
rect 130 81 137 98
rect 154 81 161 98
rect 130 69 161 81
rect 188 98 219 111
rect 188 81 195 98
rect 212 81 219 98
rect 188 69 219 81
rect 300 98 331 111
rect 300 81 307 98
rect 324 81 331 98
rect 300 69 331 81
rect 74 38 91 69
rect 188 38 205 69
rect 70 30 91 38
rect 88 12 91 30
rect 70 4 91 12
rect 166 30 205 38
rect 184 21 205 30
rect 262 30 280 38
rect 166 4 184 12
rect 262 4 280 12
<< viali >>
rect 70 428 88 446
rect 166 428 184 446
rect 262 428 280 446
rect 25 275 42 292
rect 9 178 26 195
rect 103 136 120 153
rect 273 212 290 229
rect 273 136 290 153
rect 314 136 331 153
rect 70 12 88 30
rect 166 12 184 30
rect 262 12 280 30
<< metal1 >>
rect 0 446 349 452
rect 0 428 70 446
rect 88 428 166 446
rect 184 428 262 446
rect 280 428 349 446
rect 0 422 349 428
rect 22 292 45 298
rect 22 275 25 292
rect 42 283 45 292
rect 42 275 284 283
rect 22 269 284 275
rect 270 235 284 269
rect 270 229 293 235
rect 270 212 273 229
rect 290 212 293 229
rect 270 206 293 212
rect 5 195 31 202
rect 5 192 9 195
rect 4 178 9 192
rect 26 192 31 195
rect 26 178 201 192
rect 5 170 31 178
rect 98 157 125 160
rect 98 131 99 157
rect 187 159 201 178
rect 187 153 293 159
rect 187 145 273 153
rect 98 128 125 131
rect 270 136 273 145
rect 290 136 293 153
rect 270 130 293 136
rect 309 158 335 161
rect 309 129 335 132
rect 0 30 349 36
rect 0 12 70 30
rect 88 12 166 30
rect 184 12 262 30
rect 280 12 349 30
rect 0 6 349 12
<< via1 >>
rect 99 153 125 157
rect 99 136 103 153
rect 103 136 120 153
rect 120 136 125 153
rect 99 131 125 136
rect 309 153 335 158
rect 309 136 314 153
rect 314 136 331 153
rect 331 136 335 153
rect 309 132 335 136
<< metal2 >>
rect 315 161 329 476
rect 99 157 125 160
rect 98 136 99 150
rect 99 128 125 131
rect 309 158 335 161
rect 309 129 335 132
rect 315 0 329 129
<< labels >>
flabel metal2 98 143 98 143 0 FreeSans 80 0 0 0 din
port 1 nsew
flabel metal1 124 437 124 437 0 FreeSans 80 0 0 0 vdd
port 3 nsew
flabel metal1 124 20 124 20 0 FreeSans 80 0 0 0 gnd
port 4 nsew
flabel locali 38 135 38 135 0 FreeSans 80 0 0 0 enb
flabel locali 153 158 153 158 0 FreeSans 80 0 0 0 net1
flabel pdiff 260 332 260 332 0 FreeSans 80 0 0 0 net2
flabel ndiff 258 87 258 87 0 FreeSans 80 0 0 0 net3
flabel metal1 4 184 4 184 0 FreeSans 80 0 0 0 en
port 5 nsew
flabel metal2 321 184 321 184 0 FreeSans 80 0 0 0 wbl
port 6 nsew
<< properties >>
string FIXED_BBOX 0 0 349 476
<< end >>
