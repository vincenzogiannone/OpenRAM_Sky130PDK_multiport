magic
tech sky130A
magscale 1 2
timestamp 1643671299
<< checkpaint >>
rect -1319 -1316 2441 1591
<< nwell >>
rect -54 223 1176 331
rect -59 55 1181 223
rect -54 -54 1176 55
<< scpmos >>
rect 60 0 90 277
rect 168 0 198 277
rect 276 0 306 277
rect 384 0 414 277
rect 492 0 522 277
rect 600 0 630 277
rect 708 0 738 277
rect 816 0 846 277
rect 924 0 954 277
rect 1032 0 1062 277
<< pdiff >>
rect 0 156 60 277
rect 0 122 8 156
rect 42 122 60 156
rect 0 0 60 122
rect 90 156 168 277
rect 90 122 112 156
rect 146 122 168 156
rect 90 0 168 122
rect 198 156 276 277
rect 198 122 220 156
rect 254 122 276 156
rect 198 0 276 122
rect 306 156 384 277
rect 306 122 328 156
rect 362 122 384 156
rect 306 0 384 122
rect 414 156 492 277
rect 414 122 436 156
rect 470 122 492 156
rect 414 0 492 122
rect 522 156 600 277
rect 522 122 544 156
rect 578 122 600 156
rect 522 0 600 122
rect 630 156 708 277
rect 630 122 652 156
rect 686 122 708 156
rect 630 0 708 122
rect 738 156 816 277
rect 738 122 760 156
rect 794 122 816 156
rect 738 0 816 122
rect 846 156 924 277
rect 846 122 868 156
rect 902 122 924 156
rect 846 0 924 122
rect 954 156 1032 277
rect 954 122 976 156
rect 1010 122 1032 156
rect 954 0 1032 122
rect 1062 156 1122 277
rect 1062 122 1080 156
rect 1114 122 1122 156
rect 1062 0 1122 122
<< pdiffc >>
rect 8 122 42 156
rect 112 122 146 156
rect 220 122 254 156
rect 328 122 362 156
rect 436 122 470 156
rect 544 122 578 156
rect 652 122 686 156
rect 760 122 794 156
rect 868 122 902 156
rect 976 122 1010 156
rect 1080 122 1114 156
<< poly >>
rect 60 277 90 303
rect 168 277 198 303
rect 276 277 306 303
rect 384 277 414 303
rect 492 277 522 303
rect 600 277 630 303
rect 708 277 738 303
rect 816 277 846 303
rect 924 277 954 303
rect 1032 277 1062 303
rect 60 -26 90 0
rect 168 -26 198 0
rect 276 -26 306 0
rect 384 -26 414 0
rect 492 -26 522 0
rect 600 -26 630 0
rect 708 -26 738 0
rect 816 -26 846 0
rect 924 -26 954 0
rect 1032 -26 1062 0
rect 60 -56 1062 -26
<< locali >>
rect 8 156 42 172
rect 8 106 42 122
rect 112 156 146 172
rect 112 72 146 122
rect 220 156 254 172
rect 220 106 254 122
rect 328 156 362 172
rect 328 72 362 122
rect 436 156 470 172
rect 436 106 470 122
rect 544 156 578 172
rect 544 72 578 122
rect 652 156 686 172
rect 652 106 686 122
rect 760 156 794 172
rect 760 72 794 122
rect 868 156 902 172
rect 868 106 902 122
rect 976 156 1010 172
rect 976 72 1010 122
rect 1080 156 1114 172
rect 1080 106 1114 122
rect 112 38 1010 72
use contact_9  contact_9_0
timestamp 1643671299
transform 1 0 1072 0 1 98
box 0 0 2 2
use contact_9  contact_9_1
timestamp 1643671299
transform 1 0 968 0 1 98
box 0 0 2 2
use contact_9  contact_9_2
timestamp 1643671299
transform 1 0 860 0 1 98
box 0 0 2 2
use contact_9  contact_9_3
timestamp 1643671299
transform 1 0 752 0 1 98
box 0 0 2 2
use contact_9  contact_9_4
timestamp 1643671299
transform 1 0 644 0 1 98
box 0 0 2 2
use contact_9  contact_9_5
timestamp 1643671299
transform 1 0 536 0 1 98
box 0 0 2 2
use contact_9  contact_9_6
timestamp 1643671299
transform 1 0 428 0 1 98
box 0 0 2 2
use contact_9  contact_9_7
timestamp 1643671299
transform 1 0 320 0 1 98
box 0 0 2 2
use contact_9  contact_9_8
timestamp 1643671299
transform 1 0 212 0 1 98
box 0 0 2 2
use contact_9  contact_9_9
timestamp 1643671299
transform 1 0 104 0 1 98
box 0 0 2 2
use contact_9  contact_9_10
timestamp 1643671299
transform 1 0 0 0 1 98
box 0 0 2 2
<< labels >>
rlabel mvvaractor s 561 -41 561 -41 4 G
rlabel locali s 237 139 237 139 4 S
rlabel locali s 453 139 453 139 4 S
rlabel locali s 25 139 25 139 4 S
rlabel locali s 669 139 669 139 4 S
rlabel locali s 1097 139 1097 139 4 S
rlabel locali s 885 139 885 139 4 S
rlabel locali s 561 55 561 55 4 D
<< properties >>
string FIXED_BBOX -54 -56 1176 55
string GDS_FILE sram_0rw2r1w_16_32_sky130A.gds
string GDS_END 1220708
string GDS_START 1218024
<< end >>
