magic
tech sky130A
magscale 1 2
timestamp 1643671299
<< checkpaint >>
rect 3288 -1260 54316 2310
<< via1 >>
rect 4658 954 4710 1006
rect 6214 954 6266 1006
rect 7770 954 7822 1006
rect 9326 954 9378 1006
rect 10882 954 10934 1006
rect 12438 954 12490 1006
rect 13994 954 14046 1006
rect 15550 954 15602 1006
rect 17106 954 17158 1006
rect 18662 954 18714 1006
rect 20218 954 20270 1006
rect 21774 954 21826 1006
rect 23330 954 23382 1006
rect 24886 954 24938 1006
rect 26442 954 26494 1006
rect 27998 954 28050 1006
rect 29554 954 29606 1006
rect 31110 954 31162 1006
rect 32666 954 32718 1006
rect 34222 954 34274 1006
rect 35778 954 35830 1006
rect 37334 954 37386 1006
rect 38890 954 38942 1006
rect 40446 954 40498 1006
rect 42002 954 42054 1006
rect 43558 954 43610 1006
rect 45114 954 45166 1006
rect 46670 954 46722 1006
rect 48226 954 48278 1006
rect 49782 954 49834 1006
rect 51338 954 51390 1006
rect 52894 954 52946 1006
rect 4658 8 4710 60
rect 6214 8 6266 60
rect 7770 8 7822 60
rect 9326 8 9378 60
rect 10882 8 10934 60
rect 12438 8 12490 60
rect 13994 8 14046 60
rect 15550 8 15602 60
rect 17106 8 17158 60
rect 18662 8 18714 60
rect 20218 8 20270 60
rect 21774 8 21826 60
rect 23330 8 23382 60
rect 24886 8 24938 60
rect 26442 8 26494 60
rect 27998 8 28050 60
rect 29554 8 29606 60
rect 31110 8 31162 60
rect 32666 8 32718 60
rect 34222 8 34274 60
rect 35778 8 35830 60
rect 37334 8 37386 60
rect 38890 8 38942 60
rect 40446 8 40498 60
rect 42002 8 42054 60
rect 43558 8 43610 60
rect 45114 8 45166 60
rect 46670 8 46722 60
rect 48226 8 48278 60
rect 49782 8 49834 60
rect 51338 8 51390 60
rect 52894 8 52946 60
<< metal2 >>
rect 4664 1008 4704 1014
rect 6220 1008 6260 1014
rect 7776 1008 7816 1014
rect 9332 1008 9372 1014
rect 10888 1008 10928 1014
rect 12444 1008 12484 1014
rect 14000 1008 14040 1014
rect 15556 1008 15596 1014
rect 17112 1008 17152 1014
rect 18668 1008 18708 1014
rect 20224 1008 20264 1014
rect 21780 1008 21820 1014
rect 23336 1008 23376 1014
rect 24892 1008 24932 1014
rect 26448 1008 26488 1014
rect 28004 1008 28044 1014
rect 29560 1008 29600 1014
rect 31116 1008 31156 1014
rect 32672 1008 32712 1014
rect 34228 1008 34268 1014
rect 35784 1008 35824 1014
rect 37340 1008 37380 1014
rect 38896 1008 38936 1014
rect 40452 1008 40492 1014
rect 42008 1008 42048 1014
rect 43564 1008 43604 1014
rect 45120 1008 45160 1014
rect 46676 1008 46716 1014
rect 48232 1008 48272 1014
rect 49788 1008 49828 1014
rect 51344 1008 51384 1014
rect 52900 1008 52940 1014
rect 4664 946 4704 952
rect 6220 946 6260 952
rect 7776 946 7816 952
rect 9332 946 9372 952
rect 10888 946 10928 952
rect 12444 946 12484 952
rect 14000 946 14040 952
rect 15556 946 15596 952
rect 17112 946 17152 952
rect 18668 946 18708 952
rect 20224 946 20264 952
rect 21780 946 21820 952
rect 23336 946 23376 952
rect 24892 946 24932 952
rect 26448 946 26488 952
rect 28004 946 28044 952
rect 29560 946 29600 952
rect 31116 946 31156 952
rect 32672 946 32712 952
rect 34228 946 34268 952
rect 35784 946 35824 952
rect 37340 946 37380 952
rect 38896 946 38936 952
rect 40452 946 40492 952
rect 42008 946 42048 952
rect 43564 946 43604 952
rect 45120 946 45160 952
rect 46676 946 46716 952
rect 48232 946 48272 952
rect 49788 946 49828 952
rect 51344 946 51384 952
rect 52900 946 52940 952
rect 4562 0 4590 240
rect 4664 62 4704 68
rect 4664 0 4704 6
rect 4750 0 4778 240
rect 6118 0 6146 240
rect 6220 62 6260 68
rect 6220 0 6260 6
rect 6306 0 6334 240
rect 7674 0 7702 240
rect 7776 62 7816 68
rect 7776 0 7816 6
rect 7862 0 7890 240
rect 9230 0 9258 240
rect 9332 62 9372 68
rect 9332 0 9372 6
rect 9418 0 9446 240
rect 10786 0 10814 240
rect 10888 62 10928 68
rect 10888 0 10928 6
rect 10974 0 11002 240
rect 12342 0 12370 240
rect 12444 62 12484 68
rect 12444 0 12484 6
rect 12530 0 12558 240
rect 13898 0 13926 240
rect 14000 62 14040 68
rect 14000 0 14040 6
rect 14086 0 14114 240
rect 15454 0 15482 240
rect 15556 62 15596 68
rect 15556 0 15596 6
rect 15642 0 15670 240
rect 17010 0 17038 240
rect 17112 62 17152 68
rect 17112 0 17152 6
rect 17198 0 17226 240
rect 18566 0 18594 240
rect 18668 62 18708 68
rect 18668 0 18708 6
rect 18754 0 18782 240
rect 20122 0 20150 240
rect 20224 62 20264 68
rect 20224 0 20264 6
rect 20310 0 20338 240
rect 21678 0 21706 240
rect 21780 62 21820 68
rect 21780 0 21820 6
rect 21866 0 21894 240
rect 23234 0 23262 240
rect 23336 62 23376 68
rect 23336 0 23376 6
rect 23422 0 23450 240
rect 24790 0 24818 240
rect 24892 62 24932 68
rect 24892 0 24932 6
rect 24978 0 25006 240
rect 26346 0 26374 240
rect 26448 62 26488 68
rect 26448 0 26488 6
rect 26534 0 26562 240
rect 27902 0 27930 240
rect 28004 62 28044 68
rect 28004 0 28044 6
rect 28090 0 28118 240
rect 29458 0 29486 240
rect 29560 62 29600 68
rect 29560 0 29600 6
rect 29646 0 29674 240
rect 31014 0 31042 240
rect 31116 62 31156 68
rect 31116 0 31156 6
rect 31202 0 31230 240
rect 32570 0 32598 240
rect 32672 62 32712 68
rect 32672 0 32712 6
rect 32758 0 32786 240
rect 34126 0 34154 240
rect 34228 62 34268 68
rect 34228 0 34268 6
rect 34314 0 34342 240
rect 35682 0 35710 240
rect 35784 62 35824 68
rect 35784 0 35824 6
rect 35870 0 35898 240
rect 37238 0 37266 240
rect 37340 62 37380 68
rect 37340 0 37380 6
rect 37426 0 37454 240
rect 38794 0 38822 240
rect 38896 62 38936 68
rect 38896 0 38936 6
rect 38982 0 39010 240
rect 40350 0 40378 240
rect 40452 62 40492 68
rect 40452 0 40492 6
rect 40538 0 40566 240
rect 41906 0 41934 240
rect 42008 62 42048 68
rect 42008 0 42048 6
rect 42094 0 42122 240
rect 43462 0 43490 240
rect 43564 62 43604 68
rect 43564 0 43604 6
rect 43650 0 43678 240
rect 45018 0 45046 240
rect 45120 62 45160 68
rect 45120 0 45160 6
rect 45206 0 45234 240
rect 46574 0 46602 240
rect 46676 62 46716 68
rect 46676 0 46716 6
rect 46762 0 46790 240
rect 48130 0 48158 240
rect 48232 62 48272 68
rect 48232 0 48272 6
rect 48318 0 48346 240
rect 49686 0 49714 240
rect 49788 62 49828 68
rect 49788 0 49828 6
rect 49874 0 49902 240
rect 51242 0 51270 240
rect 51344 62 51384 68
rect 51344 0 51384 6
rect 51430 0 51458 240
rect 52798 0 52826 240
rect 52900 62 52940 68
rect 52900 0 52940 6
rect 52986 0 53014 240
<< via2 >>
rect 4656 1006 4712 1008
rect 4656 954 4658 1006
rect 4658 954 4710 1006
rect 4710 954 4712 1006
rect 4656 952 4712 954
rect 6212 1006 6268 1008
rect 6212 954 6214 1006
rect 6214 954 6266 1006
rect 6266 954 6268 1006
rect 6212 952 6268 954
rect 7768 1006 7824 1008
rect 7768 954 7770 1006
rect 7770 954 7822 1006
rect 7822 954 7824 1006
rect 7768 952 7824 954
rect 9324 1006 9380 1008
rect 9324 954 9326 1006
rect 9326 954 9378 1006
rect 9378 954 9380 1006
rect 9324 952 9380 954
rect 10880 1006 10936 1008
rect 10880 954 10882 1006
rect 10882 954 10934 1006
rect 10934 954 10936 1006
rect 10880 952 10936 954
rect 12436 1006 12492 1008
rect 12436 954 12438 1006
rect 12438 954 12490 1006
rect 12490 954 12492 1006
rect 12436 952 12492 954
rect 13992 1006 14048 1008
rect 13992 954 13994 1006
rect 13994 954 14046 1006
rect 14046 954 14048 1006
rect 13992 952 14048 954
rect 15548 1006 15604 1008
rect 15548 954 15550 1006
rect 15550 954 15602 1006
rect 15602 954 15604 1006
rect 15548 952 15604 954
rect 17104 1006 17160 1008
rect 17104 954 17106 1006
rect 17106 954 17158 1006
rect 17158 954 17160 1006
rect 17104 952 17160 954
rect 18660 1006 18716 1008
rect 18660 954 18662 1006
rect 18662 954 18714 1006
rect 18714 954 18716 1006
rect 18660 952 18716 954
rect 20216 1006 20272 1008
rect 20216 954 20218 1006
rect 20218 954 20270 1006
rect 20270 954 20272 1006
rect 20216 952 20272 954
rect 21772 1006 21828 1008
rect 21772 954 21774 1006
rect 21774 954 21826 1006
rect 21826 954 21828 1006
rect 21772 952 21828 954
rect 23328 1006 23384 1008
rect 23328 954 23330 1006
rect 23330 954 23382 1006
rect 23382 954 23384 1006
rect 23328 952 23384 954
rect 24884 1006 24940 1008
rect 24884 954 24886 1006
rect 24886 954 24938 1006
rect 24938 954 24940 1006
rect 24884 952 24940 954
rect 26440 1006 26496 1008
rect 26440 954 26442 1006
rect 26442 954 26494 1006
rect 26494 954 26496 1006
rect 26440 952 26496 954
rect 27996 1006 28052 1008
rect 27996 954 27998 1006
rect 27998 954 28050 1006
rect 28050 954 28052 1006
rect 27996 952 28052 954
rect 29552 1006 29608 1008
rect 29552 954 29554 1006
rect 29554 954 29606 1006
rect 29606 954 29608 1006
rect 29552 952 29608 954
rect 31108 1006 31164 1008
rect 31108 954 31110 1006
rect 31110 954 31162 1006
rect 31162 954 31164 1006
rect 31108 952 31164 954
rect 32664 1006 32720 1008
rect 32664 954 32666 1006
rect 32666 954 32718 1006
rect 32718 954 32720 1006
rect 32664 952 32720 954
rect 34220 1006 34276 1008
rect 34220 954 34222 1006
rect 34222 954 34274 1006
rect 34274 954 34276 1006
rect 34220 952 34276 954
rect 35776 1006 35832 1008
rect 35776 954 35778 1006
rect 35778 954 35830 1006
rect 35830 954 35832 1006
rect 35776 952 35832 954
rect 37332 1006 37388 1008
rect 37332 954 37334 1006
rect 37334 954 37386 1006
rect 37386 954 37388 1006
rect 37332 952 37388 954
rect 38888 1006 38944 1008
rect 38888 954 38890 1006
rect 38890 954 38942 1006
rect 38942 954 38944 1006
rect 38888 952 38944 954
rect 40444 1006 40500 1008
rect 40444 954 40446 1006
rect 40446 954 40498 1006
rect 40498 954 40500 1006
rect 40444 952 40500 954
rect 42000 1006 42056 1008
rect 42000 954 42002 1006
rect 42002 954 42054 1006
rect 42054 954 42056 1006
rect 42000 952 42056 954
rect 43556 1006 43612 1008
rect 43556 954 43558 1006
rect 43558 954 43610 1006
rect 43610 954 43612 1006
rect 43556 952 43612 954
rect 45112 1006 45168 1008
rect 45112 954 45114 1006
rect 45114 954 45166 1006
rect 45166 954 45168 1006
rect 45112 952 45168 954
rect 46668 1006 46724 1008
rect 46668 954 46670 1006
rect 46670 954 46722 1006
rect 46722 954 46724 1006
rect 46668 952 46724 954
rect 48224 1006 48280 1008
rect 48224 954 48226 1006
rect 48226 954 48278 1006
rect 48278 954 48280 1006
rect 48224 952 48280 954
rect 49780 1006 49836 1008
rect 49780 954 49782 1006
rect 49782 954 49834 1006
rect 49834 954 49836 1006
rect 49780 952 49836 954
rect 51336 1006 51392 1008
rect 51336 954 51338 1006
rect 51338 954 51390 1006
rect 51390 954 51392 1006
rect 51336 952 51392 954
rect 52892 1006 52948 1008
rect 52892 954 52894 1006
rect 52894 954 52946 1006
rect 52946 954 52948 1006
rect 52892 952 52948 954
rect 4656 60 4712 62
rect 4656 8 4658 60
rect 4658 8 4710 60
rect 4710 8 4712 60
rect 4656 6 4712 8
rect 6212 60 6268 62
rect 6212 8 6214 60
rect 6214 8 6266 60
rect 6266 8 6268 60
rect 6212 6 6268 8
rect 7768 60 7824 62
rect 7768 8 7770 60
rect 7770 8 7822 60
rect 7822 8 7824 60
rect 7768 6 7824 8
rect 9324 60 9380 62
rect 9324 8 9326 60
rect 9326 8 9378 60
rect 9378 8 9380 60
rect 9324 6 9380 8
rect 10880 60 10936 62
rect 10880 8 10882 60
rect 10882 8 10934 60
rect 10934 8 10936 60
rect 10880 6 10936 8
rect 12436 60 12492 62
rect 12436 8 12438 60
rect 12438 8 12490 60
rect 12490 8 12492 60
rect 12436 6 12492 8
rect 13992 60 14048 62
rect 13992 8 13994 60
rect 13994 8 14046 60
rect 14046 8 14048 60
rect 13992 6 14048 8
rect 15548 60 15604 62
rect 15548 8 15550 60
rect 15550 8 15602 60
rect 15602 8 15604 60
rect 15548 6 15604 8
rect 17104 60 17160 62
rect 17104 8 17106 60
rect 17106 8 17158 60
rect 17158 8 17160 60
rect 17104 6 17160 8
rect 18660 60 18716 62
rect 18660 8 18662 60
rect 18662 8 18714 60
rect 18714 8 18716 60
rect 18660 6 18716 8
rect 20216 60 20272 62
rect 20216 8 20218 60
rect 20218 8 20270 60
rect 20270 8 20272 60
rect 20216 6 20272 8
rect 21772 60 21828 62
rect 21772 8 21774 60
rect 21774 8 21826 60
rect 21826 8 21828 60
rect 21772 6 21828 8
rect 23328 60 23384 62
rect 23328 8 23330 60
rect 23330 8 23382 60
rect 23382 8 23384 60
rect 23328 6 23384 8
rect 24884 60 24940 62
rect 24884 8 24886 60
rect 24886 8 24938 60
rect 24938 8 24940 60
rect 24884 6 24940 8
rect 26440 60 26496 62
rect 26440 8 26442 60
rect 26442 8 26494 60
rect 26494 8 26496 60
rect 26440 6 26496 8
rect 27996 60 28052 62
rect 27996 8 27998 60
rect 27998 8 28050 60
rect 28050 8 28052 60
rect 27996 6 28052 8
rect 29552 60 29608 62
rect 29552 8 29554 60
rect 29554 8 29606 60
rect 29606 8 29608 60
rect 29552 6 29608 8
rect 31108 60 31164 62
rect 31108 8 31110 60
rect 31110 8 31162 60
rect 31162 8 31164 60
rect 31108 6 31164 8
rect 32664 60 32720 62
rect 32664 8 32666 60
rect 32666 8 32718 60
rect 32718 8 32720 60
rect 32664 6 32720 8
rect 34220 60 34276 62
rect 34220 8 34222 60
rect 34222 8 34274 60
rect 34274 8 34276 60
rect 34220 6 34276 8
rect 35776 60 35832 62
rect 35776 8 35778 60
rect 35778 8 35830 60
rect 35830 8 35832 60
rect 35776 6 35832 8
rect 37332 60 37388 62
rect 37332 8 37334 60
rect 37334 8 37386 60
rect 37386 8 37388 60
rect 37332 6 37388 8
rect 38888 60 38944 62
rect 38888 8 38890 60
rect 38890 8 38942 60
rect 38942 8 38944 60
rect 38888 6 38944 8
rect 40444 60 40500 62
rect 40444 8 40446 60
rect 40446 8 40498 60
rect 40498 8 40500 60
rect 40444 6 40500 8
rect 42000 60 42056 62
rect 42000 8 42002 60
rect 42002 8 42054 60
rect 42054 8 42056 60
rect 42000 6 42056 8
rect 43556 60 43612 62
rect 43556 8 43558 60
rect 43558 8 43610 60
rect 43610 8 43612 60
rect 43556 6 43612 8
rect 45112 60 45168 62
rect 45112 8 45114 60
rect 45114 8 45166 60
rect 45166 8 45168 60
rect 45112 6 45168 8
rect 46668 60 46724 62
rect 46668 8 46670 60
rect 46670 8 46722 60
rect 46722 8 46724 60
rect 46668 6 46724 8
rect 48224 60 48280 62
rect 48224 8 48226 60
rect 48226 8 48278 60
rect 48278 8 48280 60
rect 48224 6 48280 8
rect 49780 60 49836 62
rect 49780 8 49782 60
rect 49782 8 49834 60
rect 49834 8 49836 60
rect 49780 6 49836 8
rect 51336 60 51392 62
rect 51336 8 51338 60
rect 51338 8 51390 60
rect 51390 8 51392 60
rect 51336 6 51392 8
rect 52892 60 52948 62
rect 52892 8 52894 60
rect 52894 8 52946 60
rect 52946 8 52948 60
rect 52892 6 52948 8
<< metal3 >>
rect 4654 1008 4714 1010
rect 4654 952 4656 1008
rect 4712 952 4714 1008
rect 4654 950 4714 952
rect 6210 1008 6270 1010
rect 6210 952 6212 1008
rect 6268 952 6270 1008
rect 6210 950 6270 952
rect 7766 1008 7826 1010
rect 7766 952 7768 1008
rect 7824 952 7826 1008
rect 7766 950 7826 952
rect 9322 1008 9382 1010
rect 9322 952 9324 1008
rect 9380 952 9382 1008
rect 9322 950 9382 952
rect 10878 1008 10938 1010
rect 10878 952 10880 1008
rect 10936 952 10938 1008
rect 10878 950 10938 952
rect 12434 1008 12494 1010
rect 12434 952 12436 1008
rect 12492 952 12494 1008
rect 12434 950 12494 952
rect 13990 1008 14050 1010
rect 13990 952 13992 1008
rect 14048 952 14050 1008
rect 13990 950 14050 952
rect 15546 1008 15606 1010
rect 15546 952 15548 1008
rect 15604 952 15606 1008
rect 15546 950 15606 952
rect 17102 1008 17162 1010
rect 17102 952 17104 1008
rect 17160 952 17162 1008
rect 17102 950 17162 952
rect 18658 1008 18718 1010
rect 18658 952 18660 1008
rect 18716 952 18718 1008
rect 18658 950 18718 952
rect 20214 1008 20274 1010
rect 20214 952 20216 1008
rect 20272 952 20274 1008
rect 20214 950 20274 952
rect 21770 1008 21830 1010
rect 21770 952 21772 1008
rect 21828 952 21830 1008
rect 21770 950 21830 952
rect 23326 1008 23386 1010
rect 23326 952 23328 1008
rect 23384 952 23386 1008
rect 23326 950 23386 952
rect 24882 1008 24942 1010
rect 24882 952 24884 1008
rect 24940 952 24942 1008
rect 24882 950 24942 952
rect 26438 1008 26498 1010
rect 26438 952 26440 1008
rect 26496 952 26498 1008
rect 26438 950 26498 952
rect 27994 1008 28054 1010
rect 27994 952 27996 1008
rect 28052 952 28054 1008
rect 27994 950 28054 952
rect 29550 1008 29610 1010
rect 29550 952 29552 1008
rect 29608 952 29610 1008
rect 29550 950 29610 952
rect 31106 1008 31166 1010
rect 31106 952 31108 1008
rect 31164 952 31166 1008
rect 31106 950 31166 952
rect 32662 1008 32722 1010
rect 32662 952 32664 1008
rect 32720 952 32722 1008
rect 32662 950 32722 952
rect 34218 1008 34278 1010
rect 34218 952 34220 1008
rect 34276 952 34278 1008
rect 34218 950 34278 952
rect 35774 1008 35834 1010
rect 35774 952 35776 1008
rect 35832 952 35834 1008
rect 35774 950 35834 952
rect 37330 1008 37390 1010
rect 37330 952 37332 1008
rect 37388 952 37390 1008
rect 37330 950 37390 952
rect 38886 1008 38946 1010
rect 38886 952 38888 1008
rect 38944 952 38946 1008
rect 38886 950 38946 952
rect 40442 1008 40502 1010
rect 40442 952 40444 1008
rect 40500 952 40502 1008
rect 40442 950 40502 952
rect 41998 1008 42058 1010
rect 41998 952 42000 1008
rect 42056 952 42058 1008
rect 41998 950 42058 952
rect 43554 1008 43614 1010
rect 43554 952 43556 1008
rect 43612 952 43614 1008
rect 43554 950 43614 952
rect 45110 1008 45170 1010
rect 45110 952 45112 1008
rect 45168 952 45170 1008
rect 45110 950 45170 952
rect 46666 1008 46726 1010
rect 46666 952 46668 1008
rect 46724 952 46726 1008
rect 46666 950 46726 952
rect 48222 1008 48282 1010
rect 48222 952 48224 1008
rect 48280 952 48282 1008
rect 48222 950 48282 952
rect 49778 1008 49838 1010
rect 49778 952 49780 1008
rect 49836 952 49838 1008
rect 49778 950 49838 952
rect 51334 1008 51394 1010
rect 51334 952 51336 1008
rect 51392 952 51394 1008
rect 51334 950 51394 952
rect 52890 1008 52950 1010
rect 52890 952 52892 1008
rect 52948 952 52950 1008
rect 52890 950 52950 952
rect 4654 62 4714 64
rect 4654 6 4656 62
rect 4712 6 4714 62
rect 4654 4 4714 6
rect 6210 62 6270 64
rect 6210 6 6212 62
rect 6268 6 6270 62
rect 6210 4 6270 6
rect 7766 62 7826 64
rect 7766 6 7768 62
rect 7824 6 7826 62
rect 7766 4 7826 6
rect 9322 62 9382 64
rect 9322 6 9324 62
rect 9380 6 9382 62
rect 9322 4 9382 6
rect 10878 62 10938 64
rect 10878 6 10880 62
rect 10936 6 10938 62
rect 10878 4 10938 6
rect 12434 62 12494 64
rect 12434 6 12436 62
rect 12492 6 12494 62
rect 12434 4 12494 6
rect 13990 62 14050 64
rect 13990 6 13992 62
rect 14048 6 14050 62
rect 13990 4 14050 6
rect 15546 62 15606 64
rect 15546 6 15548 62
rect 15604 6 15606 62
rect 15546 4 15606 6
rect 17102 62 17162 64
rect 17102 6 17104 62
rect 17160 6 17162 62
rect 17102 4 17162 6
rect 18658 62 18718 64
rect 18658 6 18660 62
rect 18716 6 18718 62
rect 18658 4 18718 6
rect 20214 62 20274 64
rect 20214 6 20216 62
rect 20272 6 20274 62
rect 20214 4 20274 6
rect 21770 62 21830 64
rect 21770 6 21772 62
rect 21828 6 21830 62
rect 21770 4 21830 6
rect 23326 62 23386 64
rect 23326 6 23328 62
rect 23384 6 23386 62
rect 23326 4 23386 6
rect 24882 62 24942 64
rect 24882 6 24884 62
rect 24940 6 24942 62
rect 24882 4 24942 6
rect 26438 62 26498 64
rect 26438 6 26440 62
rect 26496 6 26498 62
rect 26438 4 26498 6
rect 27994 62 28054 64
rect 27994 6 27996 62
rect 28052 6 28054 62
rect 27994 4 28054 6
rect 29550 62 29610 64
rect 29550 6 29552 62
rect 29608 6 29610 62
rect 29550 4 29610 6
rect 31106 62 31166 64
rect 31106 6 31108 62
rect 31164 6 31166 62
rect 31106 4 31166 6
rect 32662 62 32722 64
rect 32662 6 32664 62
rect 32720 6 32722 62
rect 32662 4 32722 6
rect 34218 62 34278 64
rect 34218 6 34220 62
rect 34276 6 34278 62
rect 34218 4 34278 6
rect 35774 62 35834 64
rect 35774 6 35776 62
rect 35832 6 35834 62
rect 35774 4 35834 6
rect 37330 62 37390 64
rect 37330 6 37332 62
rect 37388 6 37390 62
rect 37330 4 37390 6
rect 38886 62 38946 64
rect 38886 6 38888 62
rect 38944 6 38946 62
rect 38886 4 38946 6
rect 40442 62 40502 64
rect 40442 6 40444 62
rect 40500 6 40502 62
rect 40442 4 40502 6
rect 41998 62 42058 64
rect 41998 6 42000 62
rect 42056 6 42058 62
rect 41998 4 42058 6
rect 43554 62 43614 64
rect 43554 6 43556 62
rect 43612 6 43614 62
rect 43554 4 43614 6
rect 45110 62 45170 64
rect 45110 6 45112 62
rect 45168 6 45170 62
rect 45110 4 45170 6
rect 46666 62 46726 64
rect 46666 6 46668 62
rect 46724 6 46726 62
rect 46666 4 46726 6
rect 48222 62 48282 64
rect 48222 6 48224 62
rect 48280 6 48282 62
rect 48222 4 48282 6
rect 49778 62 49838 64
rect 49778 6 49780 62
rect 49836 6 49838 62
rect 49778 4 49838 6
rect 51334 62 51394 64
rect 51334 6 51336 62
rect 51392 6 51394 62
rect 51334 4 51394 6
rect 52890 62 52950 64
rect 52890 6 52892 62
rect 52948 6 52950 62
rect 52890 4 52950 6
use contact_18  contact_18_0
timestamp 1643671299
transform 1 0 52890 0 1 950
box 0 0 1 1
use contact_17  contact_17_0
timestamp 1643671299
transform 1 0 52905 0 1 965
box 0 0 1 1
use contact_18  contact_18_1
timestamp 1643671299
transform 1 0 52890 0 1 4
box 0 0 1 1
use contact_17  contact_17_1
timestamp 1643671299
transform 1 0 52905 0 1 19
box 0 0 1 1
use contact_18  contact_18_2
timestamp 1643671299
transform 1 0 51334 0 1 950
box 0 0 1 1
use contact_17  contact_17_2
timestamp 1643671299
transform 1 0 51349 0 1 965
box 0 0 1 1
use contact_18  contact_18_3
timestamp 1643671299
transform 1 0 51334 0 1 4
box 0 0 1 1
use contact_17  contact_17_3
timestamp 1643671299
transform 1 0 51349 0 1 19
box 0 0 1 1
use contact_18  contact_18_4
timestamp 1643671299
transform 1 0 49778 0 1 950
box 0 0 1 1
use contact_17  contact_17_4
timestamp 1643671299
transform 1 0 49793 0 1 965
box 0 0 1 1
use contact_18  contact_18_5
timestamp 1643671299
transform 1 0 49778 0 1 4
box 0 0 1 1
use contact_17  contact_17_5
timestamp 1643671299
transform 1 0 49793 0 1 19
box 0 0 1 1
use contact_18  contact_18_6
timestamp 1643671299
transform 1 0 48222 0 1 950
box 0 0 1 1
use contact_17  contact_17_6
timestamp 1643671299
transform 1 0 48237 0 1 965
box 0 0 1 1
use contact_18  contact_18_7
timestamp 1643671299
transform 1 0 48222 0 1 4
box 0 0 1 1
use contact_17  contact_17_7
timestamp 1643671299
transform 1 0 48237 0 1 19
box 0 0 1 1
use contact_18  contact_18_8
timestamp 1643671299
transform 1 0 46666 0 1 950
box 0 0 1 1
use contact_17  contact_17_8
timestamp 1643671299
transform 1 0 46681 0 1 965
box 0 0 1 1
use contact_18  contact_18_9
timestamp 1643671299
transform 1 0 46666 0 1 4
box 0 0 1 1
use contact_17  contact_17_9
timestamp 1643671299
transform 1 0 46681 0 1 19
box 0 0 1 1
use contact_18  contact_18_10
timestamp 1643671299
transform 1 0 45110 0 1 950
box 0 0 1 1
use contact_17  contact_17_10
timestamp 1643671299
transform 1 0 45125 0 1 965
box 0 0 1 1
use contact_18  contact_18_11
timestamp 1643671299
transform 1 0 45110 0 1 4
box 0 0 1 1
use contact_17  contact_17_11
timestamp 1643671299
transform 1 0 45125 0 1 19
box 0 0 1 1
use contact_18  contact_18_12
timestamp 1643671299
transform 1 0 43554 0 1 950
box 0 0 1 1
use contact_17  contact_17_12
timestamp 1643671299
transform 1 0 43569 0 1 965
box 0 0 1 1
use contact_18  contact_18_13
timestamp 1643671299
transform 1 0 43554 0 1 4
box 0 0 1 1
use contact_17  contact_17_13
timestamp 1643671299
transform 1 0 43569 0 1 19
box 0 0 1 1
use contact_18  contact_18_14
timestamp 1643671299
transform 1 0 41998 0 1 950
box 0 0 1 1
use contact_17  contact_17_14
timestamp 1643671299
transform 1 0 42013 0 1 965
box 0 0 1 1
use contact_18  contact_18_15
timestamp 1643671299
transform 1 0 41998 0 1 4
box 0 0 1 1
use contact_17  contact_17_15
timestamp 1643671299
transform 1 0 42013 0 1 19
box 0 0 1 1
use contact_18  contact_18_16
timestamp 1643671299
transform 1 0 40442 0 1 950
box 0 0 1 1
use contact_17  contact_17_16
timestamp 1643671299
transform 1 0 40457 0 1 965
box 0 0 1 1
use contact_18  contact_18_17
timestamp 1643671299
transform 1 0 40442 0 1 4
box 0 0 1 1
use contact_17  contact_17_17
timestamp 1643671299
transform 1 0 40457 0 1 19
box 0 0 1 1
use contact_18  contact_18_18
timestamp 1643671299
transform 1 0 38886 0 1 950
box 0 0 1 1
use contact_17  contact_17_18
timestamp 1643671299
transform 1 0 38901 0 1 965
box 0 0 1 1
use contact_18  contact_18_19
timestamp 1643671299
transform 1 0 38886 0 1 4
box 0 0 1 1
use contact_17  contact_17_19
timestamp 1643671299
transform 1 0 38901 0 1 19
box 0 0 1 1
use contact_18  contact_18_20
timestamp 1643671299
transform 1 0 37330 0 1 950
box 0 0 1 1
use contact_17  contact_17_20
timestamp 1643671299
transform 1 0 37345 0 1 965
box 0 0 1 1
use contact_18  contact_18_21
timestamp 1643671299
transform 1 0 37330 0 1 4
box 0 0 1 1
use contact_17  contact_17_21
timestamp 1643671299
transform 1 0 37345 0 1 19
box 0 0 1 1
use contact_18  contact_18_22
timestamp 1643671299
transform 1 0 35774 0 1 950
box 0 0 1 1
use contact_17  contact_17_22
timestamp 1643671299
transform 1 0 35789 0 1 965
box 0 0 1 1
use contact_18  contact_18_23
timestamp 1643671299
transform 1 0 35774 0 1 4
box 0 0 1 1
use contact_17  contact_17_23
timestamp 1643671299
transform 1 0 35789 0 1 19
box 0 0 1 1
use contact_18  contact_18_24
timestamp 1643671299
transform 1 0 34218 0 1 950
box 0 0 1 1
use contact_17  contact_17_24
timestamp 1643671299
transform 1 0 34233 0 1 965
box 0 0 1 1
use contact_18  contact_18_25
timestamp 1643671299
transform 1 0 34218 0 1 4
box 0 0 1 1
use contact_17  contact_17_25
timestamp 1643671299
transform 1 0 34233 0 1 19
box 0 0 1 1
use contact_18  contact_18_26
timestamp 1643671299
transform 1 0 32662 0 1 950
box 0 0 1 1
use contact_17  contact_17_26
timestamp 1643671299
transform 1 0 32677 0 1 965
box 0 0 1 1
use contact_18  contact_18_27
timestamp 1643671299
transform 1 0 32662 0 1 4
box 0 0 1 1
use contact_17  contact_17_27
timestamp 1643671299
transform 1 0 32677 0 1 19
box 0 0 1 1
use contact_18  contact_18_28
timestamp 1643671299
transform 1 0 31106 0 1 950
box 0 0 1 1
use contact_17  contact_17_28
timestamp 1643671299
transform 1 0 31121 0 1 965
box 0 0 1 1
use contact_18  contact_18_29
timestamp 1643671299
transform 1 0 31106 0 1 4
box 0 0 1 1
use contact_17  contact_17_29
timestamp 1643671299
transform 1 0 31121 0 1 19
box 0 0 1 1
use contact_18  contact_18_30
timestamp 1643671299
transform 1 0 29550 0 1 950
box 0 0 1 1
use contact_17  contact_17_30
timestamp 1643671299
transform 1 0 29565 0 1 965
box 0 0 1 1
use contact_18  contact_18_31
timestamp 1643671299
transform 1 0 29550 0 1 4
box 0 0 1 1
use contact_17  contact_17_31
timestamp 1643671299
transform 1 0 29565 0 1 19
box 0 0 1 1
use contact_18  contact_18_32
timestamp 1643671299
transform 1 0 27994 0 1 950
box 0 0 1 1
use contact_17  contact_17_32
timestamp 1643671299
transform 1 0 28009 0 1 965
box 0 0 1 1
use contact_18  contact_18_33
timestamp 1643671299
transform 1 0 27994 0 1 4
box 0 0 1 1
use contact_17  contact_17_33
timestamp 1643671299
transform 1 0 28009 0 1 19
box 0 0 1 1
use contact_18  contact_18_34
timestamp 1643671299
transform 1 0 26438 0 1 950
box 0 0 1 1
use contact_17  contact_17_34
timestamp 1643671299
transform 1 0 26453 0 1 965
box 0 0 1 1
use contact_18  contact_18_35
timestamp 1643671299
transform 1 0 26438 0 1 4
box 0 0 1 1
use contact_17  contact_17_35
timestamp 1643671299
transform 1 0 26453 0 1 19
box 0 0 1 1
use contact_18  contact_18_36
timestamp 1643671299
transform 1 0 24882 0 1 950
box 0 0 1 1
use contact_17  contact_17_36
timestamp 1643671299
transform 1 0 24897 0 1 965
box 0 0 1 1
use contact_18  contact_18_37
timestamp 1643671299
transform 1 0 24882 0 1 4
box 0 0 1 1
use contact_17  contact_17_37
timestamp 1643671299
transform 1 0 24897 0 1 19
box 0 0 1 1
use contact_18  contact_18_38
timestamp 1643671299
transform 1 0 23326 0 1 950
box 0 0 1 1
use contact_17  contact_17_38
timestamp 1643671299
transform 1 0 23341 0 1 965
box 0 0 1 1
use contact_18  contact_18_39
timestamp 1643671299
transform 1 0 23326 0 1 4
box 0 0 1 1
use contact_17  contact_17_39
timestamp 1643671299
transform 1 0 23341 0 1 19
box 0 0 1 1
use contact_18  contact_18_40
timestamp 1643671299
transform 1 0 21770 0 1 950
box 0 0 1 1
use contact_17  contact_17_40
timestamp 1643671299
transform 1 0 21785 0 1 965
box 0 0 1 1
use contact_18  contact_18_41
timestamp 1643671299
transform 1 0 21770 0 1 4
box 0 0 1 1
use contact_17  contact_17_41
timestamp 1643671299
transform 1 0 21785 0 1 19
box 0 0 1 1
use contact_18  contact_18_42
timestamp 1643671299
transform 1 0 20214 0 1 950
box 0 0 1 1
use contact_17  contact_17_42
timestamp 1643671299
transform 1 0 20229 0 1 965
box 0 0 1 1
use contact_18  contact_18_43
timestamp 1643671299
transform 1 0 20214 0 1 4
box 0 0 1 1
use contact_17  contact_17_43
timestamp 1643671299
transform 1 0 20229 0 1 19
box 0 0 1 1
use contact_18  contact_18_44
timestamp 1643671299
transform 1 0 18658 0 1 950
box 0 0 1 1
use contact_17  contact_17_44
timestamp 1643671299
transform 1 0 18673 0 1 965
box 0 0 1 1
use contact_18  contact_18_45
timestamp 1643671299
transform 1 0 18658 0 1 4
box 0 0 1 1
use contact_17  contact_17_45
timestamp 1643671299
transform 1 0 18673 0 1 19
box 0 0 1 1
use contact_18  contact_18_46
timestamp 1643671299
transform 1 0 17102 0 1 950
box 0 0 1 1
use contact_17  contact_17_46
timestamp 1643671299
transform 1 0 17117 0 1 965
box 0 0 1 1
use contact_18  contact_18_47
timestamp 1643671299
transform 1 0 17102 0 1 4
box 0 0 1 1
use contact_17  contact_17_47
timestamp 1643671299
transform 1 0 17117 0 1 19
box 0 0 1 1
use contact_18  contact_18_48
timestamp 1643671299
transform 1 0 15546 0 1 950
box 0 0 1 1
use contact_17  contact_17_48
timestamp 1643671299
transform 1 0 15561 0 1 965
box 0 0 1 1
use contact_18  contact_18_49
timestamp 1643671299
transform 1 0 15546 0 1 4
box 0 0 1 1
use contact_17  contact_17_49
timestamp 1643671299
transform 1 0 15561 0 1 19
box 0 0 1 1
use contact_18  contact_18_50
timestamp 1643671299
transform 1 0 13990 0 1 950
box 0 0 1 1
use contact_17  contact_17_50
timestamp 1643671299
transform 1 0 14005 0 1 965
box 0 0 1 1
use contact_18  contact_18_51
timestamp 1643671299
transform 1 0 13990 0 1 4
box 0 0 1 1
use contact_17  contact_17_51
timestamp 1643671299
transform 1 0 14005 0 1 19
box 0 0 1 1
use contact_18  contact_18_52
timestamp 1643671299
transform 1 0 12434 0 1 950
box 0 0 1 1
use contact_17  contact_17_52
timestamp 1643671299
transform 1 0 12449 0 1 965
box 0 0 1 1
use contact_18  contact_18_53
timestamp 1643671299
transform 1 0 12434 0 1 4
box 0 0 1 1
use contact_17  contact_17_53
timestamp 1643671299
transform 1 0 12449 0 1 19
box 0 0 1 1
use contact_18  contact_18_54
timestamp 1643671299
transform 1 0 10878 0 1 950
box 0 0 1 1
use contact_17  contact_17_54
timestamp 1643671299
transform 1 0 10893 0 1 965
box 0 0 1 1
use contact_18  contact_18_55
timestamp 1643671299
transform 1 0 10878 0 1 4
box 0 0 1 1
use contact_17  contact_17_55
timestamp 1643671299
transform 1 0 10893 0 1 19
box 0 0 1 1
use contact_18  contact_18_56
timestamp 1643671299
transform 1 0 9322 0 1 950
box 0 0 1 1
use contact_17  contact_17_56
timestamp 1643671299
transform 1 0 9337 0 1 965
box 0 0 1 1
use contact_18  contact_18_57
timestamp 1643671299
transform 1 0 9322 0 1 4
box 0 0 1 1
use contact_17  contact_17_57
timestamp 1643671299
transform 1 0 9337 0 1 19
box 0 0 1 1
use contact_18  contact_18_58
timestamp 1643671299
transform 1 0 7766 0 1 950
box 0 0 1 1
use contact_17  contact_17_58
timestamp 1643671299
transform 1 0 7781 0 1 965
box 0 0 1 1
use contact_18  contact_18_59
timestamp 1643671299
transform 1 0 7766 0 1 4
box 0 0 1 1
use contact_17  contact_17_59
timestamp 1643671299
transform 1 0 7781 0 1 19
box 0 0 1 1
use contact_18  contact_18_60
timestamp 1643671299
transform 1 0 6210 0 1 950
box 0 0 1 1
use contact_17  contact_17_60
timestamp 1643671299
transform 1 0 6225 0 1 965
box 0 0 1 1
use contact_18  contact_18_61
timestamp 1643671299
transform 1 0 6210 0 1 4
box 0 0 1 1
use contact_17  contact_17_61
timestamp 1643671299
transform 1 0 6225 0 1 19
box 0 0 1 1
use contact_18  contact_18_62
timestamp 1643671299
transform 1 0 4654 0 1 950
box 0 0 1 1
use contact_17  contact_17_62
timestamp 1643671299
transform 1 0 4669 0 1 965
box 0 0 1 1
use contact_18  contact_18_63
timestamp 1643671299
transform 1 0 4654 0 1 4
box 0 0 1 1
use contact_17  contact_17_63
timestamp 1643671299
transform 1 0 4669 0 1 19
box 0 0 1 1
use sense_amp_multiport  sense_amp_multiport_0
timestamp 1643671299
transform 1 0 52784 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_1
timestamp 1643671299
transform 1 0 51228 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_2
timestamp 1643671299
transform 1 0 49672 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_3
timestamp 1643671299
transform 1 0 48116 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_4
timestamp 1643671299
transform 1 0 46560 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_5
timestamp 1643671299
transform 1 0 45004 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_6
timestamp 1643671299
transform 1 0 43448 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_7
timestamp 1643671299
transform 1 0 41892 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_8
timestamp 1643671299
transform 1 0 40336 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_9
timestamp 1643671299
transform 1 0 38780 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_10
timestamp 1643671299
transform 1 0 37224 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_11
timestamp 1643671299
transform 1 0 35668 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_12
timestamp 1643671299
transform 1 0 34112 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_13
timestamp 1643671299
transform 1 0 32556 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_14
timestamp 1643671299
transform 1 0 31000 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_15
timestamp 1643671299
transform 1 0 29444 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_16
timestamp 1643671299
transform 1 0 27888 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_17
timestamp 1643671299
transform 1 0 26332 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_18
timestamp 1643671299
transform 1 0 24776 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_19
timestamp 1643671299
transform 1 0 23220 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_20
timestamp 1643671299
transform 1 0 21664 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_21
timestamp 1643671299
transform 1 0 20108 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_22
timestamp 1643671299
transform 1 0 18552 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_23
timestamp 1643671299
transform 1 0 16996 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_24
timestamp 1643671299
transform 1 0 15440 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_25
timestamp 1643671299
transform 1 0 13884 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_26
timestamp 1643671299
transform 1 0 12328 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_27
timestamp 1643671299
transform 1 0 10772 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_28
timestamp 1643671299
transform 1 0 9216 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_29
timestamp 1643671299
transform 1 0 7660 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_30
timestamp 1643671299
transform 1 0 6104 0 1 0
box 0 0 272 1050
use sense_amp_multiport  sense_amp_multiport_31
timestamp 1643671299
transform 1 0 4548 0 1 0
box 0 0 272 1050
<< labels >>
rlabel metal3 s 43554 4 43614 64 4 gnd
rlabel metal3 s 21770 4 21830 64 4 gnd
rlabel metal3 s 20214 4 20274 64 4 gnd
rlabel metal3 s 45110 4 45170 64 4 gnd
rlabel metal3 s 49778 4 49838 64 4 gnd
rlabel metal3 s 48222 4 48282 64 4 gnd
rlabel metal3 s 41998 4 42058 64 4 gnd
rlabel metal3 s 18658 4 18718 64 4 gnd
rlabel metal3 s 34218 4 34278 64 4 gnd
rlabel metal3 s 15546 4 15606 64 4 gnd
rlabel metal3 s 40442 4 40502 64 4 gnd
rlabel metal3 s 32662 4 32722 64 4 gnd
rlabel metal3 s 27994 4 28054 64 4 gnd
rlabel metal3 s 9322 4 9382 64 4 gnd
rlabel metal3 s 7766 4 7826 64 4 gnd
rlabel metal3 s 10878 4 10938 64 4 gnd
rlabel metal3 s 37330 4 37390 64 4 gnd
rlabel metal3 s 12434 4 12494 64 4 gnd
rlabel metal3 s 38886 4 38946 64 4 gnd
rlabel metal3 s 4654 4 4714 64 4 gnd
rlabel metal3 s 29550 4 29610 64 4 gnd
rlabel metal3 s 52890 4 52950 64 4 gnd
rlabel metal3 s 23326 4 23386 64 4 gnd
rlabel metal3 s 6210 4 6270 64 4 gnd
rlabel metal3 s 24882 4 24942 64 4 gnd
rlabel metal3 s 26438 4 26498 64 4 gnd
rlabel metal3 s 35774 4 35834 64 4 gnd
rlabel metal3 s 31106 4 31166 64 4 gnd
rlabel metal3 s 13990 4 14050 64 4 gnd
rlabel metal3 s 46666 4 46726 64 4 gnd
rlabel metal3 s 51334 4 51394 64 4 gnd
rlabel metal3 s 17102 4 17162 64 4 gnd
rlabel metal3 s 4654 950 4714 1010 4 vdd
rlabel metal3 s 40442 950 40502 1010 4 vdd
rlabel metal3 s 52890 950 52950 1010 4 vdd
rlabel metal3 s 21770 950 21830 1010 4 vdd
rlabel metal3 s 29550 950 29610 1010 4 vdd
rlabel metal3 s 37330 950 37390 1010 4 vdd
rlabel metal3 s 13990 950 14050 1010 4 vdd
rlabel metal3 s 20214 950 20274 1010 4 vdd
rlabel metal3 s 35774 950 35834 1010 4 vdd
rlabel metal3 s 9322 950 9382 1010 4 vdd
rlabel metal3 s 18658 950 18718 1010 4 vdd
rlabel metal3 s 51334 950 51394 1010 4 vdd
rlabel metal3 s 43554 950 43614 1010 4 vdd
rlabel metal3 s 41998 950 42058 1010 4 vdd
rlabel metal3 s 17102 950 17162 1010 4 vdd
rlabel metal3 s 38886 950 38946 1010 4 vdd
rlabel metal3 s 48222 950 48282 1010 4 vdd
rlabel metal3 s 32662 950 32722 1010 4 vdd
rlabel metal3 s 46666 950 46726 1010 4 vdd
rlabel metal3 s 12434 950 12494 1010 4 vdd
rlabel metal3 s 15546 950 15606 1010 4 vdd
rlabel metal3 s 23326 950 23386 1010 4 vdd
rlabel metal3 s 34218 950 34278 1010 4 vdd
rlabel metal3 s 24882 950 24942 1010 4 vdd
rlabel metal3 s 45110 950 45170 1010 4 vdd
rlabel metal3 s 10878 950 10938 1010 4 vdd
rlabel metal3 s 27994 950 28054 1010 4 vdd
rlabel metal3 s 31106 950 31166 1010 4 vdd
rlabel metal3 s 7766 950 7826 1010 4 vdd
rlabel metal3 s 26438 950 26498 1010 4 vdd
rlabel metal3 s 49778 950 49838 1010 4 vdd
rlabel metal3 s 6210 950 6270 1010 4 vdd
rlabel metal2 s 4562 0 4590 240 4 rbl_0
rlabel metal2 s 4750 0 4778 240 4 data_0
rlabel metal2 s 6118 0 6146 240 4 rbl_1
rlabel metal2 s 6306 0 6334 240 4 data_1
rlabel metal2 s 7674 0 7702 240 4 rbl_2
rlabel metal2 s 7862 0 7890 240 4 data_2
rlabel metal2 s 9230 0 9258 240 4 rbl_3
rlabel metal2 s 9418 0 9446 240 4 data_3
rlabel metal2 s 10786 0 10814 240 4 rbl_4
rlabel metal2 s 10974 0 11002 240 4 data_4
rlabel metal2 s 12342 0 12370 240 4 rbl_5
rlabel metal2 s 12530 0 12558 240 4 data_5
rlabel metal2 s 13898 0 13926 240 4 rbl_6
rlabel metal2 s 14086 0 14114 240 4 data_6
rlabel metal2 s 15454 0 15482 240 4 rbl_7
rlabel metal2 s 15642 0 15670 240 4 data_7
rlabel metal2 s 17010 0 17038 240 4 rbl_8
rlabel metal2 s 17198 0 17226 240 4 data_8
rlabel metal2 s 18566 0 18594 240 4 rbl_9
rlabel metal2 s 18754 0 18782 240 4 data_9
rlabel metal2 s 20122 0 20150 240 4 rbl_10
rlabel metal2 s 20310 0 20338 240 4 data_10
rlabel metal2 s 21678 0 21706 240 4 rbl_11
rlabel metal2 s 21866 0 21894 240 4 data_11
rlabel metal2 s 23234 0 23262 240 4 rbl_12
rlabel metal2 s 23422 0 23450 240 4 data_12
rlabel metal2 s 24790 0 24818 240 4 rbl_13
rlabel metal2 s 24978 0 25006 240 4 data_13
rlabel metal2 s 26346 0 26374 240 4 rbl_14
rlabel metal2 s 26534 0 26562 240 4 data_14
rlabel metal2 s 27902 0 27930 240 4 rbl_15
rlabel metal2 s 28090 0 28118 240 4 data_15
rlabel metal2 s 29458 0 29486 240 4 rbl_16
rlabel metal2 s 29646 0 29674 240 4 data_16
rlabel metal2 s 31014 0 31042 240 4 rbl_17
rlabel metal2 s 31202 0 31230 240 4 data_17
rlabel metal2 s 32570 0 32598 240 4 rbl_18
rlabel metal2 s 32758 0 32786 240 4 data_18
rlabel metal2 s 34126 0 34154 240 4 rbl_19
rlabel metal2 s 34314 0 34342 240 4 data_19
rlabel metal2 s 35682 0 35710 240 4 rbl_20
rlabel metal2 s 35870 0 35898 240 4 data_20
rlabel metal2 s 37238 0 37266 240 4 rbl_21
rlabel metal2 s 37426 0 37454 240 4 data_21
rlabel metal2 s 38794 0 38822 240 4 rbl_22
rlabel metal2 s 38982 0 39010 240 4 data_22
rlabel metal2 s 40350 0 40378 240 4 rbl_23
rlabel metal2 s 40538 0 40566 240 4 data_23
rlabel metal2 s 41906 0 41934 240 4 rbl_24
rlabel metal2 s 42094 0 42122 240 4 data_24
rlabel metal2 s 43462 0 43490 240 4 rbl_25
rlabel metal2 s 43650 0 43678 240 4 data_25
rlabel metal2 s 45018 0 45046 240 4 rbl_26
rlabel metal2 s 45206 0 45234 240 4 data_26
rlabel metal2 s 46574 0 46602 240 4 rbl_27
rlabel metal2 s 46762 0 46790 240 4 data_27
rlabel metal2 s 48130 0 48158 240 4 rbl_28
rlabel metal2 s 48318 0 48346 240 4 data_28
rlabel metal2 s 49686 0 49714 240 4 rbl_29
rlabel metal2 s 49874 0 49902 240 4 data_29
rlabel metal2 s 51242 0 51270 240 4 rbl_30
rlabel metal2 s 51430 0 51458 240 4 data_30
rlabel metal2 s 52798 0 52826 240 4 rbl_31
rlabel metal2 s 52986 0 53014 240 4 data_31
<< properties >>
string FIXED_BBOX 0 0 53056 1050
string GDS_FILE sram_0rw2r1w_16_32_sky130A.gds
string GDS_END 814912
string GDS_START 779984
<< end >>
