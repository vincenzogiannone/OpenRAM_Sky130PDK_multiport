magic
tech sky130A
magscale 1 2
timestamp 1643671299
<< checkpaint >>
rect -1319 -1316 2657 1608
<< nwell >>
rect -54 231 1392 348
rect -59 63 1397 231
rect -54 -54 1392 63
<< scpmos >>
rect 60 0 90 294
rect 168 0 198 294
rect 276 0 306 294
rect 384 0 414 294
rect 492 0 522 294
rect 600 0 630 294
rect 708 0 738 294
rect 816 0 846 294
rect 924 0 954 294
rect 1032 0 1062 294
rect 1140 0 1170 294
rect 1248 0 1278 294
<< pdiff >>
rect 0 164 60 294
rect 0 130 8 164
rect 42 130 60 164
rect 0 0 60 130
rect 90 164 168 294
rect 90 130 112 164
rect 146 130 168 164
rect 90 0 168 130
rect 198 164 276 294
rect 198 130 220 164
rect 254 130 276 164
rect 198 0 276 130
rect 306 164 384 294
rect 306 130 328 164
rect 362 130 384 164
rect 306 0 384 130
rect 414 164 492 294
rect 414 130 436 164
rect 470 130 492 164
rect 414 0 492 130
rect 522 164 600 294
rect 522 130 544 164
rect 578 130 600 164
rect 522 0 600 130
rect 630 164 708 294
rect 630 130 652 164
rect 686 130 708 164
rect 630 0 708 130
rect 738 164 816 294
rect 738 130 760 164
rect 794 130 816 164
rect 738 0 816 130
rect 846 164 924 294
rect 846 130 868 164
rect 902 130 924 164
rect 846 0 924 130
rect 954 164 1032 294
rect 954 130 976 164
rect 1010 130 1032 164
rect 954 0 1032 130
rect 1062 164 1140 294
rect 1062 130 1084 164
rect 1118 130 1140 164
rect 1062 0 1140 130
rect 1170 164 1248 294
rect 1170 130 1192 164
rect 1226 130 1248 164
rect 1170 0 1248 130
rect 1278 164 1338 294
rect 1278 130 1296 164
rect 1330 130 1338 164
rect 1278 0 1338 130
<< pdiffc >>
rect 8 130 42 164
rect 112 130 146 164
rect 220 130 254 164
rect 328 130 362 164
rect 436 130 470 164
rect 544 130 578 164
rect 652 130 686 164
rect 760 130 794 164
rect 868 130 902 164
rect 976 130 1010 164
rect 1084 130 1118 164
rect 1192 130 1226 164
rect 1296 130 1330 164
<< poly >>
rect 60 294 90 320
rect 168 294 198 320
rect 276 294 306 320
rect 384 294 414 320
rect 492 294 522 320
rect 600 294 630 320
rect 708 294 738 320
rect 816 294 846 320
rect 924 294 954 320
rect 1032 294 1062 320
rect 1140 294 1170 320
rect 1248 294 1278 320
rect 60 -26 90 0
rect 168 -26 198 0
rect 276 -26 306 0
rect 384 -26 414 0
rect 492 -26 522 0
rect 600 -26 630 0
rect 708 -26 738 0
rect 816 -26 846 0
rect 924 -26 954 0
rect 1032 -26 1062 0
rect 1140 -26 1170 0
rect 1248 -26 1278 0
rect 60 -56 1278 -26
<< locali >>
rect 8 164 42 180
rect 8 114 42 130
rect 112 164 146 180
rect 112 80 146 130
rect 220 164 254 180
rect 220 114 254 130
rect 328 164 362 180
rect 328 80 362 130
rect 436 164 470 180
rect 436 114 470 130
rect 544 164 578 180
rect 544 80 578 130
rect 652 164 686 180
rect 652 114 686 130
rect 760 164 794 180
rect 760 80 794 130
rect 868 164 902 180
rect 868 114 902 130
rect 976 164 1010 180
rect 976 80 1010 130
rect 1084 164 1118 180
rect 1084 114 1118 130
rect 1192 164 1226 180
rect 1192 80 1226 130
rect 1296 164 1330 180
rect 1296 114 1330 130
rect 112 46 1226 80
use contact_9  contact_9_0
timestamp 1643671299
transform 1 0 1288 0 1 106
box 0 0 2 2
use contact_9  contact_9_1
timestamp 1643671299
transform 1 0 1184 0 1 106
box 0 0 2 2
use contact_9  contact_9_2
timestamp 1643671299
transform 1 0 1076 0 1 106
box 0 0 2 2
use contact_9  contact_9_3
timestamp 1643671299
transform 1 0 968 0 1 106
box 0 0 2 2
use contact_9  contact_9_4
timestamp 1643671299
transform 1 0 860 0 1 106
box 0 0 2 2
use contact_9  contact_9_5
timestamp 1643671299
transform 1 0 752 0 1 106
box 0 0 2 2
use contact_9  contact_9_6
timestamp 1643671299
transform 1 0 644 0 1 106
box 0 0 2 2
use contact_9  contact_9_7
timestamp 1643671299
transform 1 0 536 0 1 106
box 0 0 2 2
use contact_9  contact_9_8
timestamp 1643671299
transform 1 0 428 0 1 106
box 0 0 2 2
use contact_9  contact_9_9
timestamp 1643671299
transform 1 0 320 0 1 106
box 0 0 2 2
use contact_9  contact_9_10
timestamp 1643671299
transform 1 0 212 0 1 106
box 0 0 2 2
use contact_9  contact_9_11
timestamp 1643671299
transform 1 0 104 0 1 106
box 0 0 2 2
use contact_9  contact_9_12
timestamp 1643671299
transform 1 0 0 0 1 106
box 0 0 2 2
<< labels >>
rlabel mvvaractor s 669 -41 669 -41 4 G
rlabel locali s 669 147 669 147 4 S
rlabel locali s 885 147 885 147 4 S
rlabel locali s 1101 147 1101 147 4 S
rlabel locali s 1313 147 1313 147 4 S
rlabel locali s 453 147 453 147 4 S
rlabel locali s 237 147 237 147 4 S
rlabel locali s 25 147 25 147 4 S
rlabel locali s 669 63 669 63 4 D
<< properties >>
string FIXED_BBOX -54 -56 1392 63
string GDS_FILE sram_0rw2r1w_16_32_sky130A.gds
string GDS_END 1159782
string GDS_START 1156706
<< end >>
