magic
tech sky130A
magscale 1 2
timestamp 1644951705
<< checkpaint >>
rect -1260 -1302 2754 2876
<< nwell >>
rect 0 1118 1494 1616
<< pwell >>
rect 240 -42 312 42
rect 554 -42 626 42
rect 868 -42 940 42
rect 1182 -42 1254 42
<< nmos >>
rect 94 132 124 332
rect 190 132 220 332
rect 286 132 316 332
rect 382 132 412 332
rect 478 132 508 332
rect 574 132 604 332
rect 778 132 808 332
rect 874 132 904 332
rect 970 132 1000 332
rect 1074 132 1104 216
rect 1274 132 1304 216
rect 1370 132 1400 216
<< pmos >>
rect 94 1154 124 1238
rect 190 1154 220 1238
rect 286 1154 316 1238
rect 382 1154 412 1238
rect 478 1154 508 1238
rect 574 1154 604 1238
rect 778 1154 808 1238
rect 874 1154 904 1238
rect 970 1154 1000 1238
rect 1074 1154 1104 1424
rect 1274 1154 1304 1424
rect 1370 1154 1400 1424
<< ndiff >>
rect 36 298 94 332
rect 36 264 44 298
rect 78 264 94 298
rect 36 200 94 264
rect 36 166 44 200
rect 78 166 94 200
rect 36 132 94 166
rect 124 132 190 332
rect 220 132 286 332
rect 316 298 382 332
rect 316 264 332 298
rect 366 264 382 298
rect 316 200 382 264
rect 316 166 332 200
rect 366 166 382 200
rect 316 132 382 166
rect 412 132 478 332
rect 508 132 574 332
rect 604 298 662 332
rect 604 264 620 298
rect 654 264 662 298
rect 604 200 662 264
rect 604 166 620 200
rect 654 166 662 200
rect 604 132 662 166
rect 720 298 778 332
rect 720 264 728 298
rect 762 264 778 298
rect 720 200 778 264
rect 720 166 728 200
rect 762 166 778 200
rect 720 132 778 166
rect 808 132 874 332
rect 904 132 970 332
rect 1000 298 1058 332
rect 1000 264 1016 298
rect 1050 264 1058 298
rect 1000 216 1058 264
rect 1000 200 1074 216
rect 1000 166 1016 200
rect 1050 166 1074 200
rect 1000 132 1074 166
rect 1104 190 1162 216
rect 1104 156 1120 190
rect 1154 156 1162 190
rect 1104 132 1162 156
rect 1216 190 1274 216
rect 1216 156 1224 190
rect 1258 156 1274 190
rect 1216 132 1274 156
rect 1304 190 1370 216
rect 1304 156 1320 190
rect 1354 156 1370 190
rect 1304 132 1370 156
rect 1400 190 1458 216
rect 1400 156 1416 190
rect 1450 156 1458 190
rect 1400 132 1458 156
<< pdiff >>
rect 1016 1390 1074 1424
rect 1016 1356 1024 1390
rect 1058 1356 1074 1390
rect 1016 1306 1074 1356
rect 1016 1272 1024 1306
rect 1058 1272 1074 1306
rect 1016 1238 1074 1272
rect 36 1212 94 1238
rect 36 1178 44 1212
rect 78 1178 94 1212
rect 36 1154 94 1178
rect 124 1212 190 1238
rect 124 1178 140 1212
rect 174 1178 190 1212
rect 124 1154 190 1178
rect 220 1212 286 1238
rect 220 1178 236 1212
rect 270 1178 286 1212
rect 220 1154 286 1178
rect 316 1212 382 1238
rect 316 1178 332 1212
rect 366 1178 382 1212
rect 316 1154 382 1178
rect 412 1212 478 1238
rect 412 1178 428 1212
rect 462 1178 478 1212
rect 412 1154 478 1178
rect 508 1212 574 1238
rect 508 1178 524 1212
rect 558 1178 574 1212
rect 508 1154 574 1178
rect 604 1212 662 1238
rect 604 1178 620 1212
rect 654 1178 662 1212
rect 604 1154 662 1178
rect 720 1212 778 1238
rect 720 1178 728 1212
rect 762 1178 778 1212
rect 720 1154 778 1178
rect 808 1212 874 1238
rect 808 1178 824 1212
rect 858 1178 874 1212
rect 808 1154 874 1178
rect 904 1212 970 1238
rect 904 1178 920 1212
rect 954 1178 970 1212
rect 904 1154 970 1178
rect 1000 1222 1074 1238
rect 1000 1188 1024 1222
rect 1058 1188 1074 1222
rect 1000 1154 1074 1188
rect 1104 1390 1162 1424
rect 1104 1356 1120 1390
rect 1154 1356 1162 1390
rect 1104 1306 1162 1356
rect 1104 1272 1120 1306
rect 1154 1272 1162 1306
rect 1104 1222 1162 1272
rect 1104 1188 1120 1222
rect 1154 1188 1162 1222
rect 1104 1154 1162 1188
rect 1216 1390 1274 1424
rect 1216 1356 1224 1390
rect 1258 1356 1274 1390
rect 1216 1306 1274 1356
rect 1216 1272 1224 1306
rect 1258 1272 1274 1306
rect 1216 1222 1274 1272
rect 1216 1188 1224 1222
rect 1258 1188 1274 1222
rect 1216 1154 1274 1188
rect 1304 1390 1370 1424
rect 1304 1356 1320 1390
rect 1354 1356 1370 1390
rect 1304 1306 1370 1356
rect 1304 1272 1320 1306
rect 1354 1272 1370 1306
rect 1304 1222 1370 1272
rect 1304 1188 1320 1222
rect 1354 1188 1370 1222
rect 1304 1154 1370 1188
rect 1400 1390 1458 1424
rect 1400 1356 1416 1390
rect 1450 1356 1458 1390
rect 1400 1306 1458 1356
rect 1400 1272 1416 1306
rect 1450 1272 1458 1306
rect 1400 1222 1458 1272
rect 1400 1188 1416 1222
rect 1450 1188 1458 1222
rect 1400 1154 1458 1188
<< ndiffc >>
rect 44 264 78 298
rect 44 166 78 200
rect 332 264 366 298
rect 332 166 366 200
rect 620 264 654 298
rect 620 166 654 200
rect 728 264 762 298
rect 728 166 762 200
rect 1016 264 1050 298
rect 1016 166 1050 200
rect 1120 156 1154 190
rect 1224 156 1258 190
rect 1320 156 1354 190
rect 1416 156 1450 190
<< pdiffc >>
rect 1024 1356 1058 1390
rect 1024 1272 1058 1306
rect 44 1178 78 1212
rect 140 1178 174 1212
rect 236 1178 270 1212
rect 332 1178 366 1212
rect 428 1178 462 1212
rect 524 1178 558 1212
rect 620 1178 654 1212
rect 728 1178 762 1212
rect 824 1178 858 1212
rect 920 1178 954 1212
rect 1024 1188 1058 1222
rect 1120 1356 1154 1390
rect 1120 1272 1154 1306
rect 1120 1188 1154 1222
rect 1224 1356 1258 1390
rect 1224 1272 1258 1306
rect 1224 1188 1258 1222
rect 1320 1356 1354 1390
rect 1320 1272 1354 1306
rect 1320 1188 1354 1222
rect 1416 1356 1450 1390
rect 1416 1272 1450 1306
rect 1416 1188 1450 1222
<< psubdiff >>
rect 240 17 312 42
rect 240 -17 259 17
rect 293 -17 312 17
rect 240 -42 312 -17
rect 554 17 626 42
rect 554 -17 573 17
rect 607 -17 626 17
rect 554 -42 626 -17
rect 868 17 940 42
rect 868 -17 887 17
rect 921 -17 940 17
rect 868 -42 940 -17
rect 1182 17 1254 42
rect 1182 -17 1201 17
rect 1235 -17 1254 17
rect 1182 -42 1254 -17
<< nsubdiff >>
rect 240 1555 312 1580
rect 240 1521 259 1555
rect 293 1521 312 1555
rect 240 1496 312 1521
rect 554 1555 626 1580
rect 554 1521 573 1555
rect 607 1521 626 1555
rect 554 1496 626 1521
rect 868 1555 940 1580
rect 868 1521 887 1555
rect 921 1521 940 1555
rect 868 1496 940 1521
rect 1182 1555 1254 1580
rect 1182 1521 1201 1555
rect 1235 1521 1254 1555
rect 1182 1496 1254 1521
<< psubdiffcont >>
rect 259 -17 293 17
rect 573 -17 607 17
rect 887 -17 921 17
rect 1201 -17 1235 17
<< nsubdiffcont >>
rect 259 1521 293 1555
rect 573 1521 607 1555
rect 887 1521 921 1555
rect 1201 1521 1235 1555
<< poly >>
rect 1074 1424 1104 1450
rect 1274 1424 1304 1450
rect 1370 1424 1400 1450
rect 94 1238 124 1264
rect 190 1238 220 1264
rect 286 1238 316 1264
rect 382 1238 412 1264
rect 478 1238 508 1264
rect 574 1238 604 1264
rect 778 1238 808 1264
rect 874 1238 904 1264
rect 970 1238 1000 1264
rect 94 1120 124 1154
rect 70 1104 124 1120
rect 70 1070 80 1104
rect 114 1070 124 1104
rect 70 1054 124 1070
rect 94 332 124 1054
rect 190 1034 220 1154
rect 166 1018 220 1034
rect 166 984 176 1018
rect 210 984 220 1018
rect 166 968 220 984
rect 190 332 220 968
rect 286 948 316 1154
rect 262 932 316 948
rect 262 898 272 932
rect 306 898 316 932
rect 262 882 316 898
rect 286 332 316 882
rect 382 862 412 1154
rect 358 846 412 862
rect 358 812 368 846
rect 402 812 412 846
rect 358 796 412 812
rect 382 332 412 796
rect 478 776 508 1154
rect 454 760 508 776
rect 454 726 464 760
rect 498 726 508 760
rect 454 710 508 726
rect 478 332 508 710
rect 574 690 604 1154
rect 550 674 604 690
rect 550 640 560 674
rect 594 640 604 674
rect 550 624 604 640
rect 574 332 604 624
rect 778 604 808 1154
rect 754 588 808 604
rect 754 554 764 588
rect 798 554 808 588
rect 754 538 808 554
rect 778 332 808 538
rect 874 518 904 1154
rect 850 502 904 518
rect 850 468 860 502
rect 894 468 904 502
rect 850 452 904 468
rect 874 332 904 452
rect 970 432 1000 1154
rect 1074 638 1104 1154
rect 1050 622 1104 638
rect 1050 588 1060 622
rect 1094 588 1104 622
rect 1050 572 1104 588
rect 946 416 1000 432
rect 946 382 956 416
rect 990 382 1000 416
rect 946 366 1000 382
rect 970 332 1000 366
rect 1074 216 1104 572
rect 1274 840 1304 1154
rect 1370 1120 1400 1154
rect 1346 1104 1400 1120
rect 1346 1070 1356 1104
rect 1390 1070 1400 1104
rect 1346 1054 1400 1070
rect 1274 824 1328 840
rect 1274 790 1284 824
rect 1318 790 1328 824
rect 1274 774 1328 790
rect 1274 216 1304 774
rect 1370 216 1400 1054
rect 94 106 124 132
rect 190 106 220 132
rect 286 106 316 132
rect 382 106 412 132
rect 478 106 508 132
rect 574 106 604 132
rect 778 106 808 132
rect 874 106 904 132
rect 970 106 1000 132
rect 1074 106 1104 132
rect 1274 106 1304 132
rect 1370 106 1400 132
<< polycont >>
rect 80 1070 114 1104
rect 176 984 210 1018
rect 272 898 306 932
rect 368 812 402 846
rect 464 726 498 760
rect 560 640 594 674
rect 764 554 798 588
rect 860 468 894 502
rect 1060 588 1094 622
rect 956 382 990 416
rect 1356 1070 1390 1104
rect 1284 790 1318 824
<< locali >>
rect 258 1556 294 1572
rect 572 1556 608 1572
rect 886 1556 922 1572
rect 1200 1556 1236 1572
rect 140 1555 1354 1556
rect 140 1521 259 1555
rect 293 1521 573 1555
rect 607 1521 887 1555
rect 921 1521 1201 1555
rect 1235 1521 1354 1555
rect 140 1520 1354 1521
rect 140 1238 174 1520
rect 258 1504 294 1520
rect 332 1238 366 1520
rect 524 1504 608 1520
rect 824 1504 922 1520
rect 524 1238 558 1504
rect 824 1238 858 1504
rect 1024 1424 1058 1520
rect 1200 1504 1236 1520
rect 1320 1424 1354 1520
rect 1016 1390 1064 1424
rect 1016 1356 1024 1390
rect 1058 1356 1064 1390
rect 1016 1306 1064 1356
rect 1016 1272 1024 1306
rect 1058 1272 1064 1306
rect 36 1212 84 1238
rect 36 1178 44 1212
rect 78 1178 84 1212
rect 36 1154 84 1178
rect 134 1212 180 1238
rect 134 1178 140 1212
rect 174 1178 180 1212
rect 134 1154 180 1178
rect 230 1212 276 1238
rect 230 1178 236 1212
rect 270 1178 276 1212
rect 230 1154 276 1178
rect 326 1212 372 1238
rect 326 1178 332 1212
rect 366 1178 372 1212
rect 326 1154 372 1178
rect 422 1212 468 1238
rect 422 1178 428 1212
rect 462 1178 468 1212
rect 422 1154 468 1178
rect 518 1212 564 1238
rect 518 1178 524 1212
rect 558 1178 564 1212
rect 518 1154 564 1178
rect 614 1212 662 1238
rect 614 1178 620 1212
rect 654 1178 662 1212
rect 614 1154 662 1178
rect 720 1212 768 1238
rect 720 1178 728 1212
rect 762 1178 768 1212
rect 720 1154 768 1178
rect 818 1212 864 1238
rect 818 1178 824 1212
rect 858 1178 864 1212
rect 818 1154 864 1178
rect 914 1212 960 1238
rect 914 1178 920 1212
rect 954 1178 960 1212
rect 914 1154 960 1178
rect 1016 1222 1064 1272
rect 1016 1188 1024 1222
rect 1058 1188 1064 1222
rect 1016 1154 1064 1188
rect 1114 1390 1162 1424
rect 1114 1356 1120 1390
rect 1154 1356 1162 1390
rect 1114 1306 1162 1356
rect 1114 1272 1120 1306
rect 1154 1272 1162 1306
rect 1114 1222 1162 1272
rect 1114 1188 1120 1222
rect 1154 1188 1162 1222
rect 1114 1154 1162 1188
rect 80 1104 114 1120
rect 80 1054 114 1070
rect 696 1076 728 1110
rect 176 1018 210 1034
rect 176 968 210 984
rect 272 932 306 948
rect 272 882 306 898
rect 368 846 402 862
rect 368 796 402 812
rect 464 760 498 776
rect 464 710 498 726
rect 560 674 594 690
rect 560 624 594 640
rect 628 590 662 796
rect 44 556 662 590
rect 44 332 78 556
rect 696 522 730 1076
rect 926 654 960 1154
rect 926 622 1094 654
rect 926 620 1060 622
rect 764 588 798 604
rect 1060 572 1094 588
rect 1128 608 1162 1154
rect 1216 1390 1264 1424
rect 1216 1356 1224 1390
rect 1258 1356 1264 1390
rect 1216 1306 1264 1356
rect 1216 1272 1224 1306
rect 1258 1272 1264 1306
rect 1216 1222 1264 1272
rect 1216 1188 1224 1222
rect 1258 1188 1264 1222
rect 1216 1154 1264 1188
rect 1314 1390 1360 1424
rect 1314 1356 1320 1390
rect 1354 1356 1360 1390
rect 1314 1306 1360 1356
rect 1314 1272 1320 1306
rect 1354 1272 1360 1306
rect 1314 1222 1360 1272
rect 1314 1188 1320 1222
rect 1354 1188 1360 1222
rect 1314 1154 1360 1188
rect 1410 1390 1458 1424
rect 1410 1356 1416 1390
rect 1450 1356 1458 1390
rect 1410 1306 1458 1356
rect 1410 1272 1416 1306
rect 1450 1272 1458 1306
rect 1410 1222 1458 1272
rect 1410 1188 1416 1222
rect 1450 1188 1458 1222
rect 1410 1154 1458 1188
rect 1216 730 1250 1154
rect 1356 1104 1390 1120
rect 1356 1054 1390 1070
rect 1424 876 1458 1154
rect 1284 824 1318 840
rect 1284 774 1318 790
rect 1128 574 1134 608
rect 764 538 798 554
rect 620 488 730 522
rect 860 502 894 518
rect 620 332 654 488
rect 860 452 894 468
rect 956 416 990 432
rect 956 366 990 382
rect 36 298 84 332
rect 36 264 44 298
rect 78 264 84 298
rect 36 200 84 264
rect 36 166 44 200
rect 78 166 84 200
rect 36 132 84 166
rect 326 298 372 332
rect 326 264 332 298
rect 366 264 372 298
rect 326 200 372 264
rect 326 166 332 200
rect 366 166 372 200
rect 326 132 372 166
rect 614 298 662 332
rect 614 264 620 298
rect 654 264 662 298
rect 614 200 662 264
rect 614 166 620 200
rect 654 166 662 200
rect 614 132 662 166
rect 720 298 768 332
rect 720 264 728 298
rect 762 264 768 298
rect 720 200 768 264
rect 720 166 728 200
rect 762 166 768 200
rect 720 132 768 166
rect 1010 298 1058 332
rect 1010 264 1016 298
rect 1050 264 1058 298
rect 1010 200 1058 264
rect 1128 216 1162 574
rect 1010 166 1016 200
rect 1050 166 1058 200
rect 1010 132 1058 166
rect 1114 190 1162 216
rect 1114 156 1120 190
rect 1154 156 1162 190
rect 1114 132 1162 156
rect 1216 216 1250 696
rect 1424 216 1458 842
rect 1216 190 1264 216
rect 1216 156 1224 190
rect 1258 156 1264 190
rect 1216 132 1264 156
rect 1314 190 1360 216
rect 1314 156 1320 190
rect 1354 156 1360 190
rect 1314 132 1360 156
rect 1410 190 1458 216
rect 1410 156 1416 190
rect 1450 156 1458 190
rect 1410 132 1458 156
rect 258 18 294 42
rect 332 18 366 132
rect 572 18 608 42
rect 886 18 922 42
rect 1016 18 1050 132
rect 1200 18 1236 42
rect 1320 18 1354 132
rect 140 17 1354 18
rect 140 -17 259 17
rect 293 -17 573 17
rect 607 -17 887 17
rect 921 -17 1201 17
rect 1235 -17 1354 17
rect 140 -18 1354 -17
rect 258 -42 294 -18
rect 572 -42 608 -18
rect 886 -42 922 -18
rect 1200 -42 1236 -18
<< viali >>
rect 259 1521 293 1555
rect 573 1521 607 1555
rect 887 1521 921 1555
rect 1201 1521 1235 1555
rect 44 1178 78 1212
rect 236 1178 270 1212
rect 428 1178 462 1212
rect 620 1178 654 1212
rect 728 1178 762 1212
rect 920 1178 954 1212
rect 80 1070 114 1104
rect 728 1076 762 1110
rect 176 984 210 1018
rect 272 898 306 932
rect 368 812 402 846
rect 628 796 662 830
rect 464 726 498 760
rect 560 640 594 674
rect 764 554 798 588
rect 1060 588 1094 622
rect 1356 1070 1390 1104
rect 1424 842 1458 876
rect 1284 790 1318 824
rect 1216 696 1250 730
rect 1134 574 1168 608
rect 860 468 894 502
rect 956 382 990 416
rect 728 166 762 200
rect 259 -17 293 17
rect 573 -17 607 17
rect 887 -17 921 17
rect 1201 -17 1235 17
<< metal1 >>
rect 0 1555 1494 1568
rect 0 1521 259 1555
rect 293 1521 573 1555
rect 607 1521 887 1555
rect 921 1521 1201 1555
rect 1235 1521 1494 1555
rect 0 1508 1494 1521
rect 38 1212 276 1224
rect 38 1178 44 1212
rect 78 1196 236 1212
rect 78 1178 84 1196
rect 38 1166 84 1178
rect 230 1178 236 1196
rect 270 1178 276 1212
rect 230 1166 276 1178
rect 422 1212 660 1224
rect 422 1178 428 1212
rect 462 1196 620 1212
rect 462 1178 468 1196
rect 422 1166 468 1178
rect 614 1178 620 1196
rect 654 1178 660 1212
rect 614 1166 660 1178
rect 722 1212 960 1224
rect 722 1178 728 1212
rect 762 1196 920 1212
rect 762 1178 768 1196
rect 722 1166 768 1178
rect 914 1178 920 1196
rect 954 1178 960 1212
rect 914 1166 960 1178
rect 248 1130 276 1166
rect 72 1104 126 1118
rect 72 1084 80 1104
rect 70 1070 80 1084
rect 114 1070 126 1104
rect 248 1102 506 1130
rect 70 1056 126 1070
rect 168 1018 222 1032
rect 168 998 176 1018
rect 166 984 176 998
rect 210 984 222 1018
rect 166 970 222 984
rect 264 932 318 946
rect 264 912 272 932
rect 262 898 272 912
rect 306 898 318 932
rect 478 930 506 1102
rect 632 1122 660 1166
rect 632 1116 768 1122
rect 632 1110 1396 1116
rect 632 1094 728 1110
rect 722 1076 728 1094
rect 762 1104 1396 1110
rect 762 1088 1356 1104
rect 762 1076 768 1088
rect 722 1064 768 1076
rect 1350 1070 1356 1088
rect 1390 1070 1396 1104
rect 1350 1058 1396 1070
rect 478 902 642 930
rect 262 884 318 898
rect 360 846 414 860
rect 360 826 368 846
rect 358 812 368 826
rect 402 812 414 846
rect 358 798 414 812
rect 614 836 642 902
rect 1418 876 1464 888
rect 1418 842 1424 876
rect 1458 848 1494 876
rect 1458 842 1464 848
rect 614 830 1324 836
rect 1418 830 1464 842
rect 614 796 628 830
rect 662 824 1324 830
rect 662 808 1284 824
rect 662 796 674 808
rect 614 786 674 796
rect 1278 790 1284 808
rect 1318 790 1324 824
rect 1278 778 1324 790
rect 456 760 510 774
rect 456 740 464 760
rect 454 726 464 740
rect 498 726 510 760
rect 454 712 510 726
rect 1210 730 1256 742
rect 1210 696 1216 730
rect 1250 702 1494 730
rect 1250 696 1256 702
rect 552 674 606 688
rect 1210 684 1256 696
rect 552 654 560 674
rect 550 640 560 654
rect 594 640 606 674
rect 550 626 606 640
rect 1054 622 1100 634
rect 756 588 810 602
rect 756 568 764 588
rect 754 554 764 568
rect 798 554 810 588
rect 1054 588 1060 622
rect 1094 588 1100 622
rect 1054 576 1100 588
rect 754 540 810 554
rect 852 502 906 516
rect 852 482 860 502
rect 850 468 860 482
rect 894 468 906 502
rect 850 454 906 468
rect 948 416 1002 430
rect 948 396 956 416
rect 946 382 956 396
rect 990 382 1002 416
rect 946 368 1002 382
rect 1072 212 1100 576
rect 1128 608 1174 620
rect 1128 574 1134 608
rect 1168 580 1494 608
rect 1168 574 1174 580
rect 1128 562 1174 574
rect 722 200 1100 212
rect 722 166 728 200
rect 762 184 1100 200
rect 762 166 768 184
rect 722 154 768 166
rect 0 17 1494 30
rect 0 -17 259 17
rect 293 -17 573 17
rect 607 -17 887 17
rect 921 -17 1201 17
rect 1235 -17 1494 17
rect 0 -30 1494 -17
<< labels >>
rlabel locali s 950 750 950 750 4 net9
rlabel metal1 s 652 1102 652 1102 4 net6
rlabel metal1 s 358 1106 358 1106 4 net3
rlabel mvpsubdiff s 434 218 434 218 4 net4
rlabel mvpsubdiff s 532 216 532 216 4 net5
rlabel mvpsubdiff s 252 216 252 216 4 net1
rlabel mvpsubdiff s 158 208 158 208 4 net2
rlabel mvpsubdiff s 932 242 932 242 4 net7
rlabel mvpsubdiff s 840 238 840 238 4 net8
rlabel metal1 s 70 1056 126 1084 4 A0
port 1 nsew
rlabel metal1 s 166 970 222 998 4 B0
port 2 nsew
rlabel metal1 s 262 884 318 912 4 C0
port 3 nsew
rlabel metal1 s 358 798 414 826 4 A1
port 4 nsew
rlabel metal1 s 454 712 510 740 4 B1
port 5 nsew
rlabel metal1 s 550 626 606 654 4 C1
port 6 nsew
rlabel metal1 s 754 540 810 568 4 A2
port 7 nsew
rlabel metal1 s 850 454 906 482 4 B2
port 8 nsew
rlabel metal1 s 946 368 1002 396 4 C2
port 9 nsew
rlabel metal1 s 1128 580 1494 608 4 OUT2
port 10 nsew
rlabel metal1 s 0 1508 1494 1568 4 vdd
port 11 nsew
rlabel metal1 s 0 -30 1494 30 4 gnd
port 12 nsew
rlabel metal1 s 1418 848 1494 876 4 OUT0
port 13 nsew
rlabel metal1 s 1210 702 1494 730 4 OUT1
port 14 nsew
rlabel metal1 s 98 1070 98 1070 4 A0
rlabel metal1 s 194 984 194 984 4 B0
rlabel metal1 s 290 898 290 898 4 C0
rlabel metal1 s 386 812 386 812 4 A1
rlabel metal1 s 482 726 482 726 4 B1
rlabel metal1 s 578 640 578 640 4 C1
rlabel metal1 s 782 554 782 554 4 A2
rlabel metal1 s 878 468 878 468 4 B2
rlabel metal1 s 974 382 974 382 4 C2
rlabel metal1 s 1456 862 1456 862 4 OUT0
rlabel metal1 s 1352 716 1352 716 4 OUT1
rlabel metal1 s 1311 594 1311 594 4 OUT2
rlabel metal1 s 747 1538 747 1538 4 vdd
rlabel metal1 s 747 0 747 0 4 gnd
<< properties >>
string FIXED_BBOX 0 0 1494 1538
string GDS_FILE sram_0rw2r1w_16_128_sky130A.gds
string GDS_END 1842472
string GDS_START 1817894
<< end >>
