magic
tech sky130A
magscale 1 2
timestamp 1643671299
<< checkpaint >>
rect -1260 -1302 2494 25910
<< metal1 >>
rect 536 23998 618 24026
rect 1176 23928 1204 23956
rect 234 23878 318 23906
rect 1176 23802 1204 23830
rect 56 23732 126 23760
rect 1176 23576 1204 23604
rect 1176 22536 1204 22564
rect 56 22380 126 22408
rect 1176 22310 1204 22338
rect 234 22234 318 22262
rect 1176 22184 1204 22212
rect 536 22114 618 22142
rect 536 20922 618 20950
rect 1176 20852 1204 20880
rect 234 20802 318 20830
rect 1176 20726 1204 20754
rect 56 20656 126 20684
rect 1176 20500 1204 20528
rect 1176 19460 1204 19488
rect 56 19304 126 19332
rect 1176 19234 1204 19262
rect 234 19158 318 19186
rect 1176 19108 1204 19136
rect 536 19038 618 19066
rect 536 17846 618 17874
rect 1176 17776 1204 17804
rect 234 17726 318 17754
rect 1176 17650 1204 17678
rect 56 17580 126 17608
rect 1176 17424 1204 17452
rect 1176 16384 1204 16412
rect 56 16228 126 16256
rect 1176 16158 1204 16186
rect 234 16082 318 16110
rect 1176 16032 1204 16060
rect 536 15962 618 15990
rect 536 14770 618 14798
rect 1176 14700 1204 14728
rect 234 14650 318 14678
rect 1176 14574 1204 14602
rect 56 14504 126 14532
rect 1176 14348 1204 14376
rect 1176 13308 1204 13336
rect 56 13152 126 13180
rect 1176 13082 1204 13110
rect 234 13006 318 13034
rect 1176 12956 1204 12984
rect 536 12886 618 12914
rect 536 11694 618 11722
rect 1176 11624 1204 11652
rect 234 11574 318 11602
rect 1176 11498 1204 11526
rect 56 11428 126 11456
rect 1176 11272 1204 11300
rect 1176 10232 1204 10260
rect 56 10076 126 10104
rect 1176 10006 1204 10034
rect 234 9930 318 9958
rect 1176 9880 1204 9908
rect 536 9810 618 9838
rect 536 8618 618 8646
rect 1176 8548 1204 8576
rect 234 8498 318 8526
rect 1176 8422 1204 8450
rect 56 8352 126 8380
rect 1176 8196 1204 8224
rect 1176 7156 1204 7184
rect 56 7000 126 7028
rect 1176 6930 1204 6958
rect 234 6854 318 6882
rect 1176 6804 1204 6832
rect 536 6734 618 6762
rect 536 5542 618 5570
rect 1176 5472 1204 5500
rect 234 5422 318 5450
rect 1176 5346 1204 5374
rect 56 5276 126 5304
rect 1176 5120 1204 5148
rect 1176 4080 1204 4108
rect 56 3924 126 3952
rect 1176 3854 1204 3882
rect 234 3778 318 3806
rect 1176 3728 1204 3756
rect 536 3658 618 3686
rect 536 2466 618 2494
rect 1176 2396 1204 2424
rect 234 2346 318 2374
rect 1176 2270 1204 2298
rect 56 2200 126 2228
rect 1176 2044 1204 2072
rect 1176 1004 1204 1032
rect 56 848 126 876
rect 1176 778 1204 806
rect 234 702 318 730
rect 1176 652 1204 680
rect 536 582 618 610
<< via1 >>
rect 1178 24582 1230 24634
rect 1178 23044 1230 23096
rect 1178 21506 1230 21558
rect 1178 19968 1230 20020
rect 1178 18430 1230 18482
rect 1178 16892 1230 16944
rect 1178 15354 1230 15406
rect 1178 13816 1230 13868
rect 1178 12278 1230 12330
rect 1178 10740 1230 10792
rect 1178 9202 1230 9254
rect 1178 7664 1230 7716
rect 1178 6126 1230 6178
rect 1178 4588 1230 4640
rect 1178 3050 1230 3102
rect 1178 1512 1230 1564
rect 1178 -26 1230 26
<< metal2 >>
rect 1184 24636 1224 24642
rect 0 0 28 24608
rect 1184 24574 1224 24580
rect 192 23900 220 23928
rect 1184 23098 1224 23104
rect 1184 23036 1224 23042
rect 192 22212 220 22240
rect 1184 21560 1224 21566
rect 1184 21498 1224 21504
rect 192 20824 220 20852
rect 1184 20022 1224 20028
rect 1184 19960 1224 19966
rect 192 19136 220 19164
rect 1184 18484 1224 18490
rect 1184 18422 1224 18428
rect 192 17748 220 17776
rect 1184 16946 1224 16952
rect 1184 16884 1224 16890
rect 192 16060 220 16088
rect 1184 15408 1224 15414
rect 1184 15346 1224 15352
rect 192 14672 220 14700
rect 1184 13870 1224 13876
rect 1184 13808 1224 13814
rect 192 12984 220 13012
rect 1184 12332 1224 12338
rect 1184 12270 1224 12276
rect 192 11596 220 11624
rect 1184 10794 1224 10800
rect 1184 10732 1224 10738
rect 192 9908 220 9936
rect 1184 9256 1224 9262
rect 1184 9194 1224 9200
rect 192 8520 220 8548
rect 1184 7718 1224 7724
rect 1184 7656 1224 7662
rect 192 6832 220 6860
rect 1184 6180 1224 6186
rect 1184 6118 1224 6124
rect 192 5444 220 5472
rect 1184 4642 1224 4648
rect 1184 4580 1224 4586
rect 192 3756 220 3784
rect 1184 3104 1224 3110
rect 1184 3042 1224 3048
rect 192 2368 220 2396
rect 1184 1566 1224 1572
rect 1184 1504 1224 1510
rect 192 680 220 708
rect 1184 28 1224 34
rect 1184 -34 1224 -28
<< via2 >>
rect 1176 24634 1232 24636
rect 1176 24582 1178 24634
rect 1178 24582 1230 24634
rect 1230 24582 1232 24634
rect 1176 24580 1232 24582
rect 1176 23096 1232 23098
rect 1176 23044 1178 23096
rect 1178 23044 1230 23096
rect 1230 23044 1232 23096
rect 1176 23042 1232 23044
rect 1176 21558 1232 21560
rect 1176 21506 1178 21558
rect 1178 21506 1230 21558
rect 1230 21506 1232 21558
rect 1176 21504 1232 21506
rect 1176 20020 1232 20022
rect 1176 19968 1178 20020
rect 1178 19968 1230 20020
rect 1230 19968 1232 20020
rect 1176 19966 1232 19968
rect 1176 18482 1232 18484
rect 1176 18430 1178 18482
rect 1178 18430 1230 18482
rect 1230 18430 1232 18482
rect 1176 18428 1232 18430
rect 1176 16944 1232 16946
rect 1176 16892 1178 16944
rect 1178 16892 1230 16944
rect 1230 16892 1232 16944
rect 1176 16890 1232 16892
rect 1176 15406 1232 15408
rect 1176 15354 1178 15406
rect 1178 15354 1230 15406
rect 1230 15354 1232 15406
rect 1176 15352 1232 15354
rect 1176 13868 1232 13870
rect 1176 13816 1178 13868
rect 1178 13816 1230 13868
rect 1230 13816 1232 13868
rect 1176 13814 1232 13816
rect 1176 12330 1232 12332
rect 1176 12278 1178 12330
rect 1178 12278 1230 12330
rect 1230 12278 1232 12330
rect 1176 12276 1232 12278
rect 1176 10792 1232 10794
rect 1176 10740 1178 10792
rect 1178 10740 1230 10792
rect 1230 10740 1232 10792
rect 1176 10738 1232 10740
rect 1176 9254 1232 9256
rect 1176 9202 1178 9254
rect 1178 9202 1230 9254
rect 1230 9202 1232 9254
rect 1176 9200 1232 9202
rect 1176 7716 1232 7718
rect 1176 7664 1178 7716
rect 1178 7664 1230 7716
rect 1230 7664 1232 7716
rect 1176 7662 1232 7664
rect 1176 6178 1232 6180
rect 1176 6126 1178 6178
rect 1178 6126 1230 6178
rect 1230 6126 1232 6178
rect 1176 6124 1232 6126
rect 1176 4640 1232 4642
rect 1176 4588 1178 4640
rect 1178 4588 1230 4640
rect 1230 4588 1232 4640
rect 1176 4586 1232 4588
rect 1176 3102 1232 3104
rect 1176 3050 1178 3102
rect 1178 3050 1230 3102
rect 1230 3050 1232 3102
rect 1176 3048 1232 3050
rect 1176 1564 1232 1566
rect 1176 1512 1178 1564
rect 1178 1512 1230 1564
rect 1230 1512 1232 1564
rect 1176 1510 1232 1512
rect 1176 26 1232 28
rect 1176 -26 1178 26
rect 1178 -26 1230 26
rect 1230 -26 1232 26
rect 1176 -28 1232 -26
<< metal3 >>
rect 1174 24636 1234 24638
rect 1174 24580 1176 24636
rect 1232 24580 1234 24636
rect 1174 24578 1234 24580
rect 1174 23098 1234 23100
rect 1174 23042 1176 23098
rect 1232 23042 1234 23098
rect 1174 23040 1234 23042
rect 1174 21560 1234 21562
rect 1174 21504 1176 21560
rect 1232 21504 1234 21560
rect 1174 21502 1234 21504
rect 1174 20022 1234 20024
rect 1174 19966 1176 20022
rect 1232 19966 1234 20022
rect 1174 19964 1234 19966
rect 1174 18484 1234 18486
rect 1174 18428 1176 18484
rect 1232 18428 1234 18484
rect 1174 18426 1234 18428
rect 1174 16946 1234 16948
rect 1174 16890 1176 16946
rect 1232 16890 1234 16946
rect 1174 16888 1234 16890
rect 1174 15408 1234 15410
rect 1174 15352 1176 15408
rect 1232 15352 1234 15408
rect 1174 15350 1234 15352
rect 1174 13870 1234 13872
rect 1174 13814 1176 13870
rect 1232 13814 1234 13870
rect 1174 13812 1234 13814
rect 1174 12332 1234 12334
rect 1174 12276 1176 12332
rect 1232 12276 1234 12332
rect 1174 12274 1234 12276
rect 1174 10794 1234 10796
rect 1174 10738 1176 10794
rect 1232 10738 1234 10794
rect 1174 10736 1234 10738
rect 1174 9256 1234 9258
rect 1174 9200 1176 9256
rect 1232 9200 1234 9256
rect 1174 9198 1234 9200
rect 1174 7718 1234 7720
rect 1174 7662 1176 7718
rect 1232 7662 1234 7718
rect 1174 7660 1234 7662
rect 1174 6180 1234 6182
rect 1174 6124 1176 6180
rect 1232 6124 1234 6180
rect 1174 6122 1234 6124
rect 1174 4642 1234 4644
rect 1174 4586 1176 4642
rect 1232 4586 1234 4642
rect 1174 4584 1234 4586
rect 1174 3104 1234 3106
rect 1174 3048 1176 3104
rect 1232 3048 1234 3104
rect 1174 3046 1234 3048
rect 1174 1566 1234 1568
rect 1174 1510 1176 1566
rect 1232 1510 1234 1566
rect 1174 1508 1234 1510
rect 1174 28 1234 30
rect 1174 -28 1176 28
rect 1232 -28 1234 28
rect 1174 -30 1234 -28
use contact_18  contact_18_0
timestamp 1643671299
transform 1 0 1174 0 1 24578
box 0 0 1 1
use contact_17  contact_17_0
timestamp 1643671299
transform 1 0 1189 0 1 24593
box 0 0 1 1
use contact_18  contact_18_1
timestamp 1643671299
transform 1 0 1174 0 1 23040
box 0 0 1 1
use contact_17  contact_17_1
timestamp 1643671299
transform 1 0 1189 0 1 23055
box 0 0 1 1
use contact_18  contact_18_2
timestamp 1643671299
transform 1 0 1174 0 1 21502
box 0 0 1 1
use contact_17  contact_17_2
timestamp 1643671299
transform 1 0 1189 0 1 21517
box 0 0 1 1
use contact_18  contact_18_3
timestamp 1643671299
transform 1 0 1174 0 1 23040
box 0 0 1 1
use contact_17  contact_17_3
timestamp 1643671299
transform 1 0 1189 0 1 23055
box 0 0 1 1
use contact_18  contact_18_4
timestamp 1643671299
transform 1 0 1174 0 1 21502
box 0 0 1 1
use contact_17  contact_17_4
timestamp 1643671299
transform 1 0 1189 0 1 21517
box 0 0 1 1
use contact_18  contact_18_5
timestamp 1643671299
transform 1 0 1174 0 1 19964
box 0 0 1 1
use contact_17  contact_17_5
timestamp 1643671299
transform 1 0 1189 0 1 19979
box 0 0 1 1
use contact_18  contact_18_6
timestamp 1643671299
transform 1 0 1174 0 1 18426
box 0 0 1 1
use contact_17  contact_17_6
timestamp 1643671299
transform 1 0 1189 0 1 18441
box 0 0 1 1
use contact_18  contact_18_7
timestamp 1643671299
transform 1 0 1174 0 1 19964
box 0 0 1 1
use contact_17  contact_17_7
timestamp 1643671299
transform 1 0 1189 0 1 19979
box 0 0 1 1
use contact_18  contact_18_8
timestamp 1643671299
transform 1 0 1174 0 1 18426
box 0 0 1 1
use contact_17  contact_17_8
timestamp 1643671299
transform 1 0 1189 0 1 18441
box 0 0 1 1
use contact_18  contact_18_9
timestamp 1643671299
transform 1 0 1174 0 1 16888
box 0 0 1 1
use contact_17  contact_17_9
timestamp 1643671299
transform 1 0 1189 0 1 16903
box 0 0 1 1
use contact_18  contact_18_10
timestamp 1643671299
transform 1 0 1174 0 1 15350
box 0 0 1 1
use contact_17  contact_17_10
timestamp 1643671299
transform 1 0 1189 0 1 15365
box 0 0 1 1
use contact_18  contact_18_11
timestamp 1643671299
transform 1 0 1174 0 1 16888
box 0 0 1 1
use contact_17  contact_17_11
timestamp 1643671299
transform 1 0 1189 0 1 16903
box 0 0 1 1
use contact_18  contact_18_12
timestamp 1643671299
transform 1 0 1174 0 1 15350
box 0 0 1 1
use contact_17  contact_17_12
timestamp 1643671299
transform 1 0 1189 0 1 15365
box 0 0 1 1
use contact_18  contact_18_13
timestamp 1643671299
transform 1 0 1174 0 1 13812
box 0 0 1 1
use contact_17  contact_17_13
timestamp 1643671299
transform 1 0 1189 0 1 13827
box 0 0 1 1
use contact_18  contact_18_14
timestamp 1643671299
transform 1 0 1174 0 1 12274
box 0 0 1 1
use contact_17  contact_17_14
timestamp 1643671299
transform 1 0 1189 0 1 12289
box 0 0 1 1
use contact_18  contact_18_15
timestamp 1643671299
transform 1 0 1174 0 1 13812
box 0 0 1 1
use contact_17  contact_17_15
timestamp 1643671299
transform 1 0 1189 0 1 13827
box 0 0 1 1
use contact_18  contact_18_16
timestamp 1643671299
transform 1 0 1174 0 1 12274
box 0 0 1 1
use contact_17  contact_17_16
timestamp 1643671299
transform 1 0 1189 0 1 12289
box 0 0 1 1
use contact_18  contact_18_17
timestamp 1643671299
transform 1 0 1174 0 1 10736
box 0 0 1 1
use contact_17  contact_17_17
timestamp 1643671299
transform 1 0 1189 0 1 10751
box 0 0 1 1
use contact_18  contact_18_18
timestamp 1643671299
transform 1 0 1174 0 1 9198
box 0 0 1 1
use contact_17  contact_17_18
timestamp 1643671299
transform 1 0 1189 0 1 9213
box 0 0 1 1
use contact_18  contact_18_19
timestamp 1643671299
transform 1 0 1174 0 1 10736
box 0 0 1 1
use contact_17  contact_17_19
timestamp 1643671299
transform 1 0 1189 0 1 10751
box 0 0 1 1
use contact_18  contact_18_20
timestamp 1643671299
transform 1 0 1174 0 1 9198
box 0 0 1 1
use contact_17  contact_17_20
timestamp 1643671299
transform 1 0 1189 0 1 9213
box 0 0 1 1
use contact_18  contact_18_21
timestamp 1643671299
transform 1 0 1174 0 1 7660
box 0 0 1 1
use contact_17  contact_17_21
timestamp 1643671299
transform 1 0 1189 0 1 7675
box 0 0 1 1
use contact_18  contact_18_22
timestamp 1643671299
transform 1 0 1174 0 1 6122
box 0 0 1 1
use contact_17  contact_17_22
timestamp 1643671299
transform 1 0 1189 0 1 6137
box 0 0 1 1
use contact_18  contact_18_23
timestamp 1643671299
transform 1 0 1174 0 1 7660
box 0 0 1 1
use contact_17  contact_17_23
timestamp 1643671299
transform 1 0 1189 0 1 7675
box 0 0 1 1
use contact_18  contact_18_24
timestamp 1643671299
transform 1 0 1174 0 1 6122
box 0 0 1 1
use contact_17  contact_17_24
timestamp 1643671299
transform 1 0 1189 0 1 6137
box 0 0 1 1
use contact_18  contact_18_25
timestamp 1643671299
transform 1 0 1174 0 1 4584
box 0 0 1 1
use contact_17  contact_17_25
timestamp 1643671299
transform 1 0 1189 0 1 4599
box 0 0 1 1
use contact_18  contact_18_26
timestamp 1643671299
transform 1 0 1174 0 1 3046
box 0 0 1 1
use contact_17  contact_17_26
timestamp 1643671299
transform 1 0 1189 0 1 3061
box 0 0 1 1
use contact_18  contact_18_27
timestamp 1643671299
transform 1 0 1174 0 1 4584
box 0 0 1 1
use contact_17  contact_17_27
timestamp 1643671299
transform 1 0 1189 0 1 4599
box 0 0 1 1
use contact_18  contact_18_28
timestamp 1643671299
transform 1 0 1174 0 1 3046
box 0 0 1 1
use contact_17  contact_17_28
timestamp 1643671299
transform 1 0 1189 0 1 3061
box 0 0 1 1
use contact_18  contact_18_29
timestamp 1643671299
transform 1 0 1174 0 1 1508
box 0 0 1 1
use contact_17  contact_17_29
timestamp 1643671299
transform 1 0 1189 0 1 1523
box 0 0 1 1
use contact_18  contact_18_30
timestamp 1643671299
transform 1 0 1174 0 1 -30
box 0 0 1 1
use contact_17  contact_17_30
timestamp 1643671299
transform 1 0 1189 0 1 -15
box 0 0 1 1
use contact_18  contact_18_31
timestamp 1643671299
transform 1 0 1174 0 1 1508
box 0 0 1 1
use contact_17  contact_17_31
timestamp 1643671299
transform 1 0 1189 0 1 1523
box 0 0 1 1
use wordline_driver_cell  wordline_driver_cell_0
timestamp 1643671299
transform 1 0 0 0 -1 24608
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_1
timestamp 1643671299
transform 1 0 0 0 1 21532
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_2
timestamp 1643671299
transform 1 0 0 0 -1 21532
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_3
timestamp 1643671299
transform 1 0 0 0 1 18456
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_4
timestamp 1643671299
transform 1 0 0 0 -1 18456
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_5
timestamp 1643671299
transform 1 0 0 0 1 15380
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_6
timestamp 1643671299
transform 1 0 0 0 -1 15380
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_7
timestamp 1643671299
transform 1 0 0 0 1 12304
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_8
timestamp 1643671299
transform 1 0 0 0 -1 12304
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_9
timestamp 1643671299
transform 1 0 0 0 1 9228
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_10
timestamp 1643671299
transform 1 0 0 0 -1 9228
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_11
timestamp 1643671299
transform 1 0 0 0 1 6152
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_12
timestamp 1643671299
transform 1 0 0 0 -1 6152
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_13
timestamp 1643671299
transform 1 0 0 0 1 3076
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_14
timestamp 1643671299
transform 1 0 0 0 -1 3076
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_15
timestamp 1643671299
transform 1 0 0 0 1 0
box 0 -42 1204 1616
<< labels >>
rlabel metal2 s 0 0 28 24608 4 wl_en
rlabel metal1 s 56 848 126 876 4 in0_0
rlabel metal1 s 234 702 318 730 4 in1_0
rlabel metal1 s 536 582 618 610 4 in2_0
rlabel metal1 s 1176 778 1204 806 4 rwl0_0
rlabel metal1 s 1176 1004 1204 1032 4 rwl1_0
rlabel metal1 s 1176 652 1204 680 4 wwl0_0
rlabel metal1 s 56 2200 126 2228 4 in0_1
rlabel metal1 s 234 2346 318 2374 4 in1_1
rlabel metal1 s 536 2466 618 2494 4 in2_1
rlabel metal1 s 1176 2270 1204 2298 4 rwl0_1
rlabel metal1 s 1176 2044 1204 2072 4 rwl1_1
rlabel metal1 s 1176 2396 1204 2424 4 wwl0_1
rlabel metal1 s 56 3924 126 3952 4 in0_2
rlabel metal1 s 234 3778 318 3806 4 in1_2
rlabel metal1 s 536 3658 618 3686 4 in2_2
rlabel metal1 s 1176 3854 1204 3882 4 rwl0_2
rlabel metal1 s 1176 4080 1204 4108 4 rwl1_2
rlabel metal1 s 1176 3728 1204 3756 4 wwl0_2
rlabel metal1 s 56 5276 126 5304 4 in0_3
rlabel metal1 s 234 5422 318 5450 4 in1_3
rlabel metal1 s 536 5542 618 5570 4 in2_3
rlabel metal1 s 1176 5346 1204 5374 4 rwl0_3
rlabel metal1 s 1176 5120 1204 5148 4 rwl1_3
rlabel metal1 s 1176 5472 1204 5500 4 wwl0_3
rlabel metal1 s 56 7000 126 7028 4 in0_4
rlabel metal1 s 234 6854 318 6882 4 in1_4
rlabel metal1 s 536 6734 618 6762 4 in2_4
rlabel metal1 s 1176 6930 1204 6958 4 rwl0_4
rlabel metal1 s 1176 7156 1204 7184 4 rwl1_4
rlabel metal1 s 1176 6804 1204 6832 4 wwl0_4
rlabel metal1 s 56 8352 126 8380 4 in0_5
rlabel metal1 s 234 8498 318 8526 4 in1_5
rlabel metal1 s 536 8618 618 8646 4 in2_5
rlabel metal1 s 1176 8422 1204 8450 4 rwl0_5
rlabel metal1 s 1176 8196 1204 8224 4 rwl1_5
rlabel metal1 s 1176 8548 1204 8576 4 wwl0_5
rlabel metal1 s 56 10076 126 10104 4 in0_6
rlabel metal1 s 234 9930 318 9958 4 in1_6
rlabel metal1 s 536 9810 618 9838 4 in2_6
rlabel metal1 s 1176 10006 1204 10034 4 rwl0_6
rlabel metal1 s 1176 10232 1204 10260 4 rwl1_6
rlabel metal1 s 1176 9880 1204 9908 4 wwl0_6
rlabel metal1 s 56 11428 126 11456 4 in0_7
rlabel metal1 s 234 11574 318 11602 4 in1_7
rlabel metal1 s 536 11694 618 11722 4 in2_7
rlabel metal1 s 1176 11498 1204 11526 4 rwl0_7
rlabel metal1 s 1176 11272 1204 11300 4 rwl1_7
rlabel metal1 s 1176 11624 1204 11652 4 wwl0_7
rlabel metal1 s 56 13152 126 13180 4 in0_8
rlabel metal1 s 234 13006 318 13034 4 in1_8
rlabel metal1 s 536 12886 618 12914 4 in2_8
rlabel metal1 s 1176 13082 1204 13110 4 rwl0_8
rlabel metal1 s 1176 13308 1204 13336 4 rwl1_8
rlabel metal1 s 1176 12956 1204 12984 4 wwl0_8
rlabel metal1 s 56 14504 126 14532 4 in0_9
rlabel metal1 s 234 14650 318 14678 4 in1_9
rlabel metal1 s 536 14770 618 14798 4 in2_9
rlabel metal1 s 1176 14574 1204 14602 4 rwl0_9
rlabel metal1 s 1176 14348 1204 14376 4 rwl1_9
rlabel metal1 s 1176 14700 1204 14728 4 wwl0_9
rlabel metal1 s 56 16228 126 16256 4 in0_10
rlabel metal1 s 234 16082 318 16110 4 in1_10
rlabel metal1 s 536 15962 618 15990 4 in2_10
rlabel metal1 s 1176 16158 1204 16186 4 rwl0_10
rlabel metal1 s 1176 16384 1204 16412 4 rwl1_10
rlabel metal1 s 1176 16032 1204 16060 4 wwl0_10
rlabel metal1 s 56 17580 126 17608 4 in0_11
rlabel metal1 s 234 17726 318 17754 4 in1_11
rlabel metal1 s 536 17846 618 17874 4 in2_11
rlabel metal1 s 1176 17650 1204 17678 4 rwl0_11
rlabel metal1 s 1176 17424 1204 17452 4 rwl1_11
rlabel metal1 s 1176 17776 1204 17804 4 wwl0_11
rlabel metal1 s 56 19304 126 19332 4 in0_12
rlabel metal1 s 234 19158 318 19186 4 in1_12
rlabel metal1 s 536 19038 618 19066 4 in2_12
rlabel metal1 s 1176 19234 1204 19262 4 rwl0_12
rlabel metal1 s 1176 19460 1204 19488 4 rwl1_12
rlabel metal1 s 1176 19108 1204 19136 4 wwl0_12
rlabel metal1 s 56 20656 126 20684 4 in0_13
rlabel metal1 s 234 20802 318 20830 4 in1_13
rlabel metal1 s 536 20922 618 20950 4 in2_13
rlabel metal1 s 1176 20726 1204 20754 4 rwl0_13
rlabel metal1 s 1176 20500 1204 20528 4 rwl1_13
rlabel metal1 s 1176 20852 1204 20880 4 wwl0_13
rlabel metal1 s 56 22380 126 22408 4 in0_14
rlabel metal1 s 234 22234 318 22262 4 in1_14
rlabel metal1 s 536 22114 618 22142 4 in2_14
rlabel metal1 s 1176 22310 1204 22338 4 rwl0_14
rlabel metal1 s 1176 22536 1204 22564 4 rwl1_14
rlabel metal1 s 1176 22184 1204 22212 4 wwl0_14
rlabel metal1 s 56 23732 126 23760 4 in0_15
rlabel metal1 s 234 23878 318 23906 4 in1_15
rlabel metal1 s 536 23998 618 24026 4 in2_15
rlabel metal1 s 1176 23802 1204 23830 4 rwl0_15
rlabel metal1 s 1176 23576 1204 23604 4 rwl1_15
rlabel metal1 s 1176 23928 1204 23956 4 wwl0_15
rlabel metal3 s 1174 10736 1234 10796 4 vdd
rlabel metal3 s 1204 10766 1204 10766 4 vdd
rlabel metal3 s 1174 23040 1234 23100 4 vdd
rlabel metal3 s 1174 7660 1234 7720 4 vdd
rlabel metal3 s 1174 4584 1234 4644 4 vdd
rlabel metal3 s 1174 1508 1234 1568 4 vdd
rlabel metal3 s 1174 16888 1234 16948 4 vdd
rlabel metal3 s 1174 19964 1234 20024 4 vdd
rlabel metal3 s 1204 1538 1204 1538 4 vdd
rlabel metal3 s 1174 13812 1234 13872 4 vdd
rlabel metal3 s 1174 18426 1234 18486 4 gnd
rlabel metal3 s 1174 6122 1234 6182 4 gnd
rlabel metal3 s 1174 -30 1234 30 4 gnd
rlabel metal3 s 1174 21502 1234 21562 4 gnd
rlabel metal3 s 1174 12274 1234 12334 4 gnd
rlabel metal3 s 1174 9198 1234 9258 4 gnd
rlabel metal3 s 1174 15350 1234 15410 4 gnd
rlabel metal3 s 1174 24578 1234 24638 4 gnd
rlabel metal3 s 1174 3046 1234 3106 4 gnd
<< properties >>
string FIXED_BBOX 1174 -30 1234 0
string GDS_FILE sram_0rw2r1w_16_32_sky130A.gds
string GDS_END 1077578
string GDS_START 1049208
<< end >>
