magic
tech sky130A
magscale 1 2
timestamp 1644951705
<< checkpaint >>
rect -1296 -1277 4202 2155
<< locali >>
rect 0 821 2906 855
rect 196 381 262 447
rect 330 388 364 561
rect 330 354 459 388
rect 1639 354 1673 388
rect 96 257 162 323
rect 0 -17 2906 17
use pdriver_3  pdriver_3_0
timestamp 1644951705
transform 1 0 378 0 1 0
box -36 -17 2564 895
use pnand2_0  pnand2_0_0
timestamp 1644951705
transform 1 0 0 0 1 0
box -36 -17 414 895
<< labels >>
rlabel locali s 1656 371 1656 371 4 Z
rlabel locali s 129 290 129 290 4 A
rlabel locali s 229 414 229 414 4 B
rlabel locali s 1453 0 1453 0 4 gnd
rlabel locali s 1453 838 1453 838 4 vdd
<< properties >>
string FIXED_BBOX 0 0 2906 838
string GDS_FILE sram_0rw2r1w_16_128_sky130A.gds
string GDS_END 2041634
string GDS_START 2040500
<< end >>
