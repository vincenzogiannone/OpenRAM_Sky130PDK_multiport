magic
tech sky130A
magscale 1 2
timestamp 1643593061
<< checkpaint >>
rect -1319 -1316 2765 1605
<< nwell >>
rect -54 229 1500 345
rect -59 61 1505 229
rect -54 -54 1500 61
<< scpmos >>
rect 60 0 90 291
rect 168 0 198 291
rect 276 0 306 291
rect 384 0 414 291
rect 492 0 522 291
rect 600 0 630 291
rect 708 0 738 291
rect 816 0 846 291
rect 924 0 954 291
rect 1032 0 1062 291
rect 1140 0 1170 291
rect 1248 0 1278 291
rect 1356 0 1386 291
<< pdiff >>
rect 0 162 60 291
rect 0 128 8 162
rect 42 128 60 162
rect 0 0 60 128
rect 90 162 168 291
rect 90 128 112 162
rect 146 128 168 162
rect 90 0 168 128
rect 198 162 276 291
rect 198 128 220 162
rect 254 128 276 162
rect 198 0 276 128
rect 306 162 384 291
rect 306 128 328 162
rect 362 128 384 162
rect 306 0 384 128
rect 414 162 492 291
rect 414 128 436 162
rect 470 128 492 162
rect 414 0 492 128
rect 522 162 600 291
rect 522 128 544 162
rect 578 128 600 162
rect 522 0 600 128
rect 630 162 708 291
rect 630 128 652 162
rect 686 128 708 162
rect 630 0 708 128
rect 738 162 816 291
rect 738 128 760 162
rect 794 128 816 162
rect 738 0 816 128
rect 846 162 924 291
rect 846 128 868 162
rect 902 128 924 162
rect 846 0 924 128
rect 954 162 1032 291
rect 954 128 976 162
rect 1010 128 1032 162
rect 954 0 1032 128
rect 1062 162 1140 291
rect 1062 128 1084 162
rect 1118 128 1140 162
rect 1062 0 1140 128
rect 1170 162 1248 291
rect 1170 128 1192 162
rect 1226 128 1248 162
rect 1170 0 1248 128
rect 1278 162 1356 291
rect 1278 128 1300 162
rect 1334 128 1356 162
rect 1278 0 1356 128
rect 1386 162 1446 291
rect 1386 128 1404 162
rect 1438 128 1446 162
rect 1386 0 1446 128
<< pdiffc >>
rect 8 128 42 162
rect 112 128 146 162
rect 220 128 254 162
rect 328 128 362 162
rect 436 128 470 162
rect 544 128 578 162
rect 652 128 686 162
rect 760 128 794 162
rect 868 128 902 162
rect 976 128 1010 162
rect 1084 128 1118 162
rect 1192 128 1226 162
rect 1300 128 1334 162
rect 1404 128 1438 162
<< poly >>
rect 60 291 90 317
rect 168 291 198 317
rect 276 291 306 317
rect 384 291 414 317
rect 492 291 522 317
rect 600 291 630 317
rect 708 291 738 317
rect 816 291 846 317
rect 924 291 954 317
rect 1032 291 1062 317
rect 1140 291 1170 317
rect 1248 291 1278 317
rect 1356 291 1386 317
rect 60 -26 90 0
rect 168 -26 198 0
rect 276 -26 306 0
rect 384 -26 414 0
rect 492 -26 522 0
rect 600 -26 630 0
rect 708 -26 738 0
rect 816 -26 846 0
rect 924 -26 954 0
rect 1032 -26 1062 0
rect 1140 -26 1170 0
rect 1248 -26 1278 0
rect 1356 -26 1386 0
rect 60 -56 1386 -26
<< locali >>
rect 8 162 42 178
rect 8 112 42 128
rect 112 162 146 178
rect 112 78 146 128
rect 220 162 254 178
rect 220 112 254 128
rect 328 162 362 178
rect 328 78 362 128
rect 436 162 470 178
rect 436 112 470 128
rect 544 162 578 178
rect 544 78 578 128
rect 652 162 686 178
rect 652 112 686 128
rect 760 162 794 178
rect 760 78 794 128
rect 868 162 902 178
rect 868 112 902 128
rect 976 162 1010 178
rect 976 78 1010 128
rect 1084 162 1118 178
rect 1084 112 1118 128
rect 1192 162 1226 178
rect 1192 78 1226 128
rect 1300 162 1334 178
rect 1300 112 1334 128
rect 1404 162 1438 178
rect 1404 78 1438 128
rect 112 44 1438 78
use contact_9  contact_9_0
timestamp 1643593061
transform 1 0 1396 0 1 104
box 0 0 2 2
use contact_9  contact_9_1
timestamp 1643593061
transform 1 0 1292 0 1 104
box 0 0 2 2
use contact_9  contact_9_2
timestamp 1643593061
transform 1 0 1184 0 1 104
box 0 0 2 2
use contact_9  contact_9_3
timestamp 1643593061
transform 1 0 1076 0 1 104
box 0 0 2 2
use contact_9  contact_9_4
timestamp 1643593061
transform 1 0 968 0 1 104
box 0 0 2 2
use contact_9  contact_9_5
timestamp 1643593061
transform 1 0 860 0 1 104
box 0 0 2 2
use contact_9  contact_9_6
timestamp 1643593061
transform 1 0 752 0 1 104
box 0 0 2 2
use contact_9  contact_9_7
timestamp 1643593061
transform 1 0 644 0 1 104
box 0 0 2 2
use contact_9  contact_9_8
timestamp 1643593061
transform 1 0 536 0 1 104
box 0 0 2 2
use contact_9  contact_9_9
timestamp 1643593061
transform 1 0 428 0 1 104
box 0 0 2 2
use contact_9  contact_9_10
timestamp 1643593061
transform 1 0 320 0 1 104
box 0 0 2 2
use contact_9  contact_9_11
timestamp 1643593061
transform 1 0 212 0 1 104
box 0 0 2 2
use contact_9  contact_9_12
timestamp 1643593061
transform 1 0 104 0 1 104
box 0 0 2 2
use contact_9  contact_9_13
timestamp 1643593061
transform 1 0 0 0 1 104
box 0 0 2 2
<< labels >>
rlabel mvvaractor s 723 -41 723 -41 4 G
rlabel locali s 669 145 669 145 4 S
rlabel locali s 453 145 453 145 4 S
rlabel locali s 237 145 237 145 4 S
rlabel locali s 1317 145 1317 145 4 S
rlabel locali s 25 145 25 145 4 S
rlabel locali s 1101 145 1101 145 4 S
rlabel locali s 885 145 885 145 4 S
rlabel locali s 775 61 775 61 4 D
<< properties >>
string FIXED_BBOX -54 -56 1500 61
string GDS_FILE sram_0rw2r1w_2_16_sky130A.gds
string GDS_END 539860
string GDS_START 536616
<< end >>
