magic
tech sky130A
magscale 1 2
timestamp 1644969367
<< checkpaint >>
rect -1299 -1302 2742 2176
<< metal1 >>
rect 709 812 715 864
rect 767 812 773 864
rect 709 -26 715 26
rect 767 -26 773 26
<< via1 >>
rect 715 812 767 864
rect 715 -26 767 26
<< metal2 >>
rect 713 866 769 875
rect 0 345 28 838
rect 713 801 769 810
rect -1 336 55 345
rect -1 271 55 280
rect 0 0 28 271
rect 180 232 234 260
rect 1260 228 1314 256
rect 713 28 769 37
rect 713 -37 769 -28
<< via2 >>
rect 713 864 769 866
rect 713 812 715 864
rect 715 812 767 864
rect 767 812 769 864
rect 713 810 769 812
rect -1 280 55 336
rect 713 26 769 28
rect 713 -26 715 26
rect 715 -26 767 26
rect 767 -26 769 26
rect 713 -28 769 -26
<< metal3 >>
rect 675 866 807 875
rect 675 810 713 866
rect 769 810 807 866
rect 675 801 807 810
rect -39 338 93 341
rect -39 336 1482 338
rect -39 280 -1 336
rect 55 280 1482 336
rect -39 278 1482 280
rect -39 275 93 278
rect 675 28 807 37
rect 675 -28 713 28
rect 769 -28 807 28
rect 675 -37 807 -28
use contact_18  contact_18_0
timestamp 1644969367
transform 1 0 -39 0 1 271
box 0 0 1 1
use contact_18  contact_18_1
timestamp 1644969367
transform 1 0 675 0 1 -37
box 0 0 1 1
use contact_17  contact_17_0
timestamp 1644969367
transform 1 0 709 0 1 -32
box 0 0 1 1
use contact_18  contact_18_2
timestamp 1644969367
transform 1 0 675 0 1 801
box 0 0 1 1
use contact_17  contact_17_1
timestamp 1644969367
transform 1 0 709 0 1 806
box 0 0 1 1
use dff  dff_0
timestamp 1644969367
transform 1 0 0 0 1 0
box 0 -42 1482 916
<< labels >>
rlabel metal3 s 675 801 807 875 4 vdd
rlabel metal3 s 675 -37 807 37 4 gnd
rlabel metal2 s 180 232 234 260 4 din_0
rlabel metal2 s 1260 228 1314 256 4 dout_0
rlabel metal3 s 0 278 1482 338 4 clk
<< properties >>
string FIXED_BBOX 675 -37 807 0
string GDS_FILE sram_0rw2r1w_32_128_sky130A.gds
string GDS_END 3427570
string GDS_START 3426078
<< end >>
