magic
tech sky130A
magscale 1 2
timestamp 1643671299
<< checkpaint >>
rect -1260 -1260 76562 38762
<< dnwell >>
rect 1618 1564 73966 36208
<< nwell >>
rect 1534 36124 74050 36292
rect 1534 1648 1702 36124
rect 73882 1648 74050 36124
rect 1534 1480 74050 1648
<< nsubdiff >>
rect 1929 36225 1979 36249
rect 1929 36191 1937 36225
rect 1971 36191 1979 36225
rect 1929 36167 1979 36191
rect 2265 36225 2315 36249
rect 2265 36191 2273 36225
rect 2307 36191 2315 36225
rect 2265 36167 2315 36191
rect 2601 36225 2651 36249
rect 2601 36191 2609 36225
rect 2643 36191 2651 36225
rect 2601 36167 2651 36191
rect 2937 36225 2987 36249
rect 2937 36191 2945 36225
rect 2979 36191 2987 36225
rect 2937 36167 2987 36191
rect 3273 36225 3323 36249
rect 3273 36191 3281 36225
rect 3315 36191 3323 36225
rect 3273 36167 3323 36191
rect 3609 36225 3659 36249
rect 3609 36191 3617 36225
rect 3651 36191 3659 36225
rect 3609 36167 3659 36191
rect 3945 36225 3995 36249
rect 3945 36191 3953 36225
rect 3987 36191 3995 36225
rect 3945 36167 3995 36191
rect 4281 36225 4331 36249
rect 4281 36191 4289 36225
rect 4323 36191 4331 36225
rect 4281 36167 4331 36191
rect 4617 36225 4667 36249
rect 4617 36191 4625 36225
rect 4659 36191 4667 36225
rect 4617 36167 4667 36191
rect 4953 36225 5003 36249
rect 4953 36191 4961 36225
rect 4995 36191 5003 36225
rect 4953 36167 5003 36191
rect 5289 36225 5339 36249
rect 5289 36191 5297 36225
rect 5331 36191 5339 36225
rect 5289 36167 5339 36191
rect 5625 36225 5675 36249
rect 5625 36191 5633 36225
rect 5667 36191 5675 36225
rect 5625 36167 5675 36191
rect 5961 36225 6011 36249
rect 5961 36191 5969 36225
rect 6003 36191 6011 36225
rect 5961 36167 6011 36191
rect 6297 36225 6347 36249
rect 6297 36191 6305 36225
rect 6339 36191 6347 36225
rect 6297 36167 6347 36191
rect 6633 36225 6683 36249
rect 6633 36191 6641 36225
rect 6675 36191 6683 36225
rect 6633 36167 6683 36191
rect 6969 36225 7019 36249
rect 6969 36191 6977 36225
rect 7011 36191 7019 36225
rect 6969 36167 7019 36191
rect 7305 36225 7355 36249
rect 7305 36191 7313 36225
rect 7347 36191 7355 36225
rect 7305 36167 7355 36191
rect 7641 36225 7691 36249
rect 7641 36191 7649 36225
rect 7683 36191 7691 36225
rect 7641 36167 7691 36191
rect 7977 36225 8027 36249
rect 7977 36191 7985 36225
rect 8019 36191 8027 36225
rect 7977 36167 8027 36191
rect 8313 36225 8363 36249
rect 8313 36191 8321 36225
rect 8355 36191 8363 36225
rect 8313 36167 8363 36191
rect 8649 36225 8699 36249
rect 8649 36191 8657 36225
rect 8691 36191 8699 36225
rect 8649 36167 8699 36191
rect 8985 36225 9035 36249
rect 8985 36191 8993 36225
rect 9027 36191 9035 36225
rect 8985 36167 9035 36191
rect 9321 36225 9371 36249
rect 9321 36191 9329 36225
rect 9363 36191 9371 36225
rect 9321 36167 9371 36191
rect 9657 36225 9707 36249
rect 9657 36191 9665 36225
rect 9699 36191 9707 36225
rect 9657 36167 9707 36191
rect 9993 36225 10043 36249
rect 9993 36191 10001 36225
rect 10035 36191 10043 36225
rect 9993 36167 10043 36191
rect 10329 36225 10379 36249
rect 10329 36191 10337 36225
rect 10371 36191 10379 36225
rect 10329 36167 10379 36191
rect 10665 36225 10715 36249
rect 10665 36191 10673 36225
rect 10707 36191 10715 36225
rect 10665 36167 10715 36191
rect 11001 36225 11051 36249
rect 11001 36191 11009 36225
rect 11043 36191 11051 36225
rect 11001 36167 11051 36191
rect 11337 36225 11387 36249
rect 11337 36191 11345 36225
rect 11379 36191 11387 36225
rect 11337 36167 11387 36191
rect 11673 36225 11723 36249
rect 11673 36191 11681 36225
rect 11715 36191 11723 36225
rect 11673 36167 11723 36191
rect 12009 36225 12059 36249
rect 12009 36191 12017 36225
rect 12051 36191 12059 36225
rect 12009 36167 12059 36191
rect 12345 36225 12395 36249
rect 12345 36191 12353 36225
rect 12387 36191 12395 36225
rect 12345 36167 12395 36191
rect 12681 36225 12731 36249
rect 12681 36191 12689 36225
rect 12723 36191 12731 36225
rect 12681 36167 12731 36191
rect 13017 36225 13067 36249
rect 13017 36191 13025 36225
rect 13059 36191 13067 36225
rect 13017 36167 13067 36191
rect 13353 36225 13403 36249
rect 13353 36191 13361 36225
rect 13395 36191 13403 36225
rect 13353 36167 13403 36191
rect 13689 36225 13739 36249
rect 13689 36191 13697 36225
rect 13731 36191 13739 36225
rect 13689 36167 13739 36191
rect 14025 36225 14075 36249
rect 14025 36191 14033 36225
rect 14067 36191 14075 36225
rect 14025 36167 14075 36191
rect 14361 36225 14411 36249
rect 14361 36191 14369 36225
rect 14403 36191 14411 36225
rect 14361 36167 14411 36191
rect 14697 36225 14747 36249
rect 14697 36191 14705 36225
rect 14739 36191 14747 36225
rect 14697 36167 14747 36191
rect 15033 36225 15083 36249
rect 15033 36191 15041 36225
rect 15075 36191 15083 36225
rect 15033 36167 15083 36191
rect 15369 36225 15419 36249
rect 15369 36191 15377 36225
rect 15411 36191 15419 36225
rect 15369 36167 15419 36191
rect 15705 36225 15755 36249
rect 15705 36191 15713 36225
rect 15747 36191 15755 36225
rect 15705 36167 15755 36191
rect 16041 36225 16091 36249
rect 16041 36191 16049 36225
rect 16083 36191 16091 36225
rect 16041 36167 16091 36191
rect 16377 36225 16427 36249
rect 16377 36191 16385 36225
rect 16419 36191 16427 36225
rect 16377 36167 16427 36191
rect 16713 36225 16763 36249
rect 16713 36191 16721 36225
rect 16755 36191 16763 36225
rect 16713 36167 16763 36191
rect 17049 36225 17099 36249
rect 17049 36191 17057 36225
rect 17091 36191 17099 36225
rect 17049 36167 17099 36191
rect 17385 36225 17435 36249
rect 17385 36191 17393 36225
rect 17427 36191 17435 36225
rect 17385 36167 17435 36191
rect 17721 36225 17771 36249
rect 17721 36191 17729 36225
rect 17763 36191 17771 36225
rect 17721 36167 17771 36191
rect 18057 36225 18107 36249
rect 18057 36191 18065 36225
rect 18099 36191 18107 36225
rect 18057 36167 18107 36191
rect 18393 36225 18443 36249
rect 18393 36191 18401 36225
rect 18435 36191 18443 36225
rect 18393 36167 18443 36191
rect 18729 36225 18779 36249
rect 18729 36191 18737 36225
rect 18771 36191 18779 36225
rect 18729 36167 18779 36191
rect 19065 36225 19115 36249
rect 19065 36191 19073 36225
rect 19107 36191 19115 36225
rect 19065 36167 19115 36191
rect 19401 36225 19451 36249
rect 19401 36191 19409 36225
rect 19443 36191 19451 36225
rect 19401 36167 19451 36191
rect 19737 36225 19787 36249
rect 19737 36191 19745 36225
rect 19779 36191 19787 36225
rect 19737 36167 19787 36191
rect 20073 36225 20123 36249
rect 20073 36191 20081 36225
rect 20115 36191 20123 36225
rect 20073 36167 20123 36191
rect 20409 36225 20459 36249
rect 20409 36191 20417 36225
rect 20451 36191 20459 36225
rect 20409 36167 20459 36191
rect 20745 36225 20795 36249
rect 20745 36191 20753 36225
rect 20787 36191 20795 36225
rect 20745 36167 20795 36191
rect 21081 36225 21131 36249
rect 21081 36191 21089 36225
rect 21123 36191 21131 36225
rect 21081 36167 21131 36191
rect 21417 36225 21467 36249
rect 21417 36191 21425 36225
rect 21459 36191 21467 36225
rect 21417 36167 21467 36191
rect 21753 36225 21803 36249
rect 21753 36191 21761 36225
rect 21795 36191 21803 36225
rect 21753 36167 21803 36191
rect 22089 36225 22139 36249
rect 22089 36191 22097 36225
rect 22131 36191 22139 36225
rect 22089 36167 22139 36191
rect 22425 36225 22475 36249
rect 22425 36191 22433 36225
rect 22467 36191 22475 36225
rect 22425 36167 22475 36191
rect 22761 36225 22811 36249
rect 22761 36191 22769 36225
rect 22803 36191 22811 36225
rect 22761 36167 22811 36191
rect 23097 36225 23147 36249
rect 23097 36191 23105 36225
rect 23139 36191 23147 36225
rect 23097 36167 23147 36191
rect 23433 36225 23483 36249
rect 23433 36191 23441 36225
rect 23475 36191 23483 36225
rect 23433 36167 23483 36191
rect 23769 36225 23819 36249
rect 23769 36191 23777 36225
rect 23811 36191 23819 36225
rect 23769 36167 23819 36191
rect 24105 36225 24155 36249
rect 24105 36191 24113 36225
rect 24147 36191 24155 36225
rect 24105 36167 24155 36191
rect 24441 36225 24491 36249
rect 24441 36191 24449 36225
rect 24483 36191 24491 36225
rect 24441 36167 24491 36191
rect 24777 36225 24827 36249
rect 24777 36191 24785 36225
rect 24819 36191 24827 36225
rect 24777 36167 24827 36191
rect 25113 36225 25163 36249
rect 25113 36191 25121 36225
rect 25155 36191 25163 36225
rect 25113 36167 25163 36191
rect 25449 36225 25499 36249
rect 25449 36191 25457 36225
rect 25491 36191 25499 36225
rect 25449 36167 25499 36191
rect 25785 36225 25835 36249
rect 25785 36191 25793 36225
rect 25827 36191 25835 36225
rect 25785 36167 25835 36191
rect 26121 36225 26171 36249
rect 26121 36191 26129 36225
rect 26163 36191 26171 36225
rect 26121 36167 26171 36191
rect 26457 36225 26507 36249
rect 26457 36191 26465 36225
rect 26499 36191 26507 36225
rect 26457 36167 26507 36191
rect 26793 36225 26843 36249
rect 26793 36191 26801 36225
rect 26835 36191 26843 36225
rect 26793 36167 26843 36191
rect 27129 36225 27179 36249
rect 27129 36191 27137 36225
rect 27171 36191 27179 36225
rect 27129 36167 27179 36191
rect 27465 36225 27515 36249
rect 27465 36191 27473 36225
rect 27507 36191 27515 36225
rect 27465 36167 27515 36191
rect 27801 36225 27851 36249
rect 27801 36191 27809 36225
rect 27843 36191 27851 36225
rect 27801 36167 27851 36191
rect 28137 36225 28187 36249
rect 28137 36191 28145 36225
rect 28179 36191 28187 36225
rect 28137 36167 28187 36191
rect 28473 36225 28523 36249
rect 28473 36191 28481 36225
rect 28515 36191 28523 36225
rect 28473 36167 28523 36191
rect 28809 36225 28859 36249
rect 28809 36191 28817 36225
rect 28851 36191 28859 36225
rect 28809 36167 28859 36191
rect 29145 36225 29195 36249
rect 29145 36191 29153 36225
rect 29187 36191 29195 36225
rect 29145 36167 29195 36191
rect 29481 36225 29531 36249
rect 29481 36191 29489 36225
rect 29523 36191 29531 36225
rect 29481 36167 29531 36191
rect 29817 36225 29867 36249
rect 29817 36191 29825 36225
rect 29859 36191 29867 36225
rect 29817 36167 29867 36191
rect 30153 36225 30203 36249
rect 30153 36191 30161 36225
rect 30195 36191 30203 36225
rect 30153 36167 30203 36191
rect 30489 36225 30539 36249
rect 30489 36191 30497 36225
rect 30531 36191 30539 36225
rect 30489 36167 30539 36191
rect 30825 36225 30875 36249
rect 30825 36191 30833 36225
rect 30867 36191 30875 36225
rect 30825 36167 30875 36191
rect 31161 36225 31211 36249
rect 31161 36191 31169 36225
rect 31203 36191 31211 36225
rect 31161 36167 31211 36191
rect 31497 36225 31547 36249
rect 31497 36191 31505 36225
rect 31539 36191 31547 36225
rect 31497 36167 31547 36191
rect 31833 36225 31883 36249
rect 31833 36191 31841 36225
rect 31875 36191 31883 36225
rect 31833 36167 31883 36191
rect 32169 36225 32219 36249
rect 32169 36191 32177 36225
rect 32211 36191 32219 36225
rect 32169 36167 32219 36191
rect 32505 36225 32555 36249
rect 32505 36191 32513 36225
rect 32547 36191 32555 36225
rect 32505 36167 32555 36191
rect 32841 36225 32891 36249
rect 32841 36191 32849 36225
rect 32883 36191 32891 36225
rect 32841 36167 32891 36191
rect 33177 36225 33227 36249
rect 33177 36191 33185 36225
rect 33219 36191 33227 36225
rect 33177 36167 33227 36191
rect 33513 36225 33563 36249
rect 33513 36191 33521 36225
rect 33555 36191 33563 36225
rect 33513 36167 33563 36191
rect 33849 36225 33899 36249
rect 33849 36191 33857 36225
rect 33891 36191 33899 36225
rect 33849 36167 33899 36191
rect 34185 36225 34235 36249
rect 34185 36191 34193 36225
rect 34227 36191 34235 36225
rect 34185 36167 34235 36191
rect 34521 36225 34571 36249
rect 34521 36191 34529 36225
rect 34563 36191 34571 36225
rect 34521 36167 34571 36191
rect 34857 36225 34907 36249
rect 34857 36191 34865 36225
rect 34899 36191 34907 36225
rect 34857 36167 34907 36191
rect 35193 36225 35243 36249
rect 35193 36191 35201 36225
rect 35235 36191 35243 36225
rect 35193 36167 35243 36191
rect 35529 36225 35579 36249
rect 35529 36191 35537 36225
rect 35571 36191 35579 36225
rect 35529 36167 35579 36191
rect 35865 36225 35915 36249
rect 35865 36191 35873 36225
rect 35907 36191 35915 36225
rect 35865 36167 35915 36191
rect 36201 36225 36251 36249
rect 36201 36191 36209 36225
rect 36243 36191 36251 36225
rect 36201 36167 36251 36191
rect 36537 36225 36587 36249
rect 36537 36191 36545 36225
rect 36579 36191 36587 36225
rect 36537 36167 36587 36191
rect 36873 36225 36923 36249
rect 36873 36191 36881 36225
rect 36915 36191 36923 36225
rect 36873 36167 36923 36191
rect 37209 36225 37259 36249
rect 37209 36191 37217 36225
rect 37251 36191 37259 36225
rect 37209 36167 37259 36191
rect 37545 36225 37595 36249
rect 37545 36191 37553 36225
rect 37587 36191 37595 36225
rect 37545 36167 37595 36191
rect 37881 36225 37931 36249
rect 37881 36191 37889 36225
rect 37923 36191 37931 36225
rect 37881 36167 37931 36191
rect 38217 36225 38267 36249
rect 38217 36191 38225 36225
rect 38259 36191 38267 36225
rect 38217 36167 38267 36191
rect 38553 36225 38603 36249
rect 38553 36191 38561 36225
rect 38595 36191 38603 36225
rect 38553 36167 38603 36191
rect 38889 36225 38939 36249
rect 38889 36191 38897 36225
rect 38931 36191 38939 36225
rect 38889 36167 38939 36191
rect 39225 36225 39275 36249
rect 39225 36191 39233 36225
rect 39267 36191 39275 36225
rect 39225 36167 39275 36191
rect 39561 36225 39611 36249
rect 39561 36191 39569 36225
rect 39603 36191 39611 36225
rect 39561 36167 39611 36191
rect 39897 36225 39947 36249
rect 39897 36191 39905 36225
rect 39939 36191 39947 36225
rect 39897 36167 39947 36191
rect 40233 36225 40283 36249
rect 40233 36191 40241 36225
rect 40275 36191 40283 36225
rect 40233 36167 40283 36191
rect 40569 36225 40619 36249
rect 40569 36191 40577 36225
rect 40611 36191 40619 36225
rect 40569 36167 40619 36191
rect 40905 36225 40955 36249
rect 40905 36191 40913 36225
rect 40947 36191 40955 36225
rect 40905 36167 40955 36191
rect 41241 36225 41291 36249
rect 41241 36191 41249 36225
rect 41283 36191 41291 36225
rect 41241 36167 41291 36191
rect 41577 36225 41627 36249
rect 41577 36191 41585 36225
rect 41619 36191 41627 36225
rect 41577 36167 41627 36191
rect 41913 36225 41963 36249
rect 41913 36191 41921 36225
rect 41955 36191 41963 36225
rect 41913 36167 41963 36191
rect 42249 36225 42299 36249
rect 42249 36191 42257 36225
rect 42291 36191 42299 36225
rect 42249 36167 42299 36191
rect 42585 36225 42635 36249
rect 42585 36191 42593 36225
rect 42627 36191 42635 36225
rect 42585 36167 42635 36191
rect 42921 36225 42971 36249
rect 42921 36191 42929 36225
rect 42963 36191 42971 36225
rect 42921 36167 42971 36191
rect 43257 36225 43307 36249
rect 43257 36191 43265 36225
rect 43299 36191 43307 36225
rect 43257 36167 43307 36191
rect 43593 36225 43643 36249
rect 43593 36191 43601 36225
rect 43635 36191 43643 36225
rect 43593 36167 43643 36191
rect 43929 36225 43979 36249
rect 43929 36191 43937 36225
rect 43971 36191 43979 36225
rect 43929 36167 43979 36191
rect 44265 36225 44315 36249
rect 44265 36191 44273 36225
rect 44307 36191 44315 36225
rect 44265 36167 44315 36191
rect 44601 36225 44651 36249
rect 44601 36191 44609 36225
rect 44643 36191 44651 36225
rect 44601 36167 44651 36191
rect 44937 36225 44987 36249
rect 44937 36191 44945 36225
rect 44979 36191 44987 36225
rect 44937 36167 44987 36191
rect 45273 36225 45323 36249
rect 45273 36191 45281 36225
rect 45315 36191 45323 36225
rect 45273 36167 45323 36191
rect 45609 36225 45659 36249
rect 45609 36191 45617 36225
rect 45651 36191 45659 36225
rect 45609 36167 45659 36191
rect 45945 36225 45995 36249
rect 45945 36191 45953 36225
rect 45987 36191 45995 36225
rect 45945 36167 45995 36191
rect 46281 36225 46331 36249
rect 46281 36191 46289 36225
rect 46323 36191 46331 36225
rect 46281 36167 46331 36191
rect 46617 36225 46667 36249
rect 46617 36191 46625 36225
rect 46659 36191 46667 36225
rect 46617 36167 46667 36191
rect 46953 36225 47003 36249
rect 46953 36191 46961 36225
rect 46995 36191 47003 36225
rect 46953 36167 47003 36191
rect 47289 36225 47339 36249
rect 47289 36191 47297 36225
rect 47331 36191 47339 36225
rect 47289 36167 47339 36191
rect 47625 36225 47675 36249
rect 47625 36191 47633 36225
rect 47667 36191 47675 36225
rect 47625 36167 47675 36191
rect 47961 36225 48011 36249
rect 47961 36191 47969 36225
rect 48003 36191 48011 36225
rect 47961 36167 48011 36191
rect 48297 36225 48347 36249
rect 48297 36191 48305 36225
rect 48339 36191 48347 36225
rect 48297 36167 48347 36191
rect 48633 36225 48683 36249
rect 48633 36191 48641 36225
rect 48675 36191 48683 36225
rect 48633 36167 48683 36191
rect 48969 36225 49019 36249
rect 48969 36191 48977 36225
rect 49011 36191 49019 36225
rect 48969 36167 49019 36191
rect 49305 36225 49355 36249
rect 49305 36191 49313 36225
rect 49347 36191 49355 36225
rect 49305 36167 49355 36191
rect 49641 36225 49691 36249
rect 49641 36191 49649 36225
rect 49683 36191 49691 36225
rect 49641 36167 49691 36191
rect 49977 36225 50027 36249
rect 49977 36191 49985 36225
rect 50019 36191 50027 36225
rect 49977 36167 50027 36191
rect 50313 36225 50363 36249
rect 50313 36191 50321 36225
rect 50355 36191 50363 36225
rect 50313 36167 50363 36191
rect 50649 36225 50699 36249
rect 50649 36191 50657 36225
rect 50691 36191 50699 36225
rect 50649 36167 50699 36191
rect 50985 36225 51035 36249
rect 50985 36191 50993 36225
rect 51027 36191 51035 36225
rect 50985 36167 51035 36191
rect 51321 36225 51371 36249
rect 51321 36191 51329 36225
rect 51363 36191 51371 36225
rect 51321 36167 51371 36191
rect 51657 36225 51707 36249
rect 51657 36191 51665 36225
rect 51699 36191 51707 36225
rect 51657 36167 51707 36191
rect 51993 36225 52043 36249
rect 51993 36191 52001 36225
rect 52035 36191 52043 36225
rect 51993 36167 52043 36191
rect 52329 36225 52379 36249
rect 52329 36191 52337 36225
rect 52371 36191 52379 36225
rect 52329 36167 52379 36191
rect 52665 36225 52715 36249
rect 52665 36191 52673 36225
rect 52707 36191 52715 36225
rect 52665 36167 52715 36191
rect 53001 36225 53051 36249
rect 53001 36191 53009 36225
rect 53043 36191 53051 36225
rect 53001 36167 53051 36191
rect 53337 36225 53387 36249
rect 53337 36191 53345 36225
rect 53379 36191 53387 36225
rect 53337 36167 53387 36191
rect 53673 36225 53723 36249
rect 53673 36191 53681 36225
rect 53715 36191 53723 36225
rect 53673 36167 53723 36191
rect 54009 36225 54059 36249
rect 54009 36191 54017 36225
rect 54051 36191 54059 36225
rect 54009 36167 54059 36191
rect 54345 36225 54395 36249
rect 54345 36191 54353 36225
rect 54387 36191 54395 36225
rect 54345 36167 54395 36191
rect 54681 36225 54731 36249
rect 54681 36191 54689 36225
rect 54723 36191 54731 36225
rect 54681 36167 54731 36191
rect 55017 36225 55067 36249
rect 55017 36191 55025 36225
rect 55059 36191 55067 36225
rect 55017 36167 55067 36191
rect 55353 36225 55403 36249
rect 55353 36191 55361 36225
rect 55395 36191 55403 36225
rect 55353 36167 55403 36191
rect 55689 36225 55739 36249
rect 55689 36191 55697 36225
rect 55731 36191 55739 36225
rect 55689 36167 55739 36191
rect 56025 36225 56075 36249
rect 56025 36191 56033 36225
rect 56067 36191 56075 36225
rect 56025 36167 56075 36191
rect 56361 36225 56411 36249
rect 56361 36191 56369 36225
rect 56403 36191 56411 36225
rect 56361 36167 56411 36191
rect 56697 36225 56747 36249
rect 56697 36191 56705 36225
rect 56739 36191 56747 36225
rect 56697 36167 56747 36191
rect 57033 36225 57083 36249
rect 57033 36191 57041 36225
rect 57075 36191 57083 36225
rect 57033 36167 57083 36191
rect 57369 36225 57419 36249
rect 57369 36191 57377 36225
rect 57411 36191 57419 36225
rect 57369 36167 57419 36191
rect 57705 36225 57755 36249
rect 57705 36191 57713 36225
rect 57747 36191 57755 36225
rect 57705 36167 57755 36191
rect 58041 36225 58091 36249
rect 58041 36191 58049 36225
rect 58083 36191 58091 36225
rect 58041 36167 58091 36191
rect 58377 36225 58427 36249
rect 58377 36191 58385 36225
rect 58419 36191 58427 36225
rect 58377 36167 58427 36191
rect 58713 36225 58763 36249
rect 58713 36191 58721 36225
rect 58755 36191 58763 36225
rect 58713 36167 58763 36191
rect 59049 36225 59099 36249
rect 59049 36191 59057 36225
rect 59091 36191 59099 36225
rect 59049 36167 59099 36191
rect 59385 36225 59435 36249
rect 59385 36191 59393 36225
rect 59427 36191 59435 36225
rect 59385 36167 59435 36191
rect 59721 36225 59771 36249
rect 59721 36191 59729 36225
rect 59763 36191 59771 36225
rect 59721 36167 59771 36191
rect 60057 36225 60107 36249
rect 60057 36191 60065 36225
rect 60099 36191 60107 36225
rect 60057 36167 60107 36191
rect 60393 36225 60443 36249
rect 60393 36191 60401 36225
rect 60435 36191 60443 36225
rect 60393 36167 60443 36191
rect 60729 36225 60779 36249
rect 60729 36191 60737 36225
rect 60771 36191 60779 36225
rect 60729 36167 60779 36191
rect 61065 36225 61115 36249
rect 61065 36191 61073 36225
rect 61107 36191 61115 36225
rect 61065 36167 61115 36191
rect 61401 36225 61451 36249
rect 61401 36191 61409 36225
rect 61443 36191 61451 36225
rect 61401 36167 61451 36191
rect 61737 36225 61787 36249
rect 61737 36191 61745 36225
rect 61779 36191 61787 36225
rect 61737 36167 61787 36191
rect 62073 36225 62123 36249
rect 62073 36191 62081 36225
rect 62115 36191 62123 36225
rect 62073 36167 62123 36191
rect 62409 36225 62459 36249
rect 62409 36191 62417 36225
rect 62451 36191 62459 36225
rect 62409 36167 62459 36191
rect 62745 36225 62795 36249
rect 62745 36191 62753 36225
rect 62787 36191 62795 36225
rect 62745 36167 62795 36191
rect 63081 36225 63131 36249
rect 63081 36191 63089 36225
rect 63123 36191 63131 36225
rect 63081 36167 63131 36191
rect 63417 36225 63467 36249
rect 63417 36191 63425 36225
rect 63459 36191 63467 36225
rect 63417 36167 63467 36191
rect 63753 36225 63803 36249
rect 63753 36191 63761 36225
rect 63795 36191 63803 36225
rect 63753 36167 63803 36191
rect 64089 36225 64139 36249
rect 64089 36191 64097 36225
rect 64131 36191 64139 36225
rect 64089 36167 64139 36191
rect 64425 36225 64475 36249
rect 64425 36191 64433 36225
rect 64467 36191 64475 36225
rect 64425 36167 64475 36191
rect 64761 36225 64811 36249
rect 64761 36191 64769 36225
rect 64803 36191 64811 36225
rect 64761 36167 64811 36191
rect 65097 36225 65147 36249
rect 65097 36191 65105 36225
rect 65139 36191 65147 36225
rect 65097 36167 65147 36191
rect 65433 36225 65483 36249
rect 65433 36191 65441 36225
rect 65475 36191 65483 36225
rect 65433 36167 65483 36191
rect 65769 36225 65819 36249
rect 65769 36191 65777 36225
rect 65811 36191 65819 36225
rect 65769 36167 65819 36191
rect 66105 36225 66155 36249
rect 66105 36191 66113 36225
rect 66147 36191 66155 36225
rect 66105 36167 66155 36191
rect 66441 36225 66491 36249
rect 66441 36191 66449 36225
rect 66483 36191 66491 36225
rect 66441 36167 66491 36191
rect 66777 36225 66827 36249
rect 66777 36191 66785 36225
rect 66819 36191 66827 36225
rect 66777 36167 66827 36191
rect 67113 36225 67163 36249
rect 67113 36191 67121 36225
rect 67155 36191 67163 36225
rect 67113 36167 67163 36191
rect 67449 36225 67499 36249
rect 67449 36191 67457 36225
rect 67491 36191 67499 36225
rect 67449 36167 67499 36191
rect 67785 36225 67835 36249
rect 67785 36191 67793 36225
rect 67827 36191 67835 36225
rect 67785 36167 67835 36191
rect 68121 36225 68171 36249
rect 68121 36191 68129 36225
rect 68163 36191 68171 36225
rect 68121 36167 68171 36191
rect 68457 36225 68507 36249
rect 68457 36191 68465 36225
rect 68499 36191 68507 36225
rect 68457 36167 68507 36191
rect 68793 36225 68843 36249
rect 68793 36191 68801 36225
rect 68835 36191 68843 36225
rect 68793 36167 68843 36191
rect 69129 36225 69179 36249
rect 69129 36191 69137 36225
rect 69171 36191 69179 36225
rect 69129 36167 69179 36191
rect 69465 36225 69515 36249
rect 69465 36191 69473 36225
rect 69507 36191 69515 36225
rect 69465 36167 69515 36191
rect 69801 36225 69851 36249
rect 69801 36191 69809 36225
rect 69843 36191 69851 36225
rect 69801 36167 69851 36191
rect 70137 36225 70187 36249
rect 70137 36191 70145 36225
rect 70179 36191 70187 36225
rect 70137 36167 70187 36191
rect 70473 36225 70523 36249
rect 70473 36191 70481 36225
rect 70515 36191 70523 36225
rect 70473 36167 70523 36191
rect 70809 36225 70859 36249
rect 70809 36191 70817 36225
rect 70851 36191 70859 36225
rect 70809 36167 70859 36191
rect 71145 36225 71195 36249
rect 71145 36191 71153 36225
rect 71187 36191 71195 36225
rect 71145 36167 71195 36191
rect 71481 36225 71531 36249
rect 71481 36191 71489 36225
rect 71523 36191 71531 36225
rect 71481 36167 71531 36191
rect 71817 36225 71867 36249
rect 71817 36191 71825 36225
rect 71859 36191 71867 36225
rect 71817 36167 71867 36191
rect 72153 36225 72203 36249
rect 72153 36191 72161 36225
rect 72195 36191 72203 36225
rect 72153 36167 72203 36191
rect 72489 36225 72539 36249
rect 72489 36191 72497 36225
rect 72531 36191 72539 36225
rect 72489 36167 72539 36191
rect 72825 36225 72875 36249
rect 72825 36191 72833 36225
rect 72867 36191 72875 36225
rect 72825 36167 72875 36191
rect 73161 36225 73211 36249
rect 73161 36191 73169 36225
rect 73203 36191 73211 36225
rect 73161 36167 73211 36191
rect 73497 36225 73547 36249
rect 73497 36191 73505 36225
rect 73539 36191 73547 36225
rect 73497 36167 73547 36191
rect 1593 35853 1643 35877
rect 1593 35819 1601 35853
rect 1635 35819 1643 35853
rect 1593 35795 1643 35819
rect 73941 35853 73991 35877
rect 73941 35819 73949 35853
rect 73983 35819 73991 35853
rect 73941 35795 73991 35819
rect 1593 35517 1643 35541
rect 1593 35483 1601 35517
rect 1635 35483 1643 35517
rect 1593 35459 1643 35483
rect 73941 35517 73991 35541
rect 73941 35483 73949 35517
rect 73983 35483 73991 35517
rect 73941 35459 73991 35483
rect 1593 35181 1643 35205
rect 1593 35147 1601 35181
rect 1635 35147 1643 35181
rect 1593 35123 1643 35147
rect 73941 35181 73991 35205
rect 73941 35147 73949 35181
rect 73983 35147 73991 35181
rect 73941 35123 73991 35147
rect 1593 34845 1643 34869
rect 1593 34811 1601 34845
rect 1635 34811 1643 34845
rect 1593 34787 1643 34811
rect 73941 34845 73991 34869
rect 73941 34811 73949 34845
rect 73983 34811 73991 34845
rect 73941 34787 73991 34811
rect 1593 34509 1643 34533
rect 1593 34475 1601 34509
rect 1635 34475 1643 34509
rect 1593 34451 1643 34475
rect 73941 34509 73991 34533
rect 73941 34475 73949 34509
rect 73983 34475 73991 34509
rect 73941 34451 73991 34475
rect 1593 34173 1643 34197
rect 1593 34139 1601 34173
rect 1635 34139 1643 34173
rect 1593 34115 1643 34139
rect 73941 34173 73991 34197
rect 73941 34139 73949 34173
rect 73983 34139 73991 34173
rect 73941 34115 73991 34139
rect 1593 33837 1643 33861
rect 1593 33803 1601 33837
rect 1635 33803 1643 33837
rect 1593 33779 1643 33803
rect 73941 33837 73991 33861
rect 73941 33803 73949 33837
rect 73983 33803 73991 33837
rect 73941 33779 73991 33803
rect 1593 33501 1643 33525
rect 1593 33467 1601 33501
rect 1635 33467 1643 33501
rect 1593 33443 1643 33467
rect 73941 33501 73991 33525
rect 73941 33467 73949 33501
rect 73983 33467 73991 33501
rect 73941 33443 73991 33467
rect 1593 33165 1643 33189
rect 1593 33131 1601 33165
rect 1635 33131 1643 33165
rect 1593 33107 1643 33131
rect 73941 33165 73991 33189
rect 73941 33131 73949 33165
rect 73983 33131 73991 33165
rect 73941 33107 73991 33131
rect 1593 32829 1643 32853
rect 1593 32795 1601 32829
rect 1635 32795 1643 32829
rect 1593 32771 1643 32795
rect 73941 32829 73991 32853
rect 73941 32795 73949 32829
rect 73983 32795 73991 32829
rect 73941 32771 73991 32795
rect 1593 32493 1643 32517
rect 1593 32459 1601 32493
rect 1635 32459 1643 32493
rect 1593 32435 1643 32459
rect 73941 32493 73991 32517
rect 73941 32459 73949 32493
rect 73983 32459 73991 32493
rect 73941 32435 73991 32459
rect 1593 32157 1643 32181
rect 1593 32123 1601 32157
rect 1635 32123 1643 32157
rect 1593 32099 1643 32123
rect 73941 32157 73991 32181
rect 73941 32123 73949 32157
rect 73983 32123 73991 32157
rect 73941 32099 73991 32123
rect 1593 31821 1643 31845
rect 1593 31787 1601 31821
rect 1635 31787 1643 31821
rect 1593 31763 1643 31787
rect 73941 31821 73991 31845
rect 73941 31787 73949 31821
rect 73983 31787 73991 31821
rect 73941 31763 73991 31787
rect 1593 31485 1643 31509
rect 1593 31451 1601 31485
rect 1635 31451 1643 31485
rect 1593 31427 1643 31451
rect 73941 31485 73991 31509
rect 73941 31451 73949 31485
rect 73983 31451 73991 31485
rect 73941 31427 73991 31451
rect 1593 31149 1643 31173
rect 1593 31115 1601 31149
rect 1635 31115 1643 31149
rect 1593 31091 1643 31115
rect 73941 31149 73991 31173
rect 73941 31115 73949 31149
rect 73983 31115 73991 31149
rect 73941 31091 73991 31115
rect 1593 30813 1643 30837
rect 1593 30779 1601 30813
rect 1635 30779 1643 30813
rect 1593 30755 1643 30779
rect 73941 30813 73991 30837
rect 73941 30779 73949 30813
rect 73983 30779 73991 30813
rect 73941 30755 73991 30779
rect 1593 30477 1643 30501
rect 1593 30443 1601 30477
rect 1635 30443 1643 30477
rect 1593 30419 1643 30443
rect 73941 30477 73991 30501
rect 73941 30443 73949 30477
rect 73983 30443 73991 30477
rect 73941 30419 73991 30443
rect 1593 30141 1643 30165
rect 1593 30107 1601 30141
rect 1635 30107 1643 30141
rect 1593 30083 1643 30107
rect 73941 30141 73991 30165
rect 73941 30107 73949 30141
rect 73983 30107 73991 30141
rect 73941 30083 73991 30107
rect 1593 29805 1643 29829
rect 1593 29771 1601 29805
rect 1635 29771 1643 29805
rect 1593 29747 1643 29771
rect 73941 29805 73991 29829
rect 73941 29771 73949 29805
rect 73983 29771 73991 29805
rect 73941 29747 73991 29771
rect 1593 29469 1643 29493
rect 1593 29435 1601 29469
rect 1635 29435 1643 29469
rect 1593 29411 1643 29435
rect 73941 29469 73991 29493
rect 73941 29435 73949 29469
rect 73983 29435 73991 29469
rect 73941 29411 73991 29435
rect 1593 29133 1643 29157
rect 1593 29099 1601 29133
rect 1635 29099 1643 29133
rect 1593 29075 1643 29099
rect 73941 29133 73991 29157
rect 73941 29099 73949 29133
rect 73983 29099 73991 29133
rect 73941 29075 73991 29099
rect 1593 28797 1643 28821
rect 1593 28763 1601 28797
rect 1635 28763 1643 28797
rect 1593 28739 1643 28763
rect 73941 28797 73991 28821
rect 73941 28763 73949 28797
rect 73983 28763 73991 28797
rect 73941 28739 73991 28763
rect 1593 28461 1643 28485
rect 1593 28427 1601 28461
rect 1635 28427 1643 28461
rect 1593 28403 1643 28427
rect 73941 28461 73991 28485
rect 73941 28427 73949 28461
rect 73983 28427 73991 28461
rect 73941 28403 73991 28427
rect 1593 28125 1643 28149
rect 1593 28091 1601 28125
rect 1635 28091 1643 28125
rect 1593 28067 1643 28091
rect 73941 28125 73991 28149
rect 73941 28091 73949 28125
rect 73983 28091 73991 28125
rect 73941 28067 73991 28091
rect 1593 27789 1643 27813
rect 1593 27755 1601 27789
rect 1635 27755 1643 27789
rect 1593 27731 1643 27755
rect 73941 27789 73991 27813
rect 73941 27755 73949 27789
rect 73983 27755 73991 27789
rect 73941 27731 73991 27755
rect 1593 27453 1643 27477
rect 1593 27419 1601 27453
rect 1635 27419 1643 27453
rect 1593 27395 1643 27419
rect 73941 27453 73991 27477
rect 73941 27419 73949 27453
rect 73983 27419 73991 27453
rect 73941 27395 73991 27419
rect 1593 27117 1643 27141
rect 1593 27083 1601 27117
rect 1635 27083 1643 27117
rect 1593 27059 1643 27083
rect 73941 27117 73991 27141
rect 73941 27083 73949 27117
rect 73983 27083 73991 27117
rect 73941 27059 73991 27083
rect 1593 26781 1643 26805
rect 1593 26747 1601 26781
rect 1635 26747 1643 26781
rect 1593 26723 1643 26747
rect 73941 26781 73991 26805
rect 73941 26747 73949 26781
rect 73983 26747 73991 26781
rect 73941 26723 73991 26747
rect 1593 26445 1643 26469
rect 1593 26411 1601 26445
rect 1635 26411 1643 26445
rect 1593 26387 1643 26411
rect 73941 26445 73991 26469
rect 73941 26411 73949 26445
rect 73983 26411 73991 26445
rect 73941 26387 73991 26411
rect 1593 26109 1643 26133
rect 1593 26075 1601 26109
rect 1635 26075 1643 26109
rect 1593 26051 1643 26075
rect 73941 26109 73991 26133
rect 73941 26075 73949 26109
rect 73983 26075 73991 26109
rect 73941 26051 73991 26075
rect 1593 25773 1643 25797
rect 1593 25739 1601 25773
rect 1635 25739 1643 25773
rect 1593 25715 1643 25739
rect 73941 25773 73991 25797
rect 73941 25739 73949 25773
rect 73983 25739 73991 25773
rect 73941 25715 73991 25739
rect 1593 25437 1643 25461
rect 1593 25403 1601 25437
rect 1635 25403 1643 25437
rect 1593 25379 1643 25403
rect 73941 25437 73991 25461
rect 73941 25403 73949 25437
rect 73983 25403 73991 25437
rect 73941 25379 73991 25403
rect 1593 25101 1643 25125
rect 1593 25067 1601 25101
rect 1635 25067 1643 25101
rect 1593 25043 1643 25067
rect 73941 25101 73991 25125
rect 73941 25067 73949 25101
rect 73983 25067 73991 25101
rect 73941 25043 73991 25067
rect 1593 24765 1643 24789
rect 1593 24731 1601 24765
rect 1635 24731 1643 24765
rect 1593 24707 1643 24731
rect 73941 24765 73991 24789
rect 73941 24731 73949 24765
rect 73983 24731 73991 24765
rect 73941 24707 73991 24731
rect 1593 24429 1643 24453
rect 1593 24395 1601 24429
rect 1635 24395 1643 24429
rect 1593 24371 1643 24395
rect 73941 24429 73991 24453
rect 73941 24395 73949 24429
rect 73983 24395 73991 24429
rect 73941 24371 73991 24395
rect 1593 24093 1643 24117
rect 1593 24059 1601 24093
rect 1635 24059 1643 24093
rect 1593 24035 1643 24059
rect 73941 24093 73991 24117
rect 73941 24059 73949 24093
rect 73983 24059 73991 24093
rect 73941 24035 73991 24059
rect 1593 23757 1643 23781
rect 1593 23723 1601 23757
rect 1635 23723 1643 23757
rect 1593 23699 1643 23723
rect 73941 23757 73991 23781
rect 73941 23723 73949 23757
rect 73983 23723 73991 23757
rect 73941 23699 73991 23723
rect 1593 23421 1643 23445
rect 1593 23387 1601 23421
rect 1635 23387 1643 23421
rect 1593 23363 1643 23387
rect 73941 23421 73991 23445
rect 73941 23387 73949 23421
rect 73983 23387 73991 23421
rect 73941 23363 73991 23387
rect 1593 23085 1643 23109
rect 1593 23051 1601 23085
rect 1635 23051 1643 23085
rect 1593 23027 1643 23051
rect 73941 23085 73991 23109
rect 73941 23051 73949 23085
rect 73983 23051 73991 23085
rect 73941 23027 73991 23051
rect 1593 22749 1643 22773
rect 1593 22715 1601 22749
rect 1635 22715 1643 22749
rect 1593 22691 1643 22715
rect 73941 22749 73991 22773
rect 73941 22715 73949 22749
rect 73983 22715 73991 22749
rect 73941 22691 73991 22715
rect 1593 22413 1643 22437
rect 1593 22379 1601 22413
rect 1635 22379 1643 22413
rect 1593 22355 1643 22379
rect 73941 22413 73991 22437
rect 73941 22379 73949 22413
rect 73983 22379 73991 22413
rect 73941 22355 73991 22379
rect 1593 22077 1643 22101
rect 1593 22043 1601 22077
rect 1635 22043 1643 22077
rect 1593 22019 1643 22043
rect 73941 22077 73991 22101
rect 73941 22043 73949 22077
rect 73983 22043 73991 22077
rect 73941 22019 73991 22043
rect 1593 21741 1643 21765
rect 1593 21707 1601 21741
rect 1635 21707 1643 21741
rect 1593 21683 1643 21707
rect 73941 21741 73991 21765
rect 73941 21707 73949 21741
rect 73983 21707 73991 21741
rect 73941 21683 73991 21707
rect 1593 21405 1643 21429
rect 1593 21371 1601 21405
rect 1635 21371 1643 21405
rect 1593 21347 1643 21371
rect 73941 21405 73991 21429
rect 73941 21371 73949 21405
rect 73983 21371 73991 21405
rect 73941 21347 73991 21371
rect 1593 21069 1643 21093
rect 1593 21035 1601 21069
rect 1635 21035 1643 21069
rect 1593 21011 1643 21035
rect 73941 21069 73991 21093
rect 73941 21035 73949 21069
rect 73983 21035 73991 21069
rect 73941 21011 73991 21035
rect 1593 20733 1643 20757
rect 1593 20699 1601 20733
rect 1635 20699 1643 20733
rect 1593 20675 1643 20699
rect 73941 20733 73991 20757
rect 73941 20699 73949 20733
rect 73983 20699 73991 20733
rect 73941 20675 73991 20699
rect 1593 20397 1643 20421
rect 1593 20363 1601 20397
rect 1635 20363 1643 20397
rect 1593 20339 1643 20363
rect 73941 20397 73991 20421
rect 73941 20363 73949 20397
rect 73983 20363 73991 20397
rect 73941 20339 73991 20363
rect 1593 20061 1643 20085
rect 1593 20027 1601 20061
rect 1635 20027 1643 20061
rect 1593 20003 1643 20027
rect 73941 20061 73991 20085
rect 73941 20027 73949 20061
rect 73983 20027 73991 20061
rect 73941 20003 73991 20027
rect 1593 19725 1643 19749
rect 1593 19691 1601 19725
rect 1635 19691 1643 19725
rect 1593 19667 1643 19691
rect 73941 19725 73991 19749
rect 73941 19691 73949 19725
rect 73983 19691 73991 19725
rect 73941 19667 73991 19691
rect 1593 19389 1643 19413
rect 1593 19355 1601 19389
rect 1635 19355 1643 19389
rect 1593 19331 1643 19355
rect 73941 19389 73991 19413
rect 73941 19355 73949 19389
rect 73983 19355 73991 19389
rect 73941 19331 73991 19355
rect 1593 19053 1643 19077
rect 1593 19019 1601 19053
rect 1635 19019 1643 19053
rect 1593 18995 1643 19019
rect 73941 19053 73991 19077
rect 73941 19019 73949 19053
rect 73983 19019 73991 19053
rect 73941 18995 73991 19019
rect 1593 18717 1643 18741
rect 1593 18683 1601 18717
rect 1635 18683 1643 18717
rect 1593 18659 1643 18683
rect 73941 18717 73991 18741
rect 73941 18683 73949 18717
rect 73983 18683 73991 18717
rect 73941 18659 73991 18683
rect 1593 18381 1643 18405
rect 1593 18347 1601 18381
rect 1635 18347 1643 18381
rect 1593 18323 1643 18347
rect 73941 18381 73991 18405
rect 73941 18347 73949 18381
rect 73983 18347 73991 18381
rect 73941 18323 73991 18347
rect 1593 18045 1643 18069
rect 1593 18011 1601 18045
rect 1635 18011 1643 18045
rect 1593 17987 1643 18011
rect 73941 18045 73991 18069
rect 73941 18011 73949 18045
rect 73983 18011 73991 18045
rect 73941 17987 73991 18011
rect 1593 17709 1643 17733
rect 1593 17675 1601 17709
rect 1635 17675 1643 17709
rect 1593 17651 1643 17675
rect 73941 17709 73991 17733
rect 73941 17675 73949 17709
rect 73983 17675 73991 17709
rect 73941 17651 73991 17675
rect 1593 17373 1643 17397
rect 1593 17339 1601 17373
rect 1635 17339 1643 17373
rect 1593 17315 1643 17339
rect 73941 17373 73991 17397
rect 73941 17339 73949 17373
rect 73983 17339 73991 17373
rect 73941 17315 73991 17339
rect 1593 17037 1643 17061
rect 1593 17003 1601 17037
rect 1635 17003 1643 17037
rect 1593 16979 1643 17003
rect 73941 17037 73991 17061
rect 73941 17003 73949 17037
rect 73983 17003 73991 17037
rect 73941 16979 73991 17003
rect 1593 16701 1643 16725
rect 1593 16667 1601 16701
rect 1635 16667 1643 16701
rect 1593 16643 1643 16667
rect 73941 16701 73991 16725
rect 73941 16667 73949 16701
rect 73983 16667 73991 16701
rect 73941 16643 73991 16667
rect 1593 16365 1643 16389
rect 1593 16331 1601 16365
rect 1635 16331 1643 16365
rect 1593 16307 1643 16331
rect 73941 16365 73991 16389
rect 73941 16331 73949 16365
rect 73983 16331 73991 16365
rect 73941 16307 73991 16331
rect 1593 16029 1643 16053
rect 1593 15995 1601 16029
rect 1635 15995 1643 16029
rect 1593 15971 1643 15995
rect 73941 16029 73991 16053
rect 73941 15995 73949 16029
rect 73983 15995 73991 16029
rect 73941 15971 73991 15995
rect 1593 15693 1643 15717
rect 1593 15659 1601 15693
rect 1635 15659 1643 15693
rect 1593 15635 1643 15659
rect 73941 15693 73991 15717
rect 73941 15659 73949 15693
rect 73983 15659 73991 15693
rect 73941 15635 73991 15659
rect 1593 15357 1643 15381
rect 1593 15323 1601 15357
rect 1635 15323 1643 15357
rect 1593 15299 1643 15323
rect 73941 15357 73991 15381
rect 73941 15323 73949 15357
rect 73983 15323 73991 15357
rect 73941 15299 73991 15323
rect 1593 15021 1643 15045
rect 1593 14987 1601 15021
rect 1635 14987 1643 15021
rect 1593 14963 1643 14987
rect 73941 15021 73991 15045
rect 73941 14987 73949 15021
rect 73983 14987 73991 15021
rect 73941 14963 73991 14987
rect 1593 14685 1643 14709
rect 1593 14651 1601 14685
rect 1635 14651 1643 14685
rect 1593 14627 1643 14651
rect 73941 14685 73991 14709
rect 73941 14651 73949 14685
rect 73983 14651 73991 14685
rect 73941 14627 73991 14651
rect 1593 14349 1643 14373
rect 1593 14315 1601 14349
rect 1635 14315 1643 14349
rect 1593 14291 1643 14315
rect 73941 14349 73991 14373
rect 73941 14315 73949 14349
rect 73983 14315 73991 14349
rect 73941 14291 73991 14315
rect 1593 14013 1643 14037
rect 1593 13979 1601 14013
rect 1635 13979 1643 14013
rect 1593 13955 1643 13979
rect 73941 14013 73991 14037
rect 73941 13979 73949 14013
rect 73983 13979 73991 14013
rect 73941 13955 73991 13979
rect 1593 13677 1643 13701
rect 1593 13643 1601 13677
rect 1635 13643 1643 13677
rect 1593 13619 1643 13643
rect 73941 13677 73991 13701
rect 73941 13643 73949 13677
rect 73983 13643 73991 13677
rect 73941 13619 73991 13643
rect 1593 13341 1643 13365
rect 1593 13307 1601 13341
rect 1635 13307 1643 13341
rect 1593 13283 1643 13307
rect 73941 13341 73991 13365
rect 73941 13307 73949 13341
rect 73983 13307 73991 13341
rect 73941 13283 73991 13307
rect 1593 13005 1643 13029
rect 1593 12971 1601 13005
rect 1635 12971 1643 13005
rect 1593 12947 1643 12971
rect 73941 13005 73991 13029
rect 73941 12971 73949 13005
rect 73983 12971 73991 13005
rect 73941 12947 73991 12971
rect 1593 12669 1643 12693
rect 1593 12635 1601 12669
rect 1635 12635 1643 12669
rect 1593 12611 1643 12635
rect 73941 12669 73991 12693
rect 73941 12635 73949 12669
rect 73983 12635 73991 12669
rect 73941 12611 73991 12635
rect 1593 12333 1643 12357
rect 1593 12299 1601 12333
rect 1635 12299 1643 12333
rect 1593 12275 1643 12299
rect 73941 12333 73991 12357
rect 73941 12299 73949 12333
rect 73983 12299 73991 12333
rect 73941 12275 73991 12299
rect 1593 11997 1643 12021
rect 1593 11963 1601 11997
rect 1635 11963 1643 11997
rect 1593 11939 1643 11963
rect 73941 11997 73991 12021
rect 73941 11963 73949 11997
rect 73983 11963 73991 11997
rect 73941 11939 73991 11963
rect 1593 11661 1643 11685
rect 1593 11627 1601 11661
rect 1635 11627 1643 11661
rect 1593 11603 1643 11627
rect 73941 11661 73991 11685
rect 73941 11627 73949 11661
rect 73983 11627 73991 11661
rect 73941 11603 73991 11627
rect 1593 11325 1643 11349
rect 1593 11291 1601 11325
rect 1635 11291 1643 11325
rect 1593 11267 1643 11291
rect 73941 11325 73991 11349
rect 73941 11291 73949 11325
rect 73983 11291 73991 11325
rect 73941 11267 73991 11291
rect 1593 10989 1643 11013
rect 1593 10955 1601 10989
rect 1635 10955 1643 10989
rect 1593 10931 1643 10955
rect 73941 10989 73991 11013
rect 73941 10955 73949 10989
rect 73983 10955 73991 10989
rect 73941 10931 73991 10955
rect 1593 10653 1643 10677
rect 1593 10619 1601 10653
rect 1635 10619 1643 10653
rect 1593 10595 1643 10619
rect 73941 10653 73991 10677
rect 73941 10619 73949 10653
rect 73983 10619 73991 10653
rect 73941 10595 73991 10619
rect 1593 10317 1643 10341
rect 1593 10283 1601 10317
rect 1635 10283 1643 10317
rect 1593 10259 1643 10283
rect 73941 10317 73991 10341
rect 73941 10283 73949 10317
rect 73983 10283 73991 10317
rect 73941 10259 73991 10283
rect 1593 9981 1643 10005
rect 1593 9947 1601 9981
rect 1635 9947 1643 9981
rect 1593 9923 1643 9947
rect 73941 9981 73991 10005
rect 73941 9947 73949 9981
rect 73983 9947 73991 9981
rect 73941 9923 73991 9947
rect 1593 9645 1643 9669
rect 1593 9611 1601 9645
rect 1635 9611 1643 9645
rect 1593 9587 1643 9611
rect 73941 9645 73991 9669
rect 73941 9611 73949 9645
rect 73983 9611 73991 9645
rect 73941 9587 73991 9611
rect 1593 9309 1643 9333
rect 1593 9275 1601 9309
rect 1635 9275 1643 9309
rect 1593 9251 1643 9275
rect 73941 9309 73991 9333
rect 73941 9275 73949 9309
rect 73983 9275 73991 9309
rect 73941 9251 73991 9275
rect 1593 8973 1643 8997
rect 1593 8939 1601 8973
rect 1635 8939 1643 8973
rect 1593 8915 1643 8939
rect 73941 8973 73991 8997
rect 73941 8939 73949 8973
rect 73983 8939 73991 8973
rect 73941 8915 73991 8939
rect 1593 8637 1643 8661
rect 1593 8603 1601 8637
rect 1635 8603 1643 8637
rect 1593 8579 1643 8603
rect 73941 8637 73991 8661
rect 73941 8603 73949 8637
rect 73983 8603 73991 8637
rect 73941 8579 73991 8603
rect 1593 8301 1643 8325
rect 1593 8267 1601 8301
rect 1635 8267 1643 8301
rect 1593 8243 1643 8267
rect 73941 8301 73991 8325
rect 73941 8267 73949 8301
rect 73983 8267 73991 8301
rect 73941 8243 73991 8267
rect 1593 7965 1643 7989
rect 1593 7931 1601 7965
rect 1635 7931 1643 7965
rect 1593 7907 1643 7931
rect 73941 7965 73991 7989
rect 73941 7931 73949 7965
rect 73983 7931 73991 7965
rect 73941 7907 73991 7931
rect 1593 7629 1643 7653
rect 1593 7595 1601 7629
rect 1635 7595 1643 7629
rect 1593 7571 1643 7595
rect 73941 7629 73991 7653
rect 73941 7595 73949 7629
rect 73983 7595 73991 7629
rect 73941 7571 73991 7595
rect 1593 7293 1643 7317
rect 1593 7259 1601 7293
rect 1635 7259 1643 7293
rect 1593 7235 1643 7259
rect 73941 7293 73991 7317
rect 73941 7259 73949 7293
rect 73983 7259 73991 7293
rect 73941 7235 73991 7259
rect 1593 6957 1643 6981
rect 1593 6923 1601 6957
rect 1635 6923 1643 6957
rect 1593 6899 1643 6923
rect 73941 6957 73991 6981
rect 73941 6923 73949 6957
rect 73983 6923 73991 6957
rect 73941 6899 73991 6923
rect 1593 6621 1643 6645
rect 1593 6587 1601 6621
rect 1635 6587 1643 6621
rect 1593 6563 1643 6587
rect 73941 6621 73991 6645
rect 73941 6587 73949 6621
rect 73983 6587 73991 6621
rect 73941 6563 73991 6587
rect 1593 6285 1643 6309
rect 1593 6251 1601 6285
rect 1635 6251 1643 6285
rect 1593 6227 1643 6251
rect 73941 6285 73991 6309
rect 73941 6251 73949 6285
rect 73983 6251 73991 6285
rect 73941 6227 73991 6251
rect 1593 5949 1643 5973
rect 1593 5915 1601 5949
rect 1635 5915 1643 5949
rect 1593 5891 1643 5915
rect 73941 5949 73991 5973
rect 73941 5915 73949 5949
rect 73983 5915 73991 5949
rect 73941 5891 73991 5915
rect 1593 5613 1643 5637
rect 1593 5579 1601 5613
rect 1635 5579 1643 5613
rect 1593 5555 1643 5579
rect 73941 5613 73991 5637
rect 73941 5579 73949 5613
rect 73983 5579 73991 5613
rect 73941 5555 73991 5579
rect 1593 5277 1643 5301
rect 1593 5243 1601 5277
rect 1635 5243 1643 5277
rect 1593 5219 1643 5243
rect 73941 5277 73991 5301
rect 73941 5243 73949 5277
rect 73983 5243 73991 5277
rect 73941 5219 73991 5243
rect 1593 4941 1643 4965
rect 1593 4907 1601 4941
rect 1635 4907 1643 4941
rect 1593 4883 1643 4907
rect 73941 4941 73991 4965
rect 73941 4907 73949 4941
rect 73983 4907 73991 4941
rect 73941 4883 73991 4907
rect 1593 4605 1643 4629
rect 1593 4571 1601 4605
rect 1635 4571 1643 4605
rect 1593 4547 1643 4571
rect 73941 4605 73991 4629
rect 73941 4571 73949 4605
rect 73983 4571 73991 4605
rect 73941 4547 73991 4571
rect 1593 4269 1643 4293
rect 1593 4235 1601 4269
rect 1635 4235 1643 4269
rect 1593 4211 1643 4235
rect 73941 4269 73991 4293
rect 73941 4235 73949 4269
rect 73983 4235 73991 4269
rect 73941 4211 73991 4235
rect 1593 3933 1643 3957
rect 1593 3899 1601 3933
rect 1635 3899 1643 3933
rect 1593 3875 1643 3899
rect 73941 3933 73991 3957
rect 73941 3899 73949 3933
rect 73983 3899 73991 3933
rect 73941 3875 73991 3899
rect 1593 3597 1643 3621
rect 1593 3563 1601 3597
rect 1635 3563 1643 3597
rect 1593 3539 1643 3563
rect 73941 3597 73991 3621
rect 73941 3563 73949 3597
rect 73983 3563 73991 3597
rect 73941 3539 73991 3563
rect 1593 3261 1643 3285
rect 1593 3227 1601 3261
rect 1635 3227 1643 3261
rect 1593 3203 1643 3227
rect 73941 3261 73991 3285
rect 73941 3227 73949 3261
rect 73983 3227 73991 3261
rect 73941 3203 73991 3227
rect 1593 2925 1643 2949
rect 1593 2891 1601 2925
rect 1635 2891 1643 2925
rect 1593 2867 1643 2891
rect 73941 2925 73991 2949
rect 73941 2891 73949 2925
rect 73983 2891 73991 2925
rect 73941 2867 73991 2891
rect 1593 2589 1643 2613
rect 1593 2555 1601 2589
rect 1635 2555 1643 2589
rect 1593 2531 1643 2555
rect 73941 2589 73991 2613
rect 73941 2555 73949 2589
rect 73983 2555 73991 2589
rect 73941 2531 73991 2555
rect 1593 2253 1643 2277
rect 1593 2219 1601 2253
rect 1635 2219 1643 2253
rect 1593 2195 1643 2219
rect 73941 2253 73991 2277
rect 73941 2219 73949 2253
rect 73983 2219 73991 2253
rect 73941 2195 73991 2219
rect 1593 1917 1643 1941
rect 1593 1883 1601 1917
rect 1635 1883 1643 1917
rect 1593 1859 1643 1883
rect 73941 1917 73991 1941
rect 73941 1883 73949 1917
rect 73983 1883 73991 1917
rect 73941 1859 73991 1883
rect 1929 1581 1979 1605
rect 1929 1547 1937 1581
rect 1971 1547 1979 1581
rect 1929 1523 1979 1547
rect 2265 1581 2315 1605
rect 2265 1547 2273 1581
rect 2307 1547 2315 1581
rect 2265 1523 2315 1547
rect 2601 1581 2651 1605
rect 2601 1547 2609 1581
rect 2643 1547 2651 1581
rect 2601 1523 2651 1547
rect 2937 1581 2987 1605
rect 2937 1547 2945 1581
rect 2979 1547 2987 1581
rect 2937 1523 2987 1547
rect 3273 1581 3323 1605
rect 3273 1547 3281 1581
rect 3315 1547 3323 1581
rect 3273 1523 3323 1547
rect 3609 1581 3659 1605
rect 3609 1547 3617 1581
rect 3651 1547 3659 1581
rect 3609 1523 3659 1547
rect 3945 1581 3995 1605
rect 3945 1547 3953 1581
rect 3987 1547 3995 1581
rect 3945 1523 3995 1547
rect 4281 1581 4331 1605
rect 4281 1547 4289 1581
rect 4323 1547 4331 1581
rect 4281 1523 4331 1547
rect 4617 1581 4667 1605
rect 4617 1547 4625 1581
rect 4659 1547 4667 1581
rect 4617 1523 4667 1547
rect 4953 1581 5003 1605
rect 4953 1547 4961 1581
rect 4995 1547 5003 1581
rect 4953 1523 5003 1547
rect 5289 1581 5339 1605
rect 5289 1547 5297 1581
rect 5331 1547 5339 1581
rect 5289 1523 5339 1547
rect 5625 1581 5675 1605
rect 5625 1547 5633 1581
rect 5667 1547 5675 1581
rect 5625 1523 5675 1547
rect 5961 1581 6011 1605
rect 5961 1547 5969 1581
rect 6003 1547 6011 1581
rect 5961 1523 6011 1547
rect 6297 1581 6347 1605
rect 6297 1547 6305 1581
rect 6339 1547 6347 1581
rect 6297 1523 6347 1547
rect 6633 1581 6683 1605
rect 6633 1547 6641 1581
rect 6675 1547 6683 1581
rect 6633 1523 6683 1547
rect 6969 1581 7019 1605
rect 6969 1547 6977 1581
rect 7011 1547 7019 1581
rect 6969 1523 7019 1547
rect 7305 1581 7355 1605
rect 7305 1547 7313 1581
rect 7347 1547 7355 1581
rect 7305 1523 7355 1547
rect 7641 1581 7691 1605
rect 7641 1547 7649 1581
rect 7683 1547 7691 1581
rect 7641 1523 7691 1547
rect 7977 1581 8027 1605
rect 7977 1547 7985 1581
rect 8019 1547 8027 1581
rect 7977 1523 8027 1547
rect 8313 1581 8363 1605
rect 8313 1547 8321 1581
rect 8355 1547 8363 1581
rect 8313 1523 8363 1547
rect 8649 1581 8699 1605
rect 8649 1547 8657 1581
rect 8691 1547 8699 1581
rect 8649 1523 8699 1547
rect 8985 1581 9035 1605
rect 8985 1547 8993 1581
rect 9027 1547 9035 1581
rect 8985 1523 9035 1547
rect 9321 1581 9371 1605
rect 9321 1547 9329 1581
rect 9363 1547 9371 1581
rect 9321 1523 9371 1547
rect 9657 1581 9707 1605
rect 9657 1547 9665 1581
rect 9699 1547 9707 1581
rect 9657 1523 9707 1547
rect 9993 1581 10043 1605
rect 9993 1547 10001 1581
rect 10035 1547 10043 1581
rect 9993 1523 10043 1547
rect 10329 1581 10379 1605
rect 10329 1547 10337 1581
rect 10371 1547 10379 1581
rect 10329 1523 10379 1547
rect 10665 1581 10715 1605
rect 10665 1547 10673 1581
rect 10707 1547 10715 1581
rect 10665 1523 10715 1547
rect 11001 1581 11051 1605
rect 11001 1547 11009 1581
rect 11043 1547 11051 1581
rect 11001 1523 11051 1547
rect 11337 1581 11387 1605
rect 11337 1547 11345 1581
rect 11379 1547 11387 1581
rect 11337 1523 11387 1547
rect 11673 1581 11723 1605
rect 11673 1547 11681 1581
rect 11715 1547 11723 1581
rect 11673 1523 11723 1547
rect 12009 1581 12059 1605
rect 12009 1547 12017 1581
rect 12051 1547 12059 1581
rect 12009 1523 12059 1547
rect 12345 1581 12395 1605
rect 12345 1547 12353 1581
rect 12387 1547 12395 1581
rect 12345 1523 12395 1547
rect 12681 1581 12731 1605
rect 12681 1547 12689 1581
rect 12723 1547 12731 1581
rect 12681 1523 12731 1547
rect 13017 1581 13067 1605
rect 13017 1547 13025 1581
rect 13059 1547 13067 1581
rect 13017 1523 13067 1547
rect 13353 1581 13403 1605
rect 13353 1547 13361 1581
rect 13395 1547 13403 1581
rect 13353 1523 13403 1547
rect 13689 1581 13739 1605
rect 13689 1547 13697 1581
rect 13731 1547 13739 1581
rect 13689 1523 13739 1547
rect 14025 1581 14075 1605
rect 14025 1547 14033 1581
rect 14067 1547 14075 1581
rect 14025 1523 14075 1547
rect 14361 1581 14411 1605
rect 14361 1547 14369 1581
rect 14403 1547 14411 1581
rect 14361 1523 14411 1547
rect 14697 1581 14747 1605
rect 14697 1547 14705 1581
rect 14739 1547 14747 1581
rect 14697 1523 14747 1547
rect 15033 1581 15083 1605
rect 15033 1547 15041 1581
rect 15075 1547 15083 1581
rect 15033 1523 15083 1547
rect 15369 1581 15419 1605
rect 15369 1547 15377 1581
rect 15411 1547 15419 1581
rect 15369 1523 15419 1547
rect 15705 1581 15755 1605
rect 15705 1547 15713 1581
rect 15747 1547 15755 1581
rect 15705 1523 15755 1547
rect 16041 1581 16091 1605
rect 16041 1547 16049 1581
rect 16083 1547 16091 1581
rect 16041 1523 16091 1547
rect 16377 1581 16427 1605
rect 16377 1547 16385 1581
rect 16419 1547 16427 1581
rect 16377 1523 16427 1547
rect 16713 1581 16763 1605
rect 16713 1547 16721 1581
rect 16755 1547 16763 1581
rect 16713 1523 16763 1547
rect 17049 1581 17099 1605
rect 17049 1547 17057 1581
rect 17091 1547 17099 1581
rect 17049 1523 17099 1547
rect 17385 1581 17435 1605
rect 17385 1547 17393 1581
rect 17427 1547 17435 1581
rect 17385 1523 17435 1547
rect 17721 1581 17771 1605
rect 17721 1547 17729 1581
rect 17763 1547 17771 1581
rect 17721 1523 17771 1547
rect 18057 1581 18107 1605
rect 18057 1547 18065 1581
rect 18099 1547 18107 1581
rect 18057 1523 18107 1547
rect 18393 1581 18443 1605
rect 18393 1547 18401 1581
rect 18435 1547 18443 1581
rect 18393 1523 18443 1547
rect 18729 1581 18779 1605
rect 18729 1547 18737 1581
rect 18771 1547 18779 1581
rect 18729 1523 18779 1547
rect 19065 1581 19115 1605
rect 19065 1547 19073 1581
rect 19107 1547 19115 1581
rect 19065 1523 19115 1547
rect 19401 1581 19451 1605
rect 19401 1547 19409 1581
rect 19443 1547 19451 1581
rect 19401 1523 19451 1547
rect 19737 1581 19787 1605
rect 19737 1547 19745 1581
rect 19779 1547 19787 1581
rect 19737 1523 19787 1547
rect 20073 1581 20123 1605
rect 20073 1547 20081 1581
rect 20115 1547 20123 1581
rect 20073 1523 20123 1547
rect 20409 1581 20459 1605
rect 20409 1547 20417 1581
rect 20451 1547 20459 1581
rect 20409 1523 20459 1547
rect 20745 1581 20795 1605
rect 20745 1547 20753 1581
rect 20787 1547 20795 1581
rect 20745 1523 20795 1547
rect 21081 1581 21131 1605
rect 21081 1547 21089 1581
rect 21123 1547 21131 1581
rect 21081 1523 21131 1547
rect 21417 1581 21467 1605
rect 21417 1547 21425 1581
rect 21459 1547 21467 1581
rect 21417 1523 21467 1547
rect 21753 1581 21803 1605
rect 21753 1547 21761 1581
rect 21795 1547 21803 1581
rect 21753 1523 21803 1547
rect 22089 1581 22139 1605
rect 22089 1547 22097 1581
rect 22131 1547 22139 1581
rect 22089 1523 22139 1547
rect 22425 1581 22475 1605
rect 22425 1547 22433 1581
rect 22467 1547 22475 1581
rect 22425 1523 22475 1547
rect 22761 1581 22811 1605
rect 22761 1547 22769 1581
rect 22803 1547 22811 1581
rect 22761 1523 22811 1547
rect 23097 1581 23147 1605
rect 23097 1547 23105 1581
rect 23139 1547 23147 1581
rect 23097 1523 23147 1547
rect 23433 1581 23483 1605
rect 23433 1547 23441 1581
rect 23475 1547 23483 1581
rect 23433 1523 23483 1547
rect 23769 1581 23819 1605
rect 23769 1547 23777 1581
rect 23811 1547 23819 1581
rect 23769 1523 23819 1547
rect 24105 1581 24155 1605
rect 24105 1547 24113 1581
rect 24147 1547 24155 1581
rect 24105 1523 24155 1547
rect 24441 1581 24491 1605
rect 24441 1547 24449 1581
rect 24483 1547 24491 1581
rect 24441 1523 24491 1547
rect 24777 1581 24827 1605
rect 24777 1547 24785 1581
rect 24819 1547 24827 1581
rect 24777 1523 24827 1547
rect 25113 1581 25163 1605
rect 25113 1547 25121 1581
rect 25155 1547 25163 1581
rect 25113 1523 25163 1547
rect 25449 1581 25499 1605
rect 25449 1547 25457 1581
rect 25491 1547 25499 1581
rect 25449 1523 25499 1547
rect 25785 1581 25835 1605
rect 25785 1547 25793 1581
rect 25827 1547 25835 1581
rect 25785 1523 25835 1547
rect 26121 1581 26171 1605
rect 26121 1547 26129 1581
rect 26163 1547 26171 1581
rect 26121 1523 26171 1547
rect 26457 1581 26507 1605
rect 26457 1547 26465 1581
rect 26499 1547 26507 1581
rect 26457 1523 26507 1547
rect 26793 1581 26843 1605
rect 26793 1547 26801 1581
rect 26835 1547 26843 1581
rect 26793 1523 26843 1547
rect 27129 1581 27179 1605
rect 27129 1547 27137 1581
rect 27171 1547 27179 1581
rect 27129 1523 27179 1547
rect 27465 1581 27515 1605
rect 27465 1547 27473 1581
rect 27507 1547 27515 1581
rect 27465 1523 27515 1547
rect 27801 1581 27851 1605
rect 27801 1547 27809 1581
rect 27843 1547 27851 1581
rect 27801 1523 27851 1547
rect 28137 1581 28187 1605
rect 28137 1547 28145 1581
rect 28179 1547 28187 1581
rect 28137 1523 28187 1547
rect 28473 1581 28523 1605
rect 28473 1547 28481 1581
rect 28515 1547 28523 1581
rect 28473 1523 28523 1547
rect 28809 1581 28859 1605
rect 28809 1547 28817 1581
rect 28851 1547 28859 1581
rect 28809 1523 28859 1547
rect 29145 1581 29195 1605
rect 29145 1547 29153 1581
rect 29187 1547 29195 1581
rect 29145 1523 29195 1547
rect 29481 1581 29531 1605
rect 29481 1547 29489 1581
rect 29523 1547 29531 1581
rect 29481 1523 29531 1547
rect 29817 1581 29867 1605
rect 29817 1547 29825 1581
rect 29859 1547 29867 1581
rect 29817 1523 29867 1547
rect 30153 1581 30203 1605
rect 30153 1547 30161 1581
rect 30195 1547 30203 1581
rect 30153 1523 30203 1547
rect 30489 1581 30539 1605
rect 30489 1547 30497 1581
rect 30531 1547 30539 1581
rect 30489 1523 30539 1547
rect 30825 1581 30875 1605
rect 30825 1547 30833 1581
rect 30867 1547 30875 1581
rect 30825 1523 30875 1547
rect 31161 1581 31211 1605
rect 31161 1547 31169 1581
rect 31203 1547 31211 1581
rect 31161 1523 31211 1547
rect 31497 1581 31547 1605
rect 31497 1547 31505 1581
rect 31539 1547 31547 1581
rect 31497 1523 31547 1547
rect 31833 1581 31883 1605
rect 31833 1547 31841 1581
rect 31875 1547 31883 1581
rect 31833 1523 31883 1547
rect 32169 1581 32219 1605
rect 32169 1547 32177 1581
rect 32211 1547 32219 1581
rect 32169 1523 32219 1547
rect 32505 1581 32555 1605
rect 32505 1547 32513 1581
rect 32547 1547 32555 1581
rect 32505 1523 32555 1547
rect 32841 1581 32891 1605
rect 32841 1547 32849 1581
rect 32883 1547 32891 1581
rect 32841 1523 32891 1547
rect 33177 1581 33227 1605
rect 33177 1547 33185 1581
rect 33219 1547 33227 1581
rect 33177 1523 33227 1547
rect 33513 1581 33563 1605
rect 33513 1547 33521 1581
rect 33555 1547 33563 1581
rect 33513 1523 33563 1547
rect 33849 1581 33899 1605
rect 33849 1547 33857 1581
rect 33891 1547 33899 1581
rect 33849 1523 33899 1547
rect 34185 1581 34235 1605
rect 34185 1547 34193 1581
rect 34227 1547 34235 1581
rect 34185 1523 34235 1547
rect 34521 1581 34571 1605
rect 34521 1547 34529 1581
rect 34563 1547 34571 1581
rect 34521 1523 34571 1547
rect 34857 1581 34907 1605
rect 34857 1547 34865 1581
rect 34899 1547 34907 1581
rect 34857 1523 34907 1547
rect 35193 1581 35243 1605
rect 35193 1547 35201 1581
rect 35235 1547 35243 1581
rect 35193 1523 35243 1547
rect 35529 1581 35579 1605
rect 35529 1547 35537 1581
rect 35571 1547 35579 1581
rect 35529 1523 35579 1547
rect 35865 1581 35915 1605
rect 35865 1547 35873 1581
rect 35907 1547 35915 1581
rect 35865 1523 35915 1547
rect 36201 1581 36251 1605
rect 36201 1547 36209 1581
rect 36243 1547 36251 1581
rect 36201 1523 36251 1547
rect 36537 1581 36587 1605
rect 36537 1547 36545 1581
rect 36579 1547 36587 1581
rect 36537 1523 36587 1547
rect 36873 1581 36923 1605
rect 36873 1547 36881 1581
rect 36915 1547 36923 1581
rect 36873 1523 36923 1547
rect 37209 1581 37259 1605
rect 37209 1547 37217 1581
rect 37251 1547 37259 1581
rect 37209 1523 37259 1547
rect 37545 1581 37595 1605
rect 37545 1547 37553 1581
rect 37587 1547 37595 1581
rect 37545 1523 37595 1547
rect 37881 1581 37931 1605
rect 37881 1547 37889 1581
rect 37923 1547 37931 1581
rect 37881 1523 37931 1547
rect 38217 1581 38267 1605
rect 38217 1547 38225 1581
rect 38259 1547 38267 1581
rect 38217 1523 38267 1547
rect 38553 1581 38603 1605
rect 38553 1547 38561 1581
rect 38595 1547 38603 1581
rect 38553 1523 38603 1547
rect 38889 1581 38939 1605
rect 38889 1547 38897 1581
rect 38931 1547 38939 1581
rect 38889 1523 38939 1547
rect 39225 1581 39275 1605
rect 39225 1547 39233 1581
rect 39267 1547 39275 1581
rect 39225 1523 39275 1547
rect 39561 1581 39611 1605
rect 39561 1547 39569 1581
rect 39603 1547 39611 1581
rect 39561 1523 39611 1547
rect 39897 1581 39947 1605
rect 39897 1547 39905 1581
rect 39939 1547 39947 1581
rect 39897 1523 39947 1547
rect 40233 1581 40283 1605
rect 40233 1547 40241 1581
rect 40275 1547 40283 1581
rect 40233 1523 40283 1547
rect 40569 1581 40619 1605
rect 40569 1547 40577 1581
rect 40611 1547 40619 1581
rect 40569 1523 40619 1547
rect 40905 1581 40955 1605
rect 40905 1547 40913 1581
rect 40947 1547 40955 1581
rect 40905 1523 40955 1547
rect 41241 1581 41291 1605
rect 41241 1547 41249 1581
rect 41283 1547 41291 1581
rect 41241 1523 41291 1547
rect 41577 1581 41627 1605
rect 41577 1547 41585 1581
rect 41619 1547 41627 1581
rect 41577 1523 41627 1547
rect 41913 1581 41963 1605
rect 41913 1547 41921 1581
rect 41955 1547 41963 1581
rect 41913 1523 41963 1547
rect 42249 1581 42299 1605
rect 42249 1547 42257 1581
rect 42291 1547 42299 1581
rect 42249 1523 42299 1547
rect 42585 1581 42635 1605
rect 42585 1547 42593 1581
rect 42627 1547 42635 1581
rect 42585 1523 42635 1547
rect 42921 1581 42971 1605
rect 42921 1547 42929 1581
rect 42963 1547 42971 1581
rect 42921 1523 42971 1547
rect 43257 1581 43307 1605
rect 43257 1547 43265 1581
rect 43299 1547 43307 1581
rect 43257 1523 43307 1547
rect 43593 1581 43643 1605
rect 43593 1547 43601 1581
rect 43635 1547 43643 1581
rect 43593 1523 43643 1547
rect 43929 1581 43979 1605
rect 43929 1547 43937 1581
rect 43971 1547 43979 1581
rect 43929 1523 43979 1547
rect 44265 1581 44315 1605
rect 44265 1547 44273 1581
rect 44307 1547 44315 1581
rect 44265 1523 44315 1547
rect 44601 1581 44651 1605
rect 44601 1547 44609 1581
rect 44643 1547 44651 1581
rect 44601 1523 44651 1547
rect 44937 1581 44987 1605
rect 44937 1547 44945 1581
rect 44979 1547 44987 1581
rect 44937 1523 44987 1547
rect 45273 1581 45323 1605
rect 45273 1547 45281 1581
rect 45315 1547 45323 1581
rect 45273 1523 45323 1547
rect 45609 1581 45659 1605
rect 45609 1547 45617 1581
rect 45651 1547 45659 1581
rect 45609 1523 45659 1547
rect 45945 1581 45995 1605
rect 45945 1547 45953 1581
rect 45987 1547 45995 1581
rect 45945 1523 45995 1547
rect 46281 1581 46331 1605
rect 46281 1547 46289 1581
rect 46323 1547 46331 1581
rect 46281 1523 46331 1547
rect 46617 1581 46667 1605
rect 46617 1547 46625 1581
rect 46659 1547 46667 1581
rect 46617 1523 46667 1547
rect 46953 1581 47003 1605
rect 46953 1547 46961 1581
rect 46995 1547 47003 1581
rect 46953 1523 47003 1547
rect 47289 1581 47339 1605
rect 47289 1547 47297 1581
rect 47331 1547 47339 1581
rect 47289 1523 47339 1547
rect 47625 1581 47675 1605
rect 47625 1547 47633 1581
rect 47667 1547 47675 1581
rect 47625 1523 47675 1547
rect 47961 1581 48011 1605
rect 47961 1547 47969 1581
rect 48003 1547 48011 1581
rect 47961 1523 48011 1547
rect 48297 1581 48347 1605
rect 48297 1547 48305 1581
rect 48339 1547 48347 1581
rect 48297 1523 48347 1547
rect 48633 1581 48683 1605
rect 48633 1547 48641 1581
rect 48675 1547 48683 1581
rect 48633 1523 48683 1547
rect 48969 1581 49019 1605
rect 48969 1547 48977 1581
rect 49011 1547 49019 1581
rect 48969 1523 49019 1547
rect 49305 1581 49355 1605
rect 49305 1547 49313 1581
rect 49347 1547 49355 1581
rect 49305 1523 49355 1547
rect 49641 1581 49691 1605
rect 49641 1547 49649 1581
rect 49683 1547 49691 1581
rect 49641 1523 49691 1547
rect 49977 1581 50027 1605
rect 49977 1547 49985 1581
rect 50019 1547 50027 1581
rect 49977 1523 50027 1547
rect 50313 1581 50363 1605
rect 50313 1547 50321 1581
rect 50355 1547 50363 1581
rect 50313 1523 50363 1547
rect 50649 1581 50699 1605
rect 50649 1547 50657 1581
rect 50691 1547 50699 1581
rect 50649 1523 50699 1547
rect 50985 1581 51035 1605
rect 50985 1547 50993 1581
rect 51027 1547 51035 1581
rect 50985 1523 51035 1547
rect 51321 1581 51371 1605
rect 51321 1547 51329 1581
rect 51363 1547 51371 1581
rect 51321 1523 51371 1547
rect 51657 1581 51707 1605
rect 51657 1547 51665 1581
rect 51699 1547 51707 1581
rect 51657 1523 51707 1547
rect 51993 1581 52043 1605
rect 51993 1547 52001 1581
rect 52035 1547 52043 1581
rect 51993 1523 52043 1547
rect 52329 1581 52379 1605
rect 52329 1547 52337 1581
rect 52371 1547 52379 1581
rect 52329 1523 52379 1547
rect 52665 1581 52715 1605
rect 52665 1547 52673 1581
rect 52707 1547 52715 1581
rect 52665 1523 52715 1547
rect 53001 1581 53051 1605
rect 53001 1547 53009 1581
rect 53043 1547 53051 1581
rect 53001 1523 53051 1547
rect 53337 1581 53387 1605
rect 53337 1547 53345 1581
rect 53379 1547 53387 1581
rect 53337 1523 53387 1547
rect 53673 1581 53723 1605
rect 53673 1547 53681 1581
rect 53715 1547 53723 1581
rect 53673 1523 53723 1547
rect 54009 1581 54059 1605
rect 54009 1547 54017 1581
rect 54051 1547 54059 1581
rect 54009 1523 54059 1547
rect 54345 1581 54395 1605
rect 54345 1547 54353 1581
rect 54387 1547 54395 1581
rect 54345 1523 54395 1547
rect 54681 1581 54731 1605
rect 54681 1547 54689 1581
rect 54723 1547 54731 1581
rect 54681 1523 54731 1547
rect 55017 1581 55067 1605
rect 55017 1547 55025 1581
rect 55059 1547 55067 1581
rect 55017 1523 55067 1547
rect 55353 1581 55403 1605
rect 55353 1547 55361 1581
rect 55395 1547 55403 1581
rect 55353 1523 55403 1547
rect 55689 1581 55739 1605
rect 55689 1547 55697 1581
rect 55731 1547 55739 1581
rect 55689 1523 55739 1547
rect 56025 1581 56075 1605
rect 56025 1547 56033 1581
rect 56067 1547 56075 1581
rect 56025 1523 56075 1547
rect 56361 1581 56411 1605
rect 56361 1547 56369 1581
rect 56403 1547 56411 1581
rect 56361 1523 56411 1547
rect 56697 1581 56747 1605
rect 56697 1547 56705 1581
rect 56739 1547 56747 1581
rect 56697 1523 56747 1547
rect 57033 1581 57083 1605
rect 57033 1547 57041 1581
rect 57075 1547 57083 1581
rect 57033 1523 57083 1547
rect 57369 1581 57419 1605
rect 57369 1547 57377 1581
rect 57411 1547 57419 1581
rect 57369 1523 57419 1547
rect 57705 1581 57755 1605
rect 57705 1547 57713 1581
rect 57747 1547 57755 1581
rect 57705 1523 57755 1547
rect 58041 1581 58091 1605
rect 58041 1547 58049 1581
rect 58083 1547 58091 1581
rect 58041 1523 58091 1547
rect 58377 1581 58427 1605
rect 58377 1547 58385 1581
rect 58419 1547 58427 1581
rect 58377 1523 58427 1547
rect 58713 1581 58763 1605
rect 58713 1547 58721 1581
rect 58755 1547 58763 1581
rect 58713 1523 58763 1547
rect 59049 1581 59099 1605
rect 59049 1547 59057 1581
rect 59091 1547 59099 1581
rect 59049 1523 59099 1547
rect 59385 1581 59435 1605
rect 59385 1547 59393 1581
rect 59427 1547 59435 1581
rect 59385 1523 59435 1547
rect 59721 1581 59771 1605
rect 59721 1547 59729 1581
rect 59763 1547 59771 1581
rect 59721 1523 59771 1547
rect 60057 1581 60107 1605
rect 60057 1547 60065 1581
rect 60099 1547 60107 1581
rect 60057 1523 60107 1547
rect 60393 1581 60443 1605
rect 60393 1547 60401 1581
rect 60435 1547 60443 1581
rect 60393 1523 60443 1547
rect 60729 1581 60779 1605
rect 60729 1547 60737 1581
rect 60771 1547 60779 1581
rect 60729 1523 60779 1547
rect 61065 1581 61115 1605
rect 61065 1547 61073 1581
rect 61107 1547 61115 1581
rect 61065 1523 61115 1547
rect 61401 1581 61451 1605
rect 61401 1547 61409 1581
rect 61443 1547 61451 1581
rect 61401 1523 61451 1547
rect 61737 1581 61787 1605
rect 61737 1547 61745 1581
rect 61779 1547 61787 1581
rect 61737 1523 61787 1547
rect 62073 1581 62123 1605
rect 62073 1547 62081 1581
rect 62115 1547 62123 1581
rect 62073 1523 62123 1547
rect 62409 1581 62459 1605
rect 62409 1547 62417 1581
rect 62451 1547 62459 1581
rect 62409 1523 62459 1547
rect 62745 1581 62795 1605
rect 62745 1547 62753 1581
rect 62787 1547 62795 1581
rect 62745 1523 62795 1547
rect 63081 1581 63131 1605
rect 63081 1547 63089 1581
rect 63123 1547 63131 1581
rect 63081 1523 63131 1547
rect 63417 1581 63467 1605
rect 63417 1547 63425 1581
rect 63459 1547 63467 1581
rect 63417 1523 63467 1547
rect 63753 1581 63803 1605
rect 63753 1547 63761 1581
rect 63795 1547 63803 1581
rect 63753 1523 63803 1547
rect 64089 1581 64139 1605
rect 64089 1547 64097 1581
rect 64131 1547 64139 1581
rect 64089 1523 64139 1547
rect 64425 1581 64475 1605
rect 64425 1547 64433 1581
rect 64467 1547 64475 1581
rect 64425 1523 64475 1547
rect 64761 1581 64811 1605
rect 64761 1547 64769 1581
rect 64803 1547 64811 1581
rect 64761 1523 64811 1547
rect 65097 1581 65147 1605
rect 65097 1547 65105 1581
rect 65139 1547 65147 1581
rect 65097 1523 65147 1547
rect 65433 1581 65483 1605
rect 65433 1547 65441 1581
rect 65475 1547 65483 1581
rect 65433 1523 65483 1547
rect 65769 1581 65819 1605
rect 65769 1547 65777 1581
rect 65811 1547 65819 1581
rect 65769 1523 65819 1547
rect 66105 1581 66155 1605
rect 66105 1547 66113 1581
rect 66147 1547 66155 1581
rect 66105 1523 66155 1547
rect 66441 1581 66491 1605
rect 66441 1547 66449 1581
rect 66483 1547 66491 1581
rect 66441 1523 66491 1547
rect 66777 1581 66827 1605
rect 66777 1547 66785 1581
rect 66819 1547 66827 1581
rect 66777 1523 66827 1547
rect 67113 1581 67163 1605
rect 67113 1547 67121 1581
rect 67155 1547 67163 1581
rect 67113 1523 67163 1547
rect 67449 1581 67499 1605
rect 67449 1547 67457 1581
rect 67491 1547 67499 1581
rect 67449 1523 67499 1547
rect 67785 1581 67835 1605
rect 67785 1547 67793 1581
rect 67827 1547 67835 1581
rect 67785 1523 67835 1547
rect 68121 1581 68171 1605
rect 68121 1547 68129 1581
rect 68163 1547 68171 1581
rect 68121 1523 68171 1547
rect 68457 1581 68507 1605
rect 68457 1547 68465 1581
rect 68499 1547 68507 1581
rect 68457 1523 68507 1547
rect 68793 1581 68843 1605
rect 68793 1547 68801 1581
rect 68835 1547 68843 1581
rect 68793 1523 68843 1547
rect 69129 1581 69179 1605
rect 69129 1547 69137 1581
rect 69171 1547 69179 1581
rect 69129 1523 69179 1547
rect 69465 1581 69515 1605
rect 69465 1547 69473 1581
rect 69507 1547 69515 1581
rect 69465 1523 69515 1547
rect 69801 1581 69851 1605
rect 69801 1547 69809 1581
rect 69843 1547 69851 1581
rect 69801 1523 69851 1547
rect 70137 1581 70187 1605
rect 70137 1547 70145 1581
rect 70179 1547 70187 1581
rect 70137 1523 70187 1547
rect 70473 1581 70523 1605
rect 70473 1547 70481 1581
rect 70515 1547 70523 1581
rect 70473 1523 70523 1547
rect 70809 1581 70859 1605
rect 70809 1547 70817 1581
rect 70851 1547 70859 1581
rect 70809 1523 70859 1547
rect 71145 1581 71195 1605
rect 71145 1547 71153 1581
rect 71187 1547 71195 1581
rect 71145 1523 71195 1547
rect 71481 1581 71531 1605
rect 71481 1547 71489 1581
rect 71523 1547 71531 1581
rect 71481 1523 71531 1547
rect 71817 1581 71867 1605
rect 71817 1547 71825 1581
rect 71859 1547 71867 1581
rect 71817 1523 71867 1547
rect 72153 1581 72203 1605
rect 72153 1547 72161 1581
rect 72195 1547 72203 1581
rect 72153 1523 72203 1547
rect 72489 1581 72539 1605
rect 72489 1547 72497 1581
rect 72531 1547 72539 1581
rect 72489 1523 72539 1547
rect 72825 1581 72875 1605
rect 72825 1547 72833 1581
rect 72867 1547 72875 1581
rect 72825 1523 72875 1547
rect 73161 1581 73211 1605
rect 73161 1547 73169 1581
rect 73203 1547 73211 1581
rect 73161 1523 73211 1547
rect 73497 1581 73547 1605
rect 73497 1547 73505 1581
rect 73539 1547 73547 1581
rect 73497 1523 73547 1547
<< nsubdiffcont >>
rect 1937 36191 1971 36225
rect 2273 36191 2307 36225
rect 2609 36191 2643 36225
rect 2945 36191 2979 36225
rect 3281 36191 3315 36225
rect 3617 36191 3651 36225
rect 3953 36191 3987 36225
rect 4289 36191 4323 36225
rect 4625 36191 4659 36225
rect 4961 36191 4995 36225
rect 5297 36191 5331 36225
rect 5633 36191 5667 36225
rect 5969 36191 6003 36225
rect 6305 36191 6339 36225
rect 6641 36191 6675 36225
rect 6977 36191 7011 36225
rect 7313 36191 7347 36225
rect 7649 36191 7683 36225
rect 7985 36191 8019 36225
rect 8321 36191 8355 36225
rect 8657 36191 8691 36225
rect 8993 36191 9027 36225
rect 9329 36191 9363 36225
rect 9665 36191 9699 36225
rect 10001 36191 10035 36225
rect 10337 36191 10371 36225
rect 10673 36191 10707 36225
rect 11009 36191 11043 36225
rect 11345 36191 11379 36225
rect 11681 36191 11715 36225
rect 12017 36191 12051 36225
rect 12353 36191 12387 36225
rect 12689 36191 12723 36225
rect 13025 36191 13059 36225
rect 13361 36191 13395 36225
rect 13697 36191 13731 36225
rect 14033 36191 14067 36225
rect 14369 36191 14403 36225
rect 14705 36191 14739 36225
rect 15041 36191 15075 36225
rect 15377 36191 15411 36225
rect 15713 36191 15747 36225
rect 16049 36191 16083 36225
rect 16385 36191 16419 36225
rect 16721 36191 16755 36225
rect 17057 36191 17091 36225
rect 17393 36191 17427 36225
rect 17729 36191 17763 36225
rect 18065 36191 18099 36225
rect 18401 36191 18435 36225
rect 18737 36191 18771 36225
rect 19073 36191 19107 36225
rect 19409 36191 19443 36225
rect 19745 36191 19779 36225
rect 20081 36191 20115 36225
rect 20417 36191 20451 36225
rect 20753 36191 20787 36225
rect 21089 36191 21123 36225
rect 21425 36191 21459 36225
rect 21761 36191 21795 36225
rect 22097 36191 22131 36225
rect 22433 36191 22467 36225
rect 22769 36191 22803 36225
rect 23105 36191 23139 36225
rect 23441 36191 23475 36225
rect 23777 36191 23811 36225
rect 24113 36191 24147 36225
rect 24449 36191 24483 36225
rect 24785 36191 24819 36225
rect 25121 36191 25155 36225
rect 25457 36191 25491 36225
rect 25793 36191 25827 36225
rect 26129 36191 26163 36225
rect 26465 36191 26499 36225
rect 26801 36191 26835 36225
rect 27137 36191 27171 36225
rect 27473 36191 27507 36225
rect 27809 36191 27843 36225
rect 28145 36191 28179 36225
rect 28481 36191 28515 36225
rect 28817 36191 28851 36225
rect 29153 36191 29187 36225
rect 29489 36191 29523 36225
rect 29825 36191 29859 36225
rect 30161 36191 30195 36225
rect 30497 36191 30531 36225
rect 30833 36191 30867 36225
rect 31169 36191 31203 36225
rect 31505 36191 31539 36225
rect 31841 36191 31875 36225
rect 32177 36191 32211 36225
rect 32513 36191 32547 36225
rect 32849 36191 32883 36225
rect 33185 36191 33219 36225
rect 33521 36191 33555 36225
rect 33857 36191 33891 36225
rect 34193 36191 34227 36225
rect 34529 36191 34563 36225
rect 34865 36191 34899 36225
rect 35201 36191 35235 36225
rect 35537 36191 35571 36225
rect 35873 36191 35907 36225
rect 36209 36191 36243 36225
rect 36545 36191 36579 36225
rect 36881 36191 36915 36225
rect 37217 36191 37251 36225
rect 37553 36191 37587 36225
rect 37889 36191 37923 36225
rect 38225 36191 38259 36225
rect 38561 36191 38595 36225
rect 38897 36191 38931 36225
rect 39233 36191 39267 36225
rect 39569 36191 39603 36225
rect 39905 36191 39939 36225
rect 40241 36191 40275 36225
rect 40577 36191 40611 36225
rect 40913 36191 40947 36225
rect 41249 36191 41283 36225
rect 41585 36191 41619 36225
rect 41921 36191 41955 36225
rect 42257 36191 42291 36225
rect 42593 36191 42627 36225
rect 42929 36191 42963 36225
rect 43265 36191 43299 36225
rect 43601 36191 43635 36225
rect 43937 36191 43971 36225
rect 44273 36191 44307 36225
rect 44609 36191 44643 36225
rect 44945 36191 44979 36225
rect 45281 36191 45315 36225
rect 45617 36191 45651 36225
rect 45953 36191 45987 36225
rect 46289 36191 46323 36225
rect 46625 36191 46659 36225
rect 46961 36191 46995 36225
rect 47297 36191 47331 36225
rect 47633 36191 47667 36225
rect 47969 36191 48003 36225
rect 48305 36191 48339 36225
rect 48641 36191 48675 36225
rect 48977 36191 49011 36225
rect 49313 36191 49347 36225
rect 49649 36191 49683 36225
rect 49985 36191 50019 36225
rect 50321 36191 50355 36225
rect 50657 36191 50691 36225
rect 50993 36191 51027 36225
rect 51329 36191 51363 36225
rect 51665 36191 51699 36225
rect 52001 36191 52035 36225
rect 52337 36191 52371 36225
rect 52673 36191 52707 36225
rect 53009 36191 53043 36225
rect 53345 36191 53379 36225
rect 53681 36191 53715 36225
rect 54017 36191 54051 36225
rect 54353 36191 54387 36225
rect 54689 36191 54723 36225
rect 55025 36191 55059 36225
rect 55361 36191 55395 36225
rect 55697 36191 55731 36225
rect 56033 36191 56067 36225
rect 56369 36191 56403 36225
rect 56705 36191 56739 36225
rect 57041 36191 57075 36225
rect 57377 36191 57411 36225
rect 57713 36191 57747 36225
rect 58049 36191 58083 36225
rect 58385 36191 58419 36225
rect 58721 36191 58755 36225
rect 59057 36191 59091 36225
rect 59393 36191 59427 36225
rect 59729 36191 59763 36225
rect 60065 36191 60099 36225
rect 60401 36191 60435 36225
rect 60737 36191 60771 36225
rect 61073 36191 61107 36225
rect 61409 36191 61443 36225
rect 61745 36191 61779 36225
rect 62081 36191 62115 36225
rect 62417 36191 62451 36225
rect 62753 36191 62787 36225
rect 63089 36191 63123 36225
rect 63425 36191 63459 36225
rect 63761 36191 63795 36225
rect 64097 36191 64131 36225
rect 64433 36191 64467 36225
rect 64769 36191 64803 36225
rect 65105 36191 65139 36225
rect 65441 36191 65475 36225
rect 65777 36191 65811 36225
rect 66113 36191 66147 36225
rect 66449 36191 66483 36225
rect 66785 36191 66819 36225
rect 67121 36191 67155 36225
rect 67457 36191 67491 36225
rect 67793 36191 67827 36225
rect 68129 36191 68163 36225
rect 68465 36191 68499 36225
rect 68801 36191 68835 36225
rect 69137 36191 69171 36225
rect 69473 36191 69507 36225
rect 69809 36191 69843 36225
rect 70145 36191 70179 36225
rect 70481 36191 70515 36225
rect 70817 36191 70851 36225
rect 71153 36191 71187 36225
rect 71489 36191 71523 36225
rect 71825 36191 71859 36225
rect 72161 36191 72195 36225
rect 72497 36191 72531 36225
rect 72833 36191 72867 36225
rect 73169 36191 73203 36225
rect 73505 36191 73539 36225
rect 1601 35819 1635 35853
rect 73949 35819 73983 35853
rect 1601 35483 1635 35517
rect 73949 35483 73983 35517
rect 1601 35147 1635 35181
rect 73949 35147 73983 35181
rect 1601 34811 1635 34845
rect 73949 34811 73983 34845
rect 1601 34475 1635 34509
rect 73949 34475 73983 34509
rect 1601 34139 1635 34173
rect 73949 34139 73983 34173
rect 1601 33803 1635 33837
rect 73949 33803 73983 33837
rect 1601 33467 1635 33501
rect 73949 33467 73983 33501
rect 1601 33131 1635 33165
rect 73949 33131 73983 33165
rect 1601 32795 1635 32829
rect 73949 32795 73983 32829
rect 1601 32459 1635 32493
rect 73949 32459 73983 32493
rect 1601 32123 1635 32157
rect 73949 32123 73983 32157
rect 1601 31787 1635 31821
rect 73949 31787 73983 31821
rect 1601 31451 1635 31485
rect 73949 31451 73983 31485
rect 1601 31115 1635 31149
rect 73949 31115 73983 31149
rect 1601 30779 1635 30813
rect 73949 30779 73983 30813
rect 1601 30443 1635 30477
rect 73949 30443 73983 30477
rect 1601 30107 1635 30141
rect 73949 30107 73983 30141
rect 1601 29771 1635 29805
rect 73949 29771 73983 29805
rect 1601 29435 1635 29469
rect 73949 29435 73983 29469
rect 1601 29099 1635 29133
rect 73949 29099 73983 29133
rect 1601 28763 1635 28797
rect 73949 28763 73983 28797
rect 1601 28427 1635 28461
rect 73949 28427 73983 28461
rect 1601 28091 1635 28125
rect 73949 28091 73983 28125
rect 1601 27755 1635 27789
rect 73949 27755 73983 27789
rect 1601 27419 1635 27453
rect 73949 27419 73983 27453
rect 1601 27083 1635 27117
rect 73949 27083 73983 27117
rect 1601 26747 1635 26781
rect 73949 26747 73983 26781
rect 1601 26411 1635 26445
rect 73949 26411 73983 26445
rect 1601 26075 1635 26109
rect 73949 26075 73983 26109
rect 1601 25739 1635 25773
rect 73949 25739 73983 25773
rect 1601 25403 1635 25437
rect 73949 25403 73983 25437
rect 1601 25067 1635 25101
rect 73949 25067 73983 25101
rect 1601 24731 1635 24765
rect 73949 24731 73983 24765
rect 1601 24395 1635 24429
rect 73949 24395 73983 24429
rect 1601 24059 1635 24093
rect 73949 24059 73983 24093
rect 1601 23723 1635 23757
rect 73949 23723 73983 23757
rect 1601 23387 1635 23421
rect 73949 23387 73983 23421
rect 1601 23051 1635 23085
rect 73949 23051 73983 23085
rect 1601 22715 1635 22749
rect 73949 22715 73983 22749
rect 1601 22379 1635 22413
rect 73949 22379 73983 22413
rect 1601 22043 1635 22077
rect 73949 22043 73983 22077
rect 1601 21707 1635 21741
rect 73949 21707 73983 21741
rect 1601 21371 1635 21405
rect 73949 21371 73983 21405
rect 1601 21035 1635 21069
rect 73949 21035 73983 21069
rect 1601 20699 1635 20733
rect 73949 20699 73983 20733
rect 1601 20363 1635 20397
rect 73949 20363 73983 20397
rect 1601 20027 1635 20061
rect 73949 20027 73983 20061
rect 1601 19691 1635 19725
rect 73949 19691 73983 19725
rect 1601 19355 1635 19389
rect 73949 19355 73983 19389
rect 1601 19019 1635 19053
rect 73949 19019 73983 19053
rect 1601 18683 1635 18717
rect 73949 18683 73983 18717
rect 1601 18347 1635 18381
rect 73949 18347 73983 18381
rect 1601 18011 1635 18045
rect 73949 18011 73983 18045
rect 1601 17675 1635 17709
rect 73949 17675 73983 17709
rect 1601 17339 1635 17373
rect 73949 17339 73983 17373
rect 1601 17003 1635 17037
rect 73949 17003 73983 17037
rect 1601 16667 1635 16701
rect 73949 16667 73983 16701
rect 1601 16331 1635 16365
rect 73949 16331 73983 16365
rect 1601 15995 1635 16029
rect 73949 15995 73983 16029
rect 1601 15659 1635 15693
rect 73949 15659 73983 15693
rect 1601 15323 1635 15357
rect 73949 15323 73983 15357
rect 1601 14987 1635 15021
rect 73949 14987 73983 15021
rect 1601 14651 1635 14685
rect 73949 14651 73983 14685
rect 1601 14315 1635 14349
rect 73949 14315 73983 14349
rect 1601 13979 1635 14013
rect 73949 13979 73983 14013
rect 1601 13643 1635 13677
rect 73949 13643 73983 13677
rect 1601 13307 1635 13341
rect 73949 13307 73983 13341
rect 1601 12971 1635 13005
rect 73949 12971 73983 13005
rect 1601 12635 1635 12669
rect 73949 12635 73983 12669
rect 1601 12299 1635 12333
rect 73949 12299 73983 12333
rect 1601 11963 1635 11997
rect 73949 11963 73983 11997
rect 1601 11627 1635 11661
rect 73949 11627 73983 11661
rect 1601 11291 1635 11325
rect 73949 11291 73983 11325
rect 1601 10955 1635 10989
rect 73949 10955 73983 10989
rect 1601 10619 1635 10653
rect 73949 10619 73983 10653
rect 1601 10283 1635 10317
rect 73949 10283 73983 10317
rect 1601 9947 1635 9981
rect 73949 9947 73983 9981
rect 1601 9611 1635 9645
rect 73949 9611 73983 9645
rect 1601 9275 1635 9309
rect 73949 9275 73983 9309
rect 1601 8939 1635 8973
rect 73949 8939 73983 8973
rect 1601 8603 1635 8637
rect 73949 8603 73983 8637
rect 1601 8267 1635 8301
rect 73949 8267 73983 8301
rect 1601 7931 1635 7965
rect 73949 7931 73983 7965
rect 1601 7595 1635 7629
rect 73949 7595 73983 7629
rect 1601 7259 1635 7293
rect 73949 7259 73983 7293
rect 1601 6923 1635 6957
rect 73949 6923 73983 6957
rect 1601 6587 1635 6621
rect 73949 6587 73983 6621
rect 1601 6251 1635 6285
rect 73949 6251 73983 6285
rect 1601 5915 1635 5949
rect 73949 5915 73983 5949
rect 1601 5579 1635 5613
rect 73949 5579 73983 5613
rect 1601 5243 1635 5277
rect 73949 5243 73983 5277
rect 1601 4907 1635 4941
rect 73949 4907 73983 4941
rect 1601 4571 1635 4605
rect 73949 4571 73983 4605
rect 1601 4235 1635 4269
rect 73949 4235 73983 4269
rect 1601 3899 1635 3933
rect 73949 3899 73983 3933
rect 1601 3563 1635 3597
rect 73949 3563 73983 3597
rect 1601 3227 1635 3261
rect 73949 3227 73983 3261
rect 1601 2891 1635 2925
rect 73949 2891 73983 2925
rect 1601 2555 1635 2589
rect 73949 2555 73983 2589
rect 1601 2219 1635 2253
rect 73949 2219 73983 2253
rect 1601 1883 1635 1917
rect 73949 1883 73983 1917
rect 1937 1547 1971 1581
rect 2273 1547 2307 1581
rect 2609 1547 2643 1581
rect 2945 1547 2979 1581
rect 3281 1547 3315 1581
rect 3617 1547 3651 1581
rect 3953 1547 3987 1581
rect 4289 1547 4323 1581
rect 4625 1547 4659 1581
rect 4961 1547 4995 1581
rect 5297 1547 5331 1581
rect 5633 1547 5667 1581
rect 5969 1547 6003 1581
rect 6305 1547 6339 1581
rect 6641 1547 6675 1581
rect 6977 1547 7011 1581
rect 7313 1547 7347 1581
rect 7649 1547 7683 1581
rect 7985 1547 8019 1581
rect 8321 1547 8355 1581
rect 8657 1547 8691 1581
rect 8993 1547 9027 1581
rect 9329 1547 9363 1581
rect 9665 1547 9699 1581
rect 10001 1547 10035 1581
rect 10337 1547 10371 1581
rect 10673 1547 10707 1581
rect 11009 1547 11043 1581
rect 11345 1547 11379 1581
rect 11681 1547 11715 1581
rect 12017 1547 12051 1581
rect 12353 1547 12387 1581
rect 12689 1547 12723 1581
rect 13025 1547 13059 1581
rect 13361 1547 13395 1581
rect 13697 1547 13731 1581
rect 14033 1547 14067 1581
rect 14369 1547 14403 1581
rect 14705 1547 14739 1581
rect 15041 1547 15075 1581
rect 15377 1547 15411 1581
rect 15713 1547 15747 1581
rect 16049 1547 16083 1581
rect 16385 1547 16419 1581
rect 16721 1547 16755 1581
rect 17057 1547 17091 1581
rect 17393 1547 17427 1581
rect 17729 1547 17763 1581
rect 18065 1547 18099 1581
rect 18401 1547 18435 1581
rect 18737 1547 18771 1581
rect 19073 1547 19107 1581
rect 19409 1547 19443 1581
rect 19745 1547 19779 1581
rect 20081 1547 20115 1581
rect 20417 1547 20451 1581
rect 20753 1547 20787 1581
rect 21089 1547 21123 1581
rect 21425 1547 21459 1581
rect 21761 1547 21795 1581
rect 22097 1547 22131 1581
rect 22433 1547 22467 1581
rect 22769 1547 22803 1581
rect 23105 1547 23139 1581
rect 23441 1547 23475 1581
rect 23777 1547 23811 1581
rect 24113 1547 24147 1581
rect 24449 1547 24483 1581
rect 24785 1547 24819 1581
rect 25121 1547 25155 1581
rect 25457 1547 25491 1581
rect 25793 1547 25827 1581
rect 26129 1547 26163 1581
rect 26465 1547 26499 1581
rect 26801 1547 26835 1581
rect 27137 1547 27171 1581
rect 27473 1547 27507 1581
rect 27809 1547 27843 1581
rect 28145 1547 28179 1581
rect 28481 1547 28515 1581
rect 28817 1547 28851 1581
rect 29153 1547 29187 1581
rect 29489 1547 29523 1581
rect 29825 1547 29859 1581
rect 30161 1547 30195 1581
rect 30497 1547 30531 1581
rect 30833 1547 30867 1581
rect 31169 1547 31203 1581
rect 31505 1547 31539 1581
rect 31841 1547 31875 1581
rect 32177 1547 32211 1581
rect 32513 1547 32547 1581
rect 32849 1547 32883 1581
rect 33185 1547 33219 1581
rect 33521 1547 33555 1581
rect 33857 1547 33891 1581
rect 34193 1547 34227 1581
rect 34529 1547 34563 1581
rect 34865 1547 34899 1581
rect 35201 1547 35235 1581
rect 35537 1547 35571 1581
rect 35873 1547 35907 1581
rect 36209 1547 36243 1581
rect 36545 1547 36579 1581
rect 36881 1547 36915 1581
rect 37217 1547 37251 1581
rect 37553 1547 37587 1581
rect 37889 1547 37923 1581
rect 38225 1547 38259 1581
rect 38561 1547 38595 1581
rect 38897 1547 38931 1581
rect 39233 1547 39267 1581
rect 39569 1547 39603 1581
rect 39905 1547 39939 1581
rect 40241 1547 40275 1581
rect 40577 1547 40611 1581
rect 40913 1547 40947 1581
rect 41249 1547 41283 1581
rect 41585 1547 41619 1581
rect 41921 1547 41955 1581
rect 42257 1547 42291 1581
rect 42593 1547 42627 1581
rect 42929 1547 42963 1581
rect 43265 1547 43299 1581
rect 43601 1547 43635 1581
rect 43937 1547 43971 1581
rect 44273 1547 44307 1581
rect 44609 1547 44643 1581
rect 44945 1547 44979 1581
rect 45281 1547 45315 1581
rect 45617 1547 45651 1581
rect 45953 1547 45987 1581
rect 46289 1547 46323 1581
rect 46625 1547 46659 1581
rect 46961 1547 46995 1581
rect 47297 1547 47331 1581
rect 47633 1547 47667 1581
rect 47969 1547 48003 1581
rect 48305 1547 48339 1581
rect 48641 1547 48675 1581
rect 48977 1547 49011 1581
rect 49313 1547 49347 1581
rect 49649 1547 49683 1581
rect 49985 1547 50019 1581
rect 50321 1547 50355 1581
rect 50657 1547 50691 1581
rect 50993 1547 51027 1581
rect 51329 1547 51363 1581
rect 51665 1547 51699 1581
rect 52001 1547 52035 1581
rect 52337 1547 52371 1581
rect 52673 1547 52707 1581
rect 53009 1547 53043 1581
rect 53345 1547 53379 1581
rect 53681 1547 53715 1581
rect 54017 1547 54051 1581
rect 54353 1547 54387 1581
rect 54689 1547 54723 1581
rect 55025 1547 55059 1581
rect 55361 1547 55395 1581
rect 55697 1547 55731 1581
rect 56033 1547 56067 1581
rect 56369 1547 56403 1581
rect 56705 1547 56739 1581
rect 57041 1547 57075 1581
rect 57377 1547 57411 1581
rect 57713 1547 57747 1581
rect 58049 1547 58083 1581
rect 58385 1547 58419 1581
rect 58721 1547 58755 1581
rect 59057 1547 59091 1581
rect 59393 1547 59427 1581
rect 59729 1547 59763 1581
rect 60065 1547 60099 1581
rect 60401 1547 60435 1581
rect 60737 1547 60771 1581
rect 61073 1547 61107 1581
rect 61409 1547 61443 1581
rect 61745 1547 61779 1581
rect 62081 1547 62115 1581
rect 62417 1547 62451 1581
rect 62753 1547 62787 1581
rect 63089 1547 63123 1581
rect 63425 1547 63459 1581
rect 63761 1547 63795 1581
rect 64097 1547 64131 1581
rect 64433 1547 64467 1581
rect 64769 1547 64803 1581
rect 65105 1547 65139 1581
rect 65441 1547 65475 1581
rect 65777 1547 65811 1581
rect 66113 1547 66147 1581
rect 66449 1547 66483 1581
rect 66785 1547 66819 1581
rect 67121 1547 67155 1581
rect 67457 1547 67491 1581
rect 67793 1547 67827 1581
rect 68129 1547 68163 1581
rect 68465 1547 68499 1581
rect 68801 1547 68835 1581
rect 69137 1547 69171 1581
rect 69473 1547 69507 1581
rect 69809 1547 69843 1581
rect 70145 1547 70179 1581
rect 70481 1547 70515 1581
rect 70817 1547 70851 1581
rect 71153 1547 71187 1581
rect 71489 1547 71523 1581
rect 71825 1547 71859 1581
rect 72161 1547 72195 1581
rect 72497 1547 72531 1581
rect 72833 1547 72867 1581
rect 73169 1547 73203 1581
rect 73505 1547 73539 1581
<< locali >>
rect 1937 36225 1971 36241
rect 1937 36175 1971 36191
rect 2273 36225 2307 36241
rect 2273 36175 2307 36191
rect 2609 36225 2643 36241
rect 2609 36175 2643 36191
rect 2945 36225 2979 36241
rect 2945 36175 2979 36191
rect 3281 36225 3315 36241
rect 3281 36175 3315 36191
rect 3617 36225 3651 36241
rect 3617 36175 3651 36191
rect 3953 36225 3987 36241
rect 3953 36175 3987 36191
rect 4289 36225 4323 36241
rect 4289 36175 4323 36191
rect 4625 36225 4659 36241
rect 4625 36175 4659 36191
rect 4961 36225 4995 36241
rect 4961 36175 4995 36191
rect 5297 36225 5331 36241
rect 5297 36175 5331 36191
rect 5633 36225 5667 36241
rect 5633 36175 5667 36191
rect 5969 36225 6003 36241
rect 5969 36175 6003 36191
rect 6305 36225 6339 36241
rect 6305 36175 6339 36191
rect 6641 36225 6675 36241
rect 6641 36175 6675 36191
rect 6977 36225 7011 36241
rect 6977 36175 7011 36191
rect 7313 36225 7347 36241
rect 7313 36175 7347 36191
rect 7649 36225 7683 36241
rect 7649 36175 7683 36191
rect 7985 36225 8019 36241
rect 7985 36175 8019 36191
rect 8321 36225 8355 36241
rect 8321 36175 8355 36191
rect 8657 36225 8691 36241
rect 8657 36175 8691 36191
rect 8993 36225 9027 36241
rect 8993 36175 9027 36191
rect 9329 36225 9363 36241
rect 9329 36175 9363 36191
rect 9665 36225 9699 36241
rect 9665 36175 9699 36191
rect 10001 36225 10035 36241
rect 10001 36175 10035 36191
rect 10337 36225 10371 36241
rect 10337 36175 10371 36191
rect 10673 36225 10707 36241
rect 10673 36175 10707 36191
rect 11009 36225 11043 36241
rect 11009 36175 11043 36191
rect 11345 36225 11379 36241
rect 11345 36175 11379 36191
rect 11681 36225 11715 36241
rect 11681 36175 11715 36191
rect 12017 36225 12051 36241
rect 12017 36175 12051 36191
rect 12353 36225 12387 36241
rect 12353 36175 12387 36191
rect 12689 36225 12723 36241
rect 12689 36175 12723 36191
rect 13025 36225 13059 36241
rect 13025 36175 13059 36191
rect 13361 36225 13395 36241
rect 13361 36175 13395 36191
rect 13697 36225 13731 36241
rect 13697 36175 13731 36191
rect 14033 36225 14067 36241
rect 14033 36175 14067 36191
rect 14369 36225 14403 36241
rect 14369 36175 14403 36191
rect 14705 36225 14739 36241
rect 14705 36175 14739 36191
rect 15041 36225 15075 36241
rect 15041 36175 15075 36191
rect 15377 36225 15411 36241
rect 15377 36175 15411 36191
rect 15713 36225 15747 36241
rect 15713 36175 15747 36191
rect 16049 36225 16083 36241
rect 16049 36175 16083 36191
rect 16385 36225 16419 36241
rect 16385 36175 16419 36191
rect 16721 36225 16755 36241
rect 16721 36175 16755 36191
rect 17057 36225 17091 36241
rect 17057 36175 17091 36191
rect 17393 36225 17427 36241
rect 17393 36175 17427 36191
rect 17729 36225 17763 36241
rect 17729 36175 17763 36191
rect 18065 36225 18099 36241
rect 18065 36175 18099 36191
rect 18401 36225 18435 36241
rect 18401 36175 18435 36191
rect 18737 36225 18771 36241
rect 18737 36175 18771 36191
rect 19073 36225 19107 36241
rect 19073 36175 19107 36191
rect 19409 36225 19443 36241
rect 19409 36175 19443 36191
rect 19745 36225 19779 36241
rect 19745 36175 19779 36191
rect 20081 36225 20115 36241
rect 20081 36175 20115 36191
rect 20417 36225 20451 36241
rect 20417 36175 20451 36191
rect 20753 36225 20787 36241
rect 20753 36175 20787 36191
rect 21089 36225 21123 36241
rect 21089 36175 21123 36191
rect 21425 36225 21459 36241
rect 21425 36175 21459 36191
rect 21761 36225 21795 36241
rect 21761 36175 21795 36191
rect 22097 36225 22131 36241
rect 22097 36175 22131 36191
rect 22433 36225 22467 36241
rect 22433 36175 22467 36191
rect 22769 36225 22803 36241
rect 22769 36175 22803 36191
rect 23105 36225 23139 36241
rect 23105 36175 23139 36191
rect 23441 36225 23475 36241
rect 23441 36175 23475 36191
rect 23777 36225 23811 36241
rect 23777 36175 23811 36191
rect 24113 36225 24147 36241
rect 24113 36175 24147 36191
rect 24449 36225 24483 36241
rect 24449 36175 24483 36191
rect 24785 36225 24819 36241
rect 24785 36175 24819 36191
rect 25121 36225 25155 36241
rect 25121 36175 25155 36191
rect 25457 36225 25491 36241
rect 25457 36175 25491 36191
rect 25793 36225 25827 36241
rect 25793 36175 25827 36191
rect 26129 36225 26163 36241
rect 26129 36175 26163 36191
rect 26465 36225 26499 36241
rect 26465 36175 26499 36191
rect 26801 36225 26835 36241
rect 26801 36175 26835 36191
rect 27137 36225 27171 36241
rect 27137 36175 27171 36191
rect 27473 36225 27507 36241
rect 27473 36175 27507 36191
rect 27809 36225 27843 36241
rect 27809 36175 27843 36191
rect 28145 36225 28179 36241
rect 28145 36175 28179 36191
rect 28481 36225 28515 36241
rect 28481 36175 28515 36191
rect 28817 36225 28851 36241
rect 28817 36175 28851 36191
rect 29153 36225 29187 36241
rect 29153 36175 29187 36191
rect 29489 36225 29523 36241
rect 29489 36175 29523 36191
rect 29825 36225 29859 36241
rect 29825 36175 29859 36191
rect 30161 36225 30195 36241
rect 30161 36175 30195 36191
rect 30497 36225 30531 36241
rect 30497 36175 30531 36191
rect 30833 36225 30867 36241
rect 30833 36175 30867 36191
rect 31169 36225 31203 36241
rect 31169 36175 31203 36191
rect 31505 36225 31539 36241
rect 31505 36175 31539 36191
rect 31841 36225 31875 36241
rect 31841 36175 31875 36191
rect 32177 36225 32211 36241
rect 32177 36175 32211 36191
rect 32513 36225 32547 36241
rect 32513 36175 32547 36191
rect 32849 36225 32883 36241
rect 32849 36175 32883 36191
rect 33185 36225 33219 36241
rect 33185 36175 33219 36191
rect 33521 36225 33555 36241
rect 33521 36175 33555 36191
rect 33857 36225 33891 36241
rect 33857 36175 33891 36191
rect 34193 36225 34227 36241
rect 34193 36175 34227 36191
rect 34529 36225 34563 36241
rect 34529 36175 34563 36191
rect 34865 36225 34899 36241
rect 34865 36175 34899 36191
rect 35201 36225 35235 36241
rect 35201 36175 35235 36191
rect 35537 36225 35571 36241
rect 35537 36175 35571 36191
rect 35873 36225 35907 36241
rect 35873 36175 35907 36191
rect 36209 36225 36243 36241
rect 36209 36175 36243 36191
rect 36545 36225 36579 36241
rect 36545 36175 36579 36191
rect 36881 36225 36915 36241
rect 36881 36175 36915 36191
rect 37217 36225 37251 36241
rect 37217 36175 37251 36191
rect 37553 36225 37587 36241
rect 37553 36175 37587 36191
rect 37889 36225 37923 36241
rect 37889 36175 37923 36191
rect 38225 36225 38259 36241
rect 38225 36175 38259 36191
rect 38561 36225 38595 36241
rect 38561 36175 38595 36191
rect 38897 36225 38931 36241
rect 38897 36175 38931 36191
rect 39233 36225 39267 36241
rect 39233 36175 39267 36191
rect 39569 36225 39603 36241
rect 39569 36175 39603 36191
rect 39905 36225 39939 36241
rect 39905 36175 39939 36191
rect 40241 36225 40275 36241
rect 40241 36175 40275 36191
rect 40577 36225 40611 36241
rect 40577 36175 40611 36191
rect 40913 36225 40947 36241
rect 40913 36175 40947 36191
rect 41249 36225 41283 36241
rect 41249 36175 41283 36191
rect 41585 36225 41619 36241
rect 41585 36175 41619 36191
rect 41921 36225 41955 36241
rect 41921 36175 41955 36191
rect 42257 36225 42291 36241
rect 42257 36175 42291 36191
rect 42593 36225 42627 36241
rect 42593 36175 42627 36191
rect 42929 36225 42963 36241
rect 42929 36175 42963 36191
rect 43265 36225 43299 36241
rect 43265 36175 43299 36191
rect 43601 36225 43635 36241
rect 43601 36175 43635 36191
rect 43937 36225 43971 36241
rect 43937 36175 43971 36191
rect 44273 36225 44307 36241
rect 44273 36175 44307 36191
rect 44609 36225 44643 36241
rect 44609 36175 44643 36191
rect 44945 36225 44979 36241
rect 44945 36175 44979 36191
rect 45281 36225 45315 36241
rect 45281 36175 45315 36191
rect 45617 36225 45651 36241
rect 45617 36175 45651 36191
rect 45953 36225 45987 36241
rect 45953 36175 45987 36191
rect 46289 36225 46323 36241
rect 46289 36175 46323 36191
rect 46625 36225 46659 36241
rect 46625 36175 46659 36191
rect 46961 36225 46995 36241
rect 46961 36175 46995 36191
rect 47297 36225 47331 36241
rect 47297 36175 47331 36191
rect 47633 36225 47667 36241
rect 47633 36175 47667 36191
rect 47969 36225 48003 36241
rect 47969 36175 48003 36191
rect 48305 36225 48339 36241
rect 48305 36175 48339 36191
rect 48641 36225 48675 36241
rect 48641 36175 48675 36191
rect 48977 36225 49011 36241
rect 48977 36175 49011 36191
rect 49313 36225 49347 36241
rect 49313 36175 49347 36191
rect 49649 36225 49683 36241
rect 49649 36175 49683 36191
rect 49985 36225 50019 36241
rect 49985 36175 50019 36191
rect 50321 36225 50355 36241
rect 50321 36175 50355 36191
rect 50657 36225 50691 36241
rect 50657 36175 50691 36191
rect 50993 36225 51027 36241
rect 50993 36175 51027 36191
rect 51329 36225 51363 36241
rect 51329 36175 51363 36191
rect 51665 36225 51699 36241
rect 51665 36175 51699 36191
rect 52001 36225 52035 36241
rect 52001 36175 52035 36191
rect 52337 36225 52371 36241
rect 52337 36175 52371 36191
rect 52673 36225 52707 36241
rect 52673 36175 52707 36191
rect 53009 36225 53043 36241
rect 53009 36175 53043 36191
rect 53345 36225 53379 36241
rect 53345 36175 53379 36191
rect 53681 36225 53715 36241
rect 53681 36175 53715 36191
rect 54017 36225 54051 36241
rect 54017 36175 54051 36191
rect 54353 36225 54387 36241
rect 54353 36175 54387 36191
rect 54689 36225 54723 36241
rect 54689 36175 54723 36191
rect 55025 36225 55059 36241
rect 55025 36175 55059 36191
rect 55361 36225 55395 36241
rect 55361 36175 55395 36191
rect 55697 36225 55731 36241
rect 55697 36175 55731 36191
rect 56033 36225 56067 36241
rect 56033 36175 56067 36191
rect 56369 36225 56403 36241
rect 56369 36175 56403 36191
rect 56705 36225 56739 36241
rect 56705 36175 56739 36191
rect 57041 36225 57075 36241
rect 57041 36175 57075 36191
rect 57377 36225 57411 36241
rect 57377 36175 57411 36191
rect 57713 36225 57747 36241
rect 57713 36175 57747 36191
rect 58049 36225 58083 36241
rect 58049 36175 58083 36191
rect 58385 36225 58419 36241
rect 58385 36175 58419 36191
rect 58721 36225 58755 36241
rect 58721 36175 58755 36191
rect 59057 36225 59091 36241
rect 59057 36175 59091 36191
rect 59393 36225 59427 36241
rect 59393 36175 59427 36191
rect 59729 36225 59763 36241
rect 59729 36175 59763 36191
rect 60065 36225 60099 36241
rect 60065 36175 60099 36191
rect 60401 36225 60435 36241
rect 60401 36175 60435 36191
rect 60737 36225 60771 36241
rect 60737 36175 60771 36191
rect 61073 36225 61107 36241
rect 61073 36175 61107 36191
rect 61409 36225 61443 36241
rect 61409 36175 61443 36191
rect 61745 36225 61779 36241
rect 61745 36175 61779 36191
rect 62081 36225 62115 36241
rect 62081 36175 62115 36191
rect 62417 36225 62451 36241
rect 62417 36175 62451 36191
rect 62753 36225 62787 36241
rect 62753 36175 62787 36191
rect 63089 36225 63123 36241
rect 63089 36175 63123 36191
rect 63425 36225 63459 36241
rect 63425 36175 63459 36191
rect 63761 36225 63795 36241
rect 63761 36175 63795 36191
rect 64097 36225 64131 36241
rect 64097 36175 64131 36191
rect 64433 36225 64467 36241
rect 64433 36175 64467 36191
rect 64769 36225 64803 36241
rect 64769 36175 64803 36191
rect 65105 36225 65139 36241
rect 65105 36175 65139 36191
rect 65441 36225 65475 36241
rect 65441 36175 65475 36191
rect 65777 36225 65811 36241
rect 65777 36175 65811 36191
rect 66113 36225 66147 36241
rect 66113 36175 66147 36191
rect 66449 36225 66483 36241
rect 66449 36175 66483 36191
rect 66785 36225 66819 36241
rect 66785 36175 66819 36191
rect 67121 36225 67155 36241
rect 67121 36175 67155 36191
rect 67457 36225 67491 36241
rect 67457 36175 67491 36191
rect 67793 36225 67827 36241
rect 67793 36175 67827 36191
rect 68129 36225 68163 36241
rect 68129 36175 68163 36191
rect 68465 36225 68499 36241
rect 68465 36175 68499 36191
rect 68801 36225 68835 36241
rect 68801 36175 68835 36191
rect 69137 36225 69171 36241
rect 69137 36175 69171 36191
rect 69473 36225 69507 36241
rect 69473 36175 69507 36191
rect 69809 36225 69843 36241
rect 69809 36175 69843 36191
rect 70145 36225 70179 36241
rect 70145 36175 70179 36191
rect 70481 36225 70515 36241
rect 70481 36175 70515 36191
rect 70817 36225 70851 36241
rect 70817 36175 70851 36191
rect 71153 36225 71187 36241
rect 71153 36175 71187 36191
rect 71489 36225 71523 36241
rect 71489 36175 71523 36191
rect 71825 36225 71859 36241
rect 71825 36175 71859 36191
rect 72161 36225 72195 36241
rect 72161 36175 72195 36191
rect 72497 36225 72531 36241
rect 72497 36175 72531 36191
rect 72833 36225 72867 36241
rect 72833 36175 72867 36191
rect 73169 36225 73203 36241
rect 73169 36175 73203 36191
rect 73505 36225 73539 36241
rect 73505 36175 73539 36191
rect 1601 35853 1635 35869
rect 1601 35803 1635 35819
rect 73949 35853 73983 35869
rect 73949 35803 73983 35819
rect 1601 35517 1635 35533
rect 1601 35467 1635 35483
rect 73949 35517 73983 35533
rect 73949 35467 73983 35483
rect 1601 35181 1635 35197
rect 1601 35131 1635 35147
rect 73949 35181 73983 35197
rect 73949 35131 73983 35147
rect 1601 34845 1635 34861
rect 1601 34795 1635 34811
rect 73949 34845 73983 34861
rect 73949 34795 73983 34811
rect 1601 34509 1635 34525
rect 1601 34459 1635 34475
rect 73949 34509 73983 34525
rect 73949 34459 73983 34475
rect 1601 34173 1635 34189
rect 1601 34123 1635 34139
rect 73949 34173 73983 34189
rect 73949 34123 73983 34139
rect 1601 33837 1635 33853
rect 1601 33787 1635 33803
rect 73949 33837 73983 33853
rect 73949 33787 73983 33803
rect 1601 33501 1635 33517
rect 1601 33451 1635 33467
rect 73949 33501 73983 33517
rect 73949 33451 73983 33467
rect 1601 33165 1635 33181
rect 1601 33115 1635 33131
rect 73949 33165 73983 33181
rect 73949 33115 73983 33131
rect 1601 32829 1635 32845
rect 1601 32779 1635 32795
rect 73949 32829 73983 32845
rect 73949 32779 73983 32795
rect 1601 32493 1635 32509
rect 1601 32443 1635 32459
rect 73949 32493 73983 32509
rect 73949 32443 73983 32459
rect 1601 32157 1635 32173
rect 1601 32107 1635 32123
rect 73949 32157 73983 32173
rect 73949 32107 73983 32123
rect 1601 31821 1635 31837
rect 1601 31771 1635 31787
rect 73949 31821 73983 31837
rect 73949 31771 73983 31787
rect 1601 31485 1635 31501
rect 1601 31435 1635 31451
rect 73949 31485 73983 31501
rect 73949 31435 73983 31451
rect 1601 31149 1635 31165
rect 1601 31099 1635 31115
rect 73949 31149 73983 31165
rect 73949 31099 73983 31115
rect 1601 30813 1635 30829
rect 1601 30763 1635 30779
rect 73949 30813 73983 30829
rect 73949 30763 73983 30779
rect 1601 30477 1635 30493
rect 1601 30427 1635 30443
rect 73949 30477 73983 30493
rect 73949 30427 73983 30443
rect 1601 30141 1635 30157
rect 1601 30091 1635 30107
rect 73949 30141 73983 30157
rect 73949 30091 73983 30107
rect 1601 29805 1635 29821
rect 1601 29755 1635 29771
rect 73949 29805 73983 29821
rect 73949 29755 73983 29771
rect 1601 29469 1635 29485
rect 1601 29419 1635 29435
rect 73949 29469 73983 29485
rect 73949 29419 73983 29435
rect 1601 29133 1635 29149
rect 1601 29083 1635 29099
rect 73949 29133 73983 29149
rect 73949 29083 73983 29099
rect 1601 28797 1635 28813
rect 1601 28747 1635 28763
rect 73949 28797 73983 28813
rect 73949 28747 73983 28763
rect 1601 28461 1635 28477
rect 1601 28411 1635 28427
rect 73949 28461 73983 28477
rect 73949 28411 73983 28427
rect 1601 28125 1635 28141
rect 1601 28075 1635 28091
rect 73949 28125 73983 28141
rect 73949 28075 73983 28091
rect 1601 27789 1635 27805
rect 1601 27739 1635 27755
rect 73949 27789 73983 27805
rect 73949 27739 73983 27755
rect 1601 27453 1635 27469
rect 1601 27403 1635 27419
rect 73949 27453 73983 27469
rect 73949 27403 73983 27419
rect 1601 27117 1635 27133
rect 1601 27067 1635 27083
rect 73949 27117 73983 27133
rect 73949 27067 73983 27083
rect 1601 26781 1635 26797
rect 1601 26731 1635 26747
rect 73949 26781 73983 26797
rect 73949 26731 73983 26747
rect 1601 26445 1635 26461
rect 1601 26395 1635 26411
rect 73949 26445 73983 26461
rect 73949 26395 73983 26411
rect 1601 26109 1635 26125
rect 1601 26059 1635 26075
rect 73949 26109 73983 26125
rect 73949 26059 73983 26075
rect 1601 25773 1635 25789
rect 1601 25723 1635 25739
rect 73949 25773 73983 25789
rect 73949 25723 73983 25739
rect 1601 25437 1635 25453
rect 1601 25387 1635 25403
rect 73949 25437 73983 25453
rect 73949 25387 73983 25403
rect 1601 25101 1635 25117
rect 1601 25051 1635 25067
rect 73949 25101 73983 25117
rect 73949 25051 73983 25067
rect 1601 24765 1635 24781
rect 1601 24715 1635 24731
rect 73949 24765 73983 24781
rect 73949 24715 73983 24731
rect 1601 24429 1635 24445
rect 1601 24379 1635 24395
rect 73949 24429 73983 24445
rect 73949 24379 73983 24395
rect 1601 24093 1635 24109
rect 1601 24043 1635 24059
rect 73949 24093 73983 24109
rect 73949 24043 73983 24059
rect 1601 23757 1635 23773
rect 1601 23707 1635 23723
rect 73949 23757 73983 23773
rect 73949 23707 73983 23723
rect 1601 23421 1635 23437
rect 1601 23371 1635 23387
rect 73949 23421 73983 23437
rect 73949 23371 73983 23387
rect 1601 23085 1635 23101
rect 1601 23035 1635 23051
rect 73949 23085 73983 23101
rect 73949 23035 73983 23051
rect 1601 22749 1635 22765
rect 1601 22699 1635 22715
rect 73949 22749 73983 22765
rect 73949 22699 73983 22715
rect 1601 22413 1635 22429
rect 1601 22363 1635 22379
rect 73949 22413 73983 22429
rect 73949 22363 73983 22379
rect 1601 22077 1635 22093
rect 1601 22027 1635 22043
rect 73949 22077 73983 22093
rect 73949 22027 73983 22043
rect 1601 21741 1635 21757
rect 1601 21691 1635 21707
rect 73949 21741 73983 21757
rect 73949 21691 73983 21707
rect 1601 21405 1635 21421
rect 1601 21355 1635 21371
rect 73949 21405 73983 21421
rect 73949 21355 73983 21371
rect 1601 21069 1635 21085
rect 1601 21019 1635 21035
rect 73949 21069 73983 21085
rect 73949 21019 73983 21035
rect 1601 20733 1635 20749
rect 1601 20683 1635 20699
rect 73949 20733 73983 20749
rect 73949 20683 73983 20699
rect 1601 20397 1635 20413
rect 1601 20347 1635 20363
rect 73949 20397 73983 20413
rect 73949 20347 73983 20363
rect 1601 20061 1635 20077
rect 1601 20011 1635 20027
rect 73949 20061 73983 20077
rect 73949 20011 73983 20027
rect 1601 19725 1635 19741
rect 1601 19675 1635 19691
rect 73949 19725 73983 19741
rect 73949 19675 73983 19691
rect 1601 19389 1635 19405
rect 1601 19339 1635 19355
rect 73949 19389 73983 19405
rect 73949 19339 73983 19355
rect 1601 19053 1635 19069
rect 1601 19003 1635 19019
rect 73949 19053 73983 19069
rect 73949 19003 73983 19019
rect 1601 18717 1635 18733
rect 1601 18667 1635 18683
rect 73949 18717 73983 18733
rect 73949 18667 73983 18683
rect 1601 18381 1635 18397
rect 1601 18331 1635 18347
rect 73949 18381 73983 18397
rect 73949 18331 73983 18347
rect 1601 18045 1635 18061
rect 1601 17995 1635 18011
rect 73949 18045 73983 18061
rect 73949 17995 73983 18011
rect 1601 17709 1635 17725
rect 1601 17659 1635 17675
rect 73949 17709 73983 17725
rect 73949 17659 73983 17675
rect 1601 17373 1635 17389
rect 1601 17323 1635 17339
rect 73949 17373 73983 17389
rect 73949 17323 73983 17339
rect 1601 17037 1635 17053
rect 1601 16987 1635 17003
rect 73949 17037 73983 17053
rect 73949 16987 73983 17003
rect 1601 16701 1635 16717
rect 1601 16651 1635 16667
rect 73949 16701 73983 16717
rect 73949 16651 73983 16667
rect 1601 16365 1635 16381
rect 1601 16315 1635 16331
rect 73949 16365 73983 16381
rect 73949 16315 73983 16331
rect 1601 16029 1635 16045
rect 1601 15979 1635 15995
rect 73949 16029 73983 16045
rect 73949 15979 73983 15995
rect 1601 15693 1635 15709
rect 1601 15643 1635 15659
rect 73949 15693 73983 15709
rect 73949 15643 73983 15659
rect 1601 15357 1635 15373
rect 1601 15307 1635 15323
rect 73949 15357 73983 15373
rect 73949 15307 73983 15323
rect 1601 15021 1635 15037
rect 1601 14971 1635 14987
rect 73949 15021 73983 15037
rect 73949 14971 73983 14987
rect 1601 14685 1635 14701
rect 1601 14635 1635 14651
rect 73949 14685 73983 14701
rect 73949 14635 73983 14651
rect 1601 14349 1635 14365
rect 1601 14299 1635 14315
rect 73949 14349 73983 14365
rect 73949 14299 73983 14315
rect 1601 14013 1635 14029
rect 1601 13963 1635 13979
rect 73949 14013 73983 14029
rect 73949 13963 73983 13979
rect 1601 13677 1635 13693
rect 1601 13627 1635 13643
rect 73949 13677 73983 13693
rect 73949 13627 73983 13643
rect 1601 13341 1635 13357
rect 1601 13291 1635 13307
rect 73949 13341 73983 13357
rect 73949 13291 73983 13307
rect 1601 13005 1635 13021
rect 1601 12955 1635 12971
rect 73949 13005 73983 13021
rect 73949 12955 73983 12971
rect 1601 12669 1635 12685
rect 1601 12619 1635 12635
rect 73949 12669 73983 12685
rect 73949 12619 73983 12635
rect 1601 12333 1635 12349
rect 1601 12283 1635 12299
rect 73949 12333 73983 12349
rect 73949 12283 73983 12299
rect 1601 11997 1635 12013
rect 1601 11947 1635 11963
rect 73949 11997 73983 12013
rect 73949 11947 73983 11963
rect 1601 11661 1635 11677
rect 1601 11611 1635 11627
rect 73949 11661 73983 11677
rect 73949 11611 73983 11627
rect 1601 11325 1635 11341
rect 1601 11275 1635 11291
rect 73949 11325 73983 11341
rect 73949 11275 73983 11291
rect 1601 10989 1635 11005
rect 1601 10939 1635 10955
rect 73949 10989 73983 11005
rect 73949 10939 73983 10955
rect 1601 10653 1635 10669
rect 1601 10603 1635 10619
rect 73949 10653 73983 10669
rect 73949 10603 73983 10619
rect 1601 10317 1635 10333
rect 1601 10267 1635 10283
rect 73949 10317 73983 10333
rect 73949 10267 73983 10283
rect 1601 9981 1635 9997
rect 1601 9931 1635 9947
rect 73949 9981 73983 9997
rect 73949 9931 73983 9947
rect 1601 9645 1635 9661
rect 1601 9595 1635 9611
rect 73949 9645 73983 9661
rect 73949 9595 73983 9611
rect 1601 9309 1635 9325
rect 1601 9259 1635 9275
rect 73949 9309 73983 9325
rect 73949 9259 73983 9275
rect 1601 8973 1635 8989
rect 1601 8923 1635 8939
rect 73949 8973 73983 8989
rect 73949 8923 73983 8939
rect 1601 8637 1635 8653
rect 1601 8587 1635 8603
rect 73949 8637 73983 8653
rect 73949 8587 73983 8603
rect 1601 8301 1635 8317
rect 1601 8251 1635 8267
rect 73949 8301 73983 8317
rect 73949 8251 73983 8267
rect 1601 7965 1635 7981
rect 1601 7915 1635 7931
rect 73949 7965 73983 7981
rect 73949 7915 73983 7931
rect 1601 7629 1635 7645
rect 1601 7579 1635 7595
rect 73949 7629 73983 7645
rect 73949 7579 73983 7595
rect 1601 7293 1635 7309
rect 1601 7243 1635 7259
rect 73949 7293 73983 7309
rect 73949 7243 73983 7259
rect 1601 6957 1635 6973
rect 1601 6907 1635 6923
rect 73949 6957 73983 6973
rect 73949 6907 73983 6923
rect 1601 6621 1635 6637
rect 1601 6571 1635 6587
rect 73949 6621 73983 6637
rect 73949 6571 73983 6587
rect 1601 6285 1635 6301
rect 1601 6235 1635 6251
rect 73949 6285 73983 6301
rect 73949 6235 73983 6251
rect 1601 5949 1635 5965
rect 1601 5899 1635 5915
rect 73949 5949 73983 5965
rect 73949 5899 73983 5915
rect 1601 5613 1635 5629
rect 1601 5563 1635 5579
rect 73949 5613 73983 5629
rect 73949 5563 73983 5579
rect 1601 5277 1635 5293
rect 1601 5227 1635 5243
rect 73949 5277 73983 5293
rect 73949 5227 73983 5243
rect 1601 4941 1635 4957
rect 1601 4891 1635 4907
rect 73949 4941 73983 4957
rect 73949 4891 73983 4907
rect 1601 4605 1635 4621
rect 1601 4555 1635 4571
rect 73949 4605 73983 4621
rect 73949 4555 73983 4571
rect 1601 4269 1635 4285
rect 1601 4219 1635 4235
rect 73949 4269 73983 4285
rect 73949 4219 73983 4235
rect 1601 3933 1635 3949
rect 1601 3883 1635 3899
rect 73949 3933 73983 3949
rect 73949 3883 73983 3899
rect 1601 3597 1635 3613
rect 1601 3547 1635 3563
rect 73949 3597 73983 3613
rect 73949 3547 73983 3563
rect 1601 3261 1635 3277
rect 1601 3211 1635 3227
rect 73949 3261 73983 3277
rect 73949 3211 73983 3227
rect 1601 2925 1635 2941
rect 1601 2875 1635 2891
rect 73949 2925 73983 2941
rect 73949 2875 73983 2891
rect 1601 2589 1635 2605
rect 1601 2539 1635 2555
rect 73949 2589 73983 2605
rect 73949 2539 73983 2555
rect 1601 2253 1635 2269
rect 1601 2203 1635 2219
rect 73949 2253 73983 2269
rect 73949 2203 73983 2219
rect 1601 1917 1635 1933
rect 1601 1867 1635 1883
rect 73949 1917 73983 1933
rect 73949 1867 73983 1883
rect 1937 1581 1971 1597
rect 1937 1531 1971 1547
rect 2273 1581 2307 1597
rect 2273 1531 2307 1547
rect 2609 1581 2643 1597
rect 2609 1531 2643 1547
rect 2945 1581 2979 1597
rect 2945 1531 2979 1547
rect 3281 1581 3315 1597
rect 3281 1531 3315 1547
rect 3617 1581 3651 1597
rect 3617 1531 3651 1547
rect 3953 1581 3987 1597
rect 3953 1531 3987 1547
rect 4289 1581 4323 1597
rect 4289 1531 4323 1547
rect 4625 1581 4659 1597
rect 4625 1531 4659 1547
rect 4961 1581 4995 1597
rect 4961 1531 4995 1547
rect 5297 1581 5331 1597
rect 5297 1531 5331 1547
rect 5633 1581 5667 1597
rect 5633 1531 5667 1547
rect 5969 1581 6003 1597
rect 5969 1531 6003 1547
rect 6305 1581 6339 1597
rect 6305 1531 6339 1547
rect 6641 1581 6675 1597
rect 6641 1531 6675 1547
rect 6977 1581 7011 1597
rect 6977 1531 7011 1547
rect 7313 1581 7347 1597
rect 7313 1531 7347 1547
rect 7649 1581 7683 1597
rect 7649 1531 7683 1547
rect 7985 1581 8019 1597
rect 7985 1531 8019 1547
rect 8321 1581 8355 1597
rect 8321 1531 8355 1547
rect 8657 1581 8691 1597
rect 8657 1531 8691 1547
rect 8993 1581 9027 1597
rect 8993 1531 9027 1547
rect 9329 1581 9363 1597
rect 9329 1531 9363 1547
rect 9665 1581 9699 1597
rect 9665 1531 9699 1547
rect 10001 1581 10035 1597
rect 10001 1531 10035 1547
rect 10337 1581 10371 1597
rect 10337 1531 10371 1547
rect 10673 1581 10707 1597
rect 10673 1531 10707 1547
rect 11009 1581 11043 1597
rect 11009 1531 11043 1547
rect 11345 1581 11379 1597
rect 11345 1531 11379 1547
rect 11681 1581 11715 1597
rect 11681 1531 11715 1547
rect 12017 1581 12051 1597
rect 12017 1531 12051 1547
rect 12353 1581 12387 1597
rect 12353 1531 12387 1547
rect 12689 1581 12723 1597
rect 12689 1531 12723 1547
rect 13025 1581 13059 1597
rect 13025 1531 13059 1547
rect 13361 1581 13395 1597
rect 13361 1531 13395 1547
rect 13697 1581 13731 1597
rect 13697 1531 13731 1547
rect 14033 1581 14067 1597
rect 14033 1531 14067 1547
rect 14369 1581 14403 1597
rect 14369 1531 14403 1547
rect 14705 1581 14739 1597
rect 14705 1531 14739 1547
rect 15041 1581 15075 1597
rect 15041 1531 15075 1547
rect 15377 1581 15411 1597
rect 15377 1531 15411 1547
rect 15713 1581 15747 1597
rect 15713 1531 15747 1547
rect 16049 1581 16083 1597
rect 16049 1531 16083 1547
rect 16385 1581 16419 1597
rect 16385 1531 16419 1547
rect 16721 1581 16755 1597
rect 16721 1531 16755 1547
rect 17057 1581 17091 1597
rect 17057 1531 17091 1547
rect 17393 1581 17427 1597
rect 17393 1531 17427 1547
rect 17729 1581 17763 1597
rect 17729 1531 17763 1547
rect 18065 1581 18099 1597
rect 18065 1531 18099 1547
rect 18401 1581 18435 1597
rect 18401 1531 18435 1547
rect 18737 1581 18771 1597
rect 18737 1531 18771 1547
rect 19073 1581 19107 1597
rect 19073 1531 19107 1547
rect 19409 1581 19443 1597
rect 19409 1531 19443 1547
rect 19745 1581 19779 1597
rect 19745 1531 19779 1547
rect 20081 1581 20115 1597
rect 20081 1531 20115 1547
rect 20417 1581 20451 1597
rect 20417 1531 20451 1547
rect 20753 1581 20787 1597
rect 20753 1531 20787 1547
rect 21089 1581 21123 1597
rect 21089 1531 21123 1547
rect 21425 1581 21459 1597
rect 21425 1531 21459 1547
rect 21761 1581 21795 1597
rect 21761 1531 21795 1547
rect 22097 1581 22131 1597
rect 22097 1531 22131 1547
rect 22433 1581 22467 1597
rect 22433 1531 22467 1547
rect 22769 1581 22803 1597
rect 22769 1531 22803 1547
rect 23105 1581 23139 1597
rect 23105 1531 23139 1547
rect 23441 1581 23475 1597
rect 23441 1531 23475 1547
rect 23777 1581 23811 1597
rect 23777 1531 23811 1547
rect 24113 1581 24147 1597
rect 24113 1531 24147 1547
rect 24449 1581 24483 1597
rect 24449 1531 24483 1547
rect 24785 1581 24819 1597
rect 24785 1531 24819 1547
rect 25121 1581 25155 1597
rect 25121 1531 25155 1547
rect 25457 1581 25491 1597
rect 25457 1531 25491 1547
rect 25793 1581 25827 1597
rect 25793 1531 25827 1547
rect 26129 1581 26163 1597
rect 26129 1531 26163 1547
rect 26465 1581 26499 1597
rect 26465 1531 26499 1547
rect 26801 1581 26835 1597
rect 26801 1531 26835 1547
rect 27137 1581 27171 1597
rect 27137 1531 27171 1547
rect 27473 1581 27507 1597
rect 27473 1531 27507 1547
rect 27809 1581 27843 1597
rect 27809 1531 27843 1547
rect 28145 1581 28179 1597
rect 28145 1531 28179 1547
rect 28481 1581 28515 1597
rect 28481 1531 28515 1547
rect 28817 1581 28851 1597
rect 28817 1531 28851 1547
rect 29153 1581 29187 1597
rect 29153 1531 29187 1547
rect 29489 1581 29523 1597
rect 29489 1531 29523 1547
rect 29825 1581 29859 1597
rect 29825 1531 29859 1547
rect 30161 1581 30195 1597
rect 30161 1531 30195 1547
rect 30497 1581 30531 1597
rect 30497 1531 30531 1547
rect 30833 1581 30867 1597
rect 30833 1531 30867 1547
rect 31169 1581 31203 1597
rect 31169 1531 31203 1547
rect 31505 1581 31539 1597
rect 31505 1531 31539 1547
rect 31841 1581 31875 1597
rect 31841 1531 31875 1547
rect 32177 1581 32211 1597
rect 32177 1531 32211 1547
rect 32513 1581 32547 1597
rect 32513 1531 32547 1547
rect 32849 1581 32883 1597
rect 32849 1531 32883 1547
rect 33185 1581 33219 1597
rect 33185 1531 33219 1547
rect 33521 1581 33555 1597
rect 33521 1531 33555 1547
rect 33857 1581 33891 1597
rect 33857 1531 33891 1547
rect 34193 1581 34227 1597
rect 34193 1531 34227 1547
rect 34529 1581 34563 1597
rect 34529 1531 34563 1547
rect 34865 1581 34899 1597
rect 34865 1531 34899 1547
rect 35201 1581 35235 1597
rect 35201 1531 35235 1547
rect 35537 1581 35571 1597
rect 35537 1531 35571 1547
rect 35873 1581 35907 1597
rect 35873 1531 35907 1547
rect 36209 1581 36243 1597
rect 36209 1531 36243 1547
rect 36545 1581 36579 1597
rect 36545 1531 36579 1547
rect 36881 1581 36915 1597
rect 36881 1531 36915 1547
rect 37217 1581 37251 1597
rect 37217 1531 37251 1547
rect 37553 1581 37587 1597
rect 37553 1531 37587 1547
rect 37889 1581 37923 1597
rect 37889 1531 37923 1547
rect 38225 1581 38259 1597
rect 38225 1531 38259 1547
rect 38561 1581 38595 1597
rect 38561 1531 38595 1547
rect 38897 1581 38931 1597
rect 38897 1531 38931 1547
rect 39233 1581 39267 1597
rect 39233 1531 39267 1547
rect 39569 1581 39603 1597
rect 39569 1531 39603 1547
rect 39905 1581 39939 1597
rect 39905 1531 39939 1547
rect 40241 1581 40275 1597
rect 40241 1531 40275 1547
rect 40577 1581 40611 1597
rect 40577 1531 40611 1547
rect 40913 1581 40947 1597
rect 40913 1531 40947 1547
rect 41249 1581 41283 1597
rect 41249 1531 41283 1547
rect 41585 1581 41619 1597
rect 41585 1531 41619 1547
rect 41921 1581 41955 1597
rect 41921 1531 41955 1547
rect 42257 1581 42291 1597
rect 42257 1531 42291 1547
rect 42593 1581 42627 1597
rect 42593 1531 42627 1547
rect 42929 1581 42963 1597
rect 42929 1531 42963 1547
rect 43265 1581 43299 1597
rect 43265 1531 43299 1547
rect 43601 1581 43635 1597
rect 43601 1531 43635 1547
rect 43937 1581 43971 1597
rect 43937 1531 43971 1547
rect 44273 1581 44307 1597
rect 44273 1531 44307 1547
rect 44609 1581 44643 1597
rect 44609 1531 44643 1547
rect 44945 1581 44979 1597
rect 44945 1531 44979 1547
rect 45281 1581 45315 1597
rect 45281 1531 45315 1547
rect 45617 1581 45651 1597
rect 45617 1531 45651 1547
rect 45953 1581 45987 1597
rect 45953 1531 45987 1547
rect 46289 1581 46323 1597
rect 46289 1531 46323 1547
rect 46625 1581 46659 1597
rect 46625 1531 46659 1547
rect 46961 1581 46995 1597
rect 46961 1531 46995 1547
rect 47297 1581 47331 1597
rect 47297 1531 47331 1547
rect 47633 1581 47667 1597
rect 47633 1531 47667 1547
rect 47969 1581 48003 1597
rect 47969 1531 48003 1547
rect 48305 1581 48339 1597
rect 48305 1531 48339 1547
rect 48641 1581 48675 1597
rect 48641 1531 48675 1547
rect 48977 1581 49011 1597
rect 48977 1531 49011 1547
rect 49313 1581 49347 1597
rect 49313 1531 49347 1547
rect 49649 1581 49683 1597
rect 49649 1531 49683 1547
rect 49985 1581 50019 1597
rect 49985 1531 50019 1547
rect 50321 1581 50355 1597
rect 50321 1531 50355 1547
rect 50657 1581 50691 1597
rect 50657 1531 50691 1547
rect 50993 1581 51027 1597
rect 50993 1531 51027 1547
rect 51329 1581 51363 1597
rect 51329 1531 51363 1547
rect 51665 1581 51699 1597
rect 51665 1531 51699 1547
rect 52001 1581 52035 1597
rect 52001 1531 52035 1547
rect 52337 1581 52371 1597
rect 52337 1531 52371 1547
rect 52673 1581 52707 1597
rect 52673 1531 52707 1547
rect 53009 1581 53043 1597
rect 53009 1531 53043 1547
rect 53345 1581 53379 1597
rect 53345 1531 53379 1547
rect 53681 1581 53715 1597
rect 53681 1531 53715 1547
rect 54017 1581 54051 1597
rect 54017 1531 54051 1547
rect 54353 1581 54387 1597
rect 54353 1531 54387 1547
rect 54689 1581 54723 1597
rect 54689 1531 54723 1547
rect 55025 1581 55059 1597
rect 55025 1531 55059 1547
rect 55361 1581 55395 1597
rect 55361 1531 55395 1547
rect 55697 1581 55731 1597
rect 55697 1531 55731 1547
rect 56033 1581 56067 1597
rect 56033 1531 56067 1547
rect 56369 1581 56403 1597
rect 56369 1531 56403 1547
rect 56705 1581 56739 1597
rect 56705 1531 56739 1547
rect 57041 1581 57075 1597
rect 57041 1531 57075 1547
rect 57377 1581 57411 1597
rect 57377 1531 57411 1547
rect 57713 1581 57747 1597
rect 57713 1531 57747 1547
rect 58049 1581 58083 1597
rect 58049 1531 58083 1547
rect 58385 1581 58419 1597
rect 58385 1531 58419 1547
rect 58721 1581 58755 1597
rect 58721 1531 58755 1547
rect 59057 1581 59091 1597
rect 59057 1531 59091 1547
rect 59393 1581 59427 1597
rect 59393 1531 59427 1547
rect 59729 1581 59763 1597
rect 59729 1531 59763 1547
rect 60065 1581 60099 1597
rect 60065 1531 60099 1547
rect 60401 1581 60435 1597
rect 60401 1531 60435 1547
rect 60737 1581 60771 1597
rect 60737 1531 60771 1547
rect 61073 1581 61107 1597
rect 61073 1531 61107 1547
rect 61409 1581 61443 1597
rect 61409 1531 61443 1547
rect 61745 1581 61779 1597
rect 61745 1531 61779 1547
rect 62081 1581 62115 1597
rect 62081 1531 62115 1547
rect 62417 1581 62451 1597
rect 62417 1531 62451 1547
rect 62753 1581 62787 1597
rect 62753 1531 62787 1547
rect 63089 1581 63123 1597
rect 63089 1531 63123 1547
rect 63425 1581 63459 1597
rect 63425 1531 63459 1547
rect 63761 1581 63795 1597
rect 63761 1531 63795 1547
rect 64097 1581 64131 1597
rect 64097 1531 64131 1547
rect 64433 1581 64467 1597
rect 64433 1531 64467 1547
rect 64769 1581 64803 1597
rect 64769 1531 64803 1547
rect 65105 1581 65139 1597
rect 65105 1531 65139 1547
rect 65441 1581 65475 1597
rect 65441 1531 65475 1547
rect 65777 1581 65811 1597
rect 65777 1531 65811 1547
rect 66113 1581 66147 1597
rect 66113 1531 66147 1547
rect 66449 1581 66483 1597
rect 66449 1531 66483 1547
rect 66785 1581 66819 1597
rect 66785 1531 66819 1547
rect 67121 1581 67155 1597
rect 67121 1531 67155 1547
rect 67457 1581 67491 1597
rect 67457 1531 67491 1547
rect 67793 1581 67827 1597
rect 67793 1531 67827 1547
rect 68129 1581 68163 1597
rect 68129 1531 68163 1547
rect 68465 1581 68499 1597
rect 68465 1531 68499 1547
rect 68801 1581 68835 1597
rect 68801 1531 68835 1547
rect 69137 1581 69171 1597
rect 69137 1531 69171 1547
rect 69473 1581 69507 1597
rect 69473 1531 69507 1547
rect 69809 1581 69843 1597
rect 69809 1531 69843 1547
rect 70145 1581 70179 1597
rect 70145 1531 70179 1547
rect 70481 1581 70515 1597
rect 70481 1531 70515 1547
rect 70817 1581 70851 1597
rect 70817 1531 70851 1547
rect 71153 1581 71187 1597
rect 71153 1531 71187 1547
rect 71489 1581 71523 1597
rect 71489 1531 71523 1547
rect 71825 1581 71859 1597
rect 71825 1531 71859 1547
rect 72161 1581 72195 1597
rect 72161 1531 72195 1547
rect 72497 1581 72531 1597
rect 72497 1531 72531 1547
rect 72833 1581 72867 1597
rect 72833 1531 72867 1547
rect 73169 1581 73203 1597
rect 73169 1531 73203 1547
rect 73505 1581 73539 1597
rect 73505 1531 73539 1547
<< viali >>
rect 1937 36191 1971 36225
rect 2273 36191 2307 36225
rect 2609 36191 2643 36225
rect 2945 36191 2979 36225
rect 3281 36191 3315 36225
rect 3617 36191 3651 36225
rect 3953 36191 3987 36225
rect 4289 36191 4323 36225
rect 4625 36191 4659 36225
rect 4961 36191 4995 36225
rect 5297 36191 5331 36225
rect 5633 36191 5667 36225
rect 5969 36191 6003 36225
rect 6305 36191 6339 36225
rect 6641 36191 6675 36225
rect 6977 36191 7011 36225
rect 7313 36191 7347 36225
rect 7649 36191 7683 36225
rect 7985 36191 8019 36225
rect 8321 36191 8355 36225
rect 8657 36191 8691 36225
rect 8993 36191 9027 36225
rect 9329 36191 9363 36225
rect 9665 36191 9699 36225
rect 10001 36191 10035 36225
rect 10337 36191 10371 36225
rect 10673 36191 10707 36225
rect 11009 36191 11043 36225
rect 11345 36191 11379 36225
rect 11681 36191 11715 36225
rect 12017 36191 12051 36225
rect 12353 36191 12387 36225
rect 12689 36191 12723 36225
rect 13025 36191 13059 36225
rect 13361 36191 13395 36225
rect 13697 36191 13731 36225
rect 14033 36191 14067 36225
rect 14369 36191 14403 36225
rect 14705 36191 14739 36225
rect 15041 36191 15075 36225
rect 15377 36191 15411 36225
rect 15713 36191 15747 36225
rect 16049 36191 16083 36225
rect 16385 36191 16419 36225
rect 16721 36191 16755 36225
rect 17057 36191 17091 36225
rect 17393 36191 17427 36225
rect 17729 36191 17763 36225
rect 18065 36191 18099 36225
rect 18401 36191 18435 36225
rect 18737 36191 18771 36225
rect 19073 36191 19107 36225
rect 19409 36191 19443 36225
rect 19745 36191 19779 36225
rect 20081 36191 20115 36225
rect 20417 36191 20451 36225
rect 20753 36191 20787 36225
rect 21089 36191 21123 36225
rect 21425 36191 21459 36225
rect 21761 36191 21795 36225
rect 22097 36191 22131 36225
rect 22433 36191 22467 36225
rect 22769 36191 22803 36225
rect 23105 36191 23139 36225
rect 23441 36191 23475 36225
rect 23777 36191 23811 36225
rect 24113 36191 24147 36225
rect 24449 36191 24483 36225
rect 24785 36191 24819 36225
rect 25121 36191 25155 36225
rect 25457 36191 25491 36225
rect 25793 36191 25827 36225
rect 26129 36191 26163 36225
rect 26465 36191 26499 36225
rect 26801 36191 26835 36225
rect 27137 36191 27171 36225
rect 27473 36191 27507 36225
rect 27809 36191 27843 36225
rect 28145 36191 28179 36225
rect 28481 36191 28515 36225
rect 28817 36191 28851 36225
rect 29153 36191 29187 36225
rect 29489 36191 29523 36225
rect 29825 36191 29859 36225
rect 30161 36191 30195 36225
rect 30497 36191 30531 36225
rect 30833 36191 30867 36225
rect 31169 36191 31203 36225
rect 31505 36191 31539 36225
rect 31841 36191 31875 36225
rect 32177 36191 32211 36225
rect 32513 36191 32547 36225
rect 32849 36191 32883 36225
rect 33185 36191 33219 36225
rect 33521 36191 33555 36225
rect 33857 36191 33891 36225
rect 34193 36191 34227 36225
rect 34529 36191 34563 36225
rect 34865 36191 34899 36225
rect 35201 36191 35235 36225
rect 35537 36191 35571 36225
rect 35873 36191 35907 36225
rect 36209 36191 36243 36225
rect 36545 36191 36579 36225
rect 36881 36191 36915 36225
rect 37217 36191 37251 36225
rect 37553 36191 37587 36225
rect 37889 36191 37923 36225
rect 38225 36191 38259 36225
rect 38561 36191 38595 36225
rect 38897 36191 38931 36225
rect 39233 36191 39267 36225
rect 39569 36191 39603 36225
rect 39905 36191 39939 36225
rect 40241 36191 40275 36225
rect 40577 36191 40611 36225
rect 40913 36191 40947 36225
rect 41249 36191 41283 36225
rect 41585 36191 41619 36225
rect 41921 36191 41955 36225
rect 42257 36191 42291 36225
rect 42593 36191 42627 36225
rect 42929 36191 42963 36225
rect 43265 36191 43299 36225
rect 43601 36191 43635 36225
rect 43937 36191 43971 36225
rect 44273 36191 44307 36225
rect 44609 36191 44643 36225
rect 44945 36191 44979 36225
rect 45281 36191 45315 36225
rect 45617 36191 45651 36225
rect 45953 36191 45987 36225
rect 46289 36191 46323 36225
rect 46625 36191 46659 36225
rect 46961 36191 46995 36225
rect 47297 36191 47331 36225
rect 47633 36191 47667 36225
rect 47969 36191 48003 36225
rect 48305 36191 48339 36225
rect 48641 36191 48675 36225
rect 48977 36191 49011 36225
rect 49313 36191 49347 36225
rect 49649 36191 49683 36225
rect 49985 36191 50019 36225
rect 50321 36191 50355 36225
rect 50657 36191 50691 36225
rect 50993 36191 51027 36225
rect 51329 36191 51363 36225
rect 51665 36191 51699 36225
rect 52001 36191 52035 36225
rect 52337 36191 52371 36225
rect 52673 36191 52707 36225
rect 53009 36191 53043 36225
rect 53345 36191 53379 36225
rect 53681 36191 53715 36225
rect 54017 36191 54051 36225
rect 54353 36191 54387 36225
rect 54689 36191 54723 36225
rect 55025 36191 55059 36225
rect 55361 36191 55395 36225
rect 55697 36191 55731 36225
rect 56033 36191 56067 36225
rect 56369 36191 56403 36225
rect 56705 36191 56739 36225
rect 57041 36191 57075 36225
rect 57377 36191 57411 36225
rect 57713 36191 57747 36225
rect 58049 36191 58083 36225
rect 58385 36191 58419 36225
rect 58721 36191 58755 36225
rect 59057 36191 59091 36225
rect 59393 36191 59427 36225
rect 59729 36191 59763 36225
rect 60065 36191 60099 36225
rect 60401 36191 60435 36225
rect 60737 36191 60771 36225
rect 61073 36191 61107 36225
rect 61409 36191 61443 36225
rect 61745 36191 61779 36225
rect 62081 36191 62115 36225
rect 62417 36191 62451 36225
rect 62753 36191 62787 36225
rect 63089 36191 63123 36225
rect 63425 36191 63459 36225
rect 63761 36191 63795 36225
rect 64097 36191 64131 36225
rect 64433 36191 64467 36225
rect 64769 36191 64803 36225
rect 65105 36191 65139 36225
rect 65441 36191 65475 36225
rect 65777 36191 65811 36225
rect 66113 36191 66147 36225
rect 66449 36191 66483 36225
rect 66785 36191 66819 36225
rect 67121 36191 67155 36225
rect 67457 36191 67491 36225
rect 67793 36191 67827 36225
rect 68129 36191 68163 36225
rect 68465 36191 68499 36225
rect 68801 36191 68835 36225
rect 69137 36191 69171 36225
rect 69473 36191 69507 36225
rect 69809 36191 69843 36225
rect 70145 36191 70179 36225
rect 70481 36191 70515 36225
rect 70817 36191 70851 36225
rect 71153 36191 71187 36225
rect 71489 36191 71523 36225
rect 71825 36191 71859 36225
rect 72161 36191 72195 36225
rect 72497 36191 72531 36225
rect 72833 36191 72867 36225
rect 73169 36191 73203 36225
rect 73505 36191 73539 36225
rect 1601 35819 1635 35853
rect 73949 35819 73983 35853
rect 1601 35483 1635 35517
rect 73949 35483 73983 35517
rect 1601 35147 1635 35181
rect 73949 35147 73983 35181
rect 1601 34811 1635 34845
rect 73949 34811 73983 34845
rect 1601 34475 1635 34509
rect 73949 34475 73983 34509
rect 1601 34139 1635 34173
rect 73949 34139 73983 34173
rect 1601 33803 1635 33837
rect 73949 33803 73983 33837
rect 1601 33467 1635 33501
rect 73949 33467 73983 33501
rect 1601 33131 1635 33165
rect 73949 33131 73983 33165
rect 1601 32795 1635 32829
rect 73949 32795 73983 32829
rect 1601 32459 1635 32493
rect 73949 32459 73983 32493
rect 1601 32123 1635 32157
rect 73949 32123 73983 32157
rect 1601 31787 1635 31821
rect 73949 31787 73983 31821
rect 1601 31451 1635 31485
rect 73949 31451 73983 31485
rect 1601 31115 1635 31149
rect 73949 31115 73983 31149
rect 1601 30779 1635 30813
rect 73949 30779 73983 30813
rect 1601 30443 1635 30477
rect 73949 30443 73983 30477
rect 1601 30107 1635 30141
rect 73949 30107 73983 30141
rect 1601 29771 1635 29805
rect 73949 29771 73983 29805
rect 1601 29435 1635 29469
rect 73949 29435 73983 29469
rect 1601 29099 1635 29133
rect 73949 29099 73983 29133
rect 1601 28763 1635 28797
rect 73949 28763 73983 28797
rect 1601 28427 1635 28461
rect 73949 28427 73983 28461
rect 1601 28091 1635 28125
rect 73949 28091 73983 28125
rect 1601 27755 1635 27789
rect 73949 27755 73983 27789
rect 1601 27419 1635 27453
rect 73949 27419 73983 27453
rect 1601 27083 1635 27117
rect 73949 27083 73983 27117
rect 1601 26747 1635 26781
rect 73949 26747 73983 26781
rect 1601 26411 1635 26445
rect 73949 26411 73983 26445
rect 1601 26075 1635 26109
rect 73949 26075 73983 26109
rect 1601 25739 1635 25773
rect 73949 25739 73983 25773
rect 1601 25403 1635 25437
rect 73949 25403 73983 25437
rect 1601 25067 1635 25101
rect 73949 25067 73983 25101
rect 1601 24731 1635 24765
rect 73949 24731 73983 24765
rect 1601 24395 1635 24429
rect 73949 24395 73983 24429
rect 1601 24059 1635 24093
rect 73949 24059 73983 24093
rect 1601 23723 1635 23757
rect 73949 23723 73983 23757
rect 1601 23387 1635 23421
rect 73949 23387 73983 23421
rect 1601 23051 1635 23085
rect 73949 23051 73983 23085
rect 1601 22715 1635 22749
rect 73949 22715 73983 22749
rect 1601 22379 1635 22413
rect 73949 22379 73983 22413
rect 1601 22043 1635 22077
rect 73949 22043 73983 22077
rect 1601 21707 1635 21741
rect 73949 21707 73983 21741
rect 1601 21371 1635 21405
rect 73949 21371 73983 21405
rect 1601 21035 1635 21069
rect 73949 21035 73983 21069
rect 1601 20699 1635 20733
rect 73949 20699 73983 20733
rect 1601 20363 1635 20397
rect 73949 20363 73983 20397
rect 1601 20027 1635 20061
rect 73949 20027 73983 20061
rect 1601 19691 1635 19725
rect 73949 19691 73983 19725
rect 1601 19355 1635 19389
rect 73949 19355 73983 19389
rect 1601 19019 1635 19053
rect 73949 19019 73983 19053
rect 1601 18683 1635 18717
rect 73949 18683 73983 18717
rect 1601 18347 1635 18381
rect 73949 18347 73983 18381
rect 1601 18011 1635 18045
rect 73949 18011 73983 18045
rect 1601 17675 1635 17709
rect 73949 17675 73983 17709
rect 1601 17339 1635 17373
rect 73949 17339 73983 17373
rect 1601 17003 1635 17037
rect 73949 17003 73983 17037
rect 1601 16667 1635 16701
rect 73949 16667 73983 16701
rect 1601 16331 1635 16365
rect 73949 16331 73983 16365
rect 1601 15995 1635 16029
rect 73949 15995 73983 16029
rect 1601 15659 1635 15693
rect 73949 15659 73983 15693
rect 1601 15323 1635 15357
rect 73949 15323 73983 15357
rect 1601 14987 1635 15021
rect 73949 14987 73983 15021
rect 1601 14651 1635 14685
rect 73949 14651 73983 14685
rect 1601 14315 1635 14349
rect 73949 14315 73983 14349
rect 1601 13979 1635 14013
rect 73949 13979 73983 14013
rect 1601 13643 1635 13677
rect 73949 13643 73983 13677
rect 1601 13307 1635 13341
rect 73949 13307 73983 13341
rect 1601 12971 1635 13005
rect 73949 12971 73983 13005
rect 1601 12635 1635 12669
rect 73949 12635 73983 12669
rect 1601 12299 1635 12333
rect 73949 12299 73983 12333
rect 1601 11963 1635 11997
rect 73949 11963 73983 11997
rect 1601 11627 1635 11661
rect 73949 11627 73983 11661
rect 1601 11291 1635 11325
rect 73949 11291 73983 11325
rect 1601 10955 1635 10989
rect 73949 10955 73983 10989
rect 1601 10619 1635 10653
rect 73949 10619 73983 10653
rect 1601 10283 1635 10317
rect 73949 10283 73983 10317
rect 1601 9947 1635 9981
rect 73949 9947 73983 9981
rect 1601 9611 1635 9645
rect 73949 9611 73983 9645
rect 1601 9275 1635 9309
rect 73949 9275 73983 9309
rect 1601 8939 1635 8973
rect 73949 8939 73983 8973
rect 1601 8603 1635 8637
rect 73949 8603 73983 8637
rect 1601 8267 1635 8301
rect 73949 8267 73983 8301
rect 1601 7931 1635 7965
rect 73949 7931 73983 7965
rect 1601 7595 1635 7629
rect 73949 7595 73983 7629
rect 1601 7259 1635 7293
rect 73949 7259 73983 7293
rect 1601 6923 1635 6957
rect 73949 6923 73983 6957
rect 1601 6587 1635 6621
rect 73949 6587 73983 6621
rect 1601 6251 1635 6285
rect 73949 6251 73983 6285
rect 1601 5915 1635 5949
rect 73949 5915 73983 5949
rect 1601 5579 1635 5613
rect 73949 5579 73983 5613
rect 1601 5243 1635 5277
rect 73949 5243 73983 5277
rect 1601 4907 1635 4941
rect 73949 4907 73983 4941
rect 1601 4571 1635 4605
rect 73949 4571 73983 4605
rect 1601 4235 1635 4269
rect 73949 4235 73983 4269
rect 1601 3899 1635 3933
rect 73949 3899 73983 3933
rect 1601 3563 1635 3597
rect 73949 3563 73983 3597
rect 1601 3227 1635 3261
rect 73949 3227 73983 3261
rect 1601 2891 1635 2925
rect 73949 2891 73983 2925
rect 1601 2555 1635 2589
rect 73949 2555 73983 2589
rect 1601 2219 1635 2253
rect 73949 2219 73983 2253
rect 1601 1883 1635 1917
rect 73949 1883 73983 1917
rect 1937 1547 1971 1581
rect 2273 1547 2307 1581
rect 2609 1547 2643 1581
rect 2945 1547 2979 1581
rect 3281 1547 3315 1581
rect 3617 1547 3651 1581
rect 3953 1547 3987 1581
rect 4289 1547 4323 1581
rect 4625 1547 4659 1581
rect 4961 1547 4995 1581
rect 5297 1547 5331 1581
rect 5633 1547 5667 1581
rect 5969 1547 6003 1581
rect 6305 1547 6339 1581
rect 6641 1547 6675 1581
rect 6977 1547 7011 1581
rect 7313 1547 7347 1581
rect 7649 1547 7683 1581
rect 7985 1547 8019 1581
rect 8321 1547 8355 1581
rect 8657 1547 8691 1581
rect 8993 1547 9027 1581
rect 9329 1547 9363 1581
rect 9665 1547 9699 1581
rect 10001 1547 10035 1581
rect 10337 1547 10371 1581
rect 10673 1547 10707 1581
rect 11009 1547 11043 1581
rect 11345 1547 11379 1581
rect 11681 1547 11715 1581
rect 12017 1547 12051 1581
rect 12353 1547 12387 1581
rect 12689 1547 12723 1581
rect 13025 1547 13059 1581
rect 13361 1547 13395 1581
rect 13697 1547 13731 1581
rect 14033 1547 14067 1581
rect 14369 1547 14403 1581
rect 14705 1547 14739 1581
rect 15041 1547 15075 1581
rect 15377 1547 15411 1581
rect 15713 1547 15747 1581
rect 16049 1547 16083 1581
rect 16385 1547 16419 1581
rect 16721 1547 16755 1581
rect 17057 1547 17091 1581
rect 17393 1547 17427 1581
rect 17729 1547 17763 1581
rect 18065 1547 18099 1581
rect 18401 1547 18435 1581
rect 18737 1547 18771 1581
rect 19073 1547 19107 1581
rect 19409 1547 19443 1581
rect 19745 1547 19779 1581
rect 20081 1547 20115 1581
rect 20417 1547 20451 1581
rect 20753 1547 20787 1581
rect 21089 1547 21123 1581
rect 21425 1547 21459 1581
rect 21761 1547 21795 1581
rect 22097 1547 22131 1581
rect 22433 1547 22467 1581
rect 22769 1547 22803 1581
rect 23105 1547 23139 1581
rect 23441 1547 23475 1581
rect 23777 1547 23811 1581
rect 24113 1547 24147 1581
rect 24449 1547 24483 1581
rect 24785 1547 24819 1581
rect 25121 1547 25155 1581
rect 25457 1547 25491 1581
rect 25793 1547 25827 1581
rect 26129 1547 26163 1581
rect 26465 1547 26499 1581
rect 26801 1547 26835 1581
rect 27137 1547 27171 1581
rect 27473 1547 27507 1581
rect 27809 1547 27843 1581
rect 28145 1547 28179 1581
rect 28481 1547 28515 1581
rect 28817 1547 28851 1581
rect 29153 1547 29187 1581
rect 29489 1547 29523 1581
rect 29825 1547 29859 1581
rect 30161 1547 30195 1581
rect 30497 1547 30531 1581
rect 30833 1547 30867 1581
rect 31169 1547 31203 1581
rect 31505 1547 31539 1581
rect 31841 1547 31875 1581
rect 32177 1547 32211 1581
rect 32513 1547 32547 1581
rect 32849 1547 32883 1581
rect 33185 1547 33219 1581
rect 33521 1547 33555 1581
rect 33857 1547 33891 1581
rect 34193 1547 34227 1581
rect 34529 1547 34563 1581
rect 34865 1547 34899 1581
rect 35201 1547 35235 1581
rect 35537 1547 35571 1581
rect 35873 1547 35907 1581
rect 36209 1547 36243 1581
rect 36545 1547 36579 1581
rect 36881 1547 36915 1581
rect 37217 1547 37251 1581
rect 37553 1547 37587 1581
rect 37889 1547 37923 1581
rect 38225 1547 38259 1581
rect 38561 1547 38595 1581
rect 38897 1547 38931 1581
rect 39233 1547 39267 1581
rect 39569 1547 39603 1581
rect 39905 1547 39939 1581
rect 40241 1547 40275 1581
rect 40577 1547 40611 1581
rect 40913 1547 40947 1581
rect 41249 1547 41283 1581
rect 41585 1547 41619 1581
rect 41921 1547 41955 1581
rect 42257 1547 42291 1581
rect 42593 1547 42627 1581
rect 42929 1547 42963 1581
rect 43265 1547 43299 1581
rect 43601 1547 43635 1581
rect 43937 1547 43971 1581
rect 44273 1547 44307 1581
rect 44609 1547 44643 1581
rect 44945 1547 44979 1581
rect 45281 1547 45315 1581
rect 45617 1547 45651 1581
rect 45953 1547 45987 1581
rect 46289 1547 46323 1581
rect 46625 1547 46659 1581
rect 46961 1547 46995 1581
rect 47297 1547 47331 1581
rect 47633 1547 47667 1581
rect 47969 1547 48003 1581
rect 48305 1547 48339 1581
rect 48641 1547 48675 1581
rect 48977 1547 49011 1581
rect 49313 1547 49347 1581
rect 49649 1547 49683 1581
rect 49985 1547 50019 1581
rect 50321 1547 50355 1581
rect 50657 1547 50691 1581
rect 50993 1547 51027 1581
rect 51329 1547 51363 1581
rect 51665 1547 51699 1581
rect 52001 1547 52035 1581
rect 52337 1547 52371 1581
rect 52673 1547 52707 1581
rect 53009 1547 53043 1581
rect 53345 1547 53379 1581
rect 53681 1547 53715 1581
rect 54017 1547 54051 1581
rect 54353 1547 54387 1581
rect 54689 1547 54723 1581
rect 55025 1547 55059 1581
rect 55361 1547 55395 1581
rect 55697 1547 55731 1581
rect 56033 1547 56067 1581
rect 56369 1547 56403 1581
rect 56705 1547 56739 1581
rect 57041 1547 57075 1581
rect 57377 1547 57411 1581
rect 57713 1547 57747 1581
rect 58049 1547 58083 1581
rect 58385 1547 58419 1581
rect 58721 1547 58755 1581
rect 59057 1547 59091 1581
rect 59393 1547 59427 1581
rect 59729 1547 59763 1581
rect 60065 1547 60099 1581
rect 60401 1547 60435 1581
rect 60737 1547 60771 1581
rect 61073 1547 61107 1581
rect 61409 1547 61443 1581
rect 61745 1547 61779 1581
rect 62081 1547 62115 1581
rect 62417 1547 62451 1581
rect 62753 1547 62787 1581
rect 63089 1547 63123 1581
rect 63425 1547 63459 1581
rect 63761 1547 63795 1581
rect 64097 1547 64131 1581
rect 64433 1547 64467 1581
rect 64769 1547 64803 1581
rect 65105 1547 65139 1581
rect 65441 1547 65475 1581
rect 65777 1547 65811 1581
rect 66113 1547 66147 1581
rect 66449 1547 66483 1581
rect 66785 1547 66819 1581
rect 67121 1547 67155 1581
rect 67457 1547 67491 1581
rect 67793 1547 67827 1581
rect 68129 1547 68163 1581
rect 68465 1547 68499 1581
rect 68801 1547 68835 1581
rect 69137 1547 69171 1581
rect 69473 1547 69507 1581
rect 69809 1547 69843 1581
rect 70145 1547 70179 1581
rect 70481 1547 70515 1581
rect 70817 1547 70851 1581
rect 71153 1547 71187 1581
rect 71489 1547 71523 1581
rect 71825 1547 71859 1581
rect 72161 1547 72195 1581
rect 72497 1547 72531 1581
rect 72833 1547 72867 1581
rect 73169 1547 73203 1581
rect 73505 1547 73539 1581
<< metal1 >>
rect 1506 36234 74078 36320
rect 1506 36182 1928 36234
rect 1980 36225 3608 36234
rect 3660 36225 5288 36234
rect 5340 36225 6968 36234
rect 7020 36225 8648 36234
rect 8700 36225 10328 36234
rect 10380 36225 12008 36234
rect 12060 36225 13688 36234
rect 13740 36225 15368 36234
rect 15420 36225 17048 36234
rect 17100 36225 18728 36234
rect 18780 36225 20408 36234
rect 20460 36225 22088 36234
rect 22140 36225 23768 36234
rect 23820 36225 25448 36234
rect 25500 36225 27128 36234
rect 27180 36225 28808 36234
rect 28860 36225 30488 36234
rect 30540 36225 32168 36234
rect 32220 36225 33848 36234
rect 33900 36225 35528 36234
rect 35580 36225 37208 36234
rect 37260 36225 38888 36234
rect 38940 36225 40568 36234
rect 40620 36225 42248 36234
rect 42300 36225 43928 36234
rect 43980 36225 45608 36234
rect 45660 36225 47288 36234
rect 47340 36225 48968 36234
rect 49020 36225 50648 36234
rect 50700 36225 52328 36234
rect 52380 36225 54008 36234
rect 54060 36225 55688 36234
rect 55740 36225 57368 36234
rect 57420 36225 59048 36234
rect 59100 36225 60728 36234
rect 60780 36225 62408 36234
rect 62460 36225 64088 36234
rect 64140 36225 65768 36234
rect 65820 36225 67448 36234
rect 67500 36225 69128 36234
rect 69180 36225 70808 36234
rect 70860 36225 72488 36234
rect 72540 36225 74078 36234
rect 1980 36191 2273 36225
rect 2307 36191 2609 36225
rect 2643 36191 2945 36225
rect 2979 36191 3281 36225
rect 3315 36191 3608 36225
rect 3660 36191 3953 36225
rect 3987 36191 4289 36225
rect 4323 36191 4625 36225
rect 4659 36191 4961 36225
rect 4995 36191 5288 36225
rect 5340 36191 5633 36225
rect 5667 36191 5969 36225
rect 6003 36191 6305 36225
rect 6339 36191 6641 36225
rect 6675 36191 6968 36225
rect 7020 36191 7313 36225
rect 7347 36191 7649 36225
rect 7683 36191 7985 36225
rect 8019 36191 8321 36225
rect 8355 36191 8648 36225
rect 8700 36191 8993 36225
rect 9027 36191 9329 36225
rect 9363 36191 9665 36225
rect 9699 36191 10001 36225
rect 10035 36191 10328 36225
rect 10380 36191 10673 36225
rect 10707 36191 11009 36225
rect 11043 36191 11345 36225
rect 11379 36191 11681 36225
rect 11715 36191 12008 36225
rect 12060 36191 12353 36225
rect 12387 36191 12689 36225
rect 12723 36191 13025 36225
rect 13059 36191 13361 36225
rect 13395 36191 13688 36225
rect 13740 36191 14033 36225
rect 14067 36191 14369 36225
rect 14403 36191 14705 36225
rect 14739 36191 15041 36225
rect 15075 36191 15368 36225
rect 15420 36191 15713 36225
rect 15747 36191 16049 36225
rect 16083 36191 16385 36225
rect 16419 36191 16721 36225
rect 16755 36191 17048 36225
rect 17100 36191 17393 36225
rect 17427 36191 17729 36225
rect 17763 36191 18065 36225
rect 18099 36191 18401 36225
rect 18435 36191 18728 36225
rect 18780 36191 19073 36225
rect 19107 36191 19409 36225
rect 19443 36191 19745 36225
rect 19779 36191 20081 36225
rect 20115 36191 20408 36225
rect 20460 36191 20753 36225
rect 20787 36191 21089 36225
rect 21123 36191 21425 36225
rect 21459 36191 21761 36225
rect 21795 36191 22088 36225
rect 22140 36191 22433 36225
rect 22467 36191 22769 36225
rect 22803 36191 23105 36225
rect 23139 36191 23441 36225
rect 23475 36191 23768 36225
rect 23820 36191 24113 36225
rect 24147 36191 24449 36225
rect 24483 36191 24785 36225
rect 24819 36191 25121 36225
rect 25155 36191 25448 36225
rect 25500 36191 25793 36225
rect 25827 36191 26129 36225
rect 26163 36191 26465 36225
rect 26499 36191 26801 36225
rect 26835 36191 27128 36225
rect 27180 36191 27473 36225
rect 27507 36191 27809 36225
rect 27843 36191 28145 36225
rect 28179 36191 28481 36225
rect 28515 36191 28808 36225
rect 28860 36191 29153 36225
rect 29187 36191 29489 36225
rect 29523 36191 29825 36225
rect 29859 36191 30161 36225
rect 30195 36191 30488 36225
rect 30540 36191 30833 36225
rect 30867 36191 31169 36225
rect 31203 36191 31505 36225
rect 31539 36191 31841 36225
rect 31875 36191 32168 36225
rect 32220 36191 32513 36225
rect 32547 36191 32849 36225
rect 32883 36191 33185 36225
rect 33219 36191 33521 36225
rect 33555 36191 33848 36225
rect 33900 36191 34193 36225
rect 34227 36191 34529 36225
rect 34563 36191 34865 36225
rect 34899 36191 35201 36225
rect 35235 36191 35528 36225
rect 35580 36191 35873 36225
rect 35907 36191 36209 36225
rect 36243 36191 36545 36225
rect 36579 36191 36881 36225
rect 36915 36191 37208 36225
rect 37260 36191 37553 36225
rect 37587 36191 37889 36225
rect 37923 36191 38225 36225
rect 38259 36191 38561 36225
rect 38595 36191 38888 36225
rect 38940 36191 39233 36225
rect 39267 36191 39569 36225
rect 39603 36191 39905 36225
rect 39939 36191 40241 36225
rect 40275 36191 40568 36225
rect 40620 36191 40913 36225
rect 40947 36191 41249 36225
rect 41283 36191 41585 36225
rect 41619 36191 41921 36225
rect 41955 36191 42248 36225
rect 42300 36191 42593 36225
rect 42627 36191 42929 36225
rect 42963 36191 43265 36225
rect 43299 36191 43601 36225
rect 43635 36191 43928 36225
rect 43980 36191 44273 36225
rect 44307 36191 44609 36225
rect 44643 36191 44945 36225
rect 44979 36191 45281 36225
rect 45315 36191 45608 36225
rect 45660 36191 45953 36225
rect 45987 36191 46289 36225
rect 46323 36191 46625 36225
rect 46659 36191 46961 36225
rect 46995 36191 47288 36225
rect 47340 36191 47633 36225
rect 47667 36191 47969 36225
rect 48003 36191 48305 36225
rect 48339 36191 48641 36225
rect 48675 36191 48968 36225
rect 49020 36191 49313 36225
rect 49347 36191 49649 36225
rect 49683 36191 49985 36225
rect 50019 36191 50321 36225
rect 50355 36191 50648 36225
rect 50700 36191 50993 36225
rect 51027 36191 51329 36225
rect 51363 36191 51665 36225
rect 51699 36191 52001 36225
rect 52035 36191 52328 36225
rect 52380 36191 52673 36225
rect 52707 36191 53009 36225
rect 53043 36191 53345 36225
rect 53379 36191 53681 36225
rect 53715 36191 54008 36225
rect 54060 36191 54353 36225
rect 54387 36191 54689 36225
rect 54723 36191 55025 36225
rect 55059 36191 55361 36225
rect 55395 36191 55688 36225
rect 55740 36191 56033 36225
rect 56067 36191 56369 36225
rect 56403 36191 56705 36225
rect 56739 36191 57041 36225
rect 57075 36191 57368 36225
rect 57420 36191 57713 36225
rect 57747 36191 58049 36225
rect 58083 36191 58385 36225
rect 58419 36191 58721 36225
rect 58755 36191 59048 36225
rect 59100 36191 59393 36225
rect 59427 36191 59729 36225
rect 59763 36191 60065 36225
rect 60099 36191 60401 36225
rect 60435 36191 60728 36225
rect 60780 36191 61073 36225
rect 61107 36191 61409 36225
rect 61443 36191 61745 36225
rect 61779 36191 62081 36225
rect 62115 36191 62408 36225
rect 62460 36191 62753 36225
rect 62787 36191 63089 36225
rect 63123 36191 63425 36225
rect 63459 36191 63761 36225
rect 63795 36191 64088 36225
rect 64140 36191 64433 36225
rect 64467 36191 64769 36225
rect 64803 36191 65105 36225
rect 65139 36191 65441 36225
rect 65475 36191 65768 36225
rect 65820 36191 66113 36225
rect 66147 36191 66449 36225
rect 66483 36191 66785 36225
rect 66819 36191 67121 36225
rect 67155 36191 67448 36225
rect 67500 36191 67793 36225
rect 67827 36191 68129 36225
rect 68163 36191 68465 36225
rect 68499 36191 68801 36225
rect 68835 36191 69128 36225
rect 69180 36191 69473 36225
rect 69507 36191 69809 36225
rect 69843 36191 70145 36225
rect 70179 36191 70481 36225
rect 70515 36191 70808 36225
rect 70860 36191 71153 36225
rect 71187 36191 71489 36225
rect 71523 36191 71825 36225
rect 71859 36191 72161 36225
rect 72195 36191 72488 36225
rect 72540 36191 72833 36225
rect 72867 36191 73169 36225
rect 73203 36191 73505 36225
rect 73539 36191 74078 36225
rect 1980 36182 3608 36191
rect 3660 36182 5288 36191
rect 5340 36182 6968 36191
rect 7020 36182 8648 36191
rect 8700 36182 10328 36191
rect 10380 36182 12008 36191
rect 12060 36182 13688 36191
rect 13740 36182 15368 36191
rect 15420 36182 17048 36191
rect 17100 36182 18728 36191
rect 18780 36182 20408 36191
rect 20460 36182 22088 36191
rect 22140 36182 23768 36191
rect 23820 36182 25448 36191
rect 25500 36182 27128 36191
rect 27180 36182 28808 36191
rect 28860 36182 30488 36191
rect 30540 36182 32168 36191
rect 32220 36182 33848 36191
rect 33900 36182 35528 36191
rect 35580 36182 37208 36191
rect 37260 36182 38888 36191
rect 38940 36182 40568 36191
rect 40620 36182 42248 36191
rect 42300 36182 43928 36191
rect 43980 36182 45608 36191
rect 45660 36182 47288 36191
rect 47340 36182 48968 36191
rect 49020 36182 50648 36191
rect 50700 36182 52328 36191
rect 52380 36182 54008 36191
rect 54060 36182 55688 36191
rect 55740 36182 57368 36191
rect 57420 36182 59048 36191
rect 59100 36182 60728 36191
rect 60780 36182 62408 36191
rect 62460 36182 64088 36191
rect 64140 36182 65768 36191
rect 65820 36182 67448 36191
rect 67500 36182 69128 36191
rect 69180 36182 70808 36191
rect 70860 36182 72488 36191
rect 72540 36182 74078 36191
rect 1506 36096 74078 36182
rect 1589 35851 1592 35859
rect 1563 35821 1592 35851
rect 1589 35813 1592 35821
rect 1644 35851 1647 35859
rect 73937 35851 73940 35859
rect 1644 35821 1674 35851
rect 73911 35821 73940 35851
rect 1644 35813 1647 35821
rect 73937 35813 73940 35821
rect 73992 35851 73995 35859
rect 73992 35821 74022 35851
rect 73992 35813 73995 35821
rect 1589 35515 1592 35523
rect 1563 35485 1592 35515
rect 1589 35477 1592 35485
rect 1644 35515 1647 35523
rect 73937 35515 73940 35523
rect 1644 35485 1674 35515
rect 73911 35485 73940 35515
rect 1644 35477 1647 35485
rect 73937 35477 73940 35485
rect 73992 35515 73995 35523
rect 73992 35485 74022 35515
rect 73992 35477 73995 35485
rect 1589 35179 1592 35187
rect 1563 35149 1592 35179
rect 1589 35141 1592 35149
rect 1644 35179 1647 35187
rect 73937 35179 73940 35187
rect 1644 35149 1674 35179
rect 73911 35149 73940 35179
rect 1644 35141 1647 35149
rect 73937 35141 73940 35149
rect 73992 35179 73995 35187
rect 73992 35149 74022 35179
rect 73992 35141 73995 35149
rect 1589 34843 1592 34851
rect 1563 34813 1592 34843
rect 1589 34805 1592 34813
rect 1644 34843 1647 34851
rect 73937 34843 73940 34851
rect 1644 34813 1674 34843
rect 73911 34813 73940 34843
rect 1644 34805 1647 34813
rect 73937 34805 73940 34813
rect 73992 34843 73995 34851
rect 73992 34813 74022 34843
rect 73992 34805 73995 34813
rect 1589 34507 1592 34515
rect 1563 34477 1592 34507
rect 1589 34469 1592 34477
rect 1644 34507 1647 34515
rect 73937 34507 73940 34515
rect 1644 34477 1674 34507
rect 73911 34477 73940 34507
rect 1644 34469 1647 34477
rect 73937 34469 73940 34477
rect 73992 34507 73995 34515
rect 73992 34477 74022 34507
rect 73992 34469 73995 34477
rect 1589 34171 1592 34179
rect 1563 34141 1592 34171
rect 1589 34133 1592 34141
rect 1644 34171 1647 34179
rect 73937 34171 73940 34179
rect 1644 34141 1674 34171
rect 73911 34141 73940 34171
rect 1644 34133 1647 34141
rect 73937 34133 73940 34141
rect 73992 34171 73995 34179
rect 73992 34141 74022 34171
rect 73992 34133 73995 34141
rect 1589 33835 1592 33843
rect 1563 33805 1592 33835
rect 1589 33797 1592 33805
rect 1644 33835 1647 33843
rect 73937 33835 73940 33843
rect 1644 33805 1674 33835
rect 73911 33805 73940 33835
rect 1644 33797 1647 33805
rect 73937 33797 73940 33805
rect 73992 33835 73995 33843
rect 73992 33805 74022 33835
rect 73992 33797 73995 33805
rect 1589 33499 1592 33507
rect 1563 33469 1592 33499
rect 1589 33461 1592 33469
rect 1644 33499 1647 33507
rect 73937 33499 73940 33507
rect 1644 33469 1674 33499
rect 73911 33469 73940 33499
rect 1644 33461 1647 33469
rect 73937 33461 73940 33469
rect 73992 33499 73995 33507
rect 73992 33469 74022 33499
rect 73992 33461 73995 33469
rect 1589 33163 1592 33171
rect 1563 33133 1592 33163
rect 1589 33125 1592 33133
rect 1644 33163 1647 33171
rect 73937 33163 73940 33171
rect 1644 33133 1674 33163
rect 73911 33133 73940 33163
rect 1644 33125 1647 33133
rect 73937 33125 73940 33133
rect 73992 33163 73995 33171
rect 73992 33133 74022 33163
rect 73992 33125 73995 33133
rect 1589 32827 1592 32835
rect 1563 32797 1592 32827
rect 1589 32789 1592 32797
rect 1644 32827 1647 32835
rect 73937 32827 73940 32835
rect 1644 32797 1674 32827
rect 73911 32797 73940 32827
rect 1644 32789 1647 32797
rect 73937 32789 73940 32797
rect 73992 32827 73995 32835
rect 73992 32797 74022 32827
rect 73992 32789 73995 32797
rect 1589 32491 1592 32499
rect 1563 32461 1592 32491
rect 1589 32453 1592 32461
rect 1644 32491 1647 32499
rect 73937 32491 73940 32499
rect 1644 32461 1674 32491
rect 73911 32461 73940 32491
rect 1644 32453 1647 32461
rect 73937 32453 73940 32461
rect 73992 32491 73995 32499
rect 73992 32461 74022 32491
rect 73992 32453 73995 32461
rect 1589 32155 1592 32163
rect 1563 32125 1592 32155
rect 1589 32117 1592 32125
rect 1644 32155 1647 32163
rect 73937 32155 73940 32163
rect 1644 32125 1674 32155
rect 73911 32125 73940 32155
rect 1644 32117 1647 32125
rect 73937 32117 73940 32125
rect 73992 32155 73995 32163
rect 73992 32125 74022 32155
rect 73992 32117 73995 32125
rect 1589 31819 1592 31827
rect 1563 31789 1592 31819
rect 1589 31781 1592 31789
rect 1644 31819 1647 31827
rect 73937 31819 73940 31827
rect 1644 31789 1674 31819
rect 73911 31789 73940 31819
rect 1644 31781 1647 31789
rect 73937 31781 73940 31789
rect 73992 31819 73995 31827
rect 73992 31789 74022 31819
rect 73992 31781 73995 31789
rect 1589 31483 1592 31491
rect 1563 31453 1592 31483
rect 1589 31445 1592 31453
rect 1644 31483 1647 31491
rect 73937 31483 73940 31491
rect 1644 31453 1674 31483
rect 73911 31453 73940 31483
rect 1644 31445 1647 31453
rect 73937 31445 73940 31453
rect 73992 31483 73995 31491
rect 73992 31453 74022 31483
rect 73992 31445 73995 31453
rect 1589 31147 1592 31155
rect 1563 31117 1592 31147
rect 1589 31109 1592 31117
rect 1644 31147 1647 31155
rect 73937 31147 73940 31155
rect 1644 31117 1674 31147
rect 73911 31117 73940 31147
rect 1644 31109 1647 31117
rect 73937 31109 73940 31117
rect 73992 31147 73995 31155
rect 73992 31117 74022 31147
rect 73992 31109 73995 31117
rect 1589 30811 1592 30819
rect 1563 30781 1592 30811
rect 1589 30773 1592 30781
rect 1644 30811 1647 30819
rect 73937 30811 73940 30819
rect 1644 30781 1674 30811
rect 73911 30781 73940 30811
rect 1644 30773 1647 30781
rect 73937 30773 73940 30781
rect 73992 30811 73995 30819
rect 73992 30781 74022 30811
rect 73992 30773 73995 30781
rect 1589 30475 1592 30483
rect 1563 30445 1592 30475
rect 1589 30437 1592 30445
rect 1644 30475 1647 30483
rect 73937 30475 73940 30483
rect 1644 30445 1674 30475
rect 73911 30445 73940 30475
rect 1644 30437 1647 30445
rect 73937 30437 73940 30445
rect 73992 30475 73995 30483
rect 73992 30445 74022 30475
rect 73992 30437 73995 30445
rect 1589 30139 1592 30147
rect 1563 30109 1592 30139
rect 1589 30101 1592 30109
rect 1644 30139 1647 30147
rect 73937 30139 73940 30147
rect 1644 30109 1674 30139
rect 73911 30109 73940 30139
rect 1644 30101 1647 30109
rect 73937 30101 73940 30109
rect 73992 30139 73995 30147
rect 73992 30109 74022 30139
rect 73992 30101 73995 30109
rect 1589 29803 1592 29811
rect 1563 29773 1592 29803
rect 1589 29765 1592 29773
rect 1644 29803 1647 29811
rect 73937 29803 73940 29811
rect 1644 29773 1674 29803
rect 73911 29773 73940 29803
rect 1644 29765 1647 29773
rect 73937 29765 73940 29773
rect 73992 29803 73995 29811
rect 73992 29773 74022 29803
rect 73992 29765 73995 29773
rect 1589 29467 1592 29475
rect 1563 29437 1592 29467
rect 1589 29429 1592 29437
rect 1644 29467 1647 29475
rect 73937 29467 73940 29475
rect 1644 29437 1674 29467
rect 73911 29437 73940 29467
rect 1644 29429 1647 29437
rect 73937 29429 73940 29437
rect 73992 29467 73995 29475
rect 73992 29437 74022 29467
rect 73992 29429 73995 29437
rect 1589 29131 1592 29139
rect 1563 29101 1592 29131
rect 1589 29093 1592 29101
rect 1644 29131 1647 29139
rect 73937 29131 73940 29139
rect 1644 29101 1674 29131
rect 73911 29101 73940 29131
rect 1644 29093 1647 29101
rect 73937 29093 73940 29101
rect 73992 29131 73995 29139
rect 73992 29101 74022 29131
rect 73992 29093 73995 29101
rect 1589 28795 1592 28803
rect 1563 28765 1592 28795
rect 1589 28757 1592 28765
rect 1644 28795 1647 28803
rect 73937 28795 73940 28803
rect 1644 28765 1674 28795
rect 73911 28765 73940 28795
rect 1644 28757 1647 28765
rect 73937 28757 73940 28765
rect 73992 28795 73995 28803
rect 73992 28765 74022 28795
rect 73992 28757 73995 28765
rect 1589 28459 1592 28467
rect 1563 28429 1592 28459
rect 1589 28421 1592 28429
rect 1644 28459 1647 28467
rect 73937 28459 73940 28467
rect 1644 28429 1674 28459
rect 73911 28429 73940 28459
rect 1644 28421 1647 28429
rect 73937 28421 73940 28429
rect 73992 28459 73995 28467
rect 73992 28429 74022 28459
rect 73992 28421 73995 28429
rect 1589 28123 1592 28131
rect 1563 28093 1592 28123
rect 1589 28085 1592 28093
rect 1644 28123 1647 28131
rect 73937 28123 73940 28131
rect 1644 28093 1674 28123
rect 73911 28093 73940 28123
rect 1644 28085 1647 28093
rect 73937 28085 73940 28093
rect 73992 28123 73995 28131
rect 73992 28093 74022 28123
rect 73992 28085 73995 28093
rect 1589 27787 1592 27795
rect 1563 27757 1592 27787
rect 1589 27749 1592 27757
rect 1644 27787 1647 27795
rect 73937 27787 73940 27795
rect 1644 27757 1674 27787
rect 73911 27757 73940 27787
rect 1644 27749 1647 27757
rect 73937 27749 73940 27757
rect 73992 27787 73995 27795
rect 73992 27757 74022 27787
rect 73992 27749 73995 27757
rect 1589 27451 1592 27459
rect 1563 27421 1592 27451
rect 1589 27413 1592 27421
rect 1644 27451 1647 27459
rect 73937 27451 73940 27459
rect 1644 27421 1674 27451
rect 73911 27421 73940 27451
rect 1644 27413 1647 27421
rect 73937 27413 73940 27421
rect 73992 27451 73995 27459
rect 73992 27421 74022 27451
rect 73992 27413 73995 27421
rect 1589 27115 1592 27123
rect 1563 27085 1592 27115
rect 1589 27077 1592 27085
rect 1644 27115 1647 27123
rect 73937 27115 73940 27123
rect 1644 27085 1674 27115
rect 73911 27085 73940 27115
rect 1644 27077 1647 27085
rect 73937 27077 73940 27085
rect 73992 27115 73995 27123
rect 73992 27085 74022 27115
rect 73992 27077 73995 27085
rect 1589 26779 1592 26787
rect 1563 26749 1592 26779
rect 1589 26741 1592 26749
rect 1644 26779 1647 26787
rect 73937 26779 73940 26787
rect 1644 26749 1674 26779
rect 73911 26749 73940 26779
rect 1644 26741 1647 26749
rect 73937 26741 73940 26749
rect 73992 26779 73995 26787
rect 73992 26749 74022 26779
rect 73992 26741 73995 26749
rect 1589 26443 1592 26451
rect 1563 26413 1592 26443
rect 1589 26405 1592 26413
rect 1644 26443 1647 26451
rect 73937 26443 73940 26451
rect 1644 26413 1674 26443
rect 73911 26413 73940 26443
rect 1644 26405 1647 26413
rect 73937 26405 73940 26413
rect 73992 26443 73995 26451
rect 73992 26413 74022 26443
rect 73992 26405 73995 26413
rect 1589 26107 1592 26115
rect 1563 26077 1592 26107
rect 1589 26069 1592 26077
rect 1644 26107 1647 26115
rect 73937 26107 73940 26115
rect 1644 26077 1674 26107
rect 73911 26077 73940 26107
rect 1644 26069 1647 26077
rect 73937 26069 73940 26077
rect 73992 26107 73995 26115
rect 73992 26077 74022 26107
rect 73992 26069 73995 26077
rect 1589 25771 1592 25779
rect 1563 25741 1592 25771
rect 1589 25733 1592 25741
rect 1644 25771 1647 25779
rect 73937 25771 73940 25779
rect 1644 25741 1674 25771
rect 73911 25741 73940 25771
rect 1644 25733 1647 25741
rect 73937 25733 73940 25741
rect 73992 25771 73995 25779
rect 73992 25741 74022 25771
rect 73992 25733 73995 25741
rect 1589 25435 1592 25443
rect 1563 25405 1592 25435
rect 1589 25397 1592 25405
rect 1644 25435 1647 25443
rect 73937 25435 73940 25443
rect 1644 25405 1674 25435
rect 73911 25405 73940 25435
rect 1644 25397 1647 25405
rect 73937 25397 73940 25405
rect 73992 25435 73995 25443
rect 73992 25405 74022 25435
rect 73992 25397 73995 25405
rect 1589 25099 1592 25107
rect 1563 25069 1592 25099
rect 1589 25061 1592 25069
rect 1644 25099 1647 25107
rect 73937 25099 73940 25107
rect 1644 25069 1674 25099
rect 73911 25069 73940 25099
rect 1644 25061 1647 25069
rect 73937 25061 73940 25069
rect 73992 25099 73995 25107
rect 73992 25069 74022 25099
rect 73992 25061 73995 25069
rect 1589 24763 1592 24771
rect 1563 24733 1592 24763
rect 1589 24725 1592 24733
rect 1644 24763 1647 24771
rect 73937 24763 73940 24771
rect 1644 24733 1674 24763
rect 73911 24733 73940 24763
rect 1644 24725 1647 24733
rect 73937 24725 73940 24733
rect 73992 24763 73995 24771
rect 73992 24733 74022 24763
rect 73992 24725 73995 24733
rect 1589 24427 1592 24435
rect 1563 24397 1592 24427
rect 1589 24389 1592 24397
rect 1644 24427 1647 24435
rect 73937 24427 73940 24435
rect 1644 24397 1674 24427
rect 73911 24397 73940 24427
rect 1644 24389 1647 24397
rect 73937 24389 73940 24397
rect 73992 24427 73995 24435
rect 73992 24397 74022 24427
rect 73992 24389 73995 24397
rect 1589 24091 1592 24099
rect 1563 24061 1592 24091
rect 1589 24053 1592 24061
rect 1644 24091 1647 24099
rect 73937 24091 73940 24099
rect 1644 24061 1674 24091
rect 73911 24061 73940 24091
rect 1644 24053 1647 24061
rect 73937 24053 73940 24061
rect 73992 24091 73995 24099
rect 73992 24061 74022 24091
rect 73992 24053 73995 24061
rect 1589 23755 1592 23763
rect 1563 23725 1592 23755
rect 1589 23717 1592 23725
rect 1644 23755 1647 23763
rect 73937 23755 73940 23763
rect 1644 23725 1674 23755
rect 73911 23725 73940 23755
rect 1644 23717 1647 23725
rect 73937 23717 73940 23725
rect 73992 23755 73995 23763
rect 73992 23725 74022 23755
rect 73992 23717 73995 23725
rect 1589 23419 1592 23427
rect 1563 23389 1592 23419
rect 1589 23381 1592 23389
rect 1644 23419 1647 23427
rect 73937 23419 73940 23427
rect 1644 23389 1674 23419
rect 73911 23389 73940 23419
rect 1644 23381 1647 23389
rect 73937 23381 73940 23389
rect 73992 23419 73995 23427
rect 73992 23389 74022 23419
rect 73992 23381 73995 23389
rect 1589 23083 1592 23091
rect 1563 23053 1592 23083
rect 1589 23045 1592 23053
rect 1644 23083 1647 23091
rect 73937 23083 73940 23091
rect 1644 23053 1674 23083
rect 73911 23053 73940 23083
rect 1644 23045 1647 23053
rect 73937 23045 73940 23053
rect 73992 23083 73995 23091
rect 73992 23053 74022 23083
rect 73992 23045 73995 23053
rect 1589 22747 1592 22755
rect 1563 22717 1592 22747
rect 1589 22709 1592 22717
rect 1644 22747 1647 22755
rect 73937 22747 73940 22755
rect 1644 22717 1674 22747
rect 73911 22717 73940 22747
rect 1644 22709 1647 22717
rect 73937 22709 73940 22717
rect 73992 22747 73995 22755
rect 73992 22717 74022 22747
rect 73992 22709 73995 22717
rect 1589 22411 1592 22419
rect 1563 22381 1592 22411
rect 1589 22373 1592 22381
rect 1644 22411 1647 22419
rect 73937 22411 73940 22419
rect 1644 22381 1674 22411
rect 73911 22381 73940 22411
rect 1644 22373 1647 22381
rect 73937 22373 73940 22381
rect 73992 22411 73995 22419
rect 73992 22381 74022 22411
rect 73992 22373 73995 22381
rect 1589 22075 1592 22083
rect 1563 22045 1592 22075
rect 1589 22037 1592 22045
rect 1644 22075 1647 22083
rect 73937 22075 73940 22083
rect 1644 22045 1674 22075
rect 73911 22045 73940 22075
rect 1644 22037 1647 22045
rect 73937 22037 73940 22045
rect 73992 22075 73995 22083
rect 73992 22045 74022 22075
rect 73992 22037 73995 22045
rect 1589 21739 1592 21747
rect 1563 21709 1592 21739
rect 1589 21701 1592 21709
rect 1644 21739 1647 21747
rect 73937 21739 73940 21747
rect 1644 21709 1674 21739
rect 73911 21709 73940 21739
rect 1644 21701 1647 21709
rect 73937 21701 73940 21709
rect 73992 21739 73995 21747
rect 73992 21709 74022 21739
rect 73992 21701 73995 21709
rect 1589 21403 1592 21411
rect 1563 21373 1592 21403
rect 1589 21365 1592 21373
rect 1644 21403 1647 21411
rect 73937 21403 73940 21411
rect 1644 21373 1674 21403
rect 73911 21373 73940 21403
rect 1644 21365 1647 21373
rect 73937 21365 73940 21373
rect 73992 21403 73995 21411
rect 73992 21373 74022 21403
rect 73992 21365 73995 21373
rect 1589 21067 1592 21075
rect 1563 21037 1592 21067
rect 1589 21029 1592 21037
rect 1644 21067 1647 21075
rect 73937 21067 73940 21075
rect 1644 21037 1674 21067
rect 73911 21037 73940 21067
rect 1644 21029 1647 21037
rect 73937 21029 73940 21037
rect 73992 21067 73995 21075
rect 73992 21037 74022 21067
rect 73992 21029 73995 21037
rect 1589 20731 1592 20739
rect 1563 20701 1592 20731
rect 1589 20693 1592 20701
rect 1644 20731 1647 20739
rect 73937 20731 73940 20739
rect 1644 20701 1674 20731
rect 73911 20701 73940 20731
rect 1644 20693 1647 20701
rect 73937 20693 73940 20701
rect 73992 20731 73995 20739
rect 73992 20701 74022 20731
rect 73992 20693 73995 20701
rect 1589 20395 1592 20403
rect 1563 20365 1592 20395
rect 1589 20357 1592 20365
rect 1644 20395 1647 20403
rect 73937 20395 73940 20403
rect 1644 20365 1674 20395
rect 73911 20365 73940 20395
rect 1644 20357 1647 20365
rect 73937 20357 73940 20365
rect 73992 20395 73995 20403
rect 73992 20365 74022 20395
rect 73992 20357 73995 20365
rect 1589 20059 1592 20067
rect 1563 20029 1592 20059
rect 1589 20021 1592 20029
rect 1644 20059 1647 20067
rect 73937 20059 73940 20067
rect 1644 20029 1674 20059
rect 73911 20029 73940 20059
rect 1644 20021 1647 20029
rect 73937 20021 73940 20029
rect 73992 20059 73995 20067
rect 73992 20029 74022 20059
rect 73992 20021 73995 20029
rect 1589 19723 1592 19731
rect 1563 19693 1592 19723
rect 1589 19685 1592 19693
rect 1644 19723 1647 19731
rect 73937 19723 73940 19731
rect 1644 19693 1674 19723
rect 73911 19693 73940 19723
rect 1644 19685 1647 19693
rect 73937 19685 73940 19693
rect 73992 19723 73995 19731
rect 73992 19693 74022 19723
rect 73992 19685 73995 19693
rect 1589 19387 1592 19395
rect 1563 19357 1592 19387
rect 1589 19349 1592 19357
rect 1644 19387 1647 19395
rect 73937 19387 73940 19395
rect 1644 19357 1674 19387
rect 73911 19357 73940 19387
rect 1644 19349 1647 19357
rect 73937 19349 73940 19357
rect 73992 19387 73995 19395
rect 73992 19357 74022 19387
rect 73992 19349 73995 19357
rect 1589 19051 1592 19059
rect 1563 19021 1592 19051
rect 1589 19013 1592 19021
rect 1644 19051 1647 19059
rect 73937 19051 73940 19059
rect 1644 19021 1674 19051
rect 73911 19021 73940 19051
rect 1644 19013 1647 19021
rect 73937 19013 73940 19021
rect 73992 19051 73995 19059
rect 73992 19021 74022 19051
rect 73992 19013 73995 19021
rect 1589 18715 1592 18723
rect 1563 18685 1592 18715
rect 1589 18677 1592 18685
rect 1644 18715 1647 18723
rect 73937 18715 73940 18723
rect 1644 18685 1674 18715
rect 73911 18685 73940 18715
rect 1644 18677 1647 18685
rect 73937 18677 73940 18685
rect 73992 18715 73995 18723
rect 73992 18685 74022 18715
rect 73992 18677 73995 18685
rect 1589 18379 1592 18387
rect 1563 18349 1592 18379
rect 1589 18341 1592 18349
rect 1644 18379 1647 18387
rect 73937 18379 73940 18387
rect 1644 18349 1674 18379
rect 73911 18349 73940 18379
rect 1644 18341 1647 18349
rect 73937 18341 73940 18349
rect 73992 18379 73995 18387
rect 73992 18349 74022 18379
rect 73992 18341 73995 18349
rect 1589 18043 1592 18051
rect 1563 18013 1592 18043
rect 1589 18005 1592 18013
rect 1644 18043 1647 18051
rect 73937 18043 73940 18051
rect 1644 18013 1674 18043
rect 73911 18013 73940 18043
rect 1644 18005 1647 18013
rect 73937 18005 73940 18013
rect 73992 18043 73995 18051
rect 73992 18013 74022 18043
rect 73992 18005 73995 18013
rect 1589 17707 1592 17715
rect 1563 17677 1592 17707
rect 1589 17669 1592 17677
rect 1644 17707 1647 17715
rect 73937 17707 73940 17715
rect 1644 17677 1674 17707
rect 73911 17677 73940 17707
rect 1644 17669 1647 17677
rect 73937 17669 73940 17677
rect 73992 17707 73995 17715
rect 73992 17677 74022 17707
rect 73992 17669 73995 17677
rect 1589 17371 1592 17379
rect 1563 17341 1592 17371
rect 1589 17333 1592 17341
rect 1644 17371 1647 17379
rect 73937 17371 73940 17379
rect 1644 17341 1674 17371
rect 73911 17341 73940 17371
rect 1644 17333 1647 17341
rect 73937 17333 73940 17341
rect 73992 17371 73995 17379
rect 73992 17341 74022 17371
rect 73992 17333 73995 17341
rect 1589 17035 1592 17043
rect 1563 17005 1592 17035
rect 1589 16997 1592 17005
rect 1644 17035 1647 17043
rect 73937 17035 73940 17043
rect 1644 17005 1674 17035
rect 73911 17005 73940 17035
rect 1644 16997 1647 17005
rect 73937 16997 73940 17005
rect 73992 17035 73995 17043
rect 73992 17005 74022 17035
rect 73992 16997 73995 17005
rect 1589 16699 1592 16707
rect 1563 16669 1592 16699
rect 1589 16661 1592 16669
rect 1644 16699 1647 16707
rect 73937 16699 73940 16707
rect 1644 16669 1674 16699
rect 73911 16669 73940 16699
rect 1644 16661 1647 16669
rect 73937 16661 73940 16669
rect 73992 16699 73995 16707
rect 73992 16669 74022 16699
rect 73992 16661 73995 16669
rect 1589 16363 1592 16371
rect 1563 16333 1592 16363
rect 1589 16325 1592 16333
rect 1644 16363 1647 16371
rect 73937 16363 73940 16371
rect 1644 16333 1674 16363
rect 73911 16333 73940 16363
rect 1644 16325 1647 16333
rect 73937 16325 73940 16333
rect 73992 16363 73995 16371
rect 73992 16333 74022 16363
rect 73992 16325 73995 16333
rect 1589 16027 1592 16035
rect 1563 15997 1592 16027
rect 1589 15989 1592 15997
rect 1644 16027 1647 16035
rect 73937 16027 73940 16035
rect 1644 15997 1674 16027
rect 73911 15997 73940 16027
rect 1644 15989 1647 15997
rect 73937 15989 73940 15997
rect 73992 16027 73995 16035
rect 73992 15997 74022 16027
rect 73992 15989 73995 15997
rect 1589 15691 1592 15699
rect 1563 15661 1592 15691
rect 1589 15653 1592 15661
rect 1644 15691 1647 15699
rect 73937 15691 73940 15699
rect 1644 15661 1674 15691
rect 73911 15661 73940 15691
rect 1644 15653 1647 15661
rect 73937 15653 73940 15661
rect 73992 15691 73995 15699
rect 73992 15661 74022 15691
rect 73992 15653 73995 15661
rect 1589 15355 1592 15363
rect 1563 15325 1592 15355
rect 1589 15317 1592 15325
rect 1644 15355 1647 15363
rect 73937 15355 73940 15363
rect 1644 15325 1674 15355
rect 73911 15325 73940 15355
rect 1644 15317 1647 15325
rect 73937 15317 73940 15325
rect 73992 15355 73995 15363
rect 73992 15325 74022 15355
rect 73992 15317 73995 15325
rect 1589 15019 1592 15027
rect 1563 14989 1592 15019
rect 1589 14981 1592 14989
rect 1644 15019 1647 15027
rect 73937 15019 73940 15027
rect 1644 14989 1674 15019
rect 73911 14989 73940 15019
rect 1644 14981 1647 14989
rect 73937 14981 73940 14989
rect 73992 15019 73995 15027
rect 73992 14989 74022 15019
rect 73992 14981 73995 14989
rect 1589 14683 1592 14691
rect 1563 14653 1592 14683
rect 1589 14645 1592 14653
rect 1644 14683 1647 14691
rect 73937 14683 73940 14691
rect 1644 14653 1674 14683
rect 73911 14653 73940 14683
rect 1644 14645 1647 14653
rect 73937 14645 73940 14653
rect 73992 14683 73995 14691
rect 73992 14653 74022 14683
rect 73992 14645 73995 14653
rect 1589 14347 1592 14355
rect 1563 14317 1592 14347
rect 1589 14309 1592 14317
rect 1644 14347 1647 14355
rect 73937 14347 73940 14355
rect 1644 14317 1674 14347
rect 73911 14317 73940 14347
rect 1644 14309 1647 14317
rect 73937 14309 73940 14317
rect 73992 14347 73995 14355
rect 73992 14317 74022 14347
rect 73992 14309 73995 14317
rect 1589 14011 1592 14019
rect 1563 13981 1592 14011
rect 1589 13973 1592 13981
rect 1644 14011 1647 14019
rect 73937 14011 73940 14019
rect 1644 13981 1674 14011
rect 73911 13981 73940 14011
rect 1644 13973 1647 13981
rect 73937 13973 73940 13981
rect 73992 14011 73995 14019
rect 73992 13981 74022 14011
rect 73992 13973 73995 13981
rect 1589 13675 1592 13683
rect 1563 13645 1592 13675
rect 1589 13637 1592 13645
rect 1644 13675 1647 13683
rect 73937 13675 73940 13683
rect 1644 13645 1674 13675
rect 73911 13645 73940 13675
rect 1644 13637 1647 13645
rect 73937 13637 73940 13645
rect 73992 13675 73995 13683
rect 73992 13645 74022 13675
rect 73992 13637 73995 13645
rect 1589 13339 1592 13347
rect 1563 13309 1592 13339
rect 1589 13301 1592 13309
rect 1644 13339 1647 13347
rect 73937 13339 73940 13347
rect 1644 13309 1674 13339
rect 73911 13309 73940 13339
rect 1644 13301 1647 13309
rect 73937 13301 73940 13309
rect 73992 13339 73995 13347
rect 73992 13309 74022 13339
rect 73992 13301 73995 13309
rect 1589 13003 1592 13011
rect 1563 12973 1592 13003
rect 1589 12965 1592 12973
rect 1644 13003 1647 13011
rect 73937 13003 73940 13011
rect 1644 12973 1674 13003
rect 73911 12973 73940 13003
rect 1644 12965 1647 12973
rect 73937 12965 73940 12973
rect 73992 13003 73995 13011
rect 73992 12973 74022 13003
rect 73992 12965 73995 12973
rect 1589 12667 1592 12675
rect 1563 12637 1592 12667
rect 1589 12629 1592 12637
rect 1644 12667 1647 12675
rect 73937 12667 73940 12675
rect 1644 12637 1674 12667
rect 73911 12637 73940 12667
rect 1644 12629 1647 12637
rect 73937 12629 73940 12637
rect 73992 12667 73995 12675
rect 73992 12637 74022 12667
rect 73992 12629 73995 12637
rect 1589 12331 1592 12339
rect 1563 12301 1592 12331
rect 1589 12293 1592 12301
rect 1644 12331 1647 12339
rect 73937 12331 73940 12339
rect 1644 12301 1674 12331
rect 73911 12301 73940 12331
rect 1644 12293 1647 12301
rect 73937 12293 73940 12301
rect 73992 12331 73995 12339
rect 73992 12301 74022 12331
rect 73992 12293 73995 12301
rect 1589 11995 1592 12003
rect 1563 11965 1592 11995
rect 1589 11957 1592 11965
rect 1644 11995 1647 12003
rect 73937 11995 73940 12003
rect 1644 11965 1674 11995
rect 73911 11965 73940 11995
rect 1644 11957 1647 11965
rect 73937 11957 73940 11965
rect 73992 11995 73995 12003
rect 73992 11965 74022 11995
rect 73992 11957 73995 11965
rect 1589 11659 1592 11667
rect 1563 11629 1592 11659
rect 1589 11621 1592 11629
rect 1644 11659 1647 11667
rect 73937 11659 73940 11667
rect 1644 11629 1674 11659
rect 73911 11629 73940 11659
rect 1644 11621 1647 11629
rect 73937 11621 73940 11629
rect 73992 11659 73995 11667
rect 73992 11629 74022 11659
rect 73992 11621 73995 11629
rect 1589 11323 1592 11331
rect 1563 11293 1592 11323
rect 1589 11285 1592 11293
rect 1644 11323 1647 11331
rect 73937 11323 73940 11331
rect 1644 11293 1674 11323
rect 73911 11293 73940 11323
rect 1644 11285 1647 11293
rect 73937 11285 73940 11293
rect 73992 11323 73995 11331
rect 73992 11293 74022 11323
rect 73992 11285 73995 11293
rect 1589 10987 1592 10995
rect 1563 10957 1592 10987
rect 1589 10949 1592 10957
rect 1644 10987 1647 10995
rect 73937 10987 73940 10995
rect 1644 10957 1674 10987
rect 73911 10957 73940 10987
rect 1644 10949 1647 10957
rect 73937 10949 73940 10957
rect 73992 10987 73995 10995
rect 73992 10957 74022 10987
rect 73992 10949 73995 10957
rect 1589 10651 1592 10659
rect 1563 10621 1592 10651
rect 1589 10613 1592 10621
rect 1644 10651 1647 10659
rect 73937 10651 73940 10659
rect 1644 10621 1674 10651
rect 73911 10621 73940 10651
rect 1644 10613 1647 10621
rect 73937 10613 73940 10621
rect 73992 10651 73995 10659
rect 73992 10621 74022 10651
rect 73992 10613 73995 10621
rect 1589 10315 1592 10323
rect 1563 10285 1592 10315
rect 1589 10277 1592 10285
rect 1644 10315 1647 10323
rect 73937 10315 73940 10323
rect 1644 10285 1674 10315
rect 73911 10285 73940 10315
rect 1644 10277 1647 10285
rect 73937 10277 73940 10285
rect 73992 10315 73995 10323
rect 73992 10285 74022 10315
rect 73992 10277 73995 10285
rect 1589 9979 1592 9987
rect 1563 9949 1592 9979
rect 1589 9941 1592 9949
rect 1644 9979 1647 9987
rect 73937 9979 73940 9987
rect 1644 9949 1674 9979
rect 73911 9949 73940 9979
rect 1644 9941 1647 9949
rect 73937 9941 73940 9949
rect 73992 9979 73995 9987
rect 73992 9949 74022 9979
rect 73992 9941 73995 9949
rect 1589 9643 1592 9651
rect 1563 9613 1592 9643
rect 1589 9605 1592 9613
rect 1644 9643 1647 9651
rect 73937 9643 73940 9651
rect 1644 9613 1674 9643
rect 73911 9613 73940 9643
rect 1644 9605 1647 9613
rect 73937 9605 73940 9613
rect 73992 9643 73995 9651
rect 73992 9613 74022 9643
rect 73992 9605 73995 9613
rect 1589 9307 1592 9315
rect 1563 9277 1592 9307
rect 1589 9269 1592 9277
rect 1644 9307 1647 9315
rect 73937 9307 73940 9315
rect 1644 9277 1674 9307
rect 73911 9277 73940 9307
rect 1644 9269 1647 9277
rect 73937 9269 73940 9277
rect 73992 9307 73995 9315
rect 73992 9277 74022 9307
rect 73992 9269 73995 9277
rect 1589 8971 1592 8979
rect 1563 8941 1592 8971
rect 1589 8933 1592 8941
rect 1644 8971 1647 8979
rect 73937 8971 73940 8979
rect 1644 8941 1674 8971
rect 73911 8941 73940 8971
rect 1644 8933 1647 8941
rect 73937 8933 73940 8941
rect 73992 8971 73995 8979
rect 73992 8941 74022 8971
rect 73992 8933 73995 8941
rect 1589 8635 1592 8643
rect 1563 8605 1592 8635
rect 1589 8597 1592 8605
rect 1644 8635 1647 8643
rect 73937 8635 73940 8643
rect 1644 8605 1674 8635
rect 73911 8605 73940 8635
rect 1644 8597 1647 8605
rect 73937 8597 73940 8605
rect 73992 8635 73995 8643
rect 73992 8605 74022 8635
rect 73992 8597 73995 8605
rect 1589 8299 1592 8307
rect 1563 8269 1592 8299
rect 1589 8261 1592 8269
rect 1644 8299 1647 8307
rect 73937 8299 73940 8307
rect 1644 8269 1674 8299
rect 73911 8269 73940 8299
rect 1644 8261 1647 8269
rect 73937 8261 73940 8269
rect 73992 8299 73995 8307
rect 73992 8269 74022 8299
rect 73992 8261 73995 8269
rect 1589 7963 1592 7971
rect 1563 7933 1592 7963
rect 1589 7925 1592 7933
rect 1644 7963 1647 7971
rect 73937 7963 73940 7971
rect 1644 7933 1674 7963
rect 73911 7933 73940 7963
rect 1644 7925 1647 7933
rect 73937 7925 73940 7933
rect 73992 7963 73995 7971
rect 73992 7933 74022 7963
rect 73992 7925 73995 7933
rect 1589 7627 1592 7635
rect 1563 7597 1592 7627
rect 1589 7589 1592 7597
rect 1644 7627 1647 7635
rect 73937 7627 73940 7635
rect 1644 7597 1674 7627
rect 73911 7597 73940 7627
rect 1644 7589 1647 7597
rect 73937 7589 73940 7597
rect 73992 7627 73995 7635
rect 73992 7597 74022 7627
rect 73992 7589 73995 7597
rect 1589 7291 1592 7299
rect 1563 7261 1592 7291
rect 1589 7253 1592 7261
rect 1644 7291 1647 7299
rect 73937 7291 73940 7299
rect 1644 7261 1674 7291
rect 73911 7261 73940 7291
rect 1644 7253 1647 7261
rect 73937 7253 73940 7261
rect 73992 7291 73995 7299
rect 73992 7261 74022 7291
rect 73992 7253 73995 7261
rect 1589 6955 1592 6963
rect 1563 6925 1592 6955
rect 1589 6917 1592 6925
rect 1644 6955 1647 6963
rect 73937 6955 73940 6963
rect 1644 6925 1674 6955
rect 73911 6925 73940 6955
rect 1644 6917 1647 6925
rect 73937 6917 73940 6925
rect 73992 6955 73995 6963
rect 73992 6925 74022 6955
rect 73992 6917 73995 6925
rect 1589 6619 1592 6627
rect 1563 6589 1592 6619
rect 1589 6581 1592 6589
rect 1644 6619 1647 6627
rect 73937 6619 73940 6627
rect 1644 6589 1674 6619
rect 73911 6589 73940 6619
rect 1644 6581 1647 6589
rect 73937 6581 73940 6589
rect 73992 6619 73995 6627
rect 73992 6589 74022 6619
rect 73992 6581 73995 6589
rect 1589 6283 1592 6291
rect 1563 6253 1592 6283
rect 1589 6245 1592 6253
rect 1644 6283 1647 6291
rect 73937 6283 73940 6291
rect 1644 6253 1674 6283
rect 73911 6253 73940 6283
rect 1644 6245 1647 6253
rect 73937 6245 73940 6253
rect 73992 6283 73995 6291
rect 73992 6253 74022 6283
rect 73992 6245 73995 6253
rect 1589 5947 1592 5955
rect 1563 5917 1592 5947
rect 1589 5909 1592 5917
rect 1644 5947 1647 5955
rect 73937 5947 73940 5955
rect 1644 5917 1674 5947
rect 73911 5917 73940 5947
rect 1644 5909 1647 5917
rect 73937 5909 73940 5917
rect 73992 5947 73995 5955
rect 73992 5917 74022 5947
rect 73992 5909 73995 5917
rect 1589 5611 1592 5619
rect 1563 5581 1592 5611
rect 1589 5573 1592 5581
rect 1644 5611 1647 5619
rect 73937 5611 73940 5619
rect 1644 5581 1674 5611
rect 73911 5581 73940 5611
rect 1644 5573 1647 5581
rect 73937 5573 73940 5581
rect 73992 5611 73995 5619
rect 73992 5581 74022 5611
rect 73992 5573 73995 5581
rect 1589 5275 1592 5283
rect 1563 5245 1592 5275
rect 1589 5237 1592 5245
rect 1644 5275 1647 5283
rect 73937 5275 73940 5283
rect 1644 5245 1674 5275
rect 73911 5245 73940 5275
rect 1644 5237 1647 5245
rect 73937 5237 73940 5245
rect 73992 5275 73995 5283
rect 73992 5245 74022 5275
rect 73992 5237 73995 5245
rect 1589 4939 1592 4947
rect 1563 4909 1592 4939
rect 1589 4901 1592 4909
rect 1644 4939 1647 4947
rect 73937 4939 73940 4947
rect 1644 4909 1674 4939
rect 73911 4909 73940 4939
rect 1644 4901 1647 4909
rect 73937 4901 73940 4909
rect 73992 4939 73995 4947
rect 73992 4909 74022 4939
rect 73992 4901 73995 4909
rect 1589 4603 1592 4611
rect 1563 4573 1592 4603
rect 1589 4565 1592 4573
rect 1644 4603 1647 4611
rect 73937 4603 73940 4611
rect 1644 4573 1674 4603
rect 73911 4573 73940 4603
rect 1644 4565 1647 4573
rect 73937 4565 73940 4573
rect 73992 4603 73995 4611
rect 73992 4573 74022 4603
rect 73992 4565 73995 4573
rect 1589 4267 1592 4275
rect 1563 4237 1592 4267
rect 1589 4229 1592 4237
rect 1644 4267 1647 4275
rect 73937 4267 73940 4275
rect 1644 4237 1674 4267
rect 73911 4237 73940 4267
rect 1644 4229 1647 4237
rect 73937 4229 73940 4237
rect 73992 4267 73995 4275
rect 73992 4237 74022 4267
rect 73992 4229 73995 4237
rect 1589 3931 1592 3939
rect 1563 3901 1592 3931
rect 1589 3893 1592 3901
rect 1644 3931 1647 3939
rect 73937 3931 73940 3939
rect 1644 3901 1674 3931
rect 73911 3901 73940 3931
rect 1644 3893 1647 3901
rect 73937 3893 73940 3901
rect 73992 3931 73995 3939
rect 73992 3901 74022 3931
rect 73992 3893 73995 3901
rect 1589 3595 1592 3603
rect 1563 3565 1592 3595
rect 1589 3557 1592 3565
rect 1644 3595 1647 3603
rect 73937 3595 73940 3603
rect 1644 3565 1674 3595
rect 73911 3565 73940 3595
rect 1644 3557 1647 3565
rect 73937 3557 73940 3565
rect 73992 3595 73995 3603
rect 73992 3565 74022 3595
rect 73992 3557 73995 3565
rect 1589 3259 1592 3267
rect 1563 3229 1592 3259
rect 1589 3221 1592 3229
rect 1644 3259 1647 3267
rect 73937 3259 73940 3267
rect 1644 3229 1674 3259
rect 73911 3229 73940 3259
rect 1644 3221 1647 3229
rect 73937 3221 73940 3229
rect 73992 3259 73995 3267
rect 73992 3229 74022 3259
rect 73992 3221 73995 3229
rect 1589 2923 1592 2931
rect 1563 2893 1592 2923
rect 1589 2885 1592 2893
rect 1644 2923 1647 2931
rect 73937 2923 73940 2931
rect 1644 2893 1674 2923
rect 73911 2893 73940 2923
rect 1644 2885 1647 2893
rect 73937 2885 73940 2893
rect 73992 2923 73995 2931
rect 73992 2893 74022 2923
rect 73992 2885 73995 2893
rect 1589 2587 1592 2595
rect 1563 2557 1592 2587
rect 1589 2549 1592 2557
rect 1644 2587 1647 2595
rect 73937 2587 73940 2595
rect 1644 2557 1674 2587
rect 73911 2557 73940 2587
rect 1644 2549 1647 2557
rect 73937 2549 73940 2557
rect 73992 2587 73995 2595
rect 73992 2557 74022 2587
rect 73992 2549 73995 2557
rect 1589 2251 1592 2259
rect 1563 2221 1592 2251
rect 1589 2213 1592 2221
rect 1644 2251 1647 2259
rect 73937 2251 73940 2259
rect 1644 2221 1674 2251
rect 73911 2221 73940 2251
rect 1644 2213 1647 2221
rect 73937 2213 73940 2221
rect 73992 2251 73995 2259
rect 73992 2221 74022 2251
rect 73992 2213 73995 2221
rect 1589 1915 1592 1923
rect 1563 1885 1592 1915
rect 1589 1877 1592 1885
rect 1644 1915 1647 1923
rect 73937 1915 73940 1923
rect 1644 1885 1674 1915
rect 73911 1885 73940 1915
rect 1644 1877 1647 1885
rect 73937 1877 73940 1885
rect 73992 1915 73995 1923
rect 73992 1885 74022 1915
rect 73992 1877 73995 1885
rect 1506 1590 74078 1676
rect 1506 1538 1928 1590
rect 1980 1581 3608 1590
rect 3660 1581 5288 1590
rect 5340 1581 6968 1590
rect 7020 1581 8648 1590
rect 8700 1581 10328 1590
rect 10380 1581 12008 1590
rect 12060 1581 13688 1590
rect 13740 1581 15368 1590
rect 15420 1581 17048 1590
rect 17100 1581 18728 1590
rect 18780 1581 20408 1590
rect 20460 1581 22088 1590
rect 22140 1581 23768 1590
rect 23820 1581 25448 1590
rect 25500 1581 27128 1590
rect 27180 1581 28808 1590
rect 28860 1581 30488 1590
rect 30540 1581 32168 1590
rect 32220 1581 33848 1590
rect 33900 1581 35528 1590
rect 35580 1581 37208 1590
rect 37260 1581 38888 1590
rect 38940 1581 40568 1590
rect 40620 1581 42248 1590
rect 42300 1581 43928 1590
rect 43980 1581 45608 1590
rect 45660 1581 47288 1590
rect 47340 1581 48968 1590
rect 49020 1581 50648 1590
rect 50700 1581 52328 1590
rect 52380 1581 54008 1590
rect 54060 1581 55688 1590
rect 55740 1581 57368 1590
rect 57420 1581 59048 1590
rect 59100 1581 60728 1590
rect 60780 1581 62408 1590
rect 62460 1581 64088 1590
rect 64140 1581 65768 1590
rect 65820 1581 67448 1590
rect 67500 1581 69128 1590
rect 69180 1581 70808 1590
rect 70860 1581 72488 1590
rect 72540 1581 74078 1590
rect 1980 1547 2273 1581
rect 2307 1547 2609 1581
rect 2643 1547 2945 1581
rect 2979 1547 3281 1581
rect 3315 1547 3608 1581
rect 3660 1547 3953 1581
rect 3987 1547 4289 1581
rect 4323 1547 4625 1581
rect 4659 1547 4961 1581
rect 4995 1547 5288 1581
rect 5340 1547 5633 1581
rect 5667 1547 5969 1581
rect 6003 1547 6305 1581
rect 6339 1547 6641 1581
rect 6675 1547 6968 1581
rect 7020 1547 7313 1581
rect 7347 1547 7649 1581
rect 7683 1547 7985 1581
rect 8019 1547 8321 1581
rect 8355 1547 8648 1581
rect 8700 1547 8993 1581
rect 9027 1547 9329 1581
rect 9363 1547 9665 1581
rect 9699 1547 10001 1581
rect 10035 1547 10328 1581
rect 10380 1547 10673 1581
rect 10707 1547 11009 1581
rect 11043 1547 11345 1581
rect 11379 1547 11681 1581
rect 11715 1547 12008 1581
rect 12060 1547 12353 1581
rect 12387 1547 12689 1581
rect 12723 1547 13025 1581
rect 13059 1547 13361 1581
rect 13395 1547 13688 1581
rect 13740 1547 14033 1581
rect 14067 1547 14369 1581
rect 14403 1547 14705 1581
rect 14739 1547 15041 1581
rect 15075 1547 15368 1581
rect 15420 1547 15713 1581
rect 15747 1547 16049 1581
rect 16083 1547 16385 1581
rect 16419 1547 16721 1581
rect 16755 1547 17048 1581
rect 17100 1547 17393 1581
rect 17427 1547 17729 1581
rect 17763 1547 18065 1581
rect 18099 1547 18401 1581
rect 18435 1547 18728 1581
rect 18780 1547 19073 1581
rect 19107 1547 19409 1581
rect 19443 1547 19745 1581
rect 19779 1547 20081 1581
rect 20115 1547 20408 1581
rect 20460 1547 20753 1581
rect 20787 1547 21089 1581
rect 21123 1547 21425 1581
rect 21459 1547 21761 1581
rect 21795 1547 22088 1581
rect 22140 1547 22433 1581
rect 22467 1547 22769 1581
rect 22803 1547 23105 1581
rect 23139 1547 23441 1581
rect 23475 1547 23768 1581
rect 23820 1547 24113 1581
rect 24147 1547 24449 1581
rect 24483 1547 24785 1581
rect 24819 1547 25121 1581
rect 25155 1547 25448 1581
rect 25500 1547 25793 1581
rect 25827 1547 26129 1581
rect 26163 1547 26465 1581
rect 26499 1547 26801 1581
rect 26835 1547 27128 1581
rect 27180 1547 27473 1581
rect 27507 1547 27809 1581
rect 27843 1547 28145 1581
rect 28179 1547 28481 1581
rect 28515 1547 28808 1581
rect 28860 1547 29153 1581
rect 29187 1547 29489 1581
rect 29523 1547 29825 1581
rect 29859 1547 30161 1581
rect 30195 1547 30488 1581
rect 30540 1547 30833 1581
rect 30867 1547 31169 1581
rect 31203 1547 31505 1581
rect 31539 1547 31841 1581
rect 31875 1547 32168 1581
rect 32220 1547 32513 1581
rect 32547 1547 32849 1581
rect 32883 1547 33185 1581
rect 33219 1547 33521 1581
rect 33555 1547 33848 1581
rect 33900 1547 34193 1581
rect 34227 1547 34529 1581
rect 34563 1547 34865 1581
rect 34899 1547 35201 1581
rect 35235 1547 35528 1581
rect 35580 1547 35873 1581
rect 35907 1547 36209 1581
rect 36243 1547 36545 1581
rect 36579 1547 36881 1581
rect 36915 1547 37208 1581
rect 37260 1547 37553 1581
rect 37587 1547 37889 1581
rect 37923 1547 38225 1581
rect 38259 1547 38561 1581
rect 38595 1547 38888 1581
rect 38940 1547 39233 1581
rect 39267 1547 39569 1581
rect 39603 1547 39905 1581
rect 39939 1547 40241 1581
rect 40275 1547 40568 1581
rect 40620 1547 40913 1581
rect 40947 1547 41249 1581
rect 41283 1547 41585 1581
rect 41619 1547 41921 1581
rect 41955 1547 42248 1581
rect 42300 1547 42593 1581
rect 42627 1547 42929 1581
rect 42963 1547 43265 1581
rect 43299 1547 43601 1581
rect 43635 1547 43928 1581
rect 43980 1547 44273 1581
rect 44307 1547 44609 1581
rect 44643 1547 44945 1581
rect 44979 1547 45281 1581
rect 45315 1547 45608 1581
rect 45660 1547 45953 1581
rect 45987 1547 46289 1581
rect 46323 1547 46625 1581
rect 46659 1547 46961 1581
rect 46995 1547 47288 1581
rect 47340 1547 47633 1581
rect 47667 1547 47969 1581
rect 48003 1547 48305 1581
rect 48339 1547 48641 1581
rect 48675 1547 48968 1581
rect 49020 1547 49313 1581
rect 49347 1547 49649 1581
rect 49683 1547 49985 1581
rect 50019 1547 50321 1581
rect 50355 1547 50648 1581
rect 50700 1547 50993 1581
rect 51027 1547 51329 1581
rect 51363 1547 51665 1581
rect 51699 1547 52001 1581
rect 52035 1547 52328 1581
rect 52380 1547 52673 1581
rect 52707 1547 53009 1581
rect 53043 1547 53345 1581
rect 53379 1547 53681 1581
rect 53715 1547 54008 1581
rect 54060 1547 54353 1581
rect 54387 1547 54689 1581
rect 54723 1547 55025 1581
rect 55059 1547 55361 1581
rect 55395 1547 55688 1581
rect 55740 1547 56033 1581
rect 56067 1547 56369 1581
rect 56403 1547 56705 1581
rect 56739 1547 57041 1581
rect 57075 1547 57368 1581
rect 57420 1547 57713 1581
rect 57747 1547 58049 1581
rect 58083 1547 58385 1581
rect 58419 1547 58721 1581
rect 58755 1547 59048 1581
rect 59100 1547 59393 1581
rect 59427 1547 59729 1581
rect 59763 1547 60065 1581
rect 60099 1547 60401 1581
rect 60435 1547 60728 1581
rect 60780 1547 61073 1581
rect 61107 1547 61409 1581
rect 61443 1547 61745 1581
rect 61779 1547 62081 1581
rect 62115 1547 62408 1581
rect 62460 1547 62753 1581
rect 62787 1547 63089 1581
rect 63123 1547 63425 1581
rect 63459 1547 63761 1581
rect 63795 1547 64088 1581
rect 64140 1547 64433 1581
rect 64467 1547 64769 1581
rect 64803 1547 65105 1581
rect 65139 1547 65441 1581
rect 65475 1547 65768 1581
rect 65820 1547 66113 1581
rect 66147 1547 66449 1581
rect 66483 1547 66785 1581
rect 66819 1547 67121 1581
rect 67155 1547 67448 1581
rect 67500 1547 67793 1581
rect 67827 1547 68129 1581
rect 68163 1547 68465 1581
rect 68499 1547 68801 1581
rect 68835 1547 69128 1581
rect 69180 1547 69473 1581
rect 69507 1547 69809 1581
rect 69843 1547 70145 1581
rect 70179 1547 70481 1581
rect 70515 1547 70808 1581
rect 70860 1547 71153 1581
rect 71187 1547 71489 1581
rect 71523 1547 71825 1581
rect 71859 1547 72161 1581
rect 72195 1547 72488 1581
rect 72540 1547 72833 1581
rect 72867 1547 73169 1581
rect 73203 1547 73505 1581
rect 73539 1547 74078 1581
rect 1980 1538 3608 1547
rect 3660 1538 5288 1547
rect 5340 1538 6968 1547
rect 7020 1538 8648 1547
rect 8700 1538 10328 1547
rect 10380 1538 12008 1547
rect 12060 1538 13688 1547
rect 13740 1538 15368 1547
rect 15420 1538 17048 1547
rect 17100 1538 18728 1547
rect 18780 1538 20408 1547
rect 20460 1538 22088 1547
rect 22140 1538 23768 1547
rect 23820 1538 25448 1547
rect 25500 1538 27128 1547
rect 27180 1538 28808 1547
rect 28860 1538 30488 1547
rect 30540 1538 32168 1547
rect 32220 1538 33848 1547
rect 33900 1538 35528 1547
rect 35580 1538 37208 1547
rect 37260 1538 38888 1547
rect 38940 1538 40568 1547
rect 40620 1538 42248 1547
rect 42300 1538 43928 1547
rect 43980 1538 45608 1547
rect 45660 1538 47288 1547
rect 47340 1538 48968 1547
rect 49020 1538 50648 1547
rect 50700 1538 52328 1547
rect 52380 1538 54008 1547
rect 54060 1538 55688 1547
rect 55740 1538 57368 1547
rect 57420 1538 59048 1547
rect 59100 1538 60728 1547
rect 60780 1538 62408 1547
rect 62460 1538 64088 1547
rect 64140 1538 65768 1547
rect 65820 1538 67448 1547
rect 67500 1538 69128 1547
rect 69180 1538 70808 1547
rect 70860 1538 72488 1547
rect 72540 1538 74078 1547
rect 1506 1452 74078 1538
<< via1 >>
rect 1928 36225 1980 36234
rect 3608 36225 3660 36234
rect 5288 36225 5340 36234
rect 6968 36225 7020 36234
rect 8648 36225 8700 36234
rect 10328 36225 10380 36234
rect 12008 36225 12060 36234
rect 13688 36225 13740 36234
rect 15368 36225 15420 36234
rect 17048 36225 17100 36234
rect 18728 36225 18780 36234
rect 20408 36225 20460 36234
rect 22088 36225 22140 36234
rect 23768 36225 23820 36234
rect 25448 36225 25500 36234
rect 27128 36225 27180 36234
rect 28808 36225 28860 36234
rect 30488 36225 30540 36234
rect 32168 36225 32220 36234
rect 33848 36225 33900 36234
rect 35528 36225 35580 36234
rect 37208 36225 37260 36234
rect 38888 36225 38940 36234
rect 40568 36225 40620 36234
rect 42248 36225 42300 36234
rect 43928 36225 43980 36234
rect 45608 36225 45660 36234
rect 47288 36225 47340 36234
rect 48968 36225 49020 36234
rect 50648 36225 50700 36234
rect 52328 36225 52380 36234
rect 54008 36225 54060 36234
rect 55688 36225 55740 36234
rect 57368 36225 57420 36234
rect 59048 36225 59100 36234
rect 60728 36225 60780 36234
rect 62408 36225 62460 36234
rect 64088 36225 64140 36234
rect 65768 36225 65820 36234
rect 67448 36225 67500 36234
rect 69128 36225 69180 36234
rect 70808 36225 70860 36234
rect 72488 36225 72540 36234
rect 1928 36191 1937 36225
rect 1937 36191 1971 36225
rect 1971 36191 1980 36225
rect 3608 36191 3617 36225
rect 3617 36191 3651 36225
rect 3651 36191 3660 36225
rect 5288 36191 5297 36225
rect 5297 36191 5331 36225
rect 5331 36191 5340 36225
rect 6968 36191 6977 36225
rect 6977 36191 7011 36225
rect 7011 36191 7020 36225
rect 8648 36191 8657 36225
rect 8657 36191 8691 36225
rect 8691 36191 8700 36225
rect 10328 36191 10337 36225
rect 10337 36191 10371 36225
rect 10371 36191 10380 36225
rect 12008 36191 12017 36225
rect 12017 36191 12051 36225
rect 12051 36191 12060 36225
rect 13688 36191 13697 36225
rect 13697 36191 13731 36225
rect 13731 36191 13740 36225
rect 15368 36191 15377 36225
rect 15377 36191 15411 36225
rect 15411 36191 15420 36225
rect 17048 36191 17057 36225
rect 17057 36191 17091 36225
rect 17091 36191 17100 36225
rect 18728 36191 18737 36225
rect 18737 36191 18771 36225
rect 18771 36191 18780 36225
rect 20408 36191 20417 36225
rect 20417 36191 20451 36225
rect 20451 36191 20460 36225
rect 22088 36191 22097 36225
rect 22097 36191 22131 36225
rect 22131 36191 22140 36225
rect 23768 36191 23777 36225
rect 23777 36191 23811 36225
rect 23811 36191 23820 36225
rect 25448 36191 25457 36225
rect 25457 36191 25491 36225
rect 25491 36191 25500 36225
rect 27128 36191 27137 36225
rect 27137 36191 27171 36225
rect 27171 36191 27180 36225
rect 28808 36191 28817 36225
rect 28817 36191 28851 36225
rect 28851 36191 28860 36225
rect 30488 36191 30497 36225
rect 30497 36191 30531 36225
rect 30531 36191 30540 36225
rect 32168 36191 32177 36225
rect 32177 36191 32211 36225
rect 32211 36191 32220 36225
rect 33848 36191 33857 36225
rect 33857 36191 33891 36225
rect 33891 36191 33900 36225
rect 35528 36191 35537 36225
rect 35537 36191 35571 36225
rect 35571 36191 35580 36225
rect 37208 36191 37217 36225
rect 37217 36191 37251 36225
rect 37251 36191 37260 36225
rect 38888 36191 38897 36225
rect 38897 36191 38931 36225
rect 38931 36191 38940 36225
rect 40568 36191 40577 36225
rect 40577 36191 40611 36225
rect 40611 36191 40620 36225
rect 42248 36191 42257 36225
rect 42257 36191 42291 36225
rect 42291 36191 42300 36225
rect 43928 36191 43937 36225
rect 43937 36191 43971 36225
rect 43971 36191 43980 36225
rect 45608 36191 45617 36225
rect 45617 36191 45651 36225
rect 45651 36191 45660 36225
rect 47288 36191 47297 36225
rect 47297 36191 47331 36225
rect 47331 36191 47340 36225
rect 48968 36191 48977 36225
rect 48977 36191 49011 36225
rect 49011 36191 49020 36225
rect 50648 36191 50657 36225
rect 50657 36191 50691 36225
rect 50691 36191 50700 36225
rect 52328 36191 52337 36225
rect 52337 36191 52371 36225
rect 52371 36191 52380 36225
rect 54008 36191 54017 36225
rect 54017 36191 54051 36225
rect 54051 36191 54060 36225
rect 55688 36191 55697 36225
rect 55697 36191 55731 36225
rect 55731 36191 55740 36225
rect 57368 36191 57377 36225
rect 57377 36191 57411 36225
rect 57411 36191 57420 36225
rect 59048 36191 59057 36225
rect 59057 36191 59091 36225
rect 59091 36191 59100 36225
rect 60728 36191 60737 36225
rect 60737 36191 60771 36225
rect 60771 36191 60780 36225
rect 62408 36191 62417 36225
rect 62417 36191 62451 36225
rect 62451 36191 62460 36225
rect 64088 36191 64097 36225
rect 64097 36191 64131 36225
rect 64131 36191 64140 36225
rect 65768 36191 65777 36225
rect 65777 36191 65811 36225
rect 65811 36191 65820 36225
rect 67448 36191 67457 36225
rect 67457 36191 67491 36225
rect 67491 36191 67500 36225
rect 69128 36191 69137 36225
rect 69137 36191 69171 36225
rect 69171 36191 69180 36225
rect 70808 36191 70817 36225
rect 70817 36191 70851 36225
rect 70851 36191 70860 36225
rect 72488 36191 72497 36225
rect 72497 36191 72531 36225
rect 72531 36191 72540 36225
rect 1928 36182 1980 36191
rect 3608 36182 3660 36191
rect 5288 36182 5340 36191
rect 6968 36182 7020 36191
rect 8648 36182 8700 36191
rect 10328 36182 10380 36191
rect 12008 36182 12060 36191
rect 13688 36182 13740 36191
rect 15368 36182 15420 36191
rect 17048 36182 17100 36191
rect 18728 36182 18780 36191
rect 20408 36182 20460 36191
rect 22088 36182 22140 36191
rect 23768 36182 23820 36191
rect 25448 36182 25500 36191
rect 27128 36182 27180 36191
rect 28808 36182 28860 36191
rect 30488 36182 30540 36191
rect 32168 36182 32220 36191
rect 33848 36182 33900 36191
rect 35528 36182 35580 36191
rect 37208 36182 37260 36191
rect 38888 36182 38940 36191
rect 40568 36182 40620 36191
rect 42248 36182 42300 36191
rect 43928 36182 43980 36191
rect 45608 36182 45660 36191
rect 47288 36182 47340 36191
rect 48968 36182 49020 36191
rect 50648 36182 50700 36191
rect 52328 36182 52380 36191
rect 54008 36182 54060 36191
rect 55688 36182 55740 36191
rect 57368 36182 57420 36191
rect 59048 36182 59100 36191
rect 60728 36182 60780 36191
rect 62408 36182 62460 36191
rect 64088 36182 64140 36191
rect 65768 36182 65820 36191
rect 67448 36182 67500 36191
rect 69128 36182 69180 36191
rect 70808 36182 70860 36191
rect 72488 36182 72540 36191
rect 1592 35853 1644 35862
rect 1592 35819 1601 35853
rect 1601 35819 1635 35853
rect 1635 35819 1644 35853
rect 73940 35853 73992 35862
rect 1592 35810 1644 35819
rect 73940 35819 73949 35853
rect 73949 35819 73983 35853
rect 73983 35819 73992 35853
rect 73940 35810 73992 35819
rect 1592 35517 1644 35526
rect 1592 35483 1601 35517
rect 1601 35483 1635 35517
rect 1635 35483 1644 35517
rect 73940 35517 73992 35526
rect 1592 35474 1644 35483
rect 73940 35483 73949 35517
rect 73949 35483 73983 35517
rect 73983 35483 73992 35517
rect 73940 35474 73992 35483
rect 1592 35181 1644 35190
rect 1592 35147 1601 35181
rect 1601 35147 1635 35181
rect 1635 35147 1644 35181
rect 73940 35181 73992 35190
rect 1592 35138 1644 35147
rect 73940 35147 73949 35181
rect 73949 35147 73983 35181
rect 73983 35147 73992 35181
rect 73940 35138 73992 35147
rect 1592 34845 1644 34854
rect 1592 34811 1601 34845
rect 1601 34811 1635 34845
rect 1635 34811 1644 34845
rect 73940 34845 73992 34854
rect 1592 34802 1644 34811
rect 73940 34811 73949 34845
rect 73949 34811 73983 34845
rect 73983 34811 73992 34845
rect 73940 34802 73992 34811
rect 1592 34509 1644 34518
rect 1592 34475 1601 34509
rect 1601 34475 1635 34509
rect 1635 34475 1644 34509
rect 73940 34509 73992 34518
rect 1592 34466 1644 34475
rect 73940 34475 73949 34509
rect 73949 34475 73983 34509
rect 73983 34475 73992 34509
rect 73940 34466 73992 34475
rect 1592 34173 1644 34182
rect 1592 34139 1601 34173
rect 1601 34139 1635 34173
rect 1635 34139 1644 34173
rect 73940 34173 73992 34182
rect 1592 34130 1644 34139
rect 73940 34139 73949 34173
rect 73949 34139 73983 34173
rect 73983 34139 73992 34173
rect 73940 34130 73992 34139
rect 1592 33837 1644 33846
rect 1592 33803 1601 33837
rect 1601 33803 1635 33837
rect 1635 33803 1644 33837
rect 73940 33837 73992 33846
rect 1592 33794 1644 33803
rect 73940 33803 73949 33837
rect 73949 33803 73983 33837
rect 73983 33803 73992 33837
rect 73940 33794 73992 33803
rect 1592 33501 1644 33510
rect 1592 33467 1601 33501
rect 1601 33467 1635 33501
rect 1635 33467 1644 33501
rect 73940 33501 73992 33510
rect 1592 33458 1644 33467
rect 73940 33467 73949 33501
rect 73949 33467 73983 33501
rect 73983 33467 73992 33501
rect 73940 33458 73992 33467
rect 1592 33165 1644 33174
rect 1592 33131 1601 33165
rect 1601 33131 1635 33165
rect 1635 33131 1644 33165
rect 73940 33165 73992 33174
rect 1592 33122 1644 33131
rect 73940 33131 73949 33165
rect 73949 33131 73983 33165
rect 73983 33131 73992 33165
rect 73940 33122 73992 33131
rect 1592 32829 1644 32838
rect 1592 32795 1601 32829
rect 1601 32795 1635 32829
rect 1635 32795 1644 32829
rect 73940 32829 73992 32838
rect 1592 32786 1644 32795
rect 73940 32795 73949 32829
rect 73949 32795 73983 32829
rect 73983 32795 73992 32829
rect 73940 32786 73992 32795
rect 1592 32493 1644 32502
rect 1592 32459 1601 32493
rect 1601 32459 1635 32493
rect 1635 32459 1644 32493
rect 73940 32493 73992 32502
rect 1592 32450 1644 32459
rect 73940 32459 73949 32493
rect 73949 32459 73983 32493
rect 73983 32459 73992 32493
rect 73940 32450 73992 32459
rect 1592 32157 1644 32166
rect 1592 32123 1601 32157
rect 1601 32123 1635 32157
rect 1635 32123 1644 32157
rect 73940 32157 73992 32166
rect 1592 32114 1644 32123
rect 73940 32123 73949 32157
rect 73949 32123 73983 32157
rect 73983 32123 73992 32157
rect 73940 32114 73992 32123
rect 1592 31821 1644 31830
rect 1592 31787 1601 31821
rect 1601 31787 1635 31821
rect 1635 31787 1644 31821
rect 73940 31821 73992 31830
rect 1592 31778 1644 31787
rect 73940 31787 73949 31821
rect 73949 31787 73983 31821
rect 73983 31787 73992 31821
rect 73940 31778 73992 31787
rect 1592 31485 1644 31494
rect 1592 31451 1601 31485
rect 1601 31451 1635 31485
rect 1635 31451 1644 31485
rect 73940 31485 73992 31494
rect 1592 31442 1644 31451
rect 73940 31451 73949 31485
rect 73949 31451 73983 31485
rect 73983 31451 73992 31485
rect 73940 31442 73992 31451
rect 1592 31149 1644 31158
rect 1592 31115 1601 31149
rect 1601 31115 1635 31149
rect 1635 31115 1644 31149
rect 73940 31149 73992 31158
rect 1592 31106 1644 31115
rect 73940 31115 73949 31149
rect 73949 31115 73983 31149
rect 73983 31115 73992 31149
rect 73940 31106 73992 31115
rect 1592 30813 1644 30822
rect 1592 30779 1601 30813
rect 1601 30779 1635 30813
rect 1635 30779 1644 30813
rect 73940 30813 73992 30822
rect 1592 30770 1644 30779
rect 73940 30779 73949 30813
rect 73949 30779 73983 30813
rect 73983 30779 73992 30813
rect 73940 30770 73992 30779
rect 1592 30477 1644 30486
rect 1592 30443 1601 30477
rect 1601 30443 1635 30477
rect 1635 30443 1644 30477
rect 73940 30477 73992 30486
rect 1592 30434 1644 30443
rect 73940 30443 73949 30477
rect 73949 30443 73983 30477
rect 73983 30443 73992 30477
rect 73940 30434 73992 30443
rect 1592 30141 1644 30150
rect 1592 30107 1601 30141
rect 1601 30107 1635 30141
rect 1635 30107 1644 30141
rect 73940 30141 73992 30150
rect 1592 30098 1644 30107
rect 73940 30107 73949 30141
rect 73949 30107 73983 30141
rect 73983 30107 73992 30141
rect 73940 30098 73992 30107
rect 1592 29805 1644 29814
rect 1592 29771 1601 29805
rect 1601 29771 1635 29805
rect 1635 29771 1644 29805
rect 73940 29805 73992 29814
rect 1592 29762 1644 29771
rect 73940 29771 73949 29805
rect 73949 29771 73983 29805
rect 73983 29771 73992 29805
rect 73940 29762 73992 29771
rect 1592 29469 1644 29478
rect 1592 29435 1601 29469
rect 1601 29435 1635 29469
rect 1635 29435 1644 29469
rect 73940 29469 73992 29478
rect 1592 29426 1644 29435
rect 73940 29435 73949 29469
rect 73949 29435 73983 29469
rect 73983 29435 73992 29469
rect 73940 29426 73992 29435
rect 1592 29133 1644 29142
rect 1592 29099 1601 29133
rect 1601 29099 1635 29133
rect 1635 29099 1644 29133
rect 73940 29133 73992 29142
rect 1592 29090 1644 29099
rect 73940 29099 73949 29133
rect 73949 29099 73983 29133
rect 73983 29099 73992 29133
rect 73940 29090 73992 29099
rect 1592 28797 1644 28806
rect 1592 28763 1601 28797
rect 1601 28763 1635 28797
rect 1635 28763 1644 28797
rect 73940 28797 73992 28806
rect 1592 28754 1644 28763
rect 73940 28763 73949 28797
rect 73949 28763 73983 28797
rect 73983 28763 73992 28797
rect 73940 28754 73992 28763
rect 1592 28461 1644 28470
rect 1592 28427 1601 28461
rect 1601 28427 1635 28461
rect 1635 28427 1644 28461
rect 73940 28461 73992 28470
rect 1592 28418 1644 28427
rect 73940 28427 73949 28461
rect 73949 28427 73983 28461
rect 73983 28427 73992 28461
rect 73940 28418 73992 28427
rect 1592 28125 1644 28134
rect 1592 28091 1601 28125
rect 1601 28091 1635 28125
rect 1635 28091 1644 28125
rect 73940 28125 73992 28134
rect 1592 28082 1644 28091
rect 73940 28091 73949 28125
rect 73949 28091 73983 28125
rect 73983 28091 73992 28125
rect 73940 28082 73992 28091
rect 1592 27789 1644 27798
rect 1592 27755 1601 27789
rect 1601 27755 1635 27789
rect 1635 27755 1644 27789
rect 73940 27789 73992 27798
rect 1592 27746 1644 27755
rect 73940 27755 73949 27789
rect 73949 27755 73983 27789
rect 73983 27755 73992 27789
rect 73940 27746 73992 27755
rect 1592 27453 1644 27462
rect 1592 27419 1601 27453
rect 1601 27419 1635 27453
rect 1635 27419 1644 27453
rect 73940 27453 73992 27462
rect 1592 27410 1644 27419
rect 73940 27419 73949 27453
rect 73949 27419 73983 27453
rect 73983 27419 73992 27453
rect 73940 27410 73992 27419
rect 1592 27117 1644 27126
rect 1592 27083 1601 27117
rect 1601 27083 1635 27117
rect 1635 27083 1644 27117
rect 73940 27117 73992 27126
rect 1592 27074 1644 27083
rect 73940 27083 73949 27117
rect 73949 27083 73983 27117
rect 73983 27083 73992 27117
rect 73940 27074 73992 27083
rect 1592 26781 1644 26790
rect 1592 26747 1601 26781
rect 1601 26747 1635 26781
rect 1635 26747 1644 26781
rect 73940 26781 73992 26790
rect 1592 26738 1644 26747
rect 73940 26747 73949 26781
rect 73949 26747 73983 26781
rect 73983 26747 73992 26781
rect 73940 26738 73992 26747
rect 1592 26445 1644 26454
rect 1592 26411 1601 26445
rect 1601 26411 1635 26445
rect 1635 26411 1644 26445
rect 73940 26445 73992 26454
rect 1592 26402 1644 26411
rect 73940 26411 73949 26445
rect 73949 26411 73983 26445
rect 73983 26411 73992 26445
rect 73940 26402 73992 26411
rect 1592 26109 1644 26118
rect 1592 26075 1601 26109
rect 1601 26075 1635 26109
rect 1635 26075 1644 26109
rect 73940 26109 73992 26118
rect 1592 26066 1644 26075
rect 73940 26075 73949 26109
rect 73949 26075 73983 26109
rect 73983 26075 73992 26109
rect 73940 26066 73992 26075
rect 1592 25773 1644 25782
rect 1592 25739 1601 25773
rect 1601 25739 1635 25773
rect 1635 25739 1644 25773
rect 73940 25773 73992 25782
rect 1592 25730 1644 25739
rect 73940 25739 73949 25773
rect 73949 25739 73983 25773
rect 73983 25739 73992 25773
rect 73940 25730 73992 25739
rect 1592 25437 1644 25446
rect 1592 25403 1601 25437
rect 1601 25403 1635 25437
rect 1635 25403 1644 25437
rect 73940 25437 73992 25446
rect 1592 25394 1644 25403
rect 73940 25403 73949 25437
rect 73949 25403 73983 25437
rect 73983 25403 73992 25437
rect 73940 25394 73992 25403
rect 1592 25101 1644 25110
rect 1592 25067 1601 25101
rect 1601 25067 1635 25101
rect 1635 25067 1644 25101
rect 73940 25101 73992 25110
rect 1592 25058 1644 25067
rect 73940 25067 73949 25101
rect 73949 25067 73983 25101
rect 73983 25067 73992 25101
rect 73940 25058 73992 25067
rect 1592 24765 1644 24774
rect 1592 24731 1601 24765
rect 1601 24731 1635 24765
rect 1635 24731 1644 24765
rect 73940 24765 73992 24774
rect 1592 24722 1644 24731
rect 73940 24731 73949 24765
rect 73949 24731 73983 24765
rect 73983 24731 73992 24765
rect 73940 24722 73992 24731
rect 1592 24429 1644 24438
rect 1592 24395 1601 24429
rect 1601 24395 1635 24429
rect 1635 24395 1644 24429
rect 73940 24429 73992 24438
rect 1592 24386 1644 24395
rect 73940 24395 73949 24429
rect 73949 24395 73983 24429
rect 73983 24395 73992 24429
rect 73940 24386 73992 24395
rect 1592 24093 1644 24102
rect 1592 24059 1601 24093
rect 1601 24059 1635 24093
rect 1635 24059 1644 24093
rect 73940 24093 73992 24102
rect 1592 24050 1644 24059
rect 73940 24059 73949 24093
rect 73949 24059 73983 24093
rect 73983 24059 73992 24093
rect 73940 24050 73992 24059
rect 1592 23757 1644 23766
rect 1592 23723 1601 23757
rect 1601 23723 1635 23757
rect 1635 23723 1644 23757
rect 73940 23757 73992 23766
rect 1592 23714 1644 23723
rect 73940 23723 73949 23757
rect 73949 23723 73983 23757
rect 73983 23723 73992 23757
rect 73940 23714 73992 23723
rect 1592 23421 1644 23430
rect 1592 23387 1601 23421
rect 1601 23387 1635 23421
rect 1635 23387 1644 23421
rect 73940 23421 73992 23430
rect 1592 23378 1644 23387
rect 73940 23387 73949 23421
rect 73949 23387 73983 23421
rect 73983 23387 73992 23421
rect 73940 23378 73992 23387
rect 1592 23085 1644 23094
rect 1592 23051 1601 23085
rect 1601 23051 1635 23085
rect 1635 23051 1644 23085
rect 73940 23085 73992 23094
rect 1592 23042 1644 23051
rect 73940 23051 73949 23085
rect 73949 23051 73983 23085
rect 73983 23051 73992 23085
rect 73940 23042 73992 23051
rect 1592 22749 1644 22758
rect 1592 22715 1601 22749
rect 1601 22715 1635 22749
rect 1635 22715 1644 22749
rect 73940 22749 73992 22758
rect 1592 22706 1644 22715
rect 73940 22715 73949 22749
rect 73949 22715 73983 22749
rect 73983 22715 73992 22749
rect 73940 22706 73992 22715
rect 1592 22413 1644 22422
rect 1592 22379 1601 22413
rect 1601 22379 1635 22413
rect 1635 22379 1644 22413
rect 73940 22413 73992 22422
rect 1592 22370 1644 22379
rect 73940 22379 73949 22413
rect 73949 22379 73983 22413
rect 73983 22379 73992 22413
rect 73940 22370 73992 22379
rect 1592 22077 1644 22086
rect 1592 22043 1601 22077
rect 1601 22043 1635 22077
rect 1635 22043 1644 22077
rect 73940 22077 73992 22086
rect 1592 22034 1644 22043
rect 73940 22043 73949 22077
rect 73949 22043 73983 22077
rect 73983 22043 73992 22077
rect 73940 22034 73992 22043
rect 1592 21741 1644 21750
rect 1592 21707 1601 21741
rect 1601 21707 1635 21741
rect 1635 21707 1644 21741
rect 73940 21741 73992 21750
rect 1592 21698 1644 21707
rect 73940 21707 73949 21741
rect 73949 21707 73983 21741
rect 73983 21707 73992 21741
rect 73940 21698 73992 21707
rect 1592 21405 1644 21414
rect 1592 21371 1601 21405
rect 1601 21371 1635 21405
rect 1635 21371 1644 21405
rect 73940 21405 73992 21414
rect 1592 21362 1644 21371
rect 73940 21371 73949 21405
rect 73949 21371 73983 21405
rect 73983 21371 73992 21405
rect 73940 21362 73992 21371
rect 1592 21069 1644 21078
rect 1592 21035 1601 21069
rect 1601 21035 1635 21069
rect 1635 21035 1644 21069
rect 73940 21069 73992 21078
rect 1592 21026 1644 21035
rect 73940 21035 73949 21069
rect 73949 21035 73983 21069
rect 73983 21035 73992 21069
rect 73940 21026 73992 21035
rect 1592 20733 1644 20742
rect 1592 20699 1601 20733
rect 1601 20699 1635 20733
rect 1635 20699 1644 20733
rect 73940 20733 73992 20742
rect 1592 20690 1644 20699
rect 73940 20699 73949 20733
rect 73949 20699 73983 20733
rect 73983 20699 73992 20733
rect 73940 20690 73992 20699
rect 1592 20397 1644 20406
rect 1592 20363 1601 20397
rect 1601 20363 1635 20397
rect 1635 20363 1644 20397
rect 73940 20397 73992 20406
rect 1592 20354 1644 20363
rect 73940 20363 73949 20397
rect 73949 20363 73983 20397
rect 73983 20363 73992 20397
rect 73940 20354 73992 20363
rect 1592 20061 1644 20070
rect 1592 20027 1601 20061
rect 1601 20027 1635 20061
rect 1635 20027 1644 20061
rect 73940 20061 73992 20070
rect 1592 20018 1644 20027
rect 73940 20027 73949 20061
rect 73949 20027 73983 20061
rect 73983 20027 73992 20061
rect 73940 20018 73992 20027
rect 1592 19725 1644 19734
rect 1592 19691 1601 19725
rect 1601 19691 1635 19725
rect 1635 19691 1644 19725
rect 73940 19725 73992 19734
rect 1592 19682 1644 19691
rect 73940 19691 73949 19725
rect 73949 19691 73983 19725
rect 73983 19691 73992 19725
rect 73940 19682 73992 19691
rect 1592 19389 1644 19398
rect 1592 19355 1601 19389
rect 1601 19355 1635 19389
rect 1635 19355 1644 19389
rect 73940 19389 73992 19398
rect 1592 19346 1644 19355
rect 73940 19355 73949 19389
rect 73949 19355 73983 19389
rect 73983 19355 73992 19389
rect 73940 19346 73992 19355
rect 1592 19053 1644 19062
rect 1592 19019 1601 19053
rect 1601 19019 1635 19053
rect 1635 19019 1644 19053
rect 73940 19053 73992 19062
rect 1592 19010 1644 19019
rect 73940 19019 73949 19053
rect 73949 19019 73983 19053
rect 73983 19019 73992 19053
rect 73940 19010 73992 19019
rect 1592 18717 1644 18726
rect 1592 18683 1601 18717
rect 1601 18683 1635 18717
rect 1635 18683 1644 18717
rect 73940 18717 73992 18726
rect 1592 18674 1644 18683
rect 73940 18683 73949 18717
rect 73949 18683 73983 18717
rect 73983 18683 73992 18717
rect 73940 18674 73992 18683
rect 1592 18381 1644 18390
rect 1592 18347 1601 18381
rect 1601 18347 1635 18381
rect 1635 18347 1644 18381
rect 73940 18381 73992 18390
rect 1592 18338 1644 18347
rect 73940 18347 73949 18381
rect 73949 18347 73983 18381
rect 73983 18347 73992 18381
rect 73940 18338 73992 18347
rect 1592 18045 1644 18054
rect 1592 18011 1601 18045
rect 1601 18011 1635 18045
rect 1635 18011 1644 18045
rect 73940 18045 73992 18054
rect 1592 18002 1644 18011
rect 73940 18011 73949 18045
rect 73949 18011 73983 18045
rect 73983 18011 73992 18045
rect 73940 18002 73992 18011
rect 1592 17709 1644 17718
rect 1592 17675 1601 17709
rect 1601 17675 1635 17709
rect 1635 17675 1644 17709
rect 73940 17709 73992 17718
rect 1592 17666 1644 17675
rect 73940 17675 73949 17709
rect 73949 17675 73983 17709
rect 73983 17675 73992 17709
rect 73940 17666 73992 17675
rect 1592 17373 1644 17382
rect 1592 17339 1601 17373
rect 1601 17339 1635 17373
rect 1635 17339 1644 17373
rect 73940 17373 73992 17382
rect 1592 17330 1644 17339
rect 73940 17339 73949 17373
rect 73949 17339 73983 17373
rect 73983 17339 73992 17373
rect 73940 17330 73992 17339
rect 1592 17037 1644 17046
rect 1592 17003 1601 17037
rect 1601 17003 1635 17037
rect 1635 17003 1644 17037
rect 73940 17037 73992 17046
rect 1592 16994 1644 17003
rect 73940 17003 73949 17037
rect 73949 17003 73983 17037
rect 73983 17003 73992 17037
rect 73940 16994 73992 17003
rect 1592 16701 1644 16710
rect 1592 16667 1601 16701
rect 1601 16667 1635 16701
rect 1635 16667 1644 16701
rect 73940 16701 73992 16710
rect 1592 16658 1644 16667
rect 73940 16667 73949 16701
rect 73949 16667 73983 16701
rect 73983 16667 73992 16701
rect 73940 16658 73992 16667
rect 1592 16365 1644 16374
rect 1592 16331 1601 16365
rect 1601 16331 1635 16365
rect 1635 16331 1644 16365
rect 73940 16365 73992 16374
rect 1592 16322 1644 16331
rect 73940 16331 73949 16365
rect 73949 16331 73983 16365
rect 73983 16331 73992 16365
rect 73940 16322 73992 16331
rect 1592 16029 1644 16038
rect 1592 15995 1601 16029
rect 1601 15995 1635 16029
rect 1635 15995 1644 16029
rect 73940 16029 73992 16038
rect 1592 15986 1644 15995
rect 73940 15995 73949 16029
rect 73949 15995 73983 16029
rect 73983 15995 73992 16029
rect 73940 15986 73992 15995
rect 1592 15693 1644 15702
rect 1592 15659 1601 15693
rect 1601 15659 1635 15693
rect 1635 15659 1644 15693
rect 73940 15693 73992 15702
rect 1592 15650 1644 15659
rect 73940 15659 73949 15693
rect 73949 15659 73983 15693
rect 73983 15659 73992 15693
rect 73940 15650 73992 15659
rect 1592 15357 1644 15366
rect 1592 15323 1601 15357
rect 1601 15323 1635 15357
rect 1635 15323 1644 15357
rect 73940 15357 73992 15366
rect 1592 15314 1644 15323
rect 73940 15323 73949 15357
rect 73949 15323 73983 15357
rect 73983 15323 73992 15357
rect 73940 15314 73992 15323
rect 1592 15021 1644 15030
rect 1592 14987 1601 15021
rect 1601 14987 1635 15021
rect 1635 14987 1644 15021
rect 73940 15021 73992 15030
rect 1592 14978 1644 14987
rect 73940 14987 73949 15021
rect 73949 14987 73983 15021
rect 73983 14987 73992 15021
rect 73940 14978 73992 14987
rect 1592 14685 1644 14694
rect 1592 14651 1601 14685
rect 1601 14651 1635 14685
rect 1635 14651 1644 14685
rect 73940 14685 73992 14694
rect 1592 14642 1644 14651
rect 73940 14651 73949 14685
rect 73949 14651 73983 14685
rect 73983 14651 73992 14685
rect 73940 14642 73992 14651
rect 1592 14349 1644 14358
rect 1592 14315 1601 14349
rect 1601 14315 1635 14349
rect 1635 14315 1644 14349
rect 73940 14349 73992 14358
rect 1592 14306 1644 14315
rect 73940 14315 73949 14349
rect 73949 14315 73983 14349
rect 73983 14315 73992 14349
rect 73940 14306 73992 14315
rect 1592 14013 1644 14022
rect 1592 13979 1601 14013
rect 1601 13979 1635 14013
rect 1635 13979 1644 14013
rect 73940 14013 73992 14022
rect 1592 13970 1644 13979
rect 73940 13979 73949 14013
rect 73949 13979 73983 14013
rect 73983 13979 73992 14013
rect 73940 13970 73992 13979
rect 1592 13677 1644 13686
rect 1592 13643 1601 13677
rect 1601 13643 1635 13677
rect 1635 13643 1644 13677
rect 73940 13677 73992 13686
rect 1592 13634 1644 13643
rect 73940 13643 73949 13677
rect 73949 13643 73983 13677
rect 73983 13643 73992 13677
rect 73940 13634 73992 13643
rect 1592 13341 1644 13350
rect 1592 13307 1601 13341
rect 1601 13307 1635 13341
rect 1635 13307 1644 13341
rect 73940 13341 73992 13350
rect 1592 13298 1644 13307
rect 73940 13307 73949 13341
rect 73949 13307 73983 13341
rect 73983 13307 73992 13341
rect 73940 13298 73992 13307
rect 1592 13005 1644 13014
rect 1592 12971 1601 13005
rect 1601 12971 1635 13005
rect 1635 12971 1644 13005
rect 73940 13005 73992 13014
rect 1592 12962 1644 12971
rect 73940 12971 73949 13005
rect 73949 12971 73983 13005
rect 73983 12971 73992 13005
rect 73940 12962 73992 12971
rect 1592 12669 1644 12678
rect 1592 12635 1601 12669
rect 1601 12635 1635 12669
rect 1635 12635 1644 12669
rect 73940 12669 73992 12678
rect 1592 12626 1644 12635
rect 73940 12635 73949 12669
rect 73949 12635 73983 12669
rect 73983 12635 73992 12669
rect 73940 12626 73992 12635
rect 1592 12333 1644 12342
rect 1592 12299 1601 12333
rect 1601 12299 1635 12333
rect 1635 12299 1644 12333
rect 73940 12333 73992 12342
rect 1592 12290 1644 12299
rect 73940 12299 73949 12333
rect 73949 12299 73983 12333
rect 73983 12299 73992 12333
rect 73940 12290 73992 12299
rect 1592 11997 1644 12006
rect 1592 11963 1601 11997
rect 1601 11963 1635 11997
rect 1635 11963 1644 11997
rect 73940 11997 73992 12006
rect 1592 11954 1644 11963
rect 73940 11963 73949 11997
rect 73949 11963 73983 11997
rect 73983 11963 73992 11997
rect 73940 11954 73992 11963
rect 1592 11661 1644 11670
rect 1592 11627 1601 11661
rect 1601 11627 1635 11661
rect 1635 11627 1644 11661
rect 73940 11661 73992 11670
rect 1592 11618 1644 11627
rect 73940 11627 73949 11661
rect 73949 11627 73983 11661
rect 73983 11627 73992 11661
rect 73940 11618 73992 11627
rect 1592 11325 1644 11334
rect 1592 11291 1601 11325
rect 1601 11291 1635 11325
rect 1635 11291 1644 11325
rect 73940 11325 73992 11334
rect 1592 11282 1644 11291
rect 73940 11291 73949 11325
rect 73949 11291 73983 11325
rect 73983 11291 73992 11325
rect 73940 11282 73992 11291
rect 1592 10989 1644 10998
rect 1592 10955 1601 10989
rect 1601 10955 1635 10989
rect 1635 10955 1644 10989
rect 73940 10989 73992 10998
rect 1592 10946 1644 10955
rect 73940 10955 73949 10989
rect 73949 10955 73983 10989
rect 73983 10955 73992 10989
rect 73940 10946 73992 10955
rect 1592 10653 1644 10662
rect 1592 10619 1601 10653
rect 1601 10619 1635 10653
rect 1635 10619 1644 10653
rect 73940 10653 73992 10662
rect 1592 10610 1644 10619
rect 73940 10619 73949 10653
rect 73949 10619 73983 10653
rect 73983 10619 73992 10653
rect 73940 10610 73992 10619
rect 1592 10317 1644 10326
rect 1592 10283 1601 10317
rect 1601 10283 1635 10317
rect 1635 10283 1644 10317
rect 73940 10317 73992 10326
rect 1592 10274 1644 10283
rect 73940 10283 73949 10317
rect 73949 10283 73983 10317
rect 73983 10283 73992 10317
rect 73940 10274 73992 10283
rect 1592 9981 1644 9990
rect 1592 9947 1601 9981
rect 1601 9947 1635 9981
rect 1635 9947 1644 9981
rect 73940 9981 73992 9990
rect 1592 9938 1644 9947
rect 73940 9947 73949 9981
rect 73949 9947 73983 9981
rect 73983 9947 73992 9981
rect 73940 9938 73992 9947
rect 1592 9645 1644 9654
rect 1592 9611 1601 9645
rect 1601 9611 1635 9645
rect 1635 9611 1644 9645
rect 73940 9645 73992 9654
rect 1592 9602 1644 9611
rect 73940 9611 73949 9645
rect 73949 9611 73983 9645
rect 73983 9611 73992 9645
rect 73940 9602 73992 9611
rect 1592 9309 1644 9318
rect 1592 9275 1601 9309
rect 1601 9275 1635 9309
rect 1635 9275 1644 9309
rect 73940 9309 73992 9318
rect 1592 9266 1644 9275
rect 73940 9275 73949 9309
rect 73949 9275 73983 9309
rect 73983 9275 73992 9309
rect 73940 9266 73992 9275
rect 1592 8973 1644 8982
rect 1592 8939 1601 8973
rect 1601 8939 1635 8973
rect 1635 8939 1644 8973
rect 73940 8973 73992 8982
rect 1592 8930 1644 8939
rect 73940 8939 73949 8973
rect 73949 8939 73983 8973
rect 73983 8939 73992 8973
rect 73940 8930 73992 8939
rect 1592 8637 1644 8646
rect 1592 8603 1601 8637
rect 1601 8603 1635 8637
rect 1635 8603 1644 8637
rect 73940 8637 73992 8646
rect 1592 8594 1644 8603
rect 73940 8603 73949 8637
rect 73949 8603 73983 8637
rect 73983 8603 73992 8637
rect 73940 8594 73992 8603
rect 1592 8301 1644 8310
rect 1592 8267 1601 8301
rect 1601 8267 1635 8301
rect 1635 8267 1644 8301
rect 73940 8301 73992 8310
rect 1592 8258 1644 8267
rect 73940 8267 73949 8301
rect 73949 8267 73983 8301
rect 73983 8267 73992 8301
rect 73940 8258 73992 8267
rect 1592 7965 1644 7974
rect 1592 7931 1601 7965
rect 1601 7931 1635 7965
rect 1635 7931 1644 7965
rect 73940 7965 73992 7974
rect 1592 7922 1644 7931
rect 73940 7931 73949 7965
rect 73949 7931 73983 7965
rect 73983 7931 73992 7965
rect 73940 7922 73992 7931
rect 1592 7629 1644 7638
rect 1592 7595 1601 7629
rect 1601 7595 1635 7629
rect 1635 7595 1644 7629
rect 73940 7629 73992 7638
rect 1592 7586 1644 7595
rect 73940 7595 73949 7629
rect 73949 7595 73983 7629
rect 73983 7595 73992 7629
rect 73940 7586 73992 7595
rect 1592 7293 1644 7302
rect 1592 7259 1601 7293
rect 1601 7259 1635 7293
rect 1635 7259 1644 7293
rect 73940 7293 73992 7302
rect 1592 7250 1644 7259
rect 73940 7259 73949 7293
rect 73949 7259 73983 7293
rect 73983 7259 73992 7293
rect 73940 7250 73992 7259
rect 1592 6957 1644 6966
rect 1592 6923 1601 6957
rect 1601 6923 1635 6957
rect 1635 6923 1644 6957
rect 73940 6957 73992 6966
rect 1592 6914 1644 6923
rect 73940 6923 73949 6957
rect 73949 6923 73983 6957
rect 73983 6923 73992 6957
rect 73940 6914 73992 6923
rect 1592 6621 1644 6630
rect 1592 6587 1601 6621
rect 1601 6587 1635 6621
rect 1635 6587 1644 6621
rect 73940 6621 73992 6630
rect 1592 6578 1644 6587
rect 73940 6587 73949 6621
rect 73949 6587 73983 6621
rect 73983 6587 73992 6621
rect 73940 6578 73992 6587
rect 1592 6285 1644 6294
rect 1592 6251 1601 6285
rect 1601 6251 1635 6285
rect 1635 6251 1644 6285
rect 73940 6285 73992 6294
rect 1592 6242 1644 6251
rect 73940 6251 73949 6285
rect 73949 6251 73983 6285
rect 73983 6251 73992 6285
rect 73940 6242 73992 6251
rect 1592 5949 1644 5958
rect 1592 5915 1601 5949
rect 1601 5915 1635 5949
rect 1635 5915 1644 5949
rect 73940 5949 73992 5958
rect 1592 5906 1644 5915
rect 73940 5915 73949 5949
rect 73949 5915 73983 5949
rect 73983 5915 73992 5949
rect 73940 5906 73992 5915
rect 1592 5613 1644 5622
rect 1592 5579 1601 5613
rect 1601 5579 1635 5613
rect 1635 5579 1644 5613
rect 73940 5613 73992 5622
rect 1592 5570 1644 5579
rect 73940 5579 73949 5613
rect 73949 5579 73983 5613
rect 73983 5579 73992 5613
rect 73940 5570 73992 5579
rect 1592 5277 1644 5286
rect 1592 5243 1601 5277
rect 1601 5243 1635 5277
rect 1635 5243 1644 5277
rect 73940 5277 73992 5286
rect 1592 5234 1644 5243
rect 73940 5243 73949 5277
rect 73949 5243 73983 5277
rect 73983 5243 73992 5277
rect 73940 5234 73992 5243
rect 1592 4941 1644 4950
rect 1592 4907 1601 4941
rect 1601 4907 1635 4941
rect 1635 4907 1644 4941
rect 73940 4941 73992 4950
rect 1592 4898 1644 4907
rect 73940 4907 73949 4941
rect 73949 4907 73983 4941
rect 73983 4907 73992 4941
rect 73940 4898 73992 4907
rect 1592 4605 1644 4614
rect 1592 4571 1601 4605
rect 1601 4571 1635 4605
rect 1635 4571 1644 4605
rect 73940 4605 73992 4614
rect 1592 4562 1644 4571
rect 73940 4571 73949 4605
rect 73949 4571 73983 4605
rect 73983 4571 73992 4605
rect 73940 4562 73992 4571
rect 1592 4269 1644 4278
rect 1592 4235 1601 4269
rect 1601 4235 1635 4269
rect 1635 4235 1644 4269
rect 73940 4269 73992 4278
rect 1592 4226 1644 4235
rect 73940 4235 73949 4269
rect 73949 4235 73983 4269
rect 73983 4235 73992 4269
rect 73940 4226 73992 4235
rect 1592 3933 1644 3942
rect 1592 3899 1601 3933
rect 1601 3899 1635 3933
rect 1635 3899 1644 3933
rect 73940 3933 73992 3942
rect 1592 3890 1644 3899
rect 73940 3899 73949 3933
rect 73949 3899 73983 3933
rect 73983 3899 73992 3933
rect 73940 3890 73992 3899
rect 1592 3597 1644 3606
rect 1592 3563 1601 3597
rect 1601 3563 1635 3597
rect 1635 3563 1644 3597
rect 73940 3597 73992 3606
rect 1592 3554 1644 3563
rect 73940 3563 73949 3597
rect 73949 3563 73983 3597
rect 73983 3563 73992 3597
rect 73940 3554 73992 3563
rect 1592 3261 1644 3270
rect 1592 3227 1601 3261
rect 1601 3227 1635 3261
rect 1635 3227 1644 3261
rect 73940 3261 73992 3270
rect 1592 3218 1644 3227
rect 73940 3227 73949 3261
rect 73949 3227 73983 3261
rect 73983 3227 73992 3261
rect 73940 3218 73992 3227
rect 1592 2925 1644 2934
rect 1592 2891 1601 2925
rect 1601 2891 1635 2925
rect 1635 2891 1644 2925
rect 73940 2925 73992 2934
rect 1592 2882 1644 2891
rect 73940 2891 73949 2925
rect 73949 2891 73983 2925
rect 73983 2891 73992 2925
rect 73940 2882 73992 2891
rect 1592 2589 1644 2598
rect 1592 2555 1601 2589
rect 1601 2555 1635 2589
rect 1635 2555 1644 2589
rect 73940 2589 73992 2598
rect 1592 2546 1644 2555
rect 73940 2555 73949 2589
rect 73949 2555 73983 2589
rect 73983 2555 73992 2589
rect 73940 2546 73992 2555
rect 1592 2253 1644 2262
rect 1592 2219 1601 2253
rect 1601 2219 1635 2253
rect 1635 2219 1644 2253
rect 73940 2253 73992 2262
rect 1592 2210 1644 2219
rect 73940 2219 73949 2253
rect 73949 2219 73983 2253
rect 73983 2219 73992 2253
rect 73940 2210 73992 2219
rect 1592 1917 1644 1926
rect 1592 1883 1601 1917
rect 1601 1883 1635 1917
rect 1635 1883 1644 1917
rect 73940 1917 73992 1926
rect 1592 1874 1644 1883
rect 73940 1883 73949 1917
rect 73949 1883 73983 1917
rect 73983 1883 73992 1917
rect 73940 1874 73992 1883
rect 1928 1581 1980 1590
rect 3608 1581 3660 1590
rect 5288 1581 5340 1590
rect 6968 1581 7020 1590
rect 8648 1581 8700 1590
rect 10328 1581 10380 1590
rect 12008 1581 12060 1590
rect 13688 1581 13740 1590
rect 15368 1581 15420 1590
rect 17048 1581 17100 1590
rect 18728 1581 18780 1590
rect 20408 1581 20460 1590
rect 22088 1581 22140 1590
rect 23768 1581 23820 1590
rect 25448 1581 25500 1590
rect 27128 1581 27180 1590
rect 28808 1581 28860 1590
rect 30488 1581 30540 1590
rect 32168 1581 32220 1590
rect 33848 1581 33900 1590
rect 35528 1581 35580 1590
rect 37208 1581 37260 1590
rect 38888 1581 38940 1590
rect 40568 1581 40620 1590
rect 42248 1581 42300 1590
rect 43928 1581 43980 1590
rect 45608 1581 45660 1590
rect 47288 1581 47340 1590
rect 48968 1581 49020 1590
rect 50648 1581 50700 1590
rect 52328 1581 52380 1590
rect 54008 1581 54060 1590
rect 55688 1581 55740 1590
rect 57368 1581 57420 1590
rect 59048 1581 59100 1590
rect 60728 1581 60780 1590
rect 62408 1581 62460 1590
rect 64088 1581 64140 1590
rect 65768 1581 65820 1590
rect 67448 1581 67500 1590
rect 69128 1581 69180 1590
rect 70808 1581 70860 1590
rect 72488 1581 72540 1590
rect 1928 1547 1937 1581
rect 1937 1547 1971 1581
rect 1971 1547 1980 1581
rect 3608 1547 3617 1581
rect 3617 1547 3651 1581
rect 3651 1547 3660 1581
rect 5288 1547 5297 1581
rect 5297 1547 5331 1581
rect 5331 1547 5340 1581
rect 6968 1547 6977 1581
rect 6977 1547 7011 1581
rect 7011 1547 7020 1581
rect 8648 1547 8657 1581
rect 8657 1547 8691 1581
rect 8691 1547 8700 1581
rect 10328 1547 10337 1581
rect 10337 1547 10371 1581
rect 10371 1547 10380 1581
rect 12008 1547 12017 1581
rect 12017 1547 12051 1581
rect 12051 1547 12060 1581
rect 13688 1547 13697 1581
rect 13697 1547 13731 1581
rect 13731 1547 13740 1581
rect 15368 1547 15377 1581
rect 15377 1547 15411 1581
rect 15411 1547 15420 1581
rect 17048 1547 17057 1581
rect 17057 1547 17091 1581
rect 17091 1547 17100 1581
rect 18728 1547 18737 1581
rect 18737 1547 18771 1581
rect 18771 1547 18780 1581
rect 20408 1547 20417 1581
rect 20417 1547 20451 1581
rect 20451 1547 20460 1581
rect 22088 1547 22097 1581
rect 22097 1547 22131 1581
rect 22131 1547 22140 1581
rect 23768 1547 23777 1581
rect 23777 1547 23811 1581
rect 23811 1547 23820 1581
rect 25448 1547 25457 1581
rect 25457 1547 25491 1581
rect 25491 1547 25500 1581
rect 27128 1547 27137 1581
rect 27137 1547 27171 1581
rect 27171 1547 27180 1581
rect 28808 1547 28817 1581
rect 28817 1547 28851 1581
rect 28851 1547 28860 1581
rect 30488 1547 30497 1581
rect 30497 1547 30531 1581
rect 30531 1547 30540 1581
rect 32168 1547 32177 1581
rect 32177 1547 32211 1581
rect 32211 1547 32220 1581
rect 33848 1547 33857 1581
rect 33857 1547 33891 1581
rect 33891 1547 33900 1581
rect 35528 1547 35537 1581
rect 35537 1547 35571 1581
rect 35571 1547 35580 1581
rect 37208 1547 37217 1581
rect 37217 1547 37251 1581
rect 37251 1547 37260 1581
rect 38888 1547 38897 1581
rect 38897 1547 38931 1581
rect 38931 1547 38940 1581
rect 40568 1547 40577 1581
rect 40577 1547 40611 1581
rect 40611 1547 40620 1581
rect 42248 1547 42257 1581
rect 42257 1547 42291 1581
rect 42291 1547 42300 1581
rect 43928 1547 43937 1581
rect 43937 1547 43971 1581
rect 43971 1547 43980 1581
rect 45608 1547 45617 1581
rect 45617 1547 45651 1581
rect 45651 1547 45660 1581
rect 47288 1547 47297 1581
rect 47297 1547 47331 1581
rect 47331 1547 47340 1581
rect 48968 1547 48977 1581
rect 48977 1547 49011 1581
rect 49011 1547 49020 1581
rect 50648 1547 50657 1581
rect 50657 1547 50691 1581
rect 50691 1547 50700 1581
rect 52328 1547 52337 1581
rect 52337 1547 52371 1581
rect 52371 1547 52380 1581
rect 54008 1547 54017 1581
rect 54017 1547 54051 1581
rect 54051 1547 54060 1581
rect 55688 1547 55697 1581
rect 55697 1547 55731 1581
rect 55731 1547 55740 1581
rect 57368 1547 57377 1581
rect 57377 1547 57411 1581
rect 57411 1547 57420 1581
rect 59048 1547 59057 1581
rect 59057 1547 59091 1581
rect 59091 1547 59100 1581
rect 60728 1547 60737 1581
rect 60737 1547 60771 1581
rect 60771 1547 60780 1581
rect 62408 1547 62417 1581
rect 62417 1547 62451 1581
rect 62451 1547 62460 1581
rect 64088 1547 64097 1581
rect 64097 1547 64131 1581
rect 64131 1547 64140 1581
rect 65768 1547 65777 1581
rect 65777 1547 65811 1581
rect 65811 1547 65820 1581
rect 67448 1547 67457 1581
rect 67457 1547 67491 1581
rect 67491 1547 67500 1581
rect 69128 1547 69137 1581
rect 69137 1547 69171 1581
rect 69171 1547 69180 1581
rect 70808 1547 70817 1581
rect 70817 1547 70851 1581
rect 70851 1547 70860 1581
rect 72488 1547 72497 1581
rect 72497 1547 72531 1581
rect 72531 1547 72540 1581
rect 1928 1538 1980 1547
rect 3608 1538 3660 1547
rect 5288 1538 5340 1547
rect 6968 1538 7020 1547
rect 8648 1538 8700 1547
rect 10328 1538 10380 1547
rect 12008 1538 12060 1547
rect 13688 1538 13740 1547
rect 15368 1538 15420 1547
rect 17048 1538 17100 1547
rect 18728 1538 18780 1547
rect 20408 1538 20460 1547
rect 22088 1538 22140 1547
rect 23768 1538 23820 1547
rect 25448 1538 25500 1547
rect 27128 1538 27180 1547
rect 28808 1538 28860 1547
rect 30488 1538 30540 1547
rect 32168 1538 32220 1547
rect 33848 1538 33900 1547
rect 35528 1538 35580 1547
rect 37208 1538 37260 1547
rect 38888 1538 38940 1547
rect 40568 1538 40620 1547
rect 42248 1538 42300 1547
rect 43928 1538 43980 1547
rect 45608 1538 45660 1547
rect 47288 1538 47340 1547
rect 48968 1538 49020 1547
rect 50648 1538 50700 1547
rect 52328 1538 52380 1547
rect 54008 1538 54060 1547
rect 55688 1538 55740 1547
rect 57368 1538 57420 1547
rect 59048 1538 59100 1547
rect 60728 1538 60780 1547
rect 62408 1538 62460 1547
rect 64088 1538 64140 1547
rect 65768 1538 65820 1547
rect 67448 1538 67500 1547
rect 69128 1538 69180 1547
rect 70808 1538 70860 1547
rect 72488 1538 72540 1547
<< metal2 >>
rect 1506 35862 1730 36320
rect 1934 36236 1974 36242
rect 3614 36236 3654 36242
rect 5294 36236 5334 36242
rect 6974 36236 7014 36242
rect 8654 36236 8694 36242
rect 10334 36236 10374 36242
rect 12014 36236 12054 36242
rect 13694 36236 13734 36242
rect 15374 36236 15414 36242
rect 17054 36236 17094 36242
rect 18734 36236 18774 36242
rect 20414 36236 20454 36242
rect 22094 36236 22134 36242
rect 23774 36236 23814 36242
rect 25454 36236 25494 36242
rect 27134 36236 27174 36242
rect 28814 36236 28854 36242
rect 30494 36236 30534 36242
rect 32174 36236 32214 36242
rect 33854 36236 33894 36242
rect 35534 36236 35574 36242
rect 37214 36236 37254 36242
rect 38894 36236 38934 36242
rect 40574 36236 40614 36242
rect 42254 36236 42294 36242
rect 43934 36236 43974 36242
rect 45614 36236 45654 36242
rect 47294 36236 47334 36242
rect 48974 36236 49014 36242
rect 50654 36236 50694 36242
rect 52334 36236 52374 36242
rect 54014 36236 54054 36242
rect 55694 36236 55734 36242
rect 57374 36236 57414 36242
rect 59054 36236 59094 36242
rect 60734 36236 60774 36242
rect 62414 36236 62454 36242
rect 64094 36236 64134 36242
rect 65774 36236 65814 36242
rect 67454 36236 67494 36242
rect 69134 36236 69174 36242
rect 70814 36236 70854 36242
rect 72494 36236 72534 36242
rect 1934 36174 1974 36180
rect 3614 36174 3654 36180
rect 5294 36174 5334 36180
rect 6974 36174 7014 36180
rect 8654 36174 8694 36180
rect 10334 36174 10374 36180
rect 12014 36174 12054 36180
rect 13694 36174 13734 36180
rect 15374 36174 15414 36180
rect 17054 36174 17094 36180
rect 18734 36174 18774 36180
rect 20414 36174 20454 36180
rect 22094 36174 22134 36180
rect 23774 36174 23814 36180
rect 25454 36174 25494 36180
rect 27134 36174 27174 36180
rect 28814 36174 28854 36180
rect 30494 36174 30534 36180
rect 32174 36174 32214 36180
rect 33854 36174 33894 36180
rect 35534 36174 35574 36180
rect 37214 36174 37254 36180
rect 38894 36174 38934 36180
rect 40574 36174 40614 36180
rect 42254 36174 42294 36180
rect 43934 36174 43974 36180
rect 45614 36174 45654 36180
rect 47294 36174 47334 36180
rect 48974 36174 49014 36180
rect 50654 36174 50694 36180
rect 52334 36174 52374 36180
rect 54014 36174 54054 36180
rect 55694 36174 55734 36180
rect 57374 36174 57414 36180
rect 59054 36174 59094 36180
rect 60734 36174 60774 36180
rect 62414 36174 62454 36180
rect 64094 36174 64134 36180
rect 65774 36174 65814 36180
rect 67454 36174 67494 36180
rect 69134 36174 69174 36180
rect 70814 36174 70854 36180
rect 72494 36174 72534 36180
rect 1506 35810 1592 35862
rect 1644 35810 1730 35862
rect 1506 35528 1730 35810
rect 1506 35472 1590 35528
rect 1646 35472 1730 35528
rect 1506 35190 1730 35472
rect 73854 35862 74078 36320
rect 73854 35810 73940 35862
rect 73992 35810 74078 35862
rect 73854 35528 74078 35810
rect 73854 35472 73938 35528
rect 73994 35472 74078 35528
rect 1506 35138 1592 35190
rect 1644 35138 1730 35190
rect 1506 34854 1730 35138
rect 1506 34802 1592 34854
rect 1644 34802 1730 34854
rect 1506 34518 1730 34802
rect 1506 34466 1592 34518
rect 1644 34466 1730 34518
rect 1506 34182 1730 34466
rect 1506 34130 1592 34182
rect 1644 34130 1730 34182
rect 1506 33848 1730 34130
rect 1506 33792 1590 33848
rect 1646 33792 1730 33848
rect 1506 33510 1730 33792
rect 1506 33458 1592 33510
rect 1644 33458 1730 33510
rect 1506 33174 1730 33458
rect 1506 33122 1592 33174
rect 1644 33122 1730 33174
rect 1506 32838 1730 33122
rect 1506 32786 1592 32838
rect 1644 32786 1730 32838
rect 1506 32502 1730 32786
rect 1506 32450 1592 32502
rect 1644 32450 1730 32502
rect 1506 32168 1730 32450
rect 1506 32112 1590 32168
rect 1646 32112 1730 32168
rect 1506 31830 1730 32112
rect 1506 31778 1592 31830
rect 1644 31778 1730 31830
rect 1506 31494 1730 31778
rect 1506 31442 1592 31494
rect 1644 31442 1730 31494
rect 1506 31158 1730 31442
rect 1506 31106 1592 31158
rect 1644 31106 1730 31158
rect 1506 30822 1730 31106
rect 1506 30770 1592 30822
rect 1644 30770 1730 30822
rect 1506 30488 1730 30770
rect 1506 30432 1590 30488
rect 1646 30432 1730 30488
rect 1506 30150 1730 30432
rect 1506 30098 1592 30150
rect 1644 30098 1730 30150
rect 1506 29814 1730 30098
rect 1506 29762 1592 29814
rect 1644 29762 1730 29814
rect 1506 29478 1730 29762
rect 1506 29426 1592 29478
rect 1644 29426 1730 29478
rect 1506 29142 1730 29426
rect 1506 29090 1592 29142
rect 1644 29090 1730 29142
rect 1506 28808 1730 29090
rect 1506 28752 1590 28808
rect 1646 28752 1730 28808
rect 1506 28470 1730 28752
rect 1506 28418 1592 28470
rect 1644 28418 1730 28470
rect 1506 28134 1730 28418
rect 1506 28082 1592 28134
rect 1644 28082 1730 28134
rect 1506 27798 1730 28082
rect 1506 27746 1592 27798
rect 1644 27746 1730 27798
rect 1506 27462 1730 27746
rect 1506 27410 1592 27462
rect 1644 27410 1730 27462
rect 1506 27128 1730 27410
rect 1506 27072 1590 27128
rect 1646 27072 1730 27128
rect 1506 26790 1730 27072
rect 1506 26738 1592 26790
rect 1644 26738 1730 26790
rect 1506 26454 1730 26738
rect 1506 26402 1592 26454
rect 1644 26402 1730 26454
rect 1506 26118 1730 26402
rect 1506 26066 1592 26118
rect 1644 26066 1730 26118
rect 1506 25782 1730 26066
rect 1506 25730 1592 25782
rect 1644 25730 1730 25782
rect 1506 25448 1730 25730
rect 1506 25392 1590 25448
rect 1646 25392 1730 25448
rect 1506 25110 1730 25392
rect 1506 25058 1592 25110
rect 1644 25058 1730 25110
rect 1506 24774 1730 25058
rect 1506 24722 1592 24774
rect 1644 24722 1730 24774
rect 1506 24438 1730 24722
rect 1506 24386 1592 24438
rect 1644 24386 1730 24438
rect 1506 24102 1730 24386
rect 1506 24050 1592 24102
rect 1644 24050 1730 24102
rect 1506 23768 1730 24050
rect 1506 23712 1590 23768
rect 1646 23712 1730 23768
rect 1506 23430 1730 23712
rect 1506 23378 1592 23430
rect 1644 23378 1730 23430
rect 1506 23094 1730 23378
rect 1506 23042 1592 23094
rect 1644 23042 1730 23094
rect 1506 22758 1730 23042
rect 1506 22706 1592 22758
rect 1644 22706 1730 22758
rect 1506 22422 1730 22706
rect 1506 22370 1592 22422
rect 1644 22370 1730 22422
rect 1506 22088 1730 22370
rect 1506 22032 1590 22088
rect 1646 22032 1730 22088
rect 1506 21750 1730 22032
rect 1506 21698 1592 21750
rect 1644 21698 1730 21750
rect 1506 21414 1730 21698
rect 1506 21362 1592 21414
rect 1644 21362 1730 21414
rect 1506 21078 1730 21362
rect 1506 21026 1592 21078
rect 1644 21026 1730 21078
rect 1506 20742 1730 21026
rect 1506 20690 1592 20742
rect 1644 20690 1730 20742
rect 1506 20408 1730 20690
rect 1506 20352 1590 20408
rect 1646 20352 1730 20408
rect 1506 20070 1730 20352
rect 1506 20018 1592 20070
rect 1644 20018 1730 20070
rect 1506 19734 1730 20018
rect 1506 19682 1592 19734
rect 1644 19682 1730 19734
rect 1506 19398 1730 19682
rect 1506 19346 1592 19398
rect 1644 19346 1730 19398
rect 1506 19062 1730 19346
rect 1506 19010 1592 19062
rect 1644 19010 1730 19062
rect 1506 18728 1730 19010
rect 1506 18672 1590 18728
rect 1646 18672 1730 18728
rect 1506 18390 1730 18672
rect 1506 18338 1592 18390
rect 1644 18338 1730 18390
rect 1506 18054 1730 18338
rect 1506 18002 1592 18054
rect 1644 18002 1730 18054
rect 1506 17718 1730 18002
rect 1506 17666 1592 17718
rect 1644 17666 1730 17718
rect 1506 17382 1730 17666
rect 1506 17330 1592 17382
rect 1644 17330 1730 17382
rect 1506 17048 1730 17330
rect 1506 16992 1590 17048
rect 1646 16992 1730 17048
rect 1506 16710 1730 16992
rect 1506 16658 1592 16710
rect 1644 16658 1730 16710
rect 1506 16374 1730 16658
rect 1506 16322 1592 16374
rect 1644 16322 1730 16374
rect 1506 16038 1730 16322
rect 1506 15986 1592 16038
rect 1644 15986 1730 16038
rect 1506 15702 1730 15986
rect 1506 15650 1592 15702
rect 1644 15650 1730 15702
rect 1506 15368 1730 15650
rect 1506 15312 1590 15368
rect 1646 15312 1730 15368
rect 1506 15030 1730 15312
rect 1506 14978 1592 15030
rect 1644 14978 1730 15030
rect 1506 14694 1730 14978
rect 1506 14642 1592 14694
rect 1644 14642 1730 14694
rect 1506 14358 1730 14642
rect 1506 14306 1592 14358
rect 1644 14306 1730 14358
rect 1506 14022 1730 14306
rect 1506 13970 1592 14022
rect 1644 13970 1730 14022
rect 1506 13688 1730 13970
rect 1506 13632 1590 13688
rect 1646 13632 1730 13688
rect 1506 13350 1730 13632
rect 1506 13298 1592 13350
rect 1644 13298 1730 13350
rect 1506 13014 1730 13298
rect 1506 12962 1592 13014
rect 1644 12962 1730 13014
rect 1506 12678 1730 12962
rect 1506 12626 1592 12678
rect 1644 12626 1730 12678
rect 1506 12342 1730 12626
rect 1506 12290 1592 12342
rect 1644 12290 1730 12342
rect 1506 12008 1730 12290
rect 1506 11952 1590 12008
rect 1646 11952 1730 12008
rect 1506 11670 1730 11952
rect 1506 11618 1592 11670
rect 1644 11618 1730 11670
rect 1506 11334 1730 11618
rect 1506 11282 1592 11334
rect 1644 11282 1730 11334
rect 1506 10998 1730 11282
rect 1506 10946 1592 10998
rect 1644 10946 1730 10998
rect 1506 10662 1730 10946
rect 1506 10610 1592 10662
rect 1644 10610 1730 10662
rect 1506 10328 1730 10610
rect 1506 10272 1590 10328
rect 1646 10272 1730 10328
rect 1506 9990 1730 10272
rect 1506 9938 1592 9990
rect 1644 9938 1730 9990
rect 1506 9654 1730 9938
rect 1506 9602 1592 9654
rect 1644 9602 1730 9654
rect 1506 9318 1730 9602
rect 1506 9266 1592 9318
rect 1644 9266 1730 9318
rect 1506 8982 1730 9266
rect 1506 8930 1592 8982
rect 1644 8930 1730 8982
rect 1506 8648 1730 8930
rect 1506 8592 1590 8648
rect 1646 8592 1730 8648
rect 1506 8310 1730 8592
rect 1506 8258 1592 8310
rect 1644 8258 1730 8310
rect 1506 7974 1730 8258
rect 1506 7922 1592 7974
rect 1644 7922 1730 7974
rect 1506 7638 1730 7922
rect 1506 7586 1592 7638
rect 1644 7586 1730 7638
rect 1506 7302 1730 7586
rect 1506 7250 1592 7302
rect 1644 7250 1730 7302
rect 1506 6968 1730 7250
rect 1506 6912 1590 6968
rect 1646 6912 1730 6968
rect 1506 6630 1730 6912
rect 1506 6578 1592 6630
rect 1644 6578 1730 6630
rect 1506 6294 1730 6578
rect 1506 6242 1592 6294
rect 1644 6242 1730 6294
rect 1506 5958 1730 6242
rect 1506 5906 1592 5958
rect 1644 5906 1730 5958
rect 1506 5622 1730 5906
rect 12130 5860 12158 11032
rect 13831 11030 13859 22940
rect 13899 12222 13927 22940
rect 13967 12706 13995 22940
rect 14035 13898 14063 22940
rect 14103 14382 14131 22940
rect 14171 15574 14199 22940
rect 18492 10155 18520 35232
rect 73854 35190 74078 35472
rect 73854 35138 73940 35190
rect 73992 35138 74078 35190
rect 73854 34854 74078 35138
rect 73854 34802 73940 34854
rect 73992 34802 74078 34854
rect 73854 34518 74078 34802
rect 73854 34466 73940 34518
rect 73992 34466 74078 34518
rect 73854 34182 74078 34466
rect 73854 34130 73940 34182
rect 73992 34130 74078 34182
rect 73854 33848 74078 34130
rect 73854 33792 73938 33848
rect 73994 33792 74078 33848
rect 73854 33510 74078 33792
rect 73854 33458 73940 33510
rect 73992 33458 74078 33510
rect 73854 33174 74078 33458
rect 73854 33122 73940 33174
rect 73992 33122 74078 33174
rect 73854 32838 74078 33122
rect 73854 32786 73940 32838
rect 73992 32786 74078 32838
rect 73854 32502 74078 32786
rect 73854 32450 73940 32502
rect 73992 32450 74078 32502
rect 73854 32168 74078 32450
rect 73854 32112 73938 32168
rect 73994 32112 74078 32168
rect 73854 31830 74078 32112
rect 73854 31778 73940 31830
rect 73992 31778 74078 31830
rect 73854 31494 74078 31778
rect 73854 31442 73940 31494
rect 73992 31442 74078 31494
rect 73854 31158 74078 31442
rect 73854 31106 73940 31158
rect 73992 31106 74078 31158
rect 73854 30822 74078 31106
rect 73854 30770 73940 30822
rect 73992 30770 74078 30822
rect 73854 30488 74078 30770
rect 73854 30432 73938 30488
rect 73994 30432 74078 30488
rect 73854 30150 74078 30432
rect 73854 30098 73940 30150
rect 73992 30098 74078 30150
rect 73854 29814 74078 30098
rect 73854 29762 73940 29814
rect 73992 29762 74078 29814
rect 73854 29478 74078 29762
rect 73854 29426 73940 29478
rect 73992 29426 74078 29478
rect 73854 29142 74078 29426
rect 73854 29090 73940 29142
rect 73992 29090 74078 29142
rect 73854 28808 74078 29090
rect 73854 28752 73938 28808
rect 73994 28752 74078 28808
rect 73854 28470 74078 28752
rect 73854 28418 73940 28470
rect 73992 28418 74078 28470
rect 73854 28134 74078 28418
rect 73854 28082 73940 28134
rect 73992 28082 74078 28134
rect 73854 27798 74078 28082
rect 73854 27746 73940 27798
rect 73992 27746 74078 27798
rect 73854 27462 74078 27746
rect 73854 27410 73940 27462
rect 73992 27410 74078 27462
rect 73854 27128 74078 27410
rect 73854 27072 73938 27128
rect 73994 27072 74078 27128
rect 73854 26790 74078 27072
rect 73854 26738 73940 26790
rect 73992 26738 74078 26790
rect 73854 26454 74078 26738
rect 73854 26402 73940 26454
rect 73992 26402 74078 26454
rect 73854 26118 74078 26402
rect 73854 26066 73940 26118
rect 73992 26066 74078 26118
rect 73854 25782 74078 26066
rect 73854 25730 73940 25782
rect 73992 25730 74078 25782
rect 73854 25448 74078 25730
rect 73854 25392 73938 25448
rect 73994 25392 74078 25448
rect 73854 25110 74078 25392
rect 73854 25058 73940 25110
rect 73992 25058 74078 25110
rect 73854 24774 74078 25058
rect 73854 24722 73940 24774
rect 73992 24722 74078 24774
rect 73854 24438 74078 24722
rect 73854 24386 73940 24438
rect 73992 24386 74078 24438
rect 73854 24102 74078 24386
rect 73854 24050 73940 24102
rect 73992 24050 74078 24102
rect 73854 23768 74078 24050
rect 73854 23712 73938 23768
rect 73994 23712 74078 23768
rect 73854 23430 74078 23712
rect 73854 23378 73940 23430
rect 73992 23378 74078 23430
rect 73854 23094 74078 23378
rect 73854 23042 73940 23094
rect 73992 23042 74078 23094
rect 73854 22758 74078 23042
rect 73854 22706 73940 22758
rect 73992 22706 74078 22758
rect 73854 22422 74078 22706
rect 73854 22370 73940 22422
rect 73992 22370 74078 22422
rect 73854 22088 74078 22370
rect 73854 22032 73938 22088
rect 73994 22032 74078 22088
rect 73854 21750 74078 22032
rect 73854 21698 73940 21750
rect 73992 21698 74078 21750
rect 73854 21414 74078 21698
rect 73854 21362 73940 21414
rect 73992 21362 74078 21414
rect 73854 21078 74078 21362
rect 73854 21026 73940 21078
rect 73992 21026 74078 21078
rect 73854 20742 74078 21026
rect 73854 20690 73940 20742
rect 73992 20690 74078 20742
rect 73854 20408 74078 20690
rect 73854 20352 73938 20408
rect 73994 20352 74078 20408
rect 73854 20070 74078 20352
rect 73854 20018 73940 20070
rect 73992 20018 74078 20070
rect 73854 19734 74078 20018
rect 73854 19682 73940 19734
rect 73992 19682 74078 19734
rect 73854 19398 74078 19682
rect 73854 19346 73940 19398
rect 73992 19346 74078 19398
rect 73854 19062 74078 19346
rect 73854 19010 73940 19062
rect 73992 19010 74078 19062
rect 73854 18728 74078 19010
rect 73854 18672 73938 18728
rect 73994 18672 74078 18728
rect 73854 18390 74078 18672
rect 73854 18338 73940 18390
rect 73992 18338 74078 18390
rect 73854 18054 74078 18338
rect 73854 18002 73940 18054
rect 73992 18002 74078 18054
rect 73854 17718 74078 18002
rect 73854 17666 73940 17718
rect 73992 17666 74078 17718
rect 73854 17382 74078 17666
rect 73854 17330 73940 17382
rect 73992 17330 74078 17382
rect 73854 17048 74078 17330
rect 73854 16992 73938 17048
rect 73994 16992 74078 17048
rect 73854 16710 74078 16992
rect 73854 16658 73940 16710
rect 73992 16658 74078 16710
rect 73854 16374 74078 16658
rect 73854 16322 73940 16374
rect 73992 16322 74078 16374
rect 73854 16038 74078 16322
rect 73854 15986 73940 16038
rect 73992 15986 74078 16038
rect 73854 15702 74078 15986
rect 73854 15650 73940 15702
rect 73992 15650 74078 15702
rect 73854 15368 74078 15650
rect 73854 15312 73938 15368
rect 73994 15312 74078 15368
rect 73854 15030 74078 15312
rect 73854 14978 73940 15030
rect 73992 14978 74078 15030
rect 73854 14694 74078 14978
rect 73854 14642 73940 14694
rect 73992 14642 74078 14694
rect 73854 14358 74078 14642
rect 73854 14306 73940 14358
rect 73992 14306 74078 14358
rect 73854 14022 74078 14306
rect 73854 13970 73940 14022
rect 73992 13970 74078 14022
rect 73854 13688 74078 13970
rect 73854 13632 73938 13688
rect 73994 13632 74078 13688
rect 73854 13350 74078 13632
rect 73854 13298 73940 13350
rect 73992 13298 74078 13350
rect 73854 13014 74078 13298
rect 73854 12962 73940 13014
rect 73992 12962 74078 13014
rect 73854 12678 74078 12962
rect 73854 12626 73940 12678
rect 73992 12626 74078 12678
rect 73854 12342 74078 12626
rect 73854 12290 73940 12342
rect 73992 12290 74078 12342
rect 73854 12008 74078 12290
rect 73854 11952 73938 12008
rect 73994 11952 74078 12008
rect 73854 11670 74078 11952
rect 73854 11618 73940 11670
rect 73992 11618 74078 11670
rect 73854 11334 74078 11618
rect 73854 11282 73940 11334
rect 73992 11282 74078 11334
rect 73854 10998 74078 11282
rect 73854 10946 73940 10998
rect 73992 10946 74078 10998
rect 73854 10662 74078 10946
rect 73854 10610 73940 10662
rect 73992 10610 74078 10662
rect 19626 8485 19654 10570
rect 73854 10328 74078 10610
rect 73854 10272 73938 10328
rect 73994 10272 74078 10328
rect 73854 9990 74078 10272
rect 73854 9938 73940 9990
rect 73992 9938 74078 9990
rect 73854 9654 74078 9938
rect 73854 9602 73940 9654
rect 73992 9602 74078 9654
rect 73854 9318 74078 9602
rect 73854 9266 73940 9318
rect 73992 9266 74078 9318
rect 11463 5846 12158 5860
rect 11463 5832 12174 5846
rect 1506 5570 1592 5622
rect 1644 5570 1730 5622
rect 1506 5288 1730 5570
rect 1506 5232 1590 5288
rect 1646 5232 1730 5288
rect 1506 4950 1730 5232
rect 1506 4898 1592 4950
rect 1644 4898 1730 4950
rect 1506 4614 1730 4898
rect 1506 4562 1592 4614
rect 1644 4562 1730 4614
rect 1506 4278 1730 4562
rect 1506 4226 1592 4278
rect 1644 4226 1730 4278
rect 1506 3942 1730 4226
rect 1506 3890 1592 3942
rect 1644 3890 1730 3942
rect 1506 3608 1730 3890
rect 1506 3552 1590 3608
rect 1646 3552 1730 3608
rect 1506 3270 1730 3552
rect 1506 3218 1592 3270
rect 1644 3218 1730 3270
rect 1506 2934 1730 3218
rect 1506 2882 1592 2934
rect 1644 2882 1730 2934
rect 1506 2598 1730 2882
rect 12114 2732 12174 5832
rect 45182 4936 45210 9173
rect 73854 8982 74078 9266
rect 73854 8930 73940 8982
rect 73992 8930 74078 8982
rect 73854 8648 74078 8930
rect 73854 8592 73938 8648
rect 73994 8592 74078 8648
rect 73854 8310 74078 8592
rect 73854 8258 73940 8310
rect 73992 8258 74078 8310
rect 73854 7974 74078 8258
rect 73854 7922 73940 7974
rect 73992 7922 74078 7974
rect 73854 7638 74078 7922
rect 73854 7586 73940 7638
rect 73992 7586 74078 7638
rect 73854 7302 74078 7586
rect 73854 7250 73940 7302
rect 73992 7250 74078 7302
rect 73854 6968 74078 7250
rect 73854 6912 73938 6968
rect 73994 6912 74078 6968
rect 73854 6630 74078 6912
rect 73854 6578 73940 6630
rect 73992 6578 74078 6630
rect 73854 6294 74078 6578
rect 73854 6242 73940 6294
rect 73992 6242 74078 6294
rect 73854 5958 74078 6242
rect 73854 5906 73940 5958
rect 73992 5906 74078 5958
rect 73854 5622 74078 5906
rect 73854 5570 73940 5622
rect 73992 5570 74078 5622
rect 73854 5288 74078 5570
rect 73854 5232 73938 5288
rect 73994 5232 74078 5288
rect 73854 4950 74078 5232
rect 12114 2704 12116 2732
rect 12172 2704 12174 2732
rect 73854 4898 73940 4950
rect 73992 4898 74078 4950
rect 73854 4614 74078 4898
rect 73854 4562 73940 4614
rect 73992 4562 74078 4614
rect 73854 4278 74078 4562
rect 73854 4226 73940 4278
rect 73992 4226 74078 4278
rect 73854 3942 74078 4226
rect 73854 3890 73940 3942
rect 73992 3890 74078 3942
rect 73854 3608 74078 3890
rect 73854 3552 73938 3608
rect 73994 3552 74078 3608
rect 73854 3270 74078 3552
rect 73854 3218 73940 3270
rect 73992 3218 74078 3270
rect 73854 2934 74078 3218
rect 73854 2882 73940 2934
rect 73992 2882 74078 2934
rect 1506 2546 1592 2598
rect 1644 2546 1730 2598
rect 1506 2262 1730 2546
rect 1506 2210 1592 2262
rect 1644 2210 1730 2262
rect 1506 1928 1730 2210
rect 1506 1872 1590 1928
rect 1646 1872 1730 1928
rect 1506 1452 1730 1872
rect 73854 2598 74078 2882
rect 73854 2546 73940 2598
rect 73992 2546 74078 2598
rect 73854 2262 74078 2546
rect 73854 2210 73940 2262
rect 73992 2210 74078 2262
rect 73854 1928 74078 2210
rect 73854 1872 73938 1928
rect 73994 1872 74078 1928
rect 1934 1592 1974 1598
rect 3614 1592 3654 1598
rect 5294 1592 5334 1598
rect 6974 1592 7014 1598
rect 8654 1592 8694 1598
rect 10334 1592 10374 1598
rect 12014 1592 12054 1598
rect 13694 1592 13734 1598
rect 15374 1592 15414 1598
rect 17054 1592 17094 1598
rect 18734 1592 18774 1598
rect 20414 1592 20454 1598
rect 22094 1592 22134 1598
rect 23774 1592 23814 1598
rect 25454 1592 25494 1598
rect 27134 1592 27174 1598
rect 28814 1592 28854 1598
rect 30494 1592 30534 1598
rect 32174 1592 32214 1598
rect 33854 1592 33894 1598
rect 35534 1592 35574 1598
rect 37214 1592 37254 1598
rect 38894 1592 38934 1598
rect 40574 1592 40614 1598
rect 42254 1592 42294 1598
rect 43934 1592 43974 1598
rect 45614 1592 45654 1598
rect 47294 1592 47334 1598
rect 48974 1592 49014 1598
rect 50654 1592 50694 1598
rect 52334 1592 52374 1598
rect 54014 1592 54054 1598
rect 55694 1592 55734 1598
rect 57374 1592 57414 1598
rect 59054 1592 59094 1598
rect 60734 1592 60774 1598
rect 62414 1592 62454 1598
rect 64094 1592 64134 1598
rect 65774 1592 65814 1598
rect 67454 1592 67494 1598
rect 69134 1592 69174 1598
rect 70814 1592 70854 1598
rect 72494 1592 72534 1598
rect 1934 1530 1974 1536
rect 3614 1530 3654 1536
rect 5294 1530 5334 1536
rect 6974 1530 7014 1536
rect 8654 1530 8694 1536
rect 10334 1530 10374 1536
rect 12014 1530 12054 1536
rect 13694 1530 13734 1536
rect 15374 1530 15414 1536
rect 17054 1530 17094 1536
rect 18734 1530 18774 1536
rect 20414 1530 20454 1536
rect 22094 1530 22134 1536
rect 23774 1530 23814 1536
rect 25454 1530 25494 1536
rect 27134 1530 27174 1536
rect 28814 1530 28854 1536
rect 30494 1530 30534 1536
rect 32174 1530 32214 1536
rect 33854 1530 33894 1536
rect 35534 1530 35574 1536
rect 37214 1530 37254 1536
rect 38894 1530 38934 1536
rect 40574 1530 40614 1536
rect 42254 1530 42294 1536
rect 43934 1530 43974 1536
rect 45614 1530 45654 1536
rect 47294 1530 47334 1536
rect 48974 1530 49014 1536
rect 50654 1530 50694 1536
rect 52334 1530 52374 1536
rect 54014 1530 54054 1536
rect 55694 1530 55734 1536
rect 57374 1530 57414 1536
rect 59054 1530 59094 1536
rect 60734 1530 60774 1536
rect 62414 1530 62454 1536
rect 64094 1530 64134 1536
rect 65774 1530 65814 1536
rect 67454 1530 67494 1536
rect 69134 1530 69174 1536
rect 70814 1530 70854 1536
rect 72494 1530 72534 1536
rect 73854 1452 74078 1872
<< via2 >>
rect 1926 36234 1982 36236
rect 1926 36182 1928 36234
rect 1928 36182 1980 36234
rect 1980 36182 1982 36234
rect 1926 36180 1982 36182
rect 3606 36234 3662 36236
rect 3606 36182 3608 36234
rect 3608 36182 3660 36234
rect 3660 36182 3662 36234
rect 3606 36180 3662 36182
rect 5286 36234 5342 36236
rect 5286 36182 5288 36234
rect 5288 36182 5340 36234
rect 5340 36182 5342 36234
rect 5286 36180 5342 36182
rect 6966 36234 7022 36236
rect 6966 36182 6968 36234
rect 6968 36182 7020 36234
rect 7020 36182 7022 36234
rect 6966 36180 7022 36182
rect 8646 36234 8702 36236
rect 8646 36182 8648 36234
rect 8648 36182 8700 36234
rect 8700 36182 8702 36234
rect 8646 36180 8702 36182
rect 10326 36234 10382 36236
rect 10326 36182 10328 36234
rect 10328 36182 10380 36234
rect 10380 36182 10382 36234
rect 10326 36180 10382 36182
rect 12006 36234 12062 36236
rect 12006 36182 12008 36234
rect 12008 36182 12060 36234
rect 12060 36182 12062 36234
rect 12006 36180 12062 36182
rect 13686 36234 13742 36236
rect 13686 36182 13688 36234
rect 13688 36182 13740 36234
rect 13740 36182 13742 36234
rect 13686 36180 13742 36182
rect 15366 36234 15422 36236
rect 15366 36182 15368 36234
rect 15368 36182 15420 36234
rect 15420 36182 15422 36234
rect 15366 36180 15422 36182
rect 17046 36234 17102 36236
rect 17046 36182 17048 36234
rect 17048 36182 17100 36234
rect 17100 36182 17102 36234
rect 17046 36180 17102 36182
rect 18726 36234 18782 36236
rect 18726 36182 18728 36234
rect 18728 36182 18780 36234
rect 18780 36182 18782 36234
rect 18726 36180 18782 36182
rect 20406 36234 20462 36236
rect 20406 36182 20408 36234
rect 20408 36182 20460 36234
rect 20460 36182 20462 36234
rect 20406 36180 20462 36182
rect 22086 36234 22142 36236
rect 22086 36182 22088 36234
rect 22088 36182 22140 36234
rect 22140 36182 22142 36234
rect 22086 36180 22142 36182
rect 23766 36234 23822 36236
rect 23766 36182 23768 36234
rect 23768 36182 23820 36234
rect 23820 36182 23822 36234
rect 23766 36180 23822 36182
rect 25446 36234 25502 36236
rect 25446 36182 25448 36234
rect 25448 36182 25500 36234
rect 25500 36182 25502 36234
rect 25446 36180 25502 36182
rect 27126 36234 27182 36236
rect 27126 36182 27128 36234
rect 27128 36182 27180 36234
rect 27180 36182 27182 36234
rect 27126 36180 27182 36182
rect 28806 36234 28862 36236
rect 28806 36182 28808 36234
rect 28808 36182 28860 36234
rect 28860 36182 28862 36234
rect 28806 36180 28862 36182
rect 30486 36234 30542 36236
rect 30486 36182 30488 36234
rect 30488 36182 30540 36234
rect 30540 36182 30542 36234
rect 30486 36180 30542 36182
rect 32166 36234 32222 36236
rect 32166 36182 32168 36234
rect 32168 36182 32220 36234
rect 32220 36182 32222 36234
rect 32166 36180 32222 36182
rect 33846 36234 33902 36236
rect 33846 36182 33848 36234
rect 33848 36182 33900 36234
rect 33900 36182 33902 36234
rect 33846 36180 33902 36182
rect 35526 36234 35582 36236
rect 35526 36182 35528 36234
rect 35528 36182 35580 36234
rect 35580 36182 35582 36234
rect 35526 36180 35582 36182
rect 37206 36234 37262 36236
rect 37206 36182 37208 36234
rect 37208 36182 37260 36234
rect 37260 36182 37262 36234
rect 37206 36180 37262 36182
rect 38886 36234 38942 36236
rect 38886 36182 38888 36234
rect 38888 36182 38940 36234
rect 38940 36182 38942 36234
rect 38886 36180 38942 36182
rect 40566 36234 40622 36236
rect 40566 36182 40568 36234
rect 40568 36182 40620 36234
rect 40620 36182 40622 36234
rect 40566 36180 40622 36182
rect 42246 36234 42302 36236
rect 42246 36182 42248 36234
rect 42248 36182 42300 36234
rect 42300 36182 42302 36234
rect 42246 36180 42302 36182
rect 43926 36234 43982 36236
rect 43926 36182 43928 36234
rect 43928 36182 43980 36234
rect 43980 36182 43982 36234
rect 43926 36180 43982 36182
rect 45606 36234 45662 36236
rect 45606 36182 45608 36234
rect 45608 36182 45660 36234
rect 45660 36182 45662 36234
rect 45606 36180 45662 36182
rect 47286 36234 47342 36236
rect 47286 36182 47288 36234
rect 47288 36182 47340 36234
rect 47340 36182 47342 36234
rect 47286 36180 47342 36182
rect 48966 36234 49022 36236
rect 48966 36182 48968 36234
rect 48968 36182 49020 36234
rect 49020 36182 49022 36234
rect 48966 36180 49022 36182
rect 50646 36234 50702 36236
rect 50646 36182 50648 36234
rect 50648 36182 50700 36234
rect 50700 36182 50702 36234
rect 50646 36180 50702 36182
rect 52326 36234 52382 36236
rect 52326 36182 52328 36234
rect 52328 36182 52380 36234
rect 52380 36182 52382 36234
rect 52326 36180 52382 36182
rect 54006 36234 54062 36236
rect 54006 36182 54008 36234
rect 54008 36182 54060 36234
rect 54060 36182 54062 36234
rect 54006 36180 54062 36182
rect 55686 36234 55742 36236
rect 55686 36182 55688 36234
rect 55688 36182 55740 36234
rect 55740 36182 55742 36234
rect 55686 36180 55742 36182
rect 57366 36234 57422 36236
rect 57366 36182 57368 36234
rect 57368 36182 57420 36234
rect 57420 36182 57422 36234
rect 57366 36180 57422 36182
rect 59046 36234 59102 36236
rect 59046 36182 59048 36234
rect 59048 36182 59100 36234
rect 59100 36182 59102 36234
rect 59046 36180 59102 36182
rect 60726 36234 60782 36236
rect 60726 36182 60728 36234
rect 60728 36182 60780 36234
rect 60780 36182 60782 36234
rect 60726 36180 60782 36182
rect 62406 36234 62462 36236
rect 62406 36182 62408 36234
rect 62408 36182 62460 36234
rect 62460 36182 62462 36234
rect 62406 36180 62462 36182
rect 64086 36234 64142 36236
rect 64086 36182 64088 36234
rect 64088 36182 64140 36234
rect 64140 36182 64142 36234
rect 64086 36180 64142 36182
rect 65766 36234 65822 36236
rect 65766 36182 65768 36234
rect 65768 36182 65820 36234
rect 65820 36182 65822 36234
rect 65766 36180 65822 36182
rect 67446 36234 67502 36236
rect 67446 36182 67448 36234
rect 67448 36182 67500 36234
rect 67500 36182 67502 36234
rect 67446 36180 67502 36182
rect 69126 36234 69182 36236
rect 69126 36182 69128 36234
rect 69128 36182 69180 36234
rect 69180 36182 69182 36234
rect 69126 36180 69182 36182
rect 70806 36234 70862 36236
rect 70806 36182 70808 36234
rect 70808 36182 70860 36234
rect 70860 36182 70862 36234
rect 70806 36180 70862 36182
rect 72486 36234 72542 36236
rect 72486 36182 72488 36234
rect 72488 36182 72540 36234
rect 72540 36182 72542 36234
rect 72486 36180 72542 36182
rect 1590 35526 1646 35528
rect 1590 35474 1592 35526
rect 1592 35474 1644 35526
rect 1644 35474 1646 35526
rect 1590 35472 1646 35474
rect 73938 35526 73994 35528
rect 73938 35474 73940 35526
rect 73940 35474 73992 35526
rect 73992 35474 73994 35526
rect 73938 35472 73994 35474
rect 1590 33846 1646 33848
rect 1590 33794 1592 33846
rect 1592 33794 1644 33846
rect 1644 33794 1646 33846
rect 1590 33792 1646 33794
rect 1590 32166 1646 32168
rect 1590 32114 1592 32166
rect 1592 32114 1644 32166
rect 1644 32114 1646 32166
rect 1590 32112 1646 32114
rect 1590 30486 1646 30488
rect 1590 30434 1592 30486
rect 1592 30434 1644 30486
rect 1644 30434 1646 30486
rect 1590 30432 1646 30434
rect 1590 28806 1646 28808
rect 1590 28754 1592 28806
rect 1592 28754 1644 28806
rect 1644 28754 1646 28806
rect 1590 28752 1646 28754
rect 1590 27126 1646 27128
rect 1590 27074 1592 27126
rect 1592 27074 1644 27126
rect 1644 27074 1646 27126
rect 1590 27072 1646 27074
rect 1590 25446 1646 25448
rect 1590 25394 1592 25446
rect 1592 25394 1644 25446
rect 1644 25394 1646 25446
rect 1590 25392 1646 25394
rect 1590 23766 1646 23768
rect 1590 23714 1592 23766
rect 1592 23714 1644 23766
rect 1644 23714 1646 23766
rect 1590 23712 1646 23714
rect 1590 22086 1646 22088
rect 1590 22034 1592 22086
rect 1592 22034 1644 22086
rect 1644 22034 1646 22086
rect 1590 22032 1646 22034
rect 1590 20406 1646 20408
rect 1590 20354 1592 20406
rect 1592 20354 1644 20406
rect 1644 20354 1646 20406
rect 1590 20352 1646 20354
rect 1590 18726 1646 18728
rect 1590 18674 1592 18726
rect 1592 18674 1644 18726
rect 1644 18674 1646 18726
rect 1590 18672 1646 18674
rect 1590 17046 1646 17048
rect 1590 16994 1592 17046
rect 1592 16994 1644 17046
rect 1644 16994 1646 17046
rect 1590 16992 1646 16994
rect 12391 15514 12447 15570
rect 13471 15518 13527 15574
rect 1590 15366 1646 15368
rect 1590 15314 1592 15366
rect 1592 15314 1644 15366
rect 1644 15314 1646 15366
rect 1590 15312 1646 15314
rect 12391 14330 12447 14386
rect 13471 14326 13527 14382
rect 12391 13838 12447 13894
rect 13471 13842 13527 13898
rect 1590 13686 1646 13688
rect 1590 13634 1592 13686
rect 1592 13634 1644 13686
rect 1644 13634 1646 13686
rect 1590 13632 1646 13634
rect 12391 12654 12447 12710
rect 13471 12650 13527 12706
rect 12391 12162 12447 12218
rect 13471 12166 13527 12222
rect 1590 12006 1646 12008
rect 1590 11954 1592 12006
rect 1592 11954 1644 12006
rect 1644 11954 1646 12006
rect 1590 11952 1646 11954
rect 12116 11032 12172 11088
rect 1590 10326 1646 10328
rect 1590 10274 1592 10326
rect 1592 10274 1644 10326
rect 1644 10274 1646 10326
rect 1590 10272 1646 10274
rect 1590 8646 1646 8648
rect 1590 8594 1592 8646
rect 1592 8594 1644 8646
rect 1644 8594 1646 8646
rect 1590 8592 1646 8594
rect 1590 6966 1646 6968
rect 1590 6914 1592 6966
rect 1592 6914 1644 6966
rect 1644 6914 1646 6966
rect 1590 6912 1646 6914
rect 2637 6040 2693 6096
rect 5997 5825 6053 5881
rect 12391 10978 12447 11034
rect 14157 15518 14213 15574
rect 14089 14326 14145 14382
rect 14021 13842 14077 13898
rect 13953 12650 14009 12706
rect 13885 12166 13941 12222
rect 13471 10974 13527 11030
rect 13817 10974 13873 11030
rect 73938 33846 73994 33848
rect 73938 33794 73940 33846
rect 73940 33794 73992 33846
rect 73992 33794 73994 33846
rect 73938 33792 73994 33794
rect 73938 32166 73994 32168
rect 73938 32114 73940 32166
rect 73940 32114 73992 32166
rect 73992 32114 73994 32166
rect 73938 32112 73994 32114
rect 73938 30486 73994 30488
rect 73938 30434 73940 30486
rect 73940 30434 73992 30486
rect 73992 30434 73994 30486
rect 73938 30432 73994 30434
rect 73938 28806 73994 28808
rect 73938 28754 73940 28806
rect 73940 28754 73992 28806
rect 73992 28754 73994 28806
rect 73938 28752 73994 28754
rect 73938 27126 73994 27128
rect 73938 27074 73940 27126
rect 73940 27074 73992 27126
rect 73992 27074 73994 27126
rect 73938 27072 73994 27074
rect 73938 25446 73994 25448
rect 73938 25394 73940 25446
rect 73940 25394 73992 25446
rect 73992 25394 73994 25446
rect 73938 25392 73994 25394
rect 73938 23766 73994 23768
rect 73938 23714 73940 23766
rect 73940 23714 73992 23766
rect 73992 23714 73994 23766
rect 73938 23712 73994 23714
rect 73938 22086 73994 22088
rect 73938 22034 73940 22086
rect 73940 22034 73992 22086
rect 73992 22034 73994 22086
rect 73938 22032 73994 22034
rect 73938 20406 73994 20408
rect 73938 20354 73940 20406
rect 73940 20354 73992 20406
rect 73992 20354 73994 20406
rect 73938 20352 73994 20354
rect 73938 18726 73994 18728
rect 73938 18674 73940 18726
rect 73940 18674 73992 18726
rect 73992 18674 73994 18726
rect 73938 18672 73994 18674
rect 73938 17046 73994 17048
rect 73938 16994 73940 17046
rect 73940 16994 73992 17046
rect 73992 16994 73994 17046
rect 73938 16992 73994 16994
rect 73938 15366 73994 15368
rect 73938 15314 73940 15366
rect 73940 15314 73992 15366
rect 73992 15314 73994 15366
rect 73938 15312 73994 15314
rect 73938 13686 73994 13688
rect 73938 13634 73940 13686
rect 73940 13634 73992 13686
rect 73992 13634 73994 13686
rect 73938 13632 73994 13634
rect 73938 12006 73994 12008
rect 73938 11954 73940 12006
rect 73940 11954 73992 12006
rect 73992 11954 73994 12006
rect 73938 11952 73994 11954
rect 13666 10099 13722 10155
rect 18478 10099 18534 10155
rect 13666 9173 13722 9229
rect 73938 10326 73994 10328
rect 73938 10274 73940 10326
rect 73940 10274 73992 10326
rect 73992 10274 73994 10326
rect 73938 10272 73994 10274
rect 24722 9252 24778 9308
rect 26278 9252 26334 9308
rect 27834 9252 27890 9308
rect 29390 9252 29446 9308
rect 30946 9252 31002 9308
rect 32502 9252 32558 9308
rect 34058 9252 34114 9308
rect 35614 9252 35670 9308
rect 37170 9252 37226 9308
rect 38726 9252 38782 9308
rect 40282 9252 40338 9308
rect 41838 9252 41894 9308
rect 43394 9252 43450 9308
rect 44950 9252 45006 9308
rect 46506 9252 46562 9308
rect 48062 9252 48118 9308
rect 45168 9173 45224 9229
rect 13666 8429 13722 8485
rect 19612 8429 19668 8485
rect 1590 5286 1646 5288
rect 1590 5234 1592 5286
rect 1592 5234 1644 5286
rect 1644 5234 1646 5286
rect 1590 5232 1646 5234
rect 2637 4856 2693 4912
rect 1590 3606 1646 3608
rect 1590 3554 1592 3606
rect 1592 3554 1644 3606
rect 1644 3554 1646 3606
rect 1590 3552 1646 3554
rect 73938 8646 73994 8648
rect 73938 8594 73940 8646
rect 73940 8594 73992 8646
rect 73992 8594 73994 8646
rect 73938 8592 73994 8594
rect 73938 6966 73994 6968
rect 73938 6914 73940 6966
rect 73940 6914 73992 6966
rect 73992 6914 73994 6966
rect 73938 6912 73994 6914
rect 73938 5286 73994 5288
rect 73938 5234 73940 5286
rect 73940 5234 73992 5286
rect 73992 5234 73994 5286
rect 73938 5232 73994 5234
rect 12116 2676 12172 2732
rect 73938 3606 73994 3608
rect 73938 3554 73940 3606
rect 73940 3554 73992 3606
rect 73992 3554 73994 3606
rect 73938 3552 73994 3554
rect 15355 2622 15411 2678
rect 16837 2622 16893 2678
rect 18319 2622 18375 2678
rect 19801 2622 19857 2678
rect 21283 2622 21339 2678
rect 22765 2622 22821 2678
rect 24247 2622 24303 2678
rect 25729 2622 25785 2678
rect 27211 2622 27267 2678
rect 28693 2622 28749 2678
rect 30175 2622 30231 2678
rect 31657 2622 31713 2678
rect 33139 2622 33195 2678
rect 34621 2622 34677 2678
rect 36103 2622 36159 2678
rect 37585 2622 37641 2678
rect 39067 2622 39123 2678
rect 1590 1926 1646 1928
rect 1590 1874 1592 1926
rect 1592 1874 1644 1926
rect 1644 1874 1646 1926
rect 1590 1872 1646 1874
rect 73938 1926 73994 1928
rect 73938 1874 73940 1926
rect 73940 1874 73992 1926
rect 73992 1874 73994 1926
rect 73938 1872 73994 1874
rect 1926 1590 1982 1592
rect 1926 1538 1928 1590
rect 1928 1538 1980 1590
rect 1980 1538 1982 1590
rect 1926 1536 1982 1538
rect 3606 1590 3662 1592
rect 3606 1538 3608 1590
rect 3608 1538 3660 1590
rect 3660 1538 3662 1590
rect 3606 1536 3662 1538
rect 5286 1590 5342 1592
rect 5286 1538 5288 1590
rect 5288 1538 5340 1590
rect 5340 1538 5342 1590
rect 5286 1536 5342 1538
rect 6966 1590 7022 1592
rect 6966 1538 6968 1590
rect 6968 1538 7020 1590
rect 7020 1538 7022 1590
rect 6966 1536 7022 1538
rect 8646 1590 8702 1592
rect 8646 1538 8648 1590
rect 8648 1538 8700 1590
rect 8700 1538 8702 1590
rect 8646 1536 8702 1538
rect 10326 1590 10382 1592
rect 10326 1538 10328 1590
rect 10328 1538 10380 1590
rect 10380 1538 10382 1590
rect 10326 1536 10382 1538
rect 12006 1590 12062 1592
rect 12006 1538 12008 1590
rect 12008 1538 12060 1590
rect 12060 1538 12062 1590
rect 12006 1536 12062 1538
rect 13686 1590 13742 1592
rect 13686 1538 13688 1590
rect 13688 1538 13740 1590
rect 13740 1538 13742 1590
rect 13686 1536 13742 1538
rect 15366 1590 15422 1592
rect 15366 1538 15368 1590
rect 15368 1538 15420 1590
rect 15420 1538 15422 1590
rect 15366 1536 15422 1538
rect 17046 1590 17102 1592
rect 17046 1538 17048 1590
rect 17048 1538 17100 1590
rect 17100 1538 17102 1590
rect 17046 1536 17102 1538
rect 18726 1590 18782 1592
rect 18726 1538 18728 1590
rect 18728 1538 18780 1590
rect 18780 1538 18782 1590
rect 18726 1536 18782 1538
rect 20406 1590 20462 1592
rect 20406 1538 20408 1590
rect 20408 1538 20460 1590
rect 20460 1538 20462 1590
rect 20406 1536 20462 1538
rect 22086 1590 22142 1592
rect 22086 1538 22088 1590
rect 22088 1538 22140 1590
rect 22140 1538 22142 1590
rect 22086 1536 22142 1538
rect 23766 1590 23822 1592
rect 23766 1538 23768 1590
rect 23768 1538 23820 1590
rect 23820 1538 23822 1590
rect 23766 1536 23822 1538
rect 25446 1590 25502 1592
rect 25446 1538 25448 1590
rect 25448 1538 25500 1590
rect 25500 1538 25502 1590
rect 25446 1536 25502 1538
rect 27126 1590 27182 1592
rect 27126 1538 27128 1590
rect 27128 1538 27180 1590
rect 27180 1538 27182 1590
rect 27126 1536 27182 1538
rect 28806 1590 28862 1592
rect 28806 1538 28808 1590
rect 28808 1538 28860 1590
rect 28860 1538 28862 1590
rect 28806 1536 28862 1538
rect 30486 1590 30542 1592
rect 30486 1538 30488 1590
rect 30488 1538 30540 1590
rect 30540 1538 30542 1590
rect 30486 1536 30542 1538
rect 32166 1590 32222 1592
rect 32166 1538 32168 1590
rect 32168 1538 32220 1590
rect 32220 1538 32222 1590
rect 32166 1536 32222 1538
rect 33846 1590 33902 1592
rect 33846 1538 33848 1590
rect 33848 1538 33900 1590
rect 33900 1538 33902 1590
rect 33846 1536 33902 1538
rect 35526 1590 35582 1592
rect 35526 1538 35528 1590
rect 35528 1538 35580 1590
rect 35580 1538 35582 1590
rect 35526 1536 35582 1538
rect 37206 1590 37262 1592
rect 37206 1538 37208 1590
rect 37208 1538 37260 1590
rect 37260 1538 37262 1590
rect 37206 1536 37262 1538
rect 38886 1590 38942 1592
rect 38886 1538 38888 1590
rect 38888 1538 38940 1590
rect 38940 1538 38942 1590
rect 38886 1536 38942 1538
rect 40566 1590 40622 1592
rect 40566 1538 40568 1590
rect 40568 1538 40620 1590
rect 40620 1538 40622 1590
rect 40566 1536 40622 1538
rect 42246 1590 42302 1592
rect 42246 1538 42248 1590
rect 42248 1538 42300 1590
rect 42300 1538 42302 1590
rect 42246 1536 42302 1538
rect 43926 1590 43982 1592
rect 43926 1538 43928 1590
rect 43928 1538 43980 1590
rect 43980 1538 43982 1590
rect 43926 1536 43982 1538
rect 45606 1590 45662 1592
rect 45606 1538 45608 1590
rect 45608 1538 45660 1590
rect 45660 1538 45662 1590
rect 45606 1536 45662 1538
rect 47286 1590 47342 1592
rect 47286 1538 47288 1590
rect 47288 1538 47340 1590
rect 47340 1538 47342 1590
rect 47286 1536 47342 1538
rect 48966 1590 49022 1592
rect 48966 1538 48968 1590
rect 48968 1538 49020 1590
rect 49020 1538 49022 1590
rect 48966 1536 49022 1538
rect 50646 1590 50702 1592
rect 50646 1538 50648 1590
rect 50648 1538 50700 1590
rect 50700 1538 50702 1590
rect 50646 1536 50702 1538
rect 52326 1590 52382 1592
rect 52326 1538 52328 1590
rect 52328 1538 52380 1590
rect 52380 1538 52382 1590
rect 52326 1536 52382 1538
rect 54006 1590 54062 1592
rect 54006 1538 54008 1590
rect 54008 1538 54060 1590
rect 54060 1538 54062 1590
rect 54006 1536 54062 1538
rect 55686 1590 55742 1592
rect 55686 1538 55688 1590
rect 55688 1538 55740 1590
rect 55740 1538 55742 1590
rect 55686 1536 55742 1538
rect 57366 1590 57422 1592
rect 57366 1538 57368 1590
rect 57368 1538 57420 1590
rect 57420 1538 57422 1590
rect 57366 1536 57422 1538
rect 59046 1590 59102 1592
rect 59046 1538 59048 1590
rect 59048 1538 59100 1590
rect 59100 1538 59102 1590
rect 59046 1536 59102 1538
rect 60726 1590 60782 1592
rect 60726 1538 60728 1590
rect 60728 1538 60780 1590
rect 60780 1538 60782 1590
rect 60726 1536 60782 1538
rect 62406 1590 62462 1592
rect 62406 1538 62408 1590
rect 62408 1538 62460 1590
rect 62460 1538 62462 1590
rect 62406 1536 62462 1538
rect 64086 1590 64142 1592
rect 64086 1538 64088 1590
rect 64088 1538 64140 1590
rect 64140 1538 64142 1590
rect 64086 1536 64142 1538
rect 65766 1590 65822 1592
rect 65766 1538 65768 1590
rect 65768 1538 65820 1590
rect 65820 1538 65822 1590
rect 65766 1536 65822 1538
rect 67446 1590 67502 1592
rect 67446 1538 67448 1590
rect 67448 1538 67500 1590
rect 67500 1538 67502 1590
rect 67446 1536 67502 1538
rect 69126 1590 69182 1592
rect 69126 1538 69128 1590
rect 69128 1538 69180 1590
rect 69180 1538 69182 1590
rect 69126 1536 69182 1538
rect 70806 1590 70862 1592
rect 70806 1538 70808 1590
rect 70808 1538 70860 1590
rect 70860 1538 70862 1590
rect 70806 1536 70862 1538
rect 72486 1590 72542 1592
rect 72486 1538 72488 1590
rect 72488 1538 72540 1590
rect 72540 1538 72542 1590
rect 72486 1536 72542 1538
<< metal3 >>
rect 302 37438 358 37500
rect 422 37438 478 37500
rect 542 37438 74998 37500
rect 75062 37438 75118 37500
rect 75182 37438 75238 37500
rect 240 37382 75300 37438
rect 302 37318 358 37382
rect 422 37318 478 37382
rect 542 37318 74998 37382
rect 75062 37318 75118 37382
rect 75182 37318 75238 37382
rect 240 37262 75300 37318
rect 302 37200 358 37262
rect 422 37200 478 37262
rect 542 37200 14518 37262
rect 14582 37200 19558 37262
rect 19622 37200 74998 37262
rect 75062 37200 75118 37262
rect 75182 37200 75238 37262
rect 902 36838 958 36900
rect 1022 36838 1078 36900
rect 1142 36838 74398 36900
rect 74462 36838 74518 36900
rect 74582 36838 74638 36900
rect 840 36782 74700 36838
rect 902 36718 958 36782
rect 1022 36718 1078 36782
rect 1142 36718 74398 36782
rect 74462 36718 74518 36782
rect 74582 36718 74638 36782
rect 840 36662 74700 36718
rect 902 36600 958 36662
rect 1022 36600 1078 36662
rect 1142 36600 1918 36662
rect 1982 36600 3718 36662
rect 3782 36600 5398 36662
rect 5462 36600 6958 36662
rect 7022 36600 8638 36662
rect 8702 36600 10438 36662
rect 10502 36600 11998 36662
rect 12062 36600 13678 36662
rect 13742 36600 15478 36662
rect 15542 36600 17158 36662
rect 17222 36600 18838 36662
rect 18902 36600 20518 36662
rect 20582 36600 22078 36662
rect 22142 36600 23758 36662
rect 23822 36600 25438 36662
rect 25502 36600 27118 36662
rect 27182 36600 28918 36662
rect 28982 36600 30478 36662
rect 30542 36600 32158 36662
rect 32222 36600 33838 36662
rect 33902 36600 35638 36662
rect 35702 36600 37318 36662
rect 37382 36600 38878 36662
rect 38942 36600 40678 36662
rect 40742 36600 42358 36662
rect 42422 36600 43918 36662
rect 43982 36600 45718 36662
rect 45782 36600 47398 36662
rect 47462 36600 48958 36662
rect 49022 36600 50638 36662
rect 50702 36600 52438 36662
rect 52502 36600 54118 36662
rect 54182 36600 55678 36662
rect 55742 36600 57358 36662
rect 57422 36600 59158 36662
rect 59222 36600 60718 36662
rect 60782 36600 62398 36662
rect 62462 36600 64198 36662
rect 64262 36600 65758 36662
rect 65822 36600 67558 36662
rect 67622 36600 69238 36662
rect 69302 36600 70798 36662
rect 70862 36600 72478 36662
rect 72542 36600 74398 36662
rect 74462 36600 74518 36662
rect 74582 36600 74638 36662
rect 1982 36238 2100 36300
rect 1920 36236 2100 36238
rect 1920 36180 1926 36236
rect 1982 36180 2100 36236
rect 1920 36120 2100 36180
rect 3600 36238 3718 36300
rect 5280 36238 5398 36300
rect 7022 36238 7140 36300
rect 8702 36238 8820 36300
rect 3600 36236 3780 36238
rect 3600 36180 3606 36236
rect 3662 36180 3780 36236
rect 3600 36120 3780 36180
rect 5280 36236 5460 36238
rect 5280 36180 5286 36236
rect 5342 36180 5460 36236
rect 5280 36120 5460 36180
rect 6960 36236 7140 36238
rect 6960 36180 6966 36236
rect 7022 36180 7140 36236
rect 6960 36120 7140 36180
rect 8640 36236 8820 36238
rect 8640 36180 8646 36236
rect 8702 36180 8820 36236
rect 8640 36120 8820 36180
rect 10320 36238 10438 36300
rect 12062 36238 12180 36300
rect 13742 36238 13860 36300
rect 10320 36236 10500 36238
rect 10320 36180 10326 36236
rect 10382 36180 10500 36236
rect 10320 36120 10500 36180
rect 12000 36236 12180 36238
rect 12000 36180 12006 36236
rect 12062 36180 12180 36236
rect 12000 36120 12180 36180
rect 13680 36236 13860 36238
rect 13680 36180 13686 36236
rect 13742 36180 13860 36236
rect 15360 36238 15478 36300
rect 17040 36238 17158 36300
rect 18720 36238 18838 36300
rect 20400 36238 20518 36300
rect 22142 36238 22260 36300
rect 23822 36238 23940 36300
rect 25502 36238 25620 36300
rect 27182 36238 27300 36300
rect 15360 36236 15540 36238
rect 13680 36120 14398 36180
rect 15360 36180 15366 36236
rect 15422 36180 15540 36236
rect 15360 36120 15540 36180
rect 17040 36236 17220 36238
rect 17040 36180 17046 36236
rect 17102 36180 17220 36236
rect 17040 36120 17220 36180
rect 18720 36236 18900 36238
rect 18720 36180 18726 36236
rect 18782 36180 18900 36236
rect 20400 36236 20580 36238
rect 20400 36182 20406 36236
rect 18720 36120 18900 36180
rect 20462 36120 20580 36236
rect 22080 36236 22260 36238
rect 22080 36180 22086 36236
rect 22142 36180 22260 36236
rect 22080 36120 22260 36180
rect 23760 36236 23940 36238
rect 23760 36180 23766 36236
rect 23822 36180 23940 36236
rect 23760 36120 23940 36180
rect 25440 36236 25620 36238
rect 25440 36180 25446 36236
rect 25502 36180 25620 36236
rect 25440 36120 25620 36180
rect 27120 36236 27300 36238
rect 27120 36180 27126 36236
rect 27182 36180 27300 36236
rect 27120 36120 27300 36180
rect 28800 36238 28918 36300
rect 30542 36238 30660 36300
rect 32222 36238 32340 36300
rect 33902 36238 34020 36300
rect 28800 36236 28980 36238
rect 28800 36180 28806 36236
rect 28862 36180 28980 36236
rect 28800 36120 28980 36180
rect 30480 36236 30660 36238
rect 30480 36180 30486 36236
rect 30542 36180 30660 36236
rect 30480 36120 30660 36180
rect 32160 36236 32340 36238
rect 32160 36180 32166 36236
rect 32222 36180 32340 36236
rect 32160 36120 32340 36180
rect 33840 36236 34020 36238
rect 33840 36180 33846 36236
rect 33902 36180 34020 36236
rect 33840 36120 34020 36180
rect 35520 36238 35638 36300
rect 37200 36238 37318 36300
rect 38942 36238 39060 36300
rect 35520 36236 35700 36238
rect 35520 36180 35526 36236
rect 35582 36180 35700 36236
rect 35520 36120 35700 36180
rect 37200 36236 37380 36238
rect 37200 36180 37206 36236
rect 37262 36180 37380 36236
rect 37200 36120 37380 36180
rect 38880 36236 39060 36238
rect 38880 36180 38886 36236
rect 38942 36180 39060 36236
rect 38880 36120 39060 36180
rect 40560 36238 40678 36300
rect 42240 36238 42358 36300
rect 43982 36238 44100 36300
rect 40560 36236 40740 36238
rect 40560 36180 40566 36236
rect 40622 36180 40740 36236
rect 40560 36120 40740 36180
rect 42240 36236 42420 36238
rect 42240 36180 42246 36236
rect 42302 36180 42420 36236
rect 42240 36120 42420 36180
rect 43920 36236 44100 36238
rect 43920 36180 43926 36236
rect 43982 36180 44100 36236
rect 43920 36120 44100 36180
rect 45600 36238 45718 36300
rect 47280 36238 47398 36300
rect 49022 36238 49140 36300
rect 50702 36238 50820 36300
rect 45600 36236 45780 36238
rect 45600 36180 45606 36236
rect 45662 36180 45780 36236
rect 45600 36120 45780 36180
rect 47280 36236 47460 36238
rect 47280 36180 47286 36236
rect 47342 36180 47460 36236
rect 47280 36120 47460 36180
rect 48960 36236 49140 36238
rect 48960 36180 48966 36236
rect 49022 36180 49140 36236
rect 48960 36120 49140 36180
rect 50640 36236 50820 36238
rect 50640 36180 50646 36236
rect 50702 36180 50820 36236
rect 50640 36120 50820 36180
rect 52320 36238 52438 36300
rect 54000 36238 54118 36300
rect 55742 36238 55860 36300
rect 57422 36238 57540 36300
rect 52320 36236 52500 36238
rect 52320 36180 52326 36236
rect 52382 36180 52500 36236
rect 52320 36120 52500 36180
rect 54000 36236 54180 36238
rect 54000 36180 54006 36236
rect 54062 36180 54180 36236
rect 54000 36120 54180 36180
rect 55680 36236 55860 36238
rect 55680 36180 55686 36236
rect 55742 36180 55860 36236
rect 55680 36120 55860 36180
rect 57360 36236 57540 36238
rect 57360 36180 57366 36236
rect 57422 36180 57540 36236
rect 57360 36120 57540 36180
rect 59040 36238 59158 36300
rect 60782 36238 60900 36300
rect 62462 36238 62580 36300
rect 59040 36236 59220 36238
rect 59040 36180 59046 36236
rect 59102 36180 59220 36236
rect 59040 36120 59220 36180
rect 60720 36236 60900 36238
rect 60720 36180 60726 36236
rect 60782 36180 60900 36236
rect 60720 36120 60900 36180
rect 62400 36236 62580 36238
rect 62400 36180 62406 36236
rect 62462 36180 62580 36236
rect 62400 36120 62580 36180
rect 64080 36238 64198 36300
rect 65822 36238 65940 36300
rect 64080 36236 64260 36238
rect 64080 36180 64086 36236
rect 64142 36180 64260 36236
rect 64080 36120 64260 36180
rect 65760 36236 65940 36238
rect 65760 36180 65766 36236
rect 65822 36180 65940 36236
rect 65760 36120 65940 36180
rect 67440 36238 67558 36300
rect 69120 36238 69238 36300
rect 70862 36238 70980 36300
rect 72542 36238 72660 36300
rect 67440 36236 67620 36238
rect 67440 36180 67446 36236
rect 67502 36180 67620 36236
rect 67440 36120 67620 36180
rect 69120 36236 69300 36238
rect 69120 36180 69126 36236
rect 69182 36180 69300 36236
rect 69120 36120 69300 36180
rect 70800 36236 70980 36238
rect 70800 36180 70806 36236
rect 70862 36180 70980 36236
rect 70800 36120 70980 36180
rect 72480 36236 72660 36238
rect 72480 36180 72486 36236
rect 72542 36180 72660 36236
rect 72480 36120 72660 36180
rect 1142 35528 1740 35580
rect 1142 35520 1590 35528
rect 1560 35472 1590 35520
rect 1646 35472 1740 35528
rect 1560 35400 1740 35472
rect 73920 35528 74100 35580
rect 73920 35472 73938 35528
rect 73994 35472 74100 35528
rect 73920 35460 74100 35472
rect 73920 35400 74398 35460
rect 14400 35278 14518 35340
rect 14582 35280 15420 35340
rect 14400 35160 14580 35278
rect 15120 35222 15420 35280
rect 19622 35278 19740 35340
rect 19560 35222 19740 35278
rect 15120 35160 15238 35222
rect 15302 35160 15420 35222
rect 19622 35160 19740 35222
rect 18360 34920 19558 34980
rect 18360 34860 18540 34920
rect 18360 34800 19678 34860
rect 1142 33848 1740 33900
rect 1142 33840 1590 33848
rect 1560 33792 1590 33840
rect 1646 33792 1740 33848
rect 1560 33720 1740 33792
rect 73920 33848 74100 33900
rect 73920 33792 73938 33848
rect 73994 33792 74100 33848
rect 14462 33720 15420 33780
rect 14462 33718 14580 33720
rect 14400 33660 14580 33718
rect 14400 33600 14998 33660
rect 15120 33600 15420 33720
rect 19560 33720 20398 33780
rect 19560 33662 19740 33720
rect 73920 33780 74100 33792
rect 73920 33720 74398 33780
rect 19622 33600 19740 33662
rect 18360 33360 19558 33420
rect 18360 33302 18540 33360
rect 18360 33240 18478 33302
rect 1560 32168 1740 32220
rect 1560 32112 1590 32168
rect 1646 32112 1740 32168
rect 1560 32100 1740 32112
rect 1142 32040 1740 32100
rect 14400 32100 14580 32220
rect 15120 32158 15238 32220
rect 15302 32158 15420 32220
rect 15120 32146 15420 32158
rect 15120 32102 15180 32146
rect 14400 32040 15118 32100
rect 15360 32040 15420 32146
rect 19560 32158 19678 32220
rect 73920 32168 74100 32220
rect 19560 32102 19740 32158
rect 19622 32040 19740 32102
rect 73920 32112 73938 32168
rect 73994 32112 74100 32168
rect 73920 32100 74100 32112
rect 73920 32040 74398 32100
rect 18360 31800 19558 31860
rect 18360 31740 18540 31800
rect 18360 31680 19678 31740
rect 14400 30660 14580 30780
rect 15062 30720 15180 30780
rect 15120 30666 15180 30720
rect 15360 30666 15420 30780
rect 15120 30660 15420 30666
rect 14400 30600 15420 30660
rect 1560 30488 1740 30540
rect 1560 30432 1590 30488
rect 1646 30432 1740 30488
rect 1560 30420 1740 30432
rect 19560 30480 19740 30660
rect 73920 30488 74398 30540
rect 1142 30360 1740 30420
rect 18360 30358 18478 30420
rect 19560 30420 19620 30480
rect 18542 30360 19620 30420
rect 73920 30432 73938 30488
rect 73994 30480 74398 30488
rect 73994 30432 74100 30480
rect 73920 30360 74100 30432
rect 18360 30300 18540 30358
rect 18360 30240 19558 30300
rect 14520 29280 15118 29340
rect 14520 29220 14580 29280
rect 14400 29160 15180 29220
rect 14400 29040 14580 29160
rect 15120 29126 15180 29160
rect 15360 29126 15420 29220
rect 15120 29040 15420 29126
rect 19560 29158 19678 29220
rect 19560 29040 19740 29158
rect 19560 28860 19620 29040
rect 1560 28808 1740 28860
rect 1560 28752 1590 28808
rect 1646 28752 1740 28808
rect 1560 28740 1740 28752
rect 1142 28680 1740 28740
rect 18360 28800 19620 28860
rect 73920 28808 74398 28860
rect 18360 28742 18540 28800
rect 73920 28752 73938 28808
rect 73994 28800 74398 28808
rect 73994 28752 74100 28800
rect 18360 28680 18478 28742
rect 73920 28680 74100 28752
rect 19622 27598 19740 27660
rect 19560 27480 19740 27598
rect 19560 27420 19620 27480
rect 18360 27360 19620 27420
rect 18360 27300 18540 27360
rect 18360 27240 19558 27300
rect 1142 27128 1740 27180
rect 1142 27120 1590 27128
rect 1560 27072 1590 27120
rect 1646 27072 1740 27128
rect 1560 27000 1740 27072
rect 73920 27128 74398 27180
rect 73920 27072 73938 27128
rect 73994 27120 74398 27128
rect 73994 27072 74100 27120
rect 73920 27000 74100 27072
rect 14400 25980 14580 26100
rect 15120 25982 15420 26100
rect 14400 25920 15118 25980
rect 15182 25920 15420 25982
rect 19560 25920 19740 26100
rect 18360 25798 18478 25860
rect 19560 25860 19620 25920
rect 18542 25800 19620 25860
rect 18360 25740 18540 25798
rect 18360 25680 19438 25740
rect 1142 25448 1740 25500
rect 1142 25440 1590 25448
rect 1560 25392 1590 25440
rect 1646 25392 1740 25448
rect 1560 25320 1740 25392
rect 73920 25448 74100 25500
rect 73920 25392 73938 25448
rect 73994 25392 74100 25448
rect 73920 25380 74100 25392
rect 73920 25320 74398 25380
rect 14400 24422 14580 24540
rect 14462 24420 14580 24422
rect 15120 24420 15420 24540
rect 19622 24478 19740 24540
rect 14462 24360 15420 24420
rect 19560 24422 19740 24478
rect 19560 24360 19678 24422
rect 19560 24300 19620 24360
rect 18360 24240 19620 24300
rect 18360 24120 18540 24240
rect 1142 23768 1740 23820
rect 1142 23760 1590 23768
rect 1560 23712 1590 23760
rect 1646 23712 1740 23768
rect 1560 23640 1740 23712
rect 73920 23768 74100 23820
rect 73920 23712 73938 23768
rect 73994 23712 74100 23768
rect 73920 23700 74100 23712
rect 73920 23640 74398 23700
rect 14520 23040 15118 23100
rect 14520 22980 14580 23040
rect 14400 22920 15420 22980
rect 14400 22800 14580 22920
rect 15120 22910 15420 22920
rect 19502 22920 19740 22980
rect 15120 22800 15180 22910
rect 15360 22862 15420 22910
rect 19560 22860 19740 22920
rect 18360 22800 19740 22860
rect 18360 22740 18540 22800
rect 18360 22680 19438 22740
rect 1560 22088 1740 22140
rect 1560 22032 1590 22088
rect 1646 22032 1740 22088
rect 1560 22020 1740 22032
rect 1142 21960 1740 22020
rect 73920 22088 74100 22140
rect 73920 22032 73938 22088
rect 73994 22032 74100 22088
rect 73920 22020 74100 22032
rect 73920 21960 74398 22020
rect 14462 21478 14580 21540
rect 14400 21420 14580 21478
rect 15120 21430 15180 21540
rect 15360 21430 15420 21540
rect 19560 21480 19678 21540
rect 15120 21420 15420 21430
rect 19666 21478 19678 21480
rect 14400 21360 15780 21420
rect 15720 21300 15780 21360
rect 15720 21240 19558 21300
rect 18360 21120 18540 21240
rect 19666 21300 19740 21478
rect 19622 21240 19740 21300
rect 1560 20408 1740 20460
rect 1560 20352 1590 20408
rect 1646 20352 1740 20408
rect 1560 20340 1740 20352
rect 1142 20280 1740 20340
rect 73920 20408 74398 20460
rect 73920 20352 73938 20408
rect 73994 20400 74398 20408
rect 73994 20352 74100 20400
rect 73920 20280 74100 20352
rect 14400 19862 14580 19980
rect 14462 19860 14580 19862
rect 15120 19918 15358 19980
rect 19502 19920 19740 19980
rect 15120 19860 15420 19918
rect 14462 19800 15420 19860
rect 19560 19800 19740 19920
rect 19560 19740 19620 19800
rect 18360 19680 19620 19740
rect 18360 19560 18540 19680
rect 1560 18728 1740 18780
rect 1560 18672 1590 18728
rect 1646 18672 1740 18728
rect 1560 18660 1740 18672
rect 1142 18600 1740 18660
rect 73920 18728 74398 18780
rect 73920 18672 73938 18728
rect 73994 18720 74398 18728
rect 73994 18672 74100 18720
rect 73920 18600 74100 18672
rect 19622 18358 19740 18420
rect 19560 18300 19740 18358
rect 18360 18240 19740 18300
rect 18360 18120 18540 18240
rect 12840 17520 14398 17580
rect 12840 17460 13020 17520
rect 12840 17400 14398 17460
rect 1142 17048 1740 17100
rect 1142 17040 1590 17048
rect 1560 16992 1590 17040
rect 1646 16992 1740 17048
rect 1560 16920 1740 16992
rect 73920 17048 74398 17100
rect 73920 16992 73938 17048
rect 73994 17040 74398 17048
rect 73994 16992 74100 17040
rect 73920 16920 74100 16992
rect 14462 16800 15420 16860
rect 14462 16798 14580 16800
rect 14400 16742 14580 16798
rect 12840 16622 13020 16740
rect 14462 16680 14580 16742
rect 15120 16680 15420 16800
rect 19560 16740 19740 16860
rect 18360 16680 19740 16740
rect 18360 16622 18540 16680
rect 12840 16560 12958 16622
rect 18360 16560 18478 16622
rect 12840 15840 14398 15900
rect 12840 15782 13020 15840
rect 12902 15720 13020 15782
rect 12360 15570 12540 15660
rect 12360 15540 12391 15570
rect 0 15514 12391 15540
rect 12447 15514 12540 15570
rect 13469 15574 14215 15576
rect 13469 15518 13471 15574
rect 13527 15518 14157 15574
rect 14213 15518 14215 15574
rect 13469 15516 14215 15518
rect 0 15480 12540 15514
rect 1142 15368 1740 15420
rect 1142 15360 1590 15368
rect 1560 15312 1590 15360
rect 1646 15312 1740 15368
rect 1560 15240 1740 15312
rect 73920 15368 74100 15420
rect 73920 15312 73938 15368
rect 73994 15312 74100 15368
rect 73920 15300 74100 15312
rect 14400 15240 15420 15300
rect 14400 15120 14580 15240
rect 15120 15214 15420 15240
rect 15120 15120 15180 15214
rect 15360 15120 15420 15214
rect 18360 15240 19740 15300
rect 73920 15240 74398 15300
rect 18360 15120 18540 15240
rect 19560 15182 19740 15240
rect 19560 15120 19678 15182
rect 12840 14998 12958 15060
rect 14400 15060 14460 15120
rect 13022 15000 14460 15060
rect 12840 14942 13020 14998
rect 12840 14880 12958 14942
rect 12360 14386 12540 14460
rect 12360 14340 12391 14386
rect 0 14330 12391 14340
rect 12447 14330 12540 14386
rect 0 14280 12540 14330
rect 13469 14382 14147 14384
rect 13469 14326 13471 14382
rect 13527 14326 14089 14382
rect 14145 14326 14147 14382
rect 13469 14324 14147 14326
rect 12902 14158 13020 14220
rect 12840 14102 13020 14158
rect 12902 14100 13020 14102
rect 12902 14040 14398 14100
rect 12360 13894 12540 13980
rect 12360 13860 12391 13894
rect 0 13838 12391 13860
rect 12447 13838 12540 13894
rect 13469 13898 14079 13900
rect 13469 13842 13471 13898
rect 13527 13842 14021 13898
rect 14077 13842 14079 13898
rect 13469 13840 14079 13842
rect 0 13800 12540 13838
rect 1142 13688 1740 13740
rect 1142 13680 1590 13688
rect 1560 13632 1590 13680
rect 1646 13632 1740 13688
rect 14462 13678 14580 13740
rect 1560 13560 1740 13632
rect 14400 13620 14580 13678
rect 15120 13674 15420 13740
rect 15120 13620 15180 13674
rect 14400 13560 15180 13620
rect 15360 13560 15420 13674
rect 18360 13678 18478 13740
rect 18360 13620 18540 13678
rect 19560 13622 19740 13740
rect 18360 13560 19558 13620
rect 19622 13560 19740 13622
rect 73920 13688 74100 13740
rect 73920 13632 73938 13688
rect 73994 13632 74100 13688
rect 73920 13620 74100 13632
rect 73920 13560 74398 13620
rect 12840 13318 12958 13380
rect 12840 13262 13020 13318
rect 12840 13200 12958 13262
rect 12360 12710 12540 12780
rect 12360 12660 12391 12710
rect 0 12654 12391 12660
rect 12447 12654 12540 12710
rect 0 12600 12540 12654
rect 13469 12706 14011 12708
rect 13469 12650 13471 12706
rect 13527 12650 13953 12706
rect 14009 12650 14011 12706
rect 13469 12648 14011 12650
rect 12902 12478 13020 12540
rect 12840 12422 13020 12478
rect 12902 12360 13020 12422
rect 12360 12218 12540 12300
rect 14400 12240 15180 12300
rect 12360 12162 12391 12218
rect 12447 12182 12540 12218
rect 13469 12222 13943 12224
rect 12447 12162 12478 12182
rect 12360 12120 12478 12162
rect 13469 12166 13471 12222
rect 13527 12166 13885 12222
rect 13941 12166 13943 12222
rect 14400 12182 14580 12240
rect 13469 12164 13943 12166
rect 14462 12120 14580 12182
rect 15120 12194 15180 12240
rect 15360 12194 15420 12300
rect 15120 12180 15420 12194
rect 19560 12238 19678 12300
rect 19560 12180 19740 12238
rect 15120 12120 15780 12180
rect 15720 12060 15780 12120
rect 18360 12120 20278 12180
rect 18360 12060 18540 12120
rect 1560 12008 1740 12060
rect 1560 11952 1590 12008
rect 1646 11952 1740 12008
rect 15720 12000 18540 12060
rect 73920 12008 74100 12060
rect 1560 11940 1740 11952
rect 1142 11880 1740 11940
rect 73920 11952 73938 12008
rect 73994 11952 74100 12008
rect 73920 11940 74100 11952
rect 73920 11880 74398 11940
rect 12840 11638 12958 11700
rect 13022 11640 14398 11700
rect 12840 11520 13020 11638
rect 12114 11088 12212 11090
rect 12114 11032 12116 11088
rect 12172 11032 12212 11088
rect 12114 11030 12212 11032
rect 12389 11034 12449 11036
rect 12389 10982 12391 11034
rect 12447 10978 12449 11034
rect 12422 10976 12449 10978
rect 13469 11030 13875 11032
rect 13469 10974 13471 11030
rect 13527 10974 13817 11030
rect 13873 10974 13875 11030
rect 13469 10972 13875 10974
rect 12902 10798 13020 10860
rect 12840 10740 13020 10798
rect 12840 10680 15420 10740
rect 14400 10560 14580 10680
rect 15120 10620 15420 10680
rect 18360 10680 19558 10740
rect 18360 10622 18540 10680
rect 19622 10678 19740 10740
rect 15120 10560 15718 10620
rect 18422 10560 18540 10622
rect 19560 10620 19740 10678
rect 19560 10560 20460 10620
rect 20280 10500 20460 10560
rect 21840 10560 23580 10620
rect 21840 10500 22020 10560
rect 20280 10440 22020 10500
rect 23400 10500 23580 10560
rect 24542 10560 25140 10620
rect 23400 10440 24598 10500
rect 24960 10500 25140 10560
rect 26222 10560 26700 10620
rect 26520 10500 26700 10560
rect 27782 10560 29820 10620
rect 28080 10500 28260 10560
rect 24960 10440 28260 10500
rect 29640 10500 29820 10560
rect 31080 10502 31260 10620
rect 32462 10560 32820 10620
rect 29342 10440 31078 10500
rect 31142 10500 31260 10502
rect 32640 10500 32820 10560
rect 34022 10560 34380 10620
rect 34200 10500 34380 10560
rect 31142 10440 34380 10500
rect 35760 10500 35940 10620
rect 37320 10502 37500 10620
rect 38702 10560 39060 10620
rect 35582 10440 37318 10500
rect 37382 10500 37500 10502
rect 38880 10500 39060 10560
rect 40142 10560 40620 10620
rect 40440 10500 40620 10560
rect 41702 10560 42180 10620
rect 42000 10500 42180 10560
rect 37382 10440 42180 10500
rect 43560 10500 43740 10620
rect 43142 10440 43740 10500
rect 1560 10328 1740 10380
rect 1560 10272 1590 10328
rect 1646 10272 1740 10328
rect 1560 10260 1740 10272
rect 1142 10200 1740 10260
rect 73920 10328 74100 10380
rect 73920 10272 73938 10328
rect 73994 10272 74100 10328
rect 73920 10260 74100 10272
rect 73920 10200 74398 10260
rect 13664 10155 18536 10157
rect 13664 10099 13666 10155
rect 13722 10099 18478 10155
rect 18534 10099 18536 10155
rect 13664 10097 18536 10099
rect 20342 9718 20460 9780
rect 20280 9662 20460 9718
rect 15782 9600 18358 9660
rect 17520 9542 17700 9600
rect 20342 9660 20460 9662
rect 21840 9660 22020 9780
rect 23400 9720 25140 9780
rect 23400 9660 23580 9720
rect 24960 9662 25140 9720
rect 26520 9662 26700 9780
rect 28080 9662 28260 9780
rect 29640 9662 29820 9780
rect 20342 9600 23580 9660
rect 25022 9600 25140 9662
rect 26582 9660 26700 9662
rect 26582 9600 28078 9660
rect 28142 9600 28260 9662
rect 29702 9660 29820 9662
rect 31080 9662 31260 9780
rect 32640 9662 32820 9780
rect 34200 9720 39060 9780
rect 34200 9662 34380 9720
rect 35760 9662 35940 9720
rect 31080 9660 31198 9662
rect 29702 9600 31198 9660
rect 32640 9660 32758 9662
rect 31262 9600 32758 9660
rect 34200 9600 34318 9662
rect 35822 9600 35940 9662
rect 37320 9662 37500 9720
rect 38880 9662 39060 9720
rect 40440 9662 40620 9780
rect 42000 9662 42180 9780
rect 43560 9662 43740 9780
rect 37320 9600 37438 9662
rect 38880 9600 38998 9662
rect 40440 9600 40558 9662
rect 42000 9600 42118 9662
rect 43560 9600 43678 9662
rect 44880 9600 46318 9660
rect 17582 9480 17700 9542
rect 30840 9480 31078 9540
rect 24542 9360 24598 9420
rect 24662 9358 24700 9396
rect 24640 9336 24700 9358
rect 24750 9358 24838 9390
rect 26222 9358 26256 9396
rect 27782 9358 27812 9396
rect 30840 9396 30900 9480
rect 33960 9480 35580 9540
rect 33960 9422 34020 9480
rect 35520 9422 35580 9480
rect 37080 9480 37318 9540
rect 29342 9358 29368 9396
rect 30840 9360 30924 9396
rect 24750 9310 24870 9358
rect 26196 9336 26256 9358
rect 27752 9336 27812 9358
rect 29308 9336 29368 9358
rect 30864 9336 30924 9360
rect 32462 9358 32480 9396
rect 34022 9358 34036 9396
rect 37080 9396 37140 9480
rect 43200 9480 43318 9540
rect 43200 9422 43260 9480
rect 44880 9540 44940 9600
rect 47942 9600 49438 9660
rect 44760 9480 44940 9540
rect 44760 9422 44820 9480
rect 35582 9358 35592 9396
rect 37080 9360 37148 9396
rect 32420 9336 32480 9358
rect 33976 9336 34036 9358
rect 35532 9336 35592 9358
rect 37088 9336 37148 9360
rect 38702 9358 38704 9396
rect 40142 9358 40260 9396
rect 41582 9360 41638 9420
rect 41702 9358 41816 9396
rect 38644 9336 38704 9358
rect 40110 9336 40260 9358
rect 41670 9336 41816 9358
rect 41836 9358 41878 9390
rect 43142 9360 43198 9420
rect 43262 9358 43372 9396
rect 24720 9308 24870 9310
rect 24720 9252 24722 9308
rect 24778 9280 24870 9308
rect 26276 9308 26336 9310
rect 24778 9252 24780 9280
rect 24720 9250 24780 9252
rect 26276 9250 26278 9308
rect 26334 9302 26336 9308
rect 27832 9308 27892 9310
rect 27832 9252 27834 9308
rect 27890 9302 27892 9308
rect 29388 9308 29448 9310
rect 27832 9250 27838 9252
rect 29388 9252 29390 9308
rect 29446 9302 29448 9308
rect 30944 9308 31004 9310
rect 29388 9250 29398 9252
rect 30944 9252 30946 9308
rect 31002 9302 31004 9308
rect 32500 9308 32560 9310
rect 30944 9250 30958 9252
rect 32500 9252 32502 9308
rect 32558 9302 32560 9308
rect 34056 9308 34116 9310
rect 32500 9250 32518 9252
rect 34056 9252 34058 9308
rect 34114 9302 34116 9308
rect 35612 9308 35672 9310
rect 34056 9250 34078 9252
rect 35612 9252 35614 9308
rect 35670 9302 35672 9308
rect 37168 9308 37228 9310
rect 35612 9250 35638 9252
rect 37168 9252 37170 9308
rect 37226 9302 37228 9308
rect 38724 9308 38784 9310
rect 37168 9250 37198 9252
rect 38724 9252 38726 9308
rect 38782 9302 38784 9308
rect 40280 9308 40340 9310
rect 38724 9250 38758 9252
rect 40280 9252 40282 9308
rect 40338 9302 40340 9308
rect 41836 9308 41896 9358
rect 43230 9336 43372 9358
rect 43392 9358 43438 9390
rect 44222 9360 44758 9420
rect 44822 9358 44928 9396
rect 40280 9250 40318 9252
rect 41836 9252 41838 9308
rect 41894 9252 41896 9308
rect 41836 9250 41896 9252
rect 43392 9308 43452 9358
rect 44790 9336 44928 9358
rect 44948 9358 44998 9390
rect 46382 9358 46484 9396
rect 43392 9252 43394 9308
rect 43450 9252 43452 9308
rect 43392 9250 43452 9252
rect 44948 9308 45008 9358
rect 44948 9252 44950 9308
rect 45006 9252 45008 9308
rect 44948 9250 45008 9252
rect 46320 9336 46484 9358
rect 13664 9229 45226 9231
rect 13664 9173 13666 9229
rect 13722 9173 45168 9229
rect 45224 9173 45226 9229
rect 13664 9171 45226 9173
rect 46320 9180 46380 9336
rect 46560 9310 46620 9420
rect 47942 9358 48040 9396
rect 46504 9308 46620 9310
rect 46504 9252 46506 9308
rect 46562 9302 46620 9308
rect 47880 9336 48040 9358
rect 46504 9250 46558 9252
rect 47880 9180 47940 9336
rect 48120 9310 48180 9420
rect 49502 9358 49620 9420
rect 48060 9308 48180 9310
rect 48060 9252 48062 9308
rect 48118 9302 48180 9308
rect 48060 9250 48118 9252
rect 49440 9300 49620 9358
rect 51000 9360 54300 9420
rect 51000 9300 51180 9360
rect 49440 9240 51180 9300
rect 52560 9240 52740 9360
rect 54120 9300 54300 9360
rect 55680 9360 57420 9420
rect 55680 9300 55860 9360
rect 54120 9240 55860 9300
rect 57240 9300 57420 9360
rect 58800 9300 58980 9420
rect 60360 9360 62100 9420
rect 60360 9300 60540 9360
rect 57240 9240 60540 9300
rect 61920 9300 62100 9360
rect 63480 9300 63660 9420
rect 65040 9300 65220 9420
rect 66600 9360 71460 9420
rect 66600 9300 66780 9360
rect 61920 9240 66780 9300
rect 68160 9240 68340 9360
rect 69720 9240 69900 9360
rect 71280 9300 71460 9360
rect 72840 9300 73020 9420
rect 71280 9240 74998 9300
rect 46320 9120 47940 9180
rect 41582 9000 43198 9060
rect 43382 9000 44758 9060
rect 17520 8760 20278 8820
rect 1560 8648 1740 8700
rect 1560 8592 1590 8648
rect 1646 8592 1740 8648
rect 17520 8640 17700 8760
rect 73920 8648 74398 8700
rect 1560 8580 1740 8592
rect 1142 8520 1740 8580
rect 73920 8592 73938 8648
rect 73994 8640 74398 8648
rect 73994 8592 74100 8640
rect 73920 8520 74100 8592
rect 13664 8485 19670 8487
rect 13664 8429 13666 8485
rect 13722 8429 19612 8485
rect 19668 8429 19670 8485
rect 13664 8427 19670 8429
rect 24600 8400 24958 8460
rect 24600 8340 24780 8400
rect 26160 8400 26518 8460
rect 26160 8340 26340 8400
rect 27720 8400 28078 8460
rect 24600 8280 26340 8340
rect 27720 8340 27900 8400
rect 29280 8400 29638 8460
rect 29280 8340 29460 8400
rect 30840 8400 31198 8460
rect 27720 8280 29460 8340
rect 30840 8280 31020 8400
rect 32400 8400 32758 8460
rect 32400 8340 32580 8400
rect 33960 8400 34318 8460
rect 33960 8340 34140 8400
rect 35520 8400 35758 8460
rect 32400 8280 34140 8340
rect 35520 8280 35700 8400
rect 37080 8400 37438 8460
rect 37080 8280 37260 8400
rect 38640 8400 38998 8460
rect 38640 8340 38820 8400
rect 40080 8400 40558 8460
rect 40080 8390 40380 8400
rect 41640 8400 42118 8460
rect 40080 8340 40140 8390
rect 38640 8280 40140 8340
rect 40320 8340 40380 8390
rect 41640 8340 41820 8400
rect 43200 8400 43678 8460
rect 43200 8340 43380 8400
rect 73920 8460 73980 8520
rect 44760 8400 48060 8460
rect 44760 8340 44940 8400
rect 40320 8280 44940 8340
rect 46320 8280 46500 8400
rect 47880 8340 48060 8400
rect 49440 8340 49620 8460
rect 51000 8400 54300 8460
rect 51000 8340 51180 8400
rect 47880 8280 51180 8340
rect 52560 8280 52740 8400
rect 54120 8340 54300 8400
rect 55680 8340 55860 8460
rect 57240 8340 57420 8460
rect 58800 8340 58980 8460
rect 60360 8400 62100 8460
rect 60360 8340 60540 8400
rect 54120 8280 60540 8340
rect 61920 8340 62100 8400
rect 63480 8340 63660 8460
rect 65040 8340 65220 8460
rect 66600 8400 71460 8460
rect 66600 8340 66780 8400
rect 61920 8280 66780 8340
rect 68160 8280 68340 8400
rect 69720 8280 69900 8400
rect 71280 8340 71460 8400
rect 72840 8400 73980 8460
rect 72840 8340 73020 8400
rect 71280 8280 73020 8340
rect 17582 7918 17700 7980
rect 17520 7800 17700 7918
rect 20640 7080 23220 7140
rect 1142 6968 1740 7020
rect 1142 6960 1590 6968
rect 1560 6912 1590 6960
rect 1646 6912 1740 6968
rect 20640 6960 20820 7080
rect 21480 6960 21660 7080
rect 22200 6960 22380 7080
rect 23040 7020 23220 7080
rect 23760 7080 24780 7140
rect 23760 7020 23940 7080
rect 23040 6960 23940 7020
rect 24600 7020 24780 7080
rect 25320 7020 25500 7140
rect 26160 7020 26340 7140
rect 26880 7080 31020 7140
rect 26880 7020 27060 7080
rect 24600 6960 27060 7020
rect 27720 6960 27900 7080
rect 28440 6960 28620 7080
rect 29280 6960 29460 7080
rect 30000 6960 30180 7080
rect 30840 7020 31020 7080
rect 31560 7020 31740 7140
rect 32400 7020 32580 7140
rect 33120 7020 33300 7140
rect 33840 7067 34140 7140
rect 33840 7020 33900 7067
rect 30840 6960 33900 7020
rect 34080 7020 34140 7067
rect 34680 7020 34860 7140
rect 35400 7080 36420 7140
rect 35400 7020 35580 7080
rect 34080 6960 35580 7020
rect 36240 7020 36420 7080
rect 36960 7080 38700 7140
rect 36960 7020 37140 7080
rect 36240 6960 37140 7020
rect 37800 6960 37980 7080
rect 38520 7020 38700 7080
rect 39360 7020 39540 7140
rect 40080 7080 41100 7140
rect 40080 7020 40260 7080
rect 38520 6960 40260 7020
rect 40920 7020 41100 7080
rect 41640 7020 41820 7140
rect 42480 7080 43380 7140
rect 42480 7020 42660 7080
rect 40920 6960 42660 7020
rect 43200 7020 43380 7080
rect 44040 7078 44158 7140
rect 44222 7080 44940 7140
rect 44040 7020 44220 7078
rect 43200 6960 44220 7020
rect 44760 6960 44940 7080
rect 73920 6968 74398 7020
rect 1560 6840 1740 6912
rect 73920 6912 73938 6968
rect 73994 6960 74398 6968
rect 73994 6912 74100 6960
rect 73920 6840 74100 6912
rect 2400 6302 2580 6420
rect 542 6240 2398 6300
rect 2462 6240 2580 6302
rect 2635 6096 2695 6098
rect 2635 6040 2637 6096
rect 2693 6040 2695 6096
rect 2635 6038 2695 6040
rect 5880 5881 6060 5940
rect 5880 5825 5997 5881
rect 6053 5825 6060 5881
rect 5880 5822 6060 5825
rect 5880 5760 5998 5822
rect 2400 5400 2580 5580
rect 2400 5340 2460 5400
rect 1142 5288 2460 5340
rect 1142 5280 1590 5288
rect 1560 5232 1590 5280
rect 1646 5280 2460 5288
rect 1646 5232 1740 5280
rect 1560 5160 1740 5232
rect 20040 5220 20220 5340
rect 20880 5280 21780 5340
rect 20880 5220 21060 5280
rect 20040 5160 21060 5220
rect 21600 5220 21780 5280
rect 22440 5220 22620 5340
rect 23160 5280 24900 5340
rect 23160 5220 23340 5280
rect 21600 5160 23340 5220
rect 24000 5160 24180 5280
rect 24720 5220 24900 5280
rect 25560 5280 27300 5340
rect 25560 5220 25740 5280
rect 24720 5160 25740 5220
rect 26280 5160 26460 5280
rect 27120 5220 27300 5280
rect 27840 5220 28020 5340
rect 28680 5220 28860 5340
rect 29400 5280 30420 5340
rect 29400 5220 29580 5280
rect 27120 5160 29580 5220
rect 30240 5220 30420 5280
rect 30960 5280 33540 5340
rect 30960 5220 31140 5280
rect 30240 5160 31140 5220
rect 31800 5160 31980 5280
rect 32520 5160 32700 5280
rect 33360 5220 33540 5280
rect 34080 5280 35100 5340
rect 34080 5220 34260 5280
rect 33360 5160 34260 5220
rect 34920 5222 35100 5280
rect 34920 5160 35038 5222
rect 35640 5220 35820 5340
rect 36480 5280 37380 5340
rect 36480 5220 36660 5280
rect 35102 5160 36660 5220
rect 37200 5220 37380 5280
rect 38040 5220 38220 5340
rect 38760 5220 38940 5340
rect 39480 5220 39660 5340
rect 40320 5220 40500 5340
rect 41040 5220 41220 5340
rect 41880 5280 42780 5340
rect 41880 5220 42060 5280
rect 37200 5160 42060 5220
rect 42600 5220 42780 5280
rect 43440 5220 43620 5340
rect 44160 5220 44340 5340
rect 45000 5220 45180 5340
rect 42600 5160 45180 5220
rect 73920 5288 74100 5340
rect 73920 5232 73938 5288
rect 73994 5232 74100 5288
rect 73920 5220 74100 5232
rect 73920 5160 74398 5220
rect 2635 4912 2695 4914
rect 2635 4856 2637 4912
rect 2693 4856 2695 4912
rect 2635 4854 2695 4856
rect 2462 4678 2580 4740
rect 2400 4560 2580 4678
rect 1142 3608 1740 3660
rect 1142 3600 1590 3608
rect 1560 3552 1590 3600
rect 1646 3552 1740 3608
rect 1560 3480 1740 3552
rect 73920 3608 74100 3660
rect 73920 3552 73938 3608
rect 73994 3552 74100 3608
rect 73920 3540 74100 3552
rect 73920 3480 74398 3540
rect 15840 3180 16020 3300
rect 17280 3180 17460 3300
rect 18840 3180 19020 3300
rect 20280 3180 20460 3300
rect 21720 3180 21900 3300
rect 23280 3240 26340 3300
rect 23280 3180 23460 3240
rect 15840 3120 23460 3180
rect 24720 3120 24900 3240
rect 26160 3180 26340 3240
rect 27720 3240 30780 3300
rect 27720 3180 27900 3240
rect 26160 3120 27900 3180
rect 29160 3120 29340 3240
rect 30600 3180 30780 3240
rect 32160 3180 32340 3300
rect 33600 3180 33780 3300
rect 35102 3240 36780 3300
rect 35102 3238 35220 3240
rect 35040 3180 35220 3238
rect 30600 3120 35518 3180
rect 36600 3180 36780 3240
rect 38040 3180 38220 3300
rect 39480 3180 39660 3300
rect 36600 3120 39660 3180
rect 12114 2732 28514 2734
rect 12114 2676 12116 2732
rect 12172 2678 28514 2732
rect 12172 2676 15355 2678
rect 12114 2674 15355 2676
rect 15353 2622 15355 2674
rect 15411 2674 16837 2678
rect 15411 2622 15413 2674
rect 15353 2580 15413 2622
rect 16835 2622 16837 2674
rect 16893 2674 18319 2678
rect 16893 2622 16895 2674
rect 16835 2580 16895 2622
rect 18317 2622 18319 2674
rect 18375 2674 19801 2678
rect 18375 2622 18377 2674
rect 15302 2520 15420 2580
rect 16800 2520 16918 2580
rect 18317 2580 18377 2622
rect 19799 2622 19801 2674
rect 19857 2674 21283 2678
rect 19857 2622 19859 2674
rect 18302 2520 18420 2580
rect 19799 2580 19859 2622
rect 21281 2622 21283 2674
rect 21339 2674 22765 2678
rect 21339 2622 21341 2674
rect 21281 2580 21341 2622
rect 22763 2622 22765 2674
rect 22821 2674 24247 2678
rect 22821 2622 22823 2674
rect 22763 2582 22823 2622
rect 24245 2622 24247 2674
rect 24303 2674 25729 2678
rect 24303 2622 24305 2674
rect 19742 2520 19860 2580
rect 21240 2520 21358 2580
rect 22763 2580 22798 2582
rect 22680 2520 22798 2580
rect 24245 2580 24305 2622
rect 25727 2622 25729 2674
rect 25785 2674 27211 2678
rect 25785 2622 25787 2674
rect 24240 2520 24358 2580
rect 25727 2580 25787 2622
rect 27209 2622 27211 2674
rect 27267 2674 28514 2678
rect 28691 2678 28751 2680
rect 27267 2622 27269 2674
rect 27209 2582 27269 2622
rect 28691 2622 28693 2678
rect 28749 2622 28751 2678
rect 25680 2520 25798 2580
rect 27209 2580 27238 2582
rect 27120 2520 27238 2580
rect 28691 2580 28751 2622
rect 30173 2678 30233 2680
rect 30173 2622 30175 2678
rect 30231 2622 30233 2678
rect 28680 2520 28798 2580
rect 30173 2580 30233 2622
rect 31655 2678 31715 2680
rect 31655 2622 31657 2678
rect 31713 2622 31715 2678
rect 31655 2582 31715 2622
rect 33137 2678 33197 2680
rect 33137 2622 33139 2678
rect 33195 2622 33197 2678
rect 33137 2582 33197 2622
rect 34619 2678 34679 2680
rect 34619 2622 34621 2678
rect 34677 2622 34679 2678
rect 34619 2582 34679 2622
rect 36101 2678 36161 2680
rect 36101 2622 36103 2678
rect 36159 2622 36161 2678
rect 30120 2520 30238 2580
rect 31655 2580 31678 2582
rect 31560 2520 31678 2580
rect 33182 2580 33197 2582
rect 33182 2520 33300 2580
rect 34622 2580 34679 2582
rect 34622 2520 34740 2580
rect 36101 2580 36161 2622
rect 37583 2678 37643 2680
rect 37583 2622 37585 2678
rect 37641 2622 37643 2678
rect 37583 2580 37643 2622
rect 39065 2678 39125 2680
rect 39065 2622 39067 2678
rect 39123 2622 39125 2678
rect 39065 2582 39125 2622
rect 36062 2520 36180 2580
rect 37560 2520 37678 2580
rect 39065 2580 39118 2582
rect 39000 2520 39118 2580
rect 15840 2340 16020 2460
rect 17280 2340 17460 2460
rect 18840 2340 19020 2460
rect 20280 2340 20460 2460
rect 21720 2340 21900 2460
rect 23280 2340 23460 2460
rect 24720 2340 24900 2460
rect 26160 2340 26340 2460
rect 27720 2340 27900 2460
rect 29160 2340 29340 2460
rect 30600 2340 30780 2460
rect 32160 2342 32340 2460
rect 32160 2340 32278 2342
rect 15840 2280 32278 2340
rect 33600 2340 33780 2460
rect 35040 2340 35220 2460
rect 36600 2340 36780 2460
rect 38040 2340 38220 2460
rect 39480 2340 39660 2460
rect 32342 2280 39660 2340
rect 1560 1928 1740 1980
rect 1560 1872 1590 1928
rect 1646 1872 1740 1928
rect 1560 1860 1740 1872
rect 73920 1928 74100 1980
rect 73920 1872 73938 1928
rect 73994 1872 74100 1928
rect 1560 1800 1918 1860
rect 73920 1860 74100 1872
rect 73920 1800 74398 1860
rect 1920 1536 1926 1558
rect 1982 1536 2100 1620
rect 1920 1502 2100 1536
rect 3600 1592 3780 1620
rect 3600 1536 3606 1592
rect 3662 1536 3780 1592
rect 3600 1502 3780 1536
rect 1920 1440 2038 1502
rect 3662 1440 3780 1502
rect 5280 1592 5460 1620
rect 5280 1536 5286 1592
rect 5342 1536 5460 1592
rect 5280 1502 5460 1536
rect 6960 1592 7140 1620
rect 6960 1536 6966 1592
rect 7022 1536 7140 1592
rect 6960 1502 7140 1536
rect 8640 1592 8820 1620
rect 8640 1536 8646 1592
rect 8702 1536 8820 1592
rect 8640 1502 8820 1536
rect 5280 1440 5398 1502
rect 7022 1440 7140 1502
rect 8702 1440 8820 1502
rect 10320 1592 10500 1620
rect 10320 1536 10326 1592
rect 10382 1536 10500 1592
rect 10320 1502 10500 1536
rect 12000 1592 12180 1620
rect 12000 1536 12006 1592
rect 12062 1536 12180 1592
rect 12000 1502 12180 1536
rect 10320 1440 10438 1502
rect 12062 1440 12180 1502
rect 13680 1592 13860 1620
rect 13680 1536 13686 1592
rect 13742 1536 13860 1592
rect 13680 1502 13860 1536
rect 15360 1592 15540 1620
rect 15360 1536 15366 1592
rect 15422 1536 15540 1592
rect 15360 1502 15540 1536
rect 13680 1440 13798 1502
rect 15422 1440 15540 1502
rect 17040 1592 17220 1620
rect 17040 1536 17046 1592
rect 17102 1536 17220 1592
rect 17040 1502 17220 1536
rect 18720 1592 18900 1620
rect 18720 1536 18726 1592
rect 18782 1536 18900 1592
rect 18720 1502 18900 1536
rect 20400 1592 20580 1620
rect 20400 1536 20406 1592
rect 20462 1536 20580 1592
rect 20400 1502 20580 1536
rect 22080 1592 22260 1620
rect 22080 1536 22086 1592
rect 22142 1536 22260 1592
rect 22080 1502 22260 1536
rect 23760 1592 23940 1620
rect 23760 1536 23766 1592
rect 23822 1536 23940 1592
rect 23760 1502 23940 1536
rect 25440 1592 25620 1620
rect 25440 1536 25446 1592
rect 25502 1536 25620 1592
rect 25440 1502 25620 1536
rect 27120 1592 27300 1620
rect 27120 1536 27126 1592
rect 27182 1536 27300 1592
rect 27120 1502 27300 1536
rect 17040 1440 17158 1502
rect 18720 1440 18838 1502
rect 20400 1440 20518 1502
rect 22080 1440 22198 1502
rect 23760 1440 23878 1502
rect 25502 1440 25620 1502
rect 27182 1440 27300 1502
rect 28800 1592 28980 1620
rect 28800 1536 28806 1592
rect 28862 1536 28980 1592
rect 28800 1500 28980 1536
rect 30480 1592 30660 1620
rect 30480 1536 30486 1592
rect 30542 1536 30660 1592
rect 30480 1502 30660 1536
rect 32160 1592 32340 1620
rect 32160 1536 32166 1592
rect 32222 1536 32340 1592
rect 32160 1502 32340 1536
rect 33840 1592 34020 1620
rect 33840 1536 33846 1592
rect 33902 1536 34020 1592
rect 33840 1502 34020 1536
rect 35520 1536 35526 1558
rect 35582 1536 35700 1620
rect 35520 1502 35700 1536
rect 28800 1440 29038 1500
rect 30542 1440 30660 1502
rect 32222 1440 32340 1502
rect 33902 1440 34020 1502
rect 35582 1440 35700 1502
rect 37200 1592 37380 1620
rect 37200 1536 37206 1592
rect 37262 1536 37380 1592
rect 37200 1500 37380 1536
rect 38880 1592 39060 1620
rect 38880 1536 38886 1592
rect 38942 1536 39060 1592
rect 37200 1440 37438 1500
rect 38880 1500 39060 1536
rect 40560 1592 40740 1620
rect 40560 1536 40566 1592
rect 40622 1536 40740 1592
rect 40560 1502 40740 1536
rect 38702 1440 39060 1500
rect 40622 1440 40740 1502
rect 42240 1592 42420 1620
rect 42240 1536 42246 1592
rect 42302 1536 42420 1592
rect 42240 1502 42420 1536
rect 43920 1592 44100 1620
rect 43920 1536 43926 1592
rect 43982 1536 44100 1592
rect 43920 1502 44100 1536
rect 45600 1592 45780 1620
rect 45600 1536 45606 1592
rect 45662 1536 45780 1592
rect 45600 1502 45780 1536
rect 47280 1592 47460 1620
rect 47280 1536 47286 1592
rect 47342 1536 47460 1592
rect 47280 1502 47460 1536
rect 48960 1592 49140 1620
rect 48960 1536 48966 1592
rect 49022 1536 49140 1592
rect 48960 1502 49140 1536
rect 50640 1592 50820 1620
rect 50640 1536 50646 1592
rect 50702 1536 50820 1592
rect 50640 1502 50820 1536
rect 42240 1440 42358 1502
rect 43920 1440 44038 1502
rect 45600 1440 45718 1502
rect 47280 1440 47398 1502
rect 49022 1440 49140 1502
rect 50702 1440 50820 1502
rect 52320 1592 52500 1620
rect 52320 1536 52326 1592
rect 52382 1536 52500 1592
rect 52320 1502 52500 1536
rect 54000 1592 54180 1620
rect 54000 1536 54006 1592
rect 54062 1536 54180 1592
rect 54000 1502 54180 1536
rect 55680 1592 55860 1620
rect 55680 1536 55686 1592
rect 55742 1536 55860 1592
rect 55680 1502 55860 1536
rect 57360 1592 57540 1620
rect 57360 1536 57366 1592
rect 57422 1536 57540 1592
rect 57360 1502 57540 1536
rect 59040 1592 59220 1620
rect 59040 1536 59046 1592
rect 59102 1536 59220 1592
rect 59040 1502 59220 1536
rect 60720 1592 60900 1620
rect 60720 1536 60726 1592
rect 60782 1536 60900 1592
rect 60720 1502 60900 1536
rect 52320 1440 52438 1502
rect 54000 1440 54118 1502
rect 55680 1440 55798 1502
rect 57422 1440 57540 1502
rect 59102 1440 59220 1502
rect 60782 1440 60900 1502
rect 62400 1592 62580 1620
rect 62400 1536 62406 1592
rect 62462 1536 62580 1592
rect 62400 1502 62580 1536
rect 64080 1592 64260 1620
rect 64080 1536 64086 1592
rect 64142 1536 64260 1592
rect 64080 1502 64260 1536
rect 65760 1592 65940 1620
rect 65760 1536 65766 1592
rect 65822 1536 65940 1592
rect 65760 1502 65940 1536
rect 62400 1440 62518 1502
rect 64142 1440 64260 1502
rect 65822 1440 65940 1502
rect 67440 1592 67620 1620
rect 67440 1536 67446 1592
rect 67502 1536 67620 1592
rect 67440 1502 67620 1536
rect 69120 1592 69300 1620
rect 69120 1536 69126 1592
rect 69182 1536 69300 1592
rect 69120 1502 69300 1536
rect 70800 1592 70980 1620
rect 70800 1536 70806 1592
rect 70862 1536 70980 1592
rect 70800 1502 70980 1536
rect 67440 1440 67558 1502
rect 69120 1440 69238 1502
rect 70862 1440 70980 1502
rect 72480 1592 72660 1620
rect 72480 1536 72486 1592
rect 72542 1536 72660 1592
rect 72480 1502 72660 1536
rect 72480 1440 72598 1502
rect 902 1078 958 1140
rect 1022 1078 1078 1140
rect 1142 1078 2038 1140
rect 2102 1078 3598 1140
rect 3662 1078 5398 1140
rect 5462 1078 6958 1140
rect 7022 1078 8638 1140
rect 8702 1078 10438 1140
rect 10502 1078 11998 1140
rect 12062 1078 13798 1140
rect 13862 1078 15358 1140
rect 15422 1078 17158 1140
rect 17222 1078 18838 1140
rect 18902 1078 20518 1140
rect 20582 1078 22198 1140
rect 22262 1078 23878 1140
rect 23942 1078 25438 1140
rect 25502 1078 27118 1140
rect 27182 1078 29038 1140
rect 29102 1078 30478 1140
rect 30542 1078 32158 1140
rect 32222 1078 33838 1140
rect 33902 1078 35518 1140
rect 35582 1078 37438 1140
rect 37502 1078 38638 1140
rect 38702 1078 40558 1140
rect 40622 1078 42358 1140
rect 42422 1078 44038 1140
rect 44102 1078 45718 1140
rect 45782 1078 47398 1140
rect 47462 1078 48958 1140
rect 49022 1078 50638 1140
rect 50702 1078 52438 1140
rect 52502 1078 54118 1140
rect 54182 1078 55798 1140
rect 55862 1078 57358 1140
rect 57422 1078 59038 1140
rect 59102 1078 60718 1140
rect 60782 1078 62518 1140
rect 62582 1078 64078 1140
rect 64142 1078 65758 1140
rect 65822 1078 67558 1140
rect 67622 1078 69238 1140
rect 69302 1078 70798 1140
rect 70862 1078 72598 1140
rect 72662 1078 74398 1140
rect 74462 1078 74518 1140
rect 74582 1078 74638 1140
rect 840 1022 74700 1078
rect 902 958 958 1022
rect 1022 958 1078 1022
rect 1142 958 74398 1022
rect 74462 958 74518 1022
rect 74582 958 74638 1022
rect 840 902 74700 958
rect 902 840 958 902
rect 1022 840 1078 902
rect 1142 840 74398 902
rect 74462 840 74518 902
rect 74582 840 74638 902
rect 302 478 358 540
rect 422 478 478 540
rect 542 478 32278 540
rect 32342 478 74998 540
rect 75062 478 75118 540
rect 75182 478 75238 540
rect 240 422 75300 478
rect 302 358 358 422
rect 422 358 478 422
rect 542 358 74998 422
rect 75062 358 75118 422
rect 75182 358 75238 422
rect 240 302 75300 358
rect 302 240 358 302
rect 422 240 478 302
rect 542 240 74998 302
rect 75062 240 75118 302
rect 75182 240 75238 302
<< via3 >>
rect 238 37438 302 37502
rect 358 37438 422 37502
rect 478 37438 542 37502
rect 74998 37438 75062 37502
rect 75118 37438 75182 37502
rect 75238 37438 75302 37502
rect 238 37318 302 37382
rect 358 37318 422 37382
rect 478 37318 542 37382
rect 74998 37318 75062 37382
rect 75118 37318 75182 37382
rect 75238 37318 75302 37382
rect 238 37198 302 37262
rect 358 37198 422 37262
rect 478 37198 542 37262
rect 14518 37198 14582 37262
rect 19558 37198 19622 37262
rect 74998 37198 75062 37262
rect 75118 37198 75182 37262
rect 75238 37198 75302 37262
rect 838 36838 902 36902
rect 958 36838 1022 36902
rect 1078 36838 1142 36902
rect 74398 36838 74462 36902
rect 74518 36838 74582 36902
rect 74638 36838 74702 36902
rect 838 36718 902 36782
rect 958 36718 1022 36782
rect 1078 36718 1142 36782
rect 74398 36718 74462 36782
rect 74518 36718 74582 36782
rect 74638 36718 74702 36782
rect 838 36598 902 36662
rect 958 36598 1022 36662
rect 1078 36598 1142 36662
rect 1918 36598 1982 36662
rect 3718 36598 3782 36662
rect 5398 36598 5462 36662
rect 6958 36598 7022 36662
rect 8638 36598 8702 36662
rect 10438 36598 10502 36662
rect 11998 36598 12062 36662
rect 13678 36598 13742 36662
rect 15478 36598 15542 36662
rect 17158 36598 17222 36662
rect 18838 36598 18902 36662
rect 20518 36598 20582 36662
rect 22078 36598 22142 36662
rect 23758 36598 23822 36662
rect 25438 36598 25502 36662
rect 27118 36598 27182 36662
rect 28918 36598 28982 36662
rect 30478 36598 30542 36662
rect 32158 36598 32222 36662
rect 33838 36598 33902 36662
rect 35638 36598 35702 36662
rect 37318 36598 37382 36662
rect 38878 36598 38942 36662
rect 40678 36598 40742 36662
rect 42358 36598 42422 36662
rect 43918 36598 43982 36662
rect 45718 36598 45782 36662
rect 47398 36598 47462 36662
rect 48958 36598 49022 36662
rect 50638 36598 50702 36662
rect 52438 36598 52502 36662
rect 54118 36598 54182 36662
rect 55678 36598 55742 36662
rect 57358 36598 57422 36662
rect 59158 36598 59222 36662
rect 60718 36598 60782 36662
rect 62398 36598 62462 36662
rect 64198 36598 64262 36662
rect 65758 36598 65822 36662
rect 67558 36598 67622 36662
rect 69238 36598 69302 36662
rect 70798 36598 70862 36662
rect 72478 36598 72542 36662
rect 74398 36598 74462 36662
rect 74518 36598 74582 36662
rect 74638 36598 74702 36662
rect 1918 36238 1982 36302
rect 3718 36238 3782 36302
rect 5398 36238 5462 36302
rect 6958 36238 7022 36302
rect 8638 36238 8702 36302
rect 10438 36238 10502 36302
rect 11998 36238 12062 36302
rect 13678 36238 13742 36302
rect 15478 36238 15542 36302
rect 17158 36238 17222 36302
rect 18838 36238 18902 36302
rect 20518 36238 20582 36302
rect 22078 36238 22142 36302
rect 23758 36238 23822 36302
rect 25438 36238 25502 36302
rect 27118 36238 27182 36302
rect 14398 36118 14462 36182
rect 20398 36180 20406 36182
rect 20406 36180 20462 36182
rect 20398 36118 20462 36180
rect 28918 36238 28982 36302
rect 30478 36238 30542 36302
rect 32158 36238 32222 36302
rect 33838 36238 33902 36302
rect 35638 36238 35702 36302
rect 37318 36238 37382 36302
rect 38878 36238 38942 36302
rect 40678 36238 40742 36302
rect 42358 36238 42422 36302
rect 43918 36238 43982 36302
rect 45718 36238 45782 36302
rect 47398 36238 47462 36302
rect 48958 36238 49022 36302
rect 50638 36238 50702 36302
rect 52438 36238 52502 36302
rect 54118 36238 54182 36302
rect 55678 36238 55742 36302
rect 57358 36238 57422 36302
rect 59158 36238 59222 36302
rect 60718 36238 60782 36302
rect 62398 36238 62462 36302
rect 64198 36238 64262 36302
rect 65758 36238 65822 36302
rect 67558 36238 67622 36302
rect 69238 36238 69302 36302
rect 70798 36238 70862 36302
rect 72478 36238 72542 36302
rect 1078 35518 1142 35582
rect 74398 35398 74462 35462
rect 14518 35278 14582 35342
rect 19558 35278 19622 35342
rect 15238 35158 15302 35222
rect 19558 35158 19622 35222
rect 19558 34918 19622 34982
rect 19678 34798 19742 34862
rect 1078 33838 1142 33902
rect 14398 33718 14462 33782
rect 14998 33598 15062 33662
rect 20398 33718 20462 33782
rect 74398 33718 74462 33782
rect 19558 33598 19622 33662
rect 19558 33358 19622 33422
rect 18478 33238 18542 33302
rect 1078 32038 1142 32102
rect 15238 32158 15302 32222
rect 15118 32038 15182 32102
rect 19678 32158 19742 32222
rect 19558 32038 19622 32102
rect 74398 32038 74462 32102
rect 19558 31798 19622 31862
rect 19678 31678 19742 31742
rect 14998 30718 15062 30782
rect 1078 30358 1142 30422
rect 18478 30358 18542 30422
rect 74398 30478 74462 30542
rect 19558 30238 19622 30302
rect 15118 29278 15182 29342
rect 19678 29158 19742 29222
rect 1078 28678 1142 28742
rect 74398 28798 74462 28862
rect 18478 28678 18542 28742
rect 19558 27598 19622 27662
rect 19558 27238 19622 27302
rect 1078 27118 1142 27182
rect 74398 27118 74462 27182
rect 15118 25918 15182 25982
rect 18478 25798 18542 25862
rect 19438 25678 19502 25742
rect 1078 25438 1142 25502
rect 74398 25318 74462 25382
rect 14398 24358 14462 24422
rect 19558 24478 19622 24542
rect 19678 24358 19742 24422
rect 1078 23758 1142 23822
rect 74398 23638 74462 23702
rect 15118 23038 15182 23102
rect 19438 22918 19502 22982
rect 15358 22798 15422 22862
rect 19438 22678 19502 22742
rect 1078 21958 1142 22022
rect 74398 21958 74462 22022
rect 14398 21478 14462 21542
rect 19678 21478 19742 21542
rect 19558 21238 19622 21302
rect 1078 20278 1142 20342
rect 74398 20398 74462 20462
rect 14398 19798 14462 19862
rect 15358 19918 15422 19982
rect 19438 19918 19502 19982
rect 1078 18598 1142 18662
rect 74398 18718 74462 18782
rect 19558 18358 19622 18422
rect 14398 17518 14462 17582
rect 14398 17398 14462 17462
rect 1078 17038 1142 17102
rect 74398 17038 74462 17102
rect 14398 16798 14462 16862
rect 14398 16678 14462 16742
rect 12958 16558 13022 16622
rect 18478 16558 18542 16622
rect 14398 15838 14462 15902
rect 12838 15718 12902 15782
rect 1078 15358 1142 15422
rect 74398 15238 74462 15302
rect 12958 14998 13022 15062
rect 19678 15118 19742 15182
rect 12958 14878 13022 14942
rect 12838 14158 12902 14222
rect 12838 14038 12902 14102
rect 14398 14038 14462 14102
rect 1078 13678 1142 13742
rect 14398 13678 14462 13742
rect 18478 13678 18542 13742
rect 19558 13558 19622 13622
rect 74398 13558 74462 13622
rect 12958 13318 13022 13382
rect 12958 13198 13022 13262
rect 12838 12478 12902 12542
rect 12838 12358 12902 12422
rect 12478 12118 12542 12182
rect 14398 12118 14462 12182
rect 19678 12238 19742 12302
rect 20278 12118 20342 12182
rect 1078 11878 1142 11942
rect 74398 11878 74462 11942
rect 12958 11638 13022 11702
rect 14398 11638 14462 11702
rect 12358 10978 12391 10982
rect 12391 10978 12422 10982
rect 12358 10918 12422 10978
rect 12838 10798 12902 10862
rect 19558 10678 19622 10742
rect 15718 10558 15782 10622
rect 18358 10558 18422 10622
rect 24478 10558 24542 10622
rect 24598 10438 24662 10502
rect 26158 10558 26222 10622
rect 27718 10558 27782 10622
rect 29278 10438 29342 10502
rect 32398 10558 32462 10622
rect 31078 10438 31142 10502
rect 33958 10558 34022 10622
rect 35518 10438 35582 10502
rect 38638 10558 38702 10622
rect 37318 10438 37382 10502
rect 40078 10558 40142 10622
rect 41638 10558 41702 10622
rect 43078 10438 43142 10502
rect 1078 10198 1142 10262
rect 74398 10198 74462 10262
rect 20278 9718 20342 9782
rect 15718 9598 15782 9662
rect 18358 9598 18422 9662
rect 20278 9598 20342 9662
rect 24958 9598 25022 9662
rect 26518 9598 26582 9662
rect 28078 9598 28142 9662
rect 29638 9598 29702 9662
rect 31198 9598 31262 9662
rect 32758 9598 32822 9662
rect 34318 9598 34382 9662
rect 35758 9598 35822 9662
rect 37438 9598 37502 9662
rect 38998 9598 39062 9662
rect 40558 9598 40622 9662
rect 42118 9598 42182 9662
rect 43678 9598 43742 9662
rect 17518 9478 17582 9542
rect 24478 9358 24542 9422
rect 24598 9358 24662 9422
rect 24838 9358 24902 9422
rect 26158 9358 26222 9422
rect 27718 9358 27782 9422
rect 29278 9358 29342 9422
rect 31078 9478 31142 9542
rect 32398 9358 32462 9422
rect 33958 9358 34022 9422
rect 35518 9358 35582 9422
rect 37318 9478 37382 9542
rect 43318 9478 43382 9542
rect 46318 9598 46382 9662
rect 47878 9598 47942 9662
rect 49438 9598 49502 9662
rect 38638 9358 38702 9422
rect 40078 9358 40142 9422
rect 41518 9358 41582 9422
rect 41638 9358 41702 9422
rect 41878 9358 41942 9422
rect 43078 9358 43142 9422
rect 43198 9358 43262 9422
rect 26278 9252 26334 9302
rect 26334 9252 26342 9302
rect 26278 9238 26342 9252
rect 27838 9252 27890 9302
rect 27890 9252 27902 9302
rect 27838 9238 27902 9252
rect 29398 9252 29446 9302
rect 29446 9252 29462 9302
rect 29398 9238 29462 9252
rect 30958 9252 31002 9302
rect 31002 9252 31022 9302
rect 30958 9238 31022 9252
rect 32518 9252 32558 9302
rect 32558 9252 32582 9302
rect 32518 9238 32582 9252
rect 34078 9252 34114 9302
rect 34114 9252 34142 9302
rect 34078 9238 34142 9252
rect 35638 9252 35670 9302
rect 35670 9252 35702 9302
rect 35638 9238 35702 9252
rect 37198 9252 37226 9302
rect 37226 9252 37262 9302
rect 37198 9238 37262 9252
rect 38758 9252 38782 9302
rect 38782 9252 38822 9302
rect 38758 9238 38822 9252
rect 43438 9358 43502 9422
rect 44158 9358 44222 9422
rect 44758 9358 44822 9422
rect 40318 9252 40338 9302
rect 40338 9252 40382 9302
rect 40318 9238 40382 9252
rect 44998 9358 45062 9422
rect 46318 9358 46382 9422
rect 47878 9358 47942 9422
rect 46558 9252 46562 9302
rect 46562 9252 46622 9302
rect 46558 9238 46622 9252
rect 49438 9358 49502 9422
rect 48118 9238 48182 9302
rect 74998 9238 75062 9302
rect 41518 8998 41582 9062
rect 43198 8998 43262 9062
rect 43318 8998 43382 9062
rect 44758 8998 44822 9062
rect 20278 8758 20342 8822
rect 1078 8518 1142 8582
rect 74398 8638 74462 8702
rect 24958 8398 25022 8462
rect 26518 8398 26582 8462
rect 28078 8398 28142 8462
rect 29638 8398 29702 8462
rect 31198 8398 31262 8462
rect 32758 8398 32822 8462
rect 34318 8398 34382 8462
rect 35758 8398 35822 8462
rect 37438 8398 37502 8462
rect 38998 8398 39062 8462
rect 40558 8398 40622 8462
rect 42118 8398 42182 8462
rect 43678 8398 43742 8462
rect 17518 7918 17582 7982
rect 1078 6958 1142 7022
rect 44158 7078 44222 7142
rect 74398 6958 74462 7022
rect 478 6238 542 6302
rect 2398 6238 2462 6302
rect 5998 5758 6062 5822
rect 1078 5278 1142 5342
rect 35038 5158 35102 5222
rect 74398 5158 74462 5222
rect 2398 4678 2462 4742
rect 1078 3598 1142 3662
rect 74398 3478 74462 3542
rect 35038 3238 35102 3302
rect 35518 3118 35582 3182
rect 15238 2518 15302 2582
rect 16918 2518 16982 2582
rect 18238 2518 18302 2582
rect 19678 2518 19742 2582
rect 21358 2518 21422 2582
rect 22798 2518 22862 2582
rect 24358 2518 24422 2582
rect 25798 2518 25862 2582
rect 27238 2518 27302 2582
rect 28798 2518 28862 2582
rect 30238 2518 30302 2582
rect 31678 2518 31742 2582
rect 33118 2518 33182 2582
rect 34558 2518 34622 2582
rect 35998 2518 36062 2582
rect 37678 2518 37742 2582
rect 39118 2518 39182 2582
rect 32278 2278 32342 2342
rect 1918 1798 1982 1862
rect 74398 1798 74462 1862
rect 1918 1592 1982 1622
rect 1918 1558 1926 1592
rect 1926 1558 1982 1592
rect 2038 1438 2102 1502
rect 3598 1438 3662 1502
rect 5398 1438 5462 1502
rect 6958 1438 7022 1502
rect 8638 1438 8702 1502
rect 10438 1438 10502 1502
rect 11998 1438 12062 1502
rect 13798 1438 13862 1502
rect 15358 1438 15422 1502
rect 17158 1438 17222 1502
rect 18838 1438 18902 1502
rect 20518 1438 20582 1502
rect 22198 1438 22262 1502
rect 23878 1438 23942 1502
rect 25438 1438 25502 1502
rect 27118 1438 27182 1502
rect 35518 1592 35582 1622
rect 35518 1558 35526 1592
rect 35526 1558 35582 1592
rect 29038 1438 29102 1502
rect 30478 1438 30542 1502
rect 32158 1438 32222 1502
rect 33838 1438 33902 1502
rect 35518 1438 35582 1502
rect 37438 1438 37502 1502
rect 38638 1438 38702 1502
rect 40558 1438 40622 1502
rect 42358 1438 42422 1502
rect 44038 1438 44102 1502
rect 45718 1438 45782 1502
rect 47398 1438 47462 1502
rect 48958 1438 49022 1502
rect 50638 1438 50702 1502
rect 52438 1438 52502 1502
rect 54118 1438 54182 1502
rect 55798 1438 55862 1502
rect 57358 1438 57422 1502
rect 59038 1438 59102 1502
rect 60718 1438 60782 1502
rect 62518 1438 62582 1502
rect 64078 1438 64142 1502
rect 65758 1438 65822 1502
rect 67558 1438 67622 1502
rect 69238 1438 69302 1502
rect 70798 1438 70862 1502
rect 72598 1438 72662 1502
rect 838 1078 902 1142
rect 958 1078 1022 1142
rect 1078 1078 1142 1142
rect 2038 1078 2102 1142
rect 3598 1078 3662 1142
rect 5398 1078 5462 1142
rect 6958 1078 7022 1142
rect 8638 1078 8702 1142
rect 10438 1078 10502 1142
rect 11998 1078 12062 1142
rect 13798 1078 13862 1142
rect 15358 1078 15422 1142
rect 17158 1078 17222 1142
rect 18838 1078 18902 1142
rect 20518 1078 20582 1142
rect 22198 1078 22262 1142
rect 23878 1078 23942 1142
rect 25438 1078 25502 1142
rect 27118 1078 27182 1142
rect 29038 1078 29102 1142
rect 30478 1078 30542 1142
rect 32158 1078 32222 1142
rect 33838 1078 33902 1142
rect 35518 1078 35582 1142
rect 37438 1078 37502 1142
rect 38638 1078 38702 1142
rect 40558 1078 40622 1142
rect 42358 1078 42422 1142
rect 44038 1078 44102 1142
rect 45718 1078 45782 1142
rect 47398 1078 47462 1142
rect 48958 1078 49022 1142
rect 50638 1078 50702 1142
rect 52438 1078 52502 1142
rect 54118 1078 54182 1142
rect 55798 1078 55862 1142
rect 57358 1078 57422 1142
rect 59038 1078 59102 1142
rect 60718 1078 60782 1142
rect 62518 1078 62582 1142
rect 64078 1078 64142 1142
rect 65758 1078 65822 1142
rect 67558 1078 67622 1142
rect 69238 1078 69302 1142
rect 70798 1078 70862 1142
rect 72598 1078 72662 1142
rect 74398 1078 74462 1142
rect 74518 1078 74582 1142
rect 74638 1078 74702 1142
rect 838 958 902 1022
rect 958 958 1022 1022
rect 1078 958 1142 1022
rect 74398 958 74462 1022
rect 74518 958 74582 1022
rect 74638 958 74702 1022
rect 838 838 902 902
rect 958 838 1022 902
rect 1078 838 1142 902
rect 74398 838 74462 902
rect 74518 838 74582 902
rect 74638 838 74702 902
rect 238 478 302 542
rect 358 478 422 542
rect 478 478 542 542
rect 32278 478 32342 542
rect 74998 478 75062 542
rect 75118 478 75182 542
rect 75238 478 75302 542
rect 238 358 302 422
rect 358 358 422 422
rect 478 358 542 422
rect 74998 358 75062 422
rect 75118 358 75182 422
rect 75238 358 75302 422
rect 238 238 302 302
rect 358 238 422 302
rect 478 238 542 302
rect 74998 238 75062 302
rect 75118 238 75182 302
rect 75238 238 75302 302
<< metal4 >>
rect 302 37438 358 37500
rect 422 37438 478 37500
rect 75062 37438 75118 37500
rect 75182 37438 75238 37500
rect 240 37382 540 37438
rect 75000 37382 75300 37438
rect 302 37318 358 37382
rect 422 37318 478 37382
rect 75062 37318 75118 37382
rect 75182 37318 75238 37382
rect 240 37262 540 37318
rect 75000 37262 75300 37318
rect 302 37198 358 37262
rect 422 37198 478 37262
rect 75062 37198 75118 37262
rect 75182 37198 75238 37262
rect 240 6302 540 37198
rect 902 36838 958 36900
rect 1022 36838 1078 36900
rect 840 36782 1140 36838
rect 902 36718 958 36782
rect 1022 36718 1078 36782
rect 840 36662 1140 36718
rect 902 36598 958 36662
rect 1022 36598 1078 36662
rect 840 35582 1140 36598
rect 1920 36302 1980 36598
rect 3720 36302 3780 36598
rect 5400 36302 5460 36598
rect 6960 36302 7020 36598
rect 8640 36302 8700 36598
rect 10440 36302 10500 36598
rect 12000 36302 12060 36598
rect 13680 36302 13740 36598
rect 840 35518 1078 35582
rect 840 33902 1140 35518
rect 840 33838 1078 33902
rect 840 32102 1140 33838
rect 14400 33782 14460 36118
rect 14520 35342 14580 37198
rect 15480 36302 15540 36598
rect 17160 36302 17220 36598
rect 18840 36302 18900 36598
rect 19560 35342 19620 37198
rect 74462 36838 74518 36900
rect 74582 36838 74638 36900
rect 74400 36782 74700 36838
rect 74462 36718 74518 36782
rect 74582 36718 74638 36782
rect 74400 36662 74700 36718
rect 74462 36598 74518 36662
rect 74582 36598 74638 36662
rect 20520 36302 20580 36598
rect 22080 36302 22140 36598
rect 23760 36302 23820 36598
rect 25440 36302 25500 36598
rect 27120 36302 27180 36598
rect 28920 36302 28980 36598
rect 30480 36302 30540 36598
rect 32160 36302 32220 36598
rect 33840 36302 33900 36598
rect 35640 36302 35700 36598
rect 37320 36302 37380 36598
rect 38880 36302 38940 36598
rect 40680 36302 40740 36598
rect 42360 36302 42420 36598
rect 43920 36302 43980 36598
rect 45720 36302 45780 36598
rect 47400 36302 47460 36598
rect 48960 36302 49020 36598
rect 50640 36302 50700 36598
rect 52440 36302 52500 36598
rect 54120 36302 54180 36598
rect 55680 36302 55740 36598
rect 57360 36302 57420 36598
rect 59160 36302 59220 36598
rect 60720 36302 60780 36598
rect 62400 36302 62460 36598
rect 64200 36302 64260 36598
rect 65760 36302 65820 36598
rect 67560 36302 67620 36598
rect 69240 36302 69300 36598
rect 70800 36302 70860 36598
rect 72480 36302 72540 36598
rect 840 32038 1078 32102
rect 840 30422 1140 32038
rect 15000 30782 15060 33598
rect 15240 32222 15300 35158
rect 19560 34982 19620 35158
rect 19560 33422 19620 33598
rect 840 30358 1078 30422
rect 840 28742 1140 30358
rect 15120 29342 15180 32038
rect 18480 30422 18540 33238
rect 19680 32222 19740 34798
rect 20400 33782 20460 36118
rect 74400 35462 74700 36598
rect 74462 35398 74700 35462
rect 74400 33782 74700 35398
rect 74462 33718 74700 33782
rect 74400 32102 74700 33718
rect 74462 32038 74700 32102
rect 19560 31862 19620 32038
rect 840 28678 1078 28742
rect 840 27182 1140 28678
rect 840 27118 1078 27182
rect 840 25502 1140 27118
rect 840 25438 1078 25502
rect 840 23822 1140 25438
rect 840 23758 1078 23822
rect 840 22022 1140 23758
rect 840 21958 1078 22022
rect 840 20342 1140 21958
rect 14400 21542 14460 24358
rect 15120 23102 15180 25918
rect 18480 25862 18540 28678
rect 19560 27662 19620 30238
rect 19680 29222 19740 31678
rect 74400 30542 74700 32038
rect 74462 30478 74700 30542
rect 74400 28862 74700 30478
rect 74462 28798 74700 28862
rect 19440 22982 19500 25678
rect 19560 24542 19620 27238
rect 74400 27182 74700 28798
rect 74462 27118 74700 27182
rect 74400 25382 74700 27118
rect 74462 25318 74700 25382
rect 840 20278 1078 20342
rect 840 18662 1140 20278
rect 15360 19982 15420 22798
rect 19440 19982 19500 22678
rect 19680 21542 19740 24358
rect 74400 23702 74700 25318
rect 74462 23638 74700 23702
rect 74400 22022 74700 23638
rect 74462 21958 74700 22022
rect 840 18598 1078 18662
rect 840 17102 1140 18598
rect 14400 17582 14460 19798
rect 19560 18422 19620 21238
rect 74400 20462 74700 21958
rect 74462 20398 74700 20462
rect 74400 18782 74700 20398
rect 74462 18718 74700 18782
rect 840 17038 1078 17102
rect 840 15422 1140 17038
rect 14400 16862 14460 17398
rect 74400 17102 74700 18718
rect 74462 17038 74700 17102
rect 840 15358 1078 15422
rect 840 13742 1140 15358
rect 12840 14222 12900 15718
rect 12960 15062 13020 16558
rect 14400 15902 14460 16678
rect 840 13678 1078 13742
rect 840 11942 1140 13678
rect 12840 12542 12900 14038
rect 12960 13382 13020 14878
rect 14400 13742 14460 14038
rect 18480 13742 18540 16558
rect 74400 15302 74700 17038
rect 74462 15238 74700 15302
rect 840 11878 1078 11942
rect 840 10262 1140 11878
rect 840 10198 1078 10262
rect 840 8582 1140 10198
rect 840 8518 1078 8582
rect 840 7022 1140 8518
rect 840 6958 1078 7022
rect 240 6238 478 6302
rect 240 542 540 6238
rect 840 5342 1140 6958
rect 840 5278 1078 5342
rect 840 3662 1140 5278
rect 2400 4742 2460 6238
rect 840 3598 1078 3662
rect 840 1142 1140 3598
rect 1920 1622 1980 1798
rect 2040 1142 2100 1438
rect 3600 1142 3660 1438
rect 5400 1142 5460 1438
rect 902 1078 958 1142
rect 1022 1078 1078 1142
rect 840 1022 1140 1078
rect 902 958 958 1022
rect 1022 958 1078 1022
rect 840 902 1140 958
rect 902 840 958 902
rect 1022 840 1078 902
rect 302 478 358 542
rect 422 478 478 542
rect 240 422 540 478
rect 302 358 358 422
rect 422 358 478 422
rect 240 302 540 358
rect 302 240 358 302
rect 422 240 478 302
rect 6000 0 6060 5758
rect 6960 1142 7020 1438
rect 8640 1142 8700 1438
rect 10440 1142 10500 1438
rect 12000 1142 12060 1438
rect 12360 0 12420 10918
rect 12480 0 12540 12118
rect 12840 10862 12900 12358
rect 12960 11702 13020 13198
rect 14400 11702 14460 12118
rect 19560 10742 19620 13558
rect 19680 12302 19740 15118
rect 74400 13622 74700 15238
rect 74462 13558 74700 13622
rect 15720 9662 15780 10558
rect 18360 9662 18420 10558
rect 20280 9782 20340 12118
rect 74400 11942 74700 13558
rect 74462 11878 74700 11942
rect 17520 7982 17580 9478
rect 20280 8822 20340 9598
rect 24480 9422 24540 10558
rect 24600 9422 24660 10438
rect 13800 1142 13860 1438
rect 15240 0 15300 2518
rect 15360 1142 15420 1438
rect 16920 0 16980 2518
rect 17160 1142 17220 1438
rect 18240 0 18300 2518
rect 18840 1142 18900 1438
rect 19680 0 19740 2518
rect 20520 1142 20580 1438
rect 21360 0 21420 2518
rect 22200 1142 22260 1438
rect 22800 0 22860 2518
rect 23880 1142 23940 1438
rect 24360 0 24420 2518
rect 24840 0 24900 9358
rect 24960 8462 25020 9598
rect 26160 9422 26220 10558
rect 25440 1142 25500 1438
rect 25800 0 25860 2518
rect 26280 0 26340 9238
rect 26520 8462 26580 9598
rect 27720 9422 27780 10558
rect 27120 1142 27180 1438
rect 27240 0 27300 2518
rect 27840 0 27900 9238
rect 28080 8462 28140 9598
rect 29280 9422 29340 10438
rect 28800 0 28860 2518
rect 29040 1142 29100 1438
rect 29400 0 29460 9238
rect 29640 8462 29700 9598
rect 31080 9542 31140 10438
rect 30240 0 30300 2518
rect 30480 1142 30540 1438
rect 30960 0 31020 9238
rect 31200 8462 31260 9598
rect 32400 9422 32460 10558
rect 31680 0 31740 2518
rect 32160 1142 32220 1438
rect 32280 542 32340 2278
rect 32520 0 32580 9238
rect 32760 8462 32820 9598
rect 33960 9422 34020 10558
rect 33120 0 33180 2518
rect 33840 1142 33900 1438
rect 34080 0 34140 9238
rect 34320 8462 34380 9598
rect 35520 9422 35580 10438
rect 35040 3302 35100 5158
rect 34560 0 34620 2518
rect 35520 1622 35580 3118
rect 35520 1142 35580 1438
rect 35640 0 35700 9238
rect 35760 8462 35820 9598
rect 37320 9542 37380 10438
rect 36000 0 36060 2518
rect 37200 0 37260 9238
rect 37440 8462 37500 9598
rect 38640 9422 38700 10558
rect 37440 1142 37500 1438
rect 37680 0 37740 2518
rect 38640 1142 38700 1438
rect 38760 0 38820 9238
rect 39000 8462 39060 9598
rect 40080 9422 40140 10558
rect 39120 0 39180 2518
rect 40320 0 40380 9238
rect 40560 8462 40620 9598
rect 41640 9422 41700 10558
rect 41520 9062 41580 9358
rect 40560 1142 40620 1438
rect 41880 0 41940 9358
rect 42120 8462 42180 9598
rect 43080 9422 43140 10438
rect 74400 10262 74700 11878
rect 74462 10198 74700 10262
rect 43200 9062 43260 9358
rect 43320 9062 43380 9478
rect 42360 1142 42420 1438
rect 43440 0 43500 9358
rect 43680 8462 43740 9598
rect 46320 9422 46380 9598
rect 47880 9422 47940 9598
rect 49440 9422 49500 9598
rect 44160 7142 44220 9358
rect 44760 9062 44820 9358
rect 44040 1142 44100 1438
rect 45000 0 45060 9358
rect 45720 1142 45780 1438
rect 46560 0 46620 9238
rect 47400 1142 47460 1438
rect 48120 0 48180 9238
rect 74400 8702 74700 10198
rect 75000 9302 75300 37198
rect 75062 9238 75300 9302
rect 74462 8638 74700 8702
rect 74400 7022 74700 8638
rect 74462 6958 74700 7022
rect 74400 5222 74700 6958
rect 74462 5158 74700 5222
rect 74400 3542 74700 5158
rect 74462 3478 74700 3542
rect 74400 1862 74700 3478
rect 74462 1798 74700 1862
rect 48960 1142 49020 1438
rect 50640 1142 50700 1438
rect 52440 1142 52500 1438
rect 54120 1142 54180 1438
rect 55800 1142 55860 1438
rect 57360 1142 57420 1438
rect 59040 1142 59100 1438
rect 60720 1142 60780 1438
rect 62520 1142 62580 1438
rect 64080 1142 64140 1438
rect 65760 1142 65820 1438
rect 67560 1142 67620 1438
rect 69240 1142 69300 1438
rect 70800 1142 70860 1438
rect 72600 1142 72660 1438
rect 74400 1142 74700 1798
rect 74462 1078 74518 1142
rect 74582 1078 74638 1142
rect 74400 1022 74700 1078
rect 74462 958 74518 1022
rect 74582 958 74638 1022
rect 74400 902 74700 958
rect 74462 840 74518 902
rect 74582 840 74638 902
rect 75000 542 75300 9238
rect 75062 478 75118 542
rect 75182 478 75238 542
rect 75000 422 75300 478
rect 75062 358 75118 422
rect 75182 358 75238 422
rect 75000 302 75300 358
rect 75062 240 75118 302
rect 75182 240 75238 302
use contact_32  contact_32_0
timestamp 1643671299
transform 1 0 75000 0 1 9240
box 0 0 1 1
use contact_32  contact_32_1
timestamp 1643671299
transform 1 0 49440 0 1 9360
box 0 0 1 1
use contact_32  contact_32_2
timestamp 1643671299
transform 1 0 49440 0 1 9600
box 0 0 1 1
use contact_32  contact_32_3
timestamp 1643671299
transform 1 0 47880 0 1 9600
box 0 0 1 1
use contact_32  contact_32_4
timestamp 1643671299
transform 1 0 47880 0 1 9360
box 0 0 1 1
use contact_32  contact_32_5
timestamp 1643671299
transform 1 0 46320 0 1 9360
box 0 0 1 1
use contact_32  contact_32_6
timestamp 1643671299
transform 1 0 46320 0 1 9600
box 0 0 1 1
use contact_32  contact_32_7
timestamp 1643671299
transform 1 0 44160 0 1 9360
box 0 0 1 1
use contact_32  contact_32_8
timestamp 1643671299
transform 1 0 44160 0 1 7080
box 0 0 1 1
use contact_32  contact_32_9
timestamp 1643671299
transform 1 0 44760 0 1 9360
box 0 0 1 1
use contact_32  contact_32_10
timestamp 1643671299
transform 1 0 44760 0 1 9000
box 0 0 1 1
use contact_32  contact_32_11
timestamp 1643671299
transform 1 0 43320 0 1 9000
box 0 0 1 1
use contact_32  contact_32_12
timestamp 1643671299
transform 1 0 43320 0 1 9480
box 0 0 1 1
use contact_32  contact_32_13
timestamp 1643671299
transform 1 0 43080 0 1 10440
box 0 0 1 1
use contact_32  contact_32_14
timestamp 1643671299
transform 1 0 43080 0 1 9360
box 0 0 1 1
use contact_32  contact_32_15
timestamp 1643671299
transform 1 0 43200 0 1 9360
box 0 0 1 1
use contact_32  contact_32_16
timestamp 1643671299
transform 1 0 43200 0 1 9000
box 0 0 1 1
use contact_32  contact_32_17
timestamp 1643671299
transform 1 0 41520 0 1 9000
box 0 0 1 1
use contact_32  contact_32_18
timestamp 1643671299
transform 1 0 41520 0 1 9360
box 0 0 1 1
use contact_32  contact_32_19
timestamp 1643671299
transform 1 0 41640 0 1 10560
box 0 0 1 1
use contact_32  contact_32_20
timestamp 1643671299
transform 1 0 41640 0 1 9360
box 0 0 1 1
use contact_32  contact_32_21
timestamp 1643671299
transform 1 0 40080 0 1 10560
box 0 0 1 1
use contact_32  contact_32_22
timestamp 1643671299
transform 1 0 40080 0 1 9360
box 0 0 1 1
use contact_32  contact_32_23
timestamp 1643671299
transform 1 0 38640 0 1 10560
box 0 0 1 1
use contact_32  contact_32_24
timestamp 1643671299
transform 1 0 38640 0 1 9360
box 0 0 1 1
use contact_32  contact_32_25
timestamp 1643671299
transform 1 0 37320 0 1 10440
box 0 0 1 1
use contact_32  contact_32_26
timestamp 1643671299
transform 1 0 37320 0 1 9480
box 0 0 1 1
use contact_32  contact_32_27
timestamp 1643671299
transform 1 0 35520 0 1 10440
box 0 0 1 1
use contact_32  contact_32_28
timestamp 1643671299
transform 1 0 35520 0 1 9360
box 0 0 1 1
use contact_32  contact_32_29
timestamp 1643671299
transform 1 0 33960 0 1 10560
box 0 0 1 1
use contact_32  contact_32_30
timestamp 1643671299
transform 1 0 33960 0 1 9360
box 0 0 1 1
use contact_32  contact_32_31
timestamp 1643671299
transform 1 0 32400 0 1 10560
box 0 0 1 1
use contact_32  contact_32_32
timestamp 1643671299
transform 1 0 32400 0 1 9360
box 0 0 1 1
use contact_32  contact_32_33
timestamp 1643671299
transform 1 0 32280 0 1 480
box 0 0 1 1
use contact_32  contact_32_34
timestamp 1643671299
transform 1 0 32280 0 1 2280
box 0 0 1 1
use contact_32  contact_32_35
timestamp 1643671299
transform 1 0 31080 0 1 10440
box 0 0 1 1
use contact_32  contact_32_36
timestamp 1643671299
transform 1 0 31080 0 1 9480
box 0 0 1 1
use contact_32  contact_32_37
timestamp 1643671299
transform 1 0 29280 0 1 10440
box 0 0 1 1
use contact_32  contact_32_38
timestamp 1643671299
transform 1 0 29280 0 1 9360
box 0 0 1 1
use contact_32  contact_32_39
timestamp 1643671299
transform 1 0 27720 0 1 10560
box 0 0 1 1
use contact_32  contact_32_40
timestamp 1643671299
transform 1 0 27720 0 1 9360
box 0 0 1 1
use contact_32  contact_32_41
timestamp 1643671299
transform 1 0 26160 0 1 10560
box 0 0 1 1
use contact_32  contact_32_42
timestamp 1643671299
transform 1 0 26160 0 1 9360
box 0 0 1 1
use contact_32  contact_32_43
timestamp 1643671299
transform 1 0 24480 0 1 10560
box 0 0 1 1
use contact_32  contact_32_44
timestamp 1643671299
transform 1 0 24480 0 1 9360
box 0 0 1 1
use contact_32  contact_32_45
timestamp 1643671299
transform 1 0 24600 0 1 9360
box 0 0 1 1
use contact_32  contact_32_46
timestamp 1643671299
transform 1 0 24600 0 1 10440
box 0 0 1 1
use contact_32  contact_32_47
timestamp 1643671299
transform 1 0 19560 0 1 13560
box 0 0 1 1
use contact_32  contact_32_48
timestamp 1643671299
transform 1 0 19560 0 1 10680
box 0 0 1 1
use contact_32  contact_32_49
timestamp 1643671299
transform 1 0 19560 0 1 37200
box 0 0 1 1
use contact_32  contact_32_50
timestamp 1643671299
transform 1 0 19560 0 1 35280
box 0 0 1 1
use contact_32  contact_32_51
timestamp 1643671299
transform 1 0 19440 0 1 22920
box 0 0 1 1
use contact_32  contact_32_52
timestamp 1643671299
transform 1 0 19440 0 1 25680
box 0 0 1 1
use contact_32  contact_32_53
timestamp 1643671299
transform 1 0 19560 0 1 32040
box 0 0 1 1
use contact_32  contact_32_54
timestamp 1643671299
transform 1 0 19560 0 1 31800
box 0 0 1 1
use contact_32  contact_32_55
timestamp 1643671299
transform 1 0 19680 0 1 29160
box 0 0 1 1
use contact_32  contact_32_56
timestamp 1643671299
transform 1 0 19680 0 1 31680
box 0 0 1 1
use contact_32  contact_32_57
timestamp 1643671299
transform 1 0 19440 0 1 19920
box 0 0 1 1
use contact_32  contact_32_58
timestamp 1643671299
transform 1 0 19440 0 1 22680
box 0 0 1 1
use contact_32  contact_32_59
timestamp 1643671299
transform 1 0 18480 0 1 13680
box 0 0 1 1
use contact_32  contact_32_60
timestamp 1643671299
transform 1 0 18480 0 1 16560
box 0 0 1 1
use contact_32  contact_32_61
timestamp 1643671299
transform 1 0 19680 0 1 32160
box 0 0 1 1
use contact_32  contact_32_62
timestamp 1643671299
transform 1 0 19680 0 1 34800
box 0 0 1 1
use contact_32  contact_32_63
timestamp 1643671299
transform 1 0 19560 0 1 35160
box 0 0 1 1
use contact_32  contact_32_64
timestamp 1643671299
transform 1 0 19560 0 1 34920
box 0 0 1 1
use contact_32  contact_32_65
timestamp 1643671299
transform 1 0 18480 0 1 25800
box 0 0 1 1
use contact_32  contact_32_66
timestamp 1643671299
transform 1 0 18480 0 1 28680
box 0 0 1 1
use contact_32  contact_32_67
timestamp 1643671299
transform 1 0 18360 0 1 10560
box 0 0 1 1
use contact_32  contact_32_68
timestamp 1643671299
transform 1 0 18360 0 1 9600
box 0 0 1 1
use contact_32  contact_32_69
timestamp 1643671299
transform 1 0 17520 0 1 9480
box 0 0 1 1
use contact_32  contact_32_70
timestamp 1643671299
transform 1 0 17520 0 1 7920
box 0 0 1 1
use contact_32  contact_32_71
timestamp 1643671299
transform 1 0 15240 0 1 35160
box 0 0 1 1
use contact_32  contact_32_72
timestamp 1643671299
transform 1 0 15240 0 1 32160
box 0 0 1 1
use contact_32  contact_32_73
timestamp 1643671299
transform 1 0 15720 0 1 9600
box 0 0 1 1
use contact_32  contact_32_74
timestamp 1643671299
transform 1 0 15720 0 1 10560
box 0 0 1 1
use contact_32  contact_32_75
timestamp 1643671299
transform 1 0 15360 0 1 19920
box 0 0 1 1
use contact_32  contact_32_76
timestamp 1643671299
transform 1 0 15360 0 1 22800
box 0 0 1 1
use contact_32  contact_32_77
timestamp 1643671299
transform 1 0 15120 0 1 25920
box 0 0 1 1
use contact_32  contact_32_78
timestamp 1643671299
transform 1 0 15120 0 1 23040
box 0 0 1 1
use contact_32  contact_32_79
timestamp 1643671299
transform 1 0 15120 0 1 32040
box 0 0 1 1
use contact_32  contact_32_80
timestamp 1643671299
transform 1 0 15120 0 1 29280
box 0 0 1 1
use contact_32  contact_32_81
timestamp 1643671299
transform 1 0 14520 0 1 37200
box 0 0 1 1
use contact_32  contact_32_82
timestamp 1643671299
transform 1 0 14520 0 1 35280
box 0 0 1 1
use contact_32  contact_32_83
timestamp 1643671299
transform 1 0 14400 0 1 13680
box 0 0 1 1
use contact_32  contact_32_84
timestamp 1643671299
transform 1 0 14400 0 1 14040
box 0 0 1 1
use contact_32  contact_32_85
timestamp 1643671299
transform 1 0 12840 0 1 14040
box 0 0 1 1
use contact_32  contact_32_86
timestamp 1643671299
transform 1 0 12840 0 1 12480
box 0 0 1 1
use contact_32  contact_32_87
timestamp 1643671299
transform 1 0 12840 0 1 12360
box 0 0 1 1
use contact_32  contact_32_88
timestamp 1643671299
transform 1 0 12840 0 1 10800
box 0 0 1 1
use contact_32  contact_32_89
timestamp 1643671299
transform 1 0 14400 0 1 16680
box 0 0 1 1
use contact_32  contact_32_90
timestamp 1643671299
transform 1 0 14400 0 1 15840
box 0 0 1 1
use contact_32  contact_32_91
timestamp 1643671299
transform 1 0 12840 0 1 14160
box 0 0 1 1
use contact_32  contact_32_92
timestamp 1643671299
transform 1 0 12840 0 1 15720
box 0 0 1 1
use contact_32  contact_32_93
timestamp 1643671299
transform 1 0 14400 0 1 16800
box 0 0 1 1
use contact_32  contact_32_94
timestamp 1643671299
transform 1 0 14400 0 1 17400
box 0 0 1 1
use contact_32  contact_32_95
timestamp 1643671299
transform 1 0 14400 0 1 19800
box 0 0 1 1
use contact_32  contact_32_96
timestamp 1643671299
transform 1 0 14400 0 1 17520
box 0 0 1 1
use contact_32  contact_32_97
timestamp 1643671299
transform 1 0 480 0 1 6240
box 0 0 1 1
use contact_32  contact_32_98
timestamp 1643671299
transform 1 0 2400 0 1 4680
box 0 0 1 1
use contact_32  contact_32_99
timestamp 1643671299
transform 1 0 2400 0 1 6240
box 0 0 1 1
use contact_32  contact_32_100
timestamp 1643671299
transform 1 0 74400 0 1 3480
box 0 0 1 1
use contact_32  contact_32_101
timestamp 1643671299
transform 1 0 74400 0 1 1800
box 0 0 1 1
use contact_32  contact_32_102
timestamp 1643671299
transform 1 0 74400 0 1 20400
box 0 0 1 1
use contact_32  contact_32_103
timestamp 1643671299
transform 1 0 74400 0 1 30480
box 0 0 1 1
use contact_32  contact_32_104
timestamp 1643671299
transform 1 0 74400 0 1 23640
box 0 0 1 1
use contact_32  contact_32_105
timestamp 1643671299
transform 1 0 74400 0 1 21960
box 0 0 1 1
use contact_32  contact_32_106
timestamp 1643671299
transform 1 0 74400 0 1 8640
box 0 0 1 1
use contact_32  contact_32_107
timestamp 1643671299
transform 1 0 74400 0 1 25320
box 0 0 1 1
use contact_32  contact_32_108
timestamp 1643671299
transform 1 0 74400 0 1 17040
box 0 0 1 1
use contact_32  contact_32_109
timestamp 1643671299
transform 1 0 74400 0 1 18720
box 0 0 1 1
use contact_32  contact_32_110
timestamp 1643671299
transform 1 0 74400 0 1 6960
box 0 0 1 1
use contact_32  contact_32_111
timestamp 1643671299
transform 1 0 74400 0 1 15240
box 0 0 1 1
use contact_32  contact_32_112
timestamp 1643671299
transform 1 0 74400 0 1 10200
box 0 0 1 1
use contact_32  contact_32_113
timestamp 1643671299
transform 1 0 74400 0 1 13560
box 0 0 1 1
use contact_32  contact_32_114
timestamp 1643671299
transform 1 0 74400 0 1 32040
box 0 0 1 1
use contact_32  contact_32_115
timestamp 1643671299
transform 1 0 74400 0 1 11880
box 0 0 1 1
use contact_32  contact_32_116
timestamp 1643671299
transform 1 0 74400 0 1 27120
box 0 0 1 1
use contact_32  contact_32_117
timestamp 1643671299
transform 1 0 74400 0 1 33720
box 0 0 1 1
use contact_32  contact_32_118
timestamp 1643671299
transform 1 0 74400 0 1 28800
box 0 0 1 1
use contact_32  contact_32_119
timestamp 1643671299
transform 1 0 74400 0 1 5160
box 0 0 1 1
use contact_32  contact_32_120
timestamp 1643671299
transform 1 0 74400 0 1 35400
box 0 0 1 1
use contact_32  contact_32_121
timestamp 1643671299
transform 1 0 72600 0 1 1080
box 0 0 1 1
use contact_32  contact_32_122
timestamp 1643671299
transform 1 0 72600 0 1 1440
box 0 0 1 1
use contact_32  contact_32_123
timestamp 1643671299
transform 1 0 72480 0 1 36600
box 0 0 1 1
use contact_32  contact_32_124
timestamp 1643671299
transform 1 0 72480 0 1 36240
box 0 0 1 1
use contact_32  contact_32_125
timestamp 1643671299
transform 1 0 70800 0 1 36600
box 0 0 1 1
use contact_32  contact_32_126
timestamp 1643671299
transform 1 0 70800 0 1 36240
box 0 0 1 1
use contact_32  contact_32_127
timestamp 1643671299
transform 1 0 70800 0 1 1080
box 0 0 1 1
use contact_32  contact_32_128
timestamp 1643671299
transform 1 0 70800 0 1 1440
box 0 0 1 1
use contact_32  contact_32_129
timestamp 1643671299
transform 1 0 69240 0 1 1080
box 0 0 1 1
use contact_32  contact_32_130
timestamp 1643671299
transform 1 0 69240 0 1 1440
box 0 0 1 1
use contact_32  contact_32_131
timestamp 1643671299
transform 1 0 69240 0 1 36600
box 0 0 1 1
use contact_32  contact_32_132
timestamp 1643671299
transform 1 0 69240 0 1 36240
box 0 0 1 1
use contact_32  contact_32_133
timestamp 1643671299
transform 1 0 67560 0 1 36600
box 0 0 1 1
use contact_32  contact_32_134
timestamp 1643671299
transform 1 0 67560 0 1 36240
box 0 0 1 1
use contact_32  contact_32_135
timestamp 1643671299
transform 1 0 67560 0 1 1080
box 0 0 1 1
use contact_32  contact_32_136
timestamp 1643671299
transform 1 0 67560 0 1 1440
box 0 0 1 1
use contact_32  contact_32_137
timestamp 1643671299
transform 1 0 65760 0 1 36600
box 0 0 1 1
use contact_32  contact_32_138
timestamp 1643671299
transform 1 0 65760 0 1 36240
box 0 0 1 1
use contact_32  contact_32_139
timestamp 1643671299
transform 1 0 65760 0 1 1080
box 0 0 1 1
use contact_32  contact_32_140
timestamp 1643671299
transform 1 0 65760 0 1 1440
box 0 0 1 1
use contact_32  contact_32_141
timestamp 1643671299
transform 1 0 64080 0 1 1080
box 0 0 1 1
use contact_32  contact_32_142
timestamp 1643671299
transform 1 0 64080 0 1 1440
box 0 0 1 1
use contact_32  contact_32_143
timestamp 1643671299
transform 1 0 64200 0 1 36600
box 0 0 1 1
use contact_32  contact_32_144
timestamp 1643671299
transform 1 0 64200 0 1 36240
box 0 0 1 1
use contact_32  contact_32_145
timestamp 1643671299
transform 1 0 62400 0 1 36600
box 0 0 1 1
use contact_32  contact_32_146
timestamp 1643671299
transform 1 0 62400 0 1 36240
box 0 0 1 1
use contact_32  contact_32_147
timestamp 1643671299
transform 1 0 62520 0 1 1080
box 0 0 1 1
use contact_32  contact_32_148
timestamp 1643671299
transform 1 0 62520 0 1 1440
box 0 0 1 1
use contact_32  contact_32_149
timestamp 1643671299
transform 1 0 60720 0 1 1080
box 0 0 1 1
use contact_32  contact_32_150
timestamp 1643671299
transform 1 0 60720 0 1 1440
box 0 0 1 1
use contact_32  contact_32_151
timestamp 1643671299
transform 1 0 60720 0 1 36600
box 0 0 1 1
use contact_32  contact_32_152
timestamp 1643671299
transform 1 0 60720 0 1 36240
box 0 0 1 1
use contact_32  contact_32_153
timestamp 1643671299
transform 1 0 59040 0 1 1080
box 0 0 1 1
use contact_32  contact_32_154
timestamp 1643671299
transform 1 0 59040 0 1 1440
box 0 0 1 1
use contact_32  contact_32_155
timestamp 1643671299
transform 1 0 59160 0 1 36600
box 0 0 1 1
use contact_32  contact_32_156
timestamp 1643671299
transform 1 0 59160 0 1 36240
box 0 0 1 1
use contact_32  contact_32_157
timestamp 1643671299
transform 1 0 57360 0 1 36600
box 0 0 1 1
use contact_32  contact_32_158
timestamp 1643671299
transform 1 0 57360 0 1 36240
box 0 0 1 1
use contact_32  contact_32_159
timestamp 1643671299
transform 1 0 57360 0 1 1080
box 0 0 1 1
use contact_32  contact_32_160
timestamp 1643671299
transform 1 0 57360 0 1 1440
box 0 0 1 1
use contact_32  contact_32_161
timestamp 1643671299
transform 1 0 55800 0 1 1080
box 0 0 1 1
use contact_32  contact_32_162
timestamp 1643671299
transform 1 0 55800 0 1 1440
box 0 0 1 1
use contact_32  contact_32_163
timestamp 1643671299
transform 1 0 55680 0 1 36600
box 0 0 1 1
use contact_32  contact_32_164
timestamp 1643671299
transform 1 0 55680 0 1 36240
box 0 0 1 1
use contact_32  contact_32_165
timestamp 1643671299
transform 1 0 54120 0 1 36600
box 0 0 1 1
use contact_32  contact_32_166
timestamp 1643671299
transform 1 0 54120 0 1 36240
box 0 0 1 1
use contact_32  contact_32_167
timestamp 1643671299
transform 1 0 54120 0 1 1080
box 0 0 1 1
use contact_32  contact_32_168
timestamp 1643671299
transform 1 0 54120 0 1 1440
box 0 0 1 1
use contact_32  contact_32_169
timestamp 1643671299
transform 1 0 52440 0 1 1080
box 0 0 1 1
use contact_32  contact_32_170
timestamp 1643671299
transform 1 0 52440 0 1 1440
box 0 0 1 1
use contact_32  contact_32_171
timestamp 1643671299
transform 1 0 52440 0 1 36600
box 0 0 1 1
use contact_32  contact_32_172
timestamp 1643671299
transform 1 0 52440 0 1 36240
box 0 0 1 1
use contact_32  contact_32_173
timestamp 1643671299
transform 1 0 50640 0 1 1080
box 0 0 1 1
use contact_32  contact_32_174
timestamp 1643671299
transform 1 0 50640 0 1 1440
box 0 0 1 1
use contact_32  contact_32_175
timestamp 1643671299
transform 1 0 50640 0 1 36600
box 0 0 1 1
use contact_32  contact_32_176
timestamp 1643671299
transform 1 0 50640 0 1 36240
box 0 0 1 1
use contact_32  contact_32_177
timestamp 1643671299
transform 1 0 48960 0 1 36600
box 0 0 1 1
use contact_32  contact_32_178
timestamp 1643671299
transform 1 0 48960 0 1 36240
box 0 0 1 1
use contact_32  contact_32_179
timestamp 1643671299
transform 1 0 48960 0 1 1080
box 0 0 1 1
use contact_32  contact_32_180
timestamp 1643671299
transform 1 0 48960 0 1 1440
box 0 0 1 1
use contact_32  contact_32_181
timestamp 1643671299
transform 1 0 47400 0 1 1080
box 0 0 1 1
use contact_32  contact_32_182
timestamp 1643671299
transform 1 0 47400 0 1 1440
box 0 0 1 1
use contact_32  contact_32_183
timestamp 1643671299
transform 1 0 47400 0 1 36600
box 0 0 1 1
use contact_32  contact_32_184
timestamp 1643671299
transform 1 0 47400 0 1 36240
box 0 0 1 1
use contact_32  contact_32_185
timestamp 1643671299
transform 1 0 45720 0 1 36600
box 0 0 1 1
use contact_32  contact_32_186
timestamp 1643671299
transform 1 0 45720 0 1 36240
box 0 0 1 1
use contact_32  contact_32_187
timestamp 1643671299
transform 1 0 45720 0 1 1080
box 0 0 1 1
use contact_32  contact_32_188
timestamp 1643671299
transform 1 0 45720 0 1 1440
box 0 0 1 1
use contact_32  contact_32_189
timestamp 1643671299
transform 1 0 44040 0 1 1080
box 0 0 1 1
use contact_32  contact_32_190
timestamp 1643671299
transform 1 0 44040 0 1 1440
box 0 0 1 1
use contact_32  contact_32_191
timestamp 1643671299
transform 1 0 43920 0 1 36600
box 0 0 1 1
use contact_32  contact_32_192
timestamp 1643671299
transform 1 0 43920 0 1 36240
box 0 0 1 1
use contact_32  contact_32_193
timestamp 1643671299
transform 1 0 43680 0 1 9600
box 0 0 1 1
use contact_32  contact_32_194
timestamp 1643671299
transform 1 0 43680 0 1 8400
box 0 0 1 1
use contact_32  contact_32_195
timestamp 1643671299
transform 1 0 42360 0 1 1080
box 0 0 1 1
use contact_32  contact_32_196
timestamp 1643671299
transform 1 0 42360 0 1 1440
box 0 0 1 1
use contact_32  contact_32_197
timestamp 1643671299
transform 1 0 42360 0 1 36600
box 0 0 1 1
use contact_32  contact_32_198
timestamp 1643671299
transform 1 0 42360 0 1 36240
box 0 0 1 1
use contact_32  contact_32_199
timestamp 1643671299
transform 1 0 42120 0 1 9600
box 0 0 1 1
use contact_32  contact_32_200
timestamp 1643671299
transform 1 0 42120 0 1 8400
box 0 0 1 1
use contact_32  contact_32_201
timestamp 1643671299
transform 1 0 40680 0 1 36600
box 0 0 1 1
use contact_32  contact_32_202
timestamp 1643671299
transform 1 0 40680 0 1 36240
box 0 0 1 1
use contact_32  contact_32_203
timestamp 1643671299
transform 1 0 40560 0 1 1080
box 0 0 1 1
use contact_32  contact_32_204
timestamp 1643671299
transform 1 0 40560 0 1 1440
box 0 0 1 1
use contact_32  contact_32_205
timestamp 1643671299
transform 1 0 40560 0 1 9600
box 0 0 1 1
use contact_32  contact_32_206
timestamp 1643671299
transform 1 0 40560 0 1 8400
box 0 0 1 1
use contact_32  contact_32_207
timestamp 1643671299
transform 1 0 38880 0 1 36600
box 0 0 1 1
use contact_32  contact_32_208
timestamp 1643671299
transform 1 0 38880 0 1 36240
box 0 0 1 1
use contact_32  contact_32_209
timestamp 1643671299
transform 1 0 38640 0 1 1080
box 0 0 1 1
use contact_32  contact_32_210
timestamp 1643671299
transform 1 0 38640 0 1 1440
box 0 0 1 1
use contact_32  contact_32_211
timestamp 1643671299
transform 1 0 39000 0 1 9600
box 0 0 1 1
use contact_32  contact_32_212
timestamp 1643671299
transform 1 0 39000 0 1 8400
box 0 0 1 1
use contact_32  contact_32_213
timestamp 1643671299
transform 1 0 37440 0 1 1080
box 0 0 1 1
use contact_32  contact_32_214
timestamp 1643671299
transform 1 0 37440 0 1 1440
box 0 0 1 1
use contact_32  contact_32_215
timestamp 1643671299
transform 1 0 37320 0 1 36600
box 0 0 1 1
use contact_32  contact_32_216
timestamp 1643671299
transform 1 0 37320 0 1 36240
box 0 0 1 1
use contact_32  contact_32_217
timestamp 1643671299
transform 1 0 37440 0 1 9600
box 0 0 1 1
use contact_32  contact_32_218
timestamp 1643671299
transform 1 0 37440 0 1 8400
box 0 0 1 1
use contact_32  contact_32_219
timestamp 1643671299
transform 1 0 35760 0 1 9600
box 0 0 1 1
use contact_32  contact_32_220
timestamp 1643671299
transform 1 0 35760 0 1 8400
box 0 0 1 1
use contact_32  contact_32_221
timestamp 1643671299
transform 1 0 35520 0 1 1080
box 0 0 1 1
use contact_32  contact_32_222
timestamp 1643671299
transform 1 0 35520 0 1 1440
box 0 0 1 1
use contact_32  contact_32_223
timestamp 1643671299
transform 1 0 35640 0 1 36600
box 0 0 1 1
use contact_32  contact_32_224
timestamp 1643671299
transform 1 0 35640 0 1 36240
box 0 0 1 1
use contact_32  contact_32_225
timestamp 1643671299
transform 1 0 35520 0 1 1560
box 0 0 1 1
use contact_32  contact_32_226
timestamp 1643671299
transform 1 0 35520 0 1 3120
box 0 0 1 1
use contact_32  contact_32_227
timestamp 1643671299
transform 1 0 35040 0 1 3240
box 0 0 1 1
use contact_32  contact_32_228
timestamp 1643671299
transform 1 0 35040 0 1 5160
box 0 0 1 1
use contact_32  contact_32_229
timestamp 1643671299
transform 1 0 34320 0 1 9600
box 0 0 1 1
use contact_32  contact_32_230
timestamp 1643671299
transform 1 0 34320 0 1 8400
box 0 0 1 1
use contact_32  contact_32_231
timestamp 1643671299
transform 1 0 33840 0 1 1080
box 0 0 1 1
use contact_32  contact_32_232
timestamp 1643671299
transform 1 0 33840 0 1 1440
box 0 0 1 1
use contact_32  contact_32_233
timestamp 1643671299
transform 1 0 33840 0 1 36600
box 0 0 1 1
use contact_32  contact_32_234
timestamp 1643671299
transform 1 0 33840 0 1 36240
box 0 0 1 1
use contact_32  contact_32_235
timestamp 1643671299
transform 1 0 32760 0 1 9600
box 0 0 1 1
use contact_32  contact_32_236
timestamp 1643671299
transform 1 0 32760 0 1 8400
box 0 0 1 1
use contact_32  contact_32_237
timestamp 1643671299
transform 1 0 32160 0 1 1080
box 0 0 1 1
use contact_32  contact_32_238
timestamp 1643671299
transform 1 0 32160 0 1 1440
box 0 0 1 1
use contact_32  contact_32_239
timestamp 1643671299
transform 1 0 32160 0 1 36600
box 0 0 1 1
use contact_32  contact_32_240
timestamp 1643671299
transform 1 0 32160 0 1 36240
box 0 0 1 1
use contact_32  contact_32_241
timestamp 1643671299
transform 1 0 31200 0 1 9600
box 0 0 1 1
use contact_32  contact_32_242
timestamp 1643671299
transform 1 0 31200 0 1 8400
box 0 0 1 1
use contact_32  contact_32_243
timestamp 1643671299
transform 1 0 30480 0 1 1080
box 0 0 1 1
use contact_32  contact_32_244
timestamp 1643671299
transform 1 0 30480 0 1 1440
box 0 0 1 1
use contact_32  contact_32_245
timestamp 1643671299
transform 1 0 30480 0 1 36600
box 0 0 1 1
use contact_32  contact_32_246
timestamp 1643671299
transform 1 0 30480 0 1 36240
box 0 0 1 1
use contact_32  contact_32_247
timestamp 1643671299
transform 1 0 29640 0 1 9600
box 0 0 1 1
use contact_32  contact_32_248
timestamp 1643671299
transform 1 0 29640 0 1 8400
box 0 0 1 1
use contact_32  contact_32_249
timestamp 1643671299
transform 1 0 28920 0 1 36600
box 0 0 1 1
use contact_32  contact_32_250
timestamp 1643671299
transform 1 0 28920 0 1 36240
box 0 0 1 1
use contact_32  contact_32_251
timestamp 1643671299
transform 1 0 29040 0 1 1080
box 0 0 1 1
use contact_32  contact_32_252
timestamp 1643671299
transform 1 0 29040 0 1 1440
box 0 0 1 1
use contact_32  contact_32_253
timestamp 1643671299
transform 1 0 28080 0 1 9600
box 0 0 1 1
use contact_32  contact_32_254
timestamp 1643671299
transform 1 0 28080 0 1 8400
box 0 0 1 1
use contact_32  contact_32_255
timestamp 1643671299
transform 1 0 27120 0 1 1080
box 0 0 1 1
use contact_32  contact_32_256
timestamp 1643671299
transform 1 0 27120 0 1 1440
box 0 0 1 1
use contact_32  contact_32_257
timestamp 1643671299
transform 1 0 27120 0 1 36600
box 0 0 1 1
use contact_32  contact_32_258
timestamp 1643671299
transform 1 0 27120 0 1 36240
box 0 0 1 1
use contact_32  contact_32_259
timestamp 1643671299
transform 1 0 26520 0 1 9600
box 0 0 1 1
use contact_32  contact_32_260
timestamp 1643671299
transform 1 0 26520 0 1 8400
box 0 0 1 1
use contact_32  contact_32_261
timestamp 1643671299
transform 1 0 25440 0 1 36600
box 0 0 1 1
use contact_32  contact_32_262
timestamp 1643671299
transform 1 0 25440 0 1 36240
box 0 0 1 1
use contact_32  contact_32_263
timestamp 1643671299
transform 1 0 25440 0 1 1080
box 0 0 1 1
use contact_32  contact_32_264
timestamp 1643671299
transform 1 0 25440 0 1 1440
box 0 0 1 1
use contact_32  contact_32_265
timestamp 1643671299
transform 1 0 24960 0 1 9600
box 0 0 1 1
use contact_32  contact_32_266
timestamp 1643671299
transform 1 0 24960 0 1 8400
box 0 0 1 1
use contact_32  contact_32_267
timestamp 1643671299
transform 1 0 23880 0 1 1080
box 0 0 1 1
use contact_32  contact_32_268
timestamp 1643671299
transform 1 0 23880 0 1 1440
box 0 0 1 1
use contact_32  contact_32_269
timestamp 1643671299
transform 1 0 23760 0 1 36600
box 0 0 1 1
use contact_32  contact_32_270
timestamp 1643671299
transform 1 0 23760 0 1 36240
box 0 0 1 1
use contact_32  contact_32_271
timestamp 1643671299
transform 1 0 22080 0 1 36600
box 0 0 1 1
use contact_32  contact_32_272
timestamp 1643671299
transform 1 0 22080 0 1 36240
box 0 0 1 1
use contact_32  contact_32_273
timestamp 1643671299
transform 1 0 22200 0 1 1080
box 0 0 1 1
use contact_32  contact_32_274
timestamp 1643671299
transform 1 0 22200 0 1 1440
box 0 0 1 1
use contact_32  contact_32_275
timestamp 1643671299
transform 1 0 20520 0 1 36600
box 0 0 1 1
use contact_32  contact_32_276
timestamp 1643671299
transform 1 0 20520 0 1 36240
box 0 0 1 1
use contact_32  contact_32_277
timestamp 1643671299
transform 1 0 20520 0 1 1080
box 0 0 1 1
use contact_32  contact_32_278
timestamp 1643671299
transform 1 0 20520 0 1 1440
box 0 0 1 1
use contact_32  contact_32_279
timestamp 1643671299
transform 1 0 19680 0 1 21480
box 0 0 1 1
use contact_32  contact_32_280
timestamp 1643671299
transform 1 0 19680 0 1 24360
box 0 0 1 1
use contact_32  contact_32_281
timestamp 1643671299
transform 1 0 20280 0 1 9720
box 0 0 1 1
use contact_32  contact_32_282
timestamp 1643671299
transform 1 0 20280 0 1 12120
box 0 0 1 1
use contact_32  contact_32_283
timestamp 1643671299
transform 1 0 19680 0 1 15120
box 0 0 1 1
use contact_32  contact_32_284
timestamp 1643671299
transform 1 0 19680 0 1 12240
box 0 0 1 1
use contact_32  contact_32_285
timestamp 1643671299
transform 1 0 20400 0 1 36120
box 0 0 1 1
use contact_32  contact_32_286
timestamp 1643671299
transform 1 0 20400 0 1 33720
box 0 0 1 1
use contact_32  contact_32_287
timestamp 1643671299
transform 1 0 19560 0 1 21240
box 0 0 1 1
use contact_32  contact_32_288
timestamp 1643671299
transform 1 0 19560 0 1 18360
box 0 0 1 1
use contact_32  contact_32_289
timestamp 1643671299
transform 1 0 18840 0 1 36600
box 0 0 1 1
use contact_32  contact_32_290
timestamp 1643671299
transform 1 0 18840 0 1 36240
box 0 0 1 1
use contact_32  contact_32_291
timestamp 1643671299
transform 1 0 18840 0 1 1080
box 0 0 1 1
use contact_32  contact_32_292
timestamp 1643671299
transform 1 0 18840 0 1 1440
box 0 0 1 1
use contact_32  contact_32_293
timestamp 1643671299
transform 1 0 19560 0 1 27600
box 0 0 1 1
use contact_32  contact_32_294
timestamp 1643671299
transform 1 0 19560 0 1 30240
box 0 0 1 1
use contact_32  contact_32_295
timestamp 1643671299
transform 1 0 19560 0 1 24480
box 0 0 1 1
use contact_32  contact_32_296
timestamp 1643671299
transform 1 0 19560 0 1 27240
box 0 0 1 1
use contact_32  contact_32_297
timestamp 1643671299
transform 1 0 19560 0 1 33600
box 0 0 1 1
use contact_32  contact_32_298
timestamp 1643671299
transform 1 0 19560 0 1 33360
box 0 0 1 1
use contact_32  contact_32_299
timestamp 1643671299
transform 1 0 18480 0 1 30360
box 0 0 1 1
use contact_32  contact_32_300
timestamp 1643671299
transform 1 0 18480 0 1 33240
box 0 0 1 1
use contact_32  contact_32_301
timestamp 1643671299
transform 1 0 20280 0 1 9600
box 0 0 1 1
use contact_32  contact_32_302
timestamp 1643671299
transform 1 0 20280 0 1 8760
box 0 0 1 1
use contact_32  contact_32_303
timestamp 1643671299
transform 1 0 17160 0 1 36600
box 0 0 1 1
use contact_32  contact_32_304
timestamp 1643671299
transform 1 0 17160 0 1 36240
box 0 0 1 1
use contact_32  contact_32_305
timestamp 1643671299
transform 1 0 17160 0 1 1080
box 0 0 1 1
use contact_32  contact_32_306
timestamp 1643671299
transform 1 0 17160 0 1 1440
box 0 0 1 1
use contact_32  contact_32_307
timestamp 1643671299
transform 1 0 15360 0 1 1080
box 0 0 1 1
use contact_32  contact_32_308
timestamp 1643671299
transform 1 0 15360 0 1 1440
box 0 0 1 1
use contact_32  contact_32_309
timestamp 1643671299
transform 1 0 15480 0 1 36600
box 0 0 1 1
use contact_32  contact_32_310
timestamp 1643671299
transform 1 0 15480 0 1 36240
box 0 0 1 1
use contact_32  contact_32_311
timestamp 1643671299
transform 1 0 15000 0 1 30720
box 0 0 1 1
use contact_32  contact_32_312
timestamp 1643671299
transform 1 0 15000 0 1 33600
box 0 0 1 1
use contact_32  contact_32_313
timestamp 1643671299
transform 1 0 14400 0 1 21480
box 0 0 1 1
use contact_32  contact_32_314
timestamp 1643671299
transform 1 0 14400 0 1 24360
box 0 0 1 1
use contact_32  contact_32_315
timestamp 1643671299
transform 1 0 13680 0 1 36600
box 0 0 1 1
use contact_32  contact_32_316
timestamp 1643671299
transform 1 0 13680 0 1 36240
box 0 0 1 1
use contact_32  contact_32_317
timestamp 1643671299
transform 1 0 14400 0 1 33720
box 0 0 1 1
use contact_32  contact_32_318
timestamp 1643671299
transform 1 0 14400 0 1 36120
box 0 0 1 1
use contact_32  contact_32_319
timestamp 1643671299
transform 1 0 13800 0 1 1080
box 0 0 1 1
use contact_32  contact_32_320
timestamp 1643671299
transform 1 0 13800 0 1 1440
box 0 0 1 1
use contact_32  contact_32_321
timestamp 1643671299
transform 1 0 12960 0 1 13320
box 0 0 1 1
use contact_32  contact_32_322
timestamp 1643671299
transform 1 0 12960 0 1 14880
box 0 0 1 1
use contact_32  contact_32_323
timestamp 1643671299
transform 1 0 12960 0 1 16560
box 0 0 1 1
use contact_32  contact_32_324
timestamp 1643671299
transform 1 0 12960 0 1 15000
box 0 0 1 1
use contact_32  contact_32_325
timestamp 1643671299
transform 1 0 14400 0 1 12120
box 0 0 1 1
use contact_32  contact_32_326
timestamp 1643671299
transform 1 0 14400 0 1 11640
box 0 0 1 1
use contact_32  contact_32_327
timestamp 1643671299
transform 1 0 12960 0 1 13200
box 0 0 1 1
use contact_32  contact_32_328
timestamp 1643671299
transform 1 0 12960 0 1 11640
box 0 0 1 1
use contact_32  contact_32_329
timestamp 1643671299
transform 1 0 12000 0 1 36600
box 0 0 1 1
use contact_32  contact_32_330
timestamp 1643671299
transform 1 0 12000 0 1 36240
box 0 0 1 1
use contact_32  contact_32_331
timestamp 1643671299
transform 1 0 12000 0 1 1080
box 0 0 1 1
use contact_32  contact_32_332
timestamp 1643671299
transform 1 0 12000 0 1 1440
box 0 0 1 1
use contact_32  contact_32_333
timestamp 1643671299
transform 1 0 10440 0 1 1080
box 0 0 1 1
use contact_32  contact_32_334
timestamp 1643671299
transform 1 0 10440 0 1 1440
box 0 0 1 1
use contact_32  contact_32_335
timestamp 1643671299
transform 1 0 10440 0 1 36600
box 0 0 1 1
use contact_32  contact_32_336
timestamp 1643671299
transform 1 0 10440 0 1 36240
box 0 0 1 1
use contact_32  contact_32_337
timestamp 1643671299
transform 1 0 8640 0 1 36600
box 0 0 1 1
use contact_32  contact_32_338
timestamp 1643671299
transform 1 0 8640 0 1 36240
box 0 0 1 1
use contact_32  contact_32_339
timestamp 1643671299
transform 1 0 8640 0 1 1080
box 0 0 1 1
use contact_32  contact_32_340
timestamp 1643671299
transform 1 0 8640 0 1 1440
box 0 0 1 1
use contact_32  contact_32_341
timestamp 1643671299
transform 1 0 6960 0 1 1080
box 0 0 1 1
use contact_32  contact_32_342
timestamp 1643671299
transform 1 0 6960 0 1 1440
box 0 0 1 1
use contact_32  contact_32_343
timestamp 1643671299
transform 1 0 6960 0 1 36600
box 0 0 1 1
use contact_32  contact_32_344
timestamp 1643671299
transform 1 0 6960 0 1 36240
box 0 0 1 1
use contact_32  contact_32_345
timestamp 1643671299
transform 1 0 5400 0 1 36600
box 0 0 1 1
use contact_32  contact_32_346
timestamp 1643671299
transform 1 0 5400 0 1 36240
box 0 0 1 1
use contact_32  contact_32_347
timestamp 1643671299
transform 1 0 5400 0 1 1080
box 0 0 1 1
use contact_32  contact_32_348
timestamp 1643671299
transform 1 0 5400 0 1 1440
box 0 0 1 1
use contact_32  contact_32_349
timestamp 1643671299
transform 1 0 3720 0 1 36600
box 0 0 1 1
use contact_32  contact_32_350
timestamp 1643671299
transform 1 0 3720 0 1 36240
box 0 0 1 1
use contact_32  contact_32_351
timestamp 1643671299
transform 1 0 3600 0 1 1080
box 0 0 1 1
use contact_32  contact_32_352
timestamp 1643671299
transform 1 0 3600 0 1 1440
box 0 0 1 1
use contact_32  contact_32_353
timestamp 1643671299
transform 1 0 1920 0 1 36600
box 0 0 1 1
use contact_32  contact_32_354
timestamp 1643671299
transform 1 0 1920 0 1 36240
box 0 0 1 1
use contact_32  contact_32_355
timestamp 1643671299
transform 1 0 2040 0 1 1080
box 0 0 1 1
use contact_32  contact_32_356
timestamp 1643671299
transform 1 0 2040 0 1 1440
box 0 0 1 1
use contact_32  contact_32_357
timestamp 1643671299
transform 1 0 1080 0 1 33840
box 0 0 1 1
use contact_32  contact_32_358
timestamp 1643671299
transform 1 0 1080 0 1 18600
box 0 0 1 1
use contact_32  contact_32_359
timestamp 1643671299
transform 1 0 1080 0 1 15360
box 0 0 1 1
use contact_32  contact_32_360
timestamp 1643671299
transform 1 0 1080 0 1 35520
box 0 0 1 1
use contact_32  contact_32_361
timestamp 1643671299
transform 1 0 1080 0 1 3600
box 0 0 1 1
use contact_32  contact_32_362
timestamp 1643671299
transform 1 0 1920 0 1 1560
box 0 0 1 1
use contact_32  contact_32_363
timestamp 1643671299
transform 1 0 1920 0 1 1800
box 0 0 1 1
use contact_32  contact_32_364
timestamp 1643671299
transform 1 0 1080 0 1 11880
box 0 0 1 1
use contact_32  contact_32_365
timestamp 1643671299
transform 1 0 1080 0 1 17040
box 0 0 1 1
use contact_32  contact_32_366
timestamp 1643671299
transform 1 0 1080 0 1 8520
box 0 0 1 1
use contact_32  contact_32_367
timestamp 1643671299
transform 1 0 1080 0 1 25440
box 0 0 1 1
use contact_32  contact_32_368
timestamp 1643671299
transform 1 0 1080 0 1 30360
box 0 0 1 1
use contact_32  contact_32_369
timestamp 1643671299
transform 1 0 1080 0 1 20280
box 0 0 1 1
use contact_32  contact_32_370
timestamp 1643671299
transform 1 0 1080 0 1 6960
box 0 0 1 1
use contact_32  contact_32_371
timestamp 1643671299
transform 1 0 1080 0 1 13680
box 0 0 1 1
use contact_32  contact_32_372
timestamp 1643671299
transform 1 0 1080 0 1 23760
box 0 0 1 1
use contact_32  contact_32_373
timestamp 1643671299
transform 1 0 1080 0 1 10200
box 0 0 1 1
use contact_32  contact_32_374
timestamp 1643671299
transform 1 0 1080 0 1 32040
box 0 0 1 1
use contact_32  contact_32_375
timestamp 1643671299
transform 1 0 1080 0 1 28680
box 0 0 1 1
use contact_32  contact_32_376
timestamp 1643671299
transform 1 0 1080 0 1 21960
box 0 0 1 1
use contact_32  contact_32_377
timestamp 1643671299
transform 1 0 1080 0 1 5280
box 0 0 1 1
use contact_32  contact_32_378
timestamp 1643671299
transform 1 0 1080 0 1 27120
box 0 0 1 1
use contact_39  contact_39_0
timestamp 1643671299
transform 1 0 75120 0 1 480
box 0 0 1 1
use contact_39  contact_39_1
timestamp 1643671299
transform 1 0 75120 0 1 37200
box 0 0 1 1
use contact_39  contact_39_2
timestamp 1643671299
transform 1 0 240 0 1 240
box 0 0 1 1
use contact_39  contact_39_3
timestamp 1643671299
transform 1 0 75240 0 1 37440
box 0 0 1 1
use contact_39  contact_39_4
timestamp 1643671299
transform 1 0 75240 0 1 480
box 0 0 1 1
use contact_39  contact_39_5
timestamp 1643671299
transform 1 0 480 0 1 37320
box 0 0 1 1
use contact_39  contact_39_6
timestamp 1643671299
transform 1 0 480 0 1 360
box 0 0 1 1
use contact_39  contact_39_7
timestamp 1643671299
transform 1 0 75120 0 1 37320
box 0 0 1 1
use contact_39  contact_39_8
timestamp 1643671299
transform 1 0 75000 0 1 37440
box 0 0 1 1
use contact_39  contact_39_9
timestamp 1643671299
transform 1 0 360 0 1 37440
box 0 0 1 1
use contact_39  contact_39_10
timestamp 1643671299
transform 1 0 75000 0 1 480
box 0 0 1 1
use contact_39  contact_39_11
timestamp 1643671299
transform 1 0 75240 0 1 37200
box 0 0 1 1
use contact_39  contact_39_12
timestamp 1643671299
transform 1 0 75240 0 1 240
box 0 0 1 1
use contact_39  contact_39_13
timestamp 1643671299
transform 1 0 75120 0 1 360
box 0 0 1 1
use contact_39  contact_39_14
timestamp 1643671299
transform 1 0 240 0 1 37320
box 0 0 1 1
use contact_39  contact_39_15
timestamp 1643671299
transform 1 0 75000 0 1 37200
box 0 0 1 1
use contact_39  contact_39_16
timestamp 1643671299
transform 1 0 360 0 1 480
box 0 0 1 1
use contact_39  contact_39_17
timestamp 1643671299
transform 1 0 360 0 1 37200
box 0 0 1 1
use contact_39  contact_39_18
timestamp 1643671299
transform 1 0 75000 0 1 240
box 0 0 1 1
use contact_39  contact_39_19
timestamp 1643671299
transform 1 0 240 0 1 360
box 0 0 1 1
use contact_39  contact_39_20
timestamp 1643671299
transform 1 0 360 0 1 240
box 0 0 1 1
use contact_39  contact_39_21
timestamp 1643671299
transform 1 0 75240 0 1 37320
box 0 0 1 1
use contact_39  contact_39_22
timestamp 1643671299
transform 1 0 480 0 1 37440
box 0 0 1 1
use contact_39  contact_39_23
timestamp 1643671299
transform 1 0 75240 0 1 360
box 0 0 1 1
use contact_39  contact_39_24
timestamp 1643671299
transform 1 0 480 0 1 480
box 0 0 1 1
use contact_39  contact_39_25
timestamp 1643671299
transform 1 0 480 0 1 37200
box 0 0 1 1
use contact_39  contact_39_26
timestamp 1643671299
transform 1 0 360 0 1 37320
box 0 0 1 1
use contact_39  contact_39_27
timestamp 1643671299
transform 1 0 360 0 1 360
box 0 0 1 1
use contact_39  contact_39_28
timestamp 1643671299
transform 1 0 75000 0 1 37320
box 0 0 1 1
use contact_39  contact_39_29
timestamp 1643671299
transform 1 0 240 0 1 37440
box 0 0 1 1
use contact_39  contact_39_30
timestamp 1643671299
transform 1 0 75000 0 1 360
box 0 0 1 1
use contact_39  contact_39_31
timestamp 1643671299
transform 1 0 240 0 1 480
box 0 0 1 1
use contact_39  contact_39_32
timestamp 1643671299
transform 1 0 240 0 1 37200
box 0 0 1 1
use contact_39  contact_39_33
timestamp 1643671299
transform 1 0 480 0 1 240
box 0 0 1 1
use contact_39  contact_39_34
timestamp 1643671299
transform 1 0 75120 0 1 37440
box 0 0 1 1
use contact_39  contact_39_35
timestamp 1643671299
transform 1 0 75120 0 1 240
box 0 0 1 1
use contact_39  contact_39_36
timestamp 1643671299
transform 1 0 74400 0 1 36720
box 0 0 1 1
use contact_39  contact_39_37
timestamp 1643671299
transform 1 0 840 0 1 36840
box 0 0 1 1
use contact_39  contact_39_38
timestamp 1643671299
transform 1 0 74640 0 1 840
box 0 0 1 1
use contact_39  contact_39_39
timestamp 1643671299
transform 1 0 1080 0 1 36600
box 0 0 1 1
use contact_39  contact_39_40
timestamp 1643671299
transform 1 0 1080 0 1 960
box 0 0 1 1
use contact_39  contact_39_41
timestamp 1643671299
transform 1 0 74520 0 1 36840
box 0 0 1 1
use contact_39  contact_39_42
timestamp 1643671299
transform 1 0 74520 0 1 36600
box 0 0 1 1
use contact_39  contact_39_43
timestamp 1643671299
transform 1 0 960 0 1 1080
box 0 0 1 1
use contact_39  contact_39_44
timestamp 1643671299
transform 1 0 74400 0 1 1080
box 0 0 1 1
use contact_39  contact_39_45
timestamp 1643671299
transform 1 0 74520 0 1 960
box 0 0 1 1
use contact_39  contact_39_46
timestamp 1643671299
transform 1 0 74400 0 1 840
box 0 0 1 1
use contact_39  contact_39_47
timestamp 1643671299
transform 1 0 840 0 1 36600
box 0 0 1 1
use contact_39  contact_39_48
timestamp 1643671299
transform 1 0 840 0 1 960
box 0 0 1 1
use contact_39  contact_39_49
timestamp 1643671299
transform 1 0 74640 0 1 36840
box 0 0 1 1
use contact_39  contact_39_50
timestamp 1643671299
transform 1 0 960 0 1 36720
box 0 0 1 1
use contact_39  contact_39_51
timestamp 1643671299
transform 1 0 960 0 1 840
box 0 0 1 1
use contact_39  contact_39_52
timestamp 1643671299
transform 1 0 74640 0 1 1080
box 0 0 1 1
use contact_39  contact_39_53
timestamp 1643671299
transform 1 0 74520 0 1 36720
box 0 0 1 1
use contact_39  contact_39_54
timestamp 1643671299
transform 1 0 74400 0 1 36840
box 0 0 1 1
use contact_39  contact_39_55
timestamp 1643671299
transform 1 0 74640 0 1 36600
box 0 0 1 1
use contact_39  contact_39_56
timestamp 1643671299
transform 1 0 74640 0 1 960
box 0 0 1 1
use contact_39  contact_39_57
timestamp 1643671299
transform 1 0 1080 0 1 36720
box 0 0 1 1
use contact_39  contact_39_58
timestamp 1643671299
transform 1 0 1080 0 1 1080
box 0 0 1 1
use contact_39  contact_39_59
timestamp 1643671299
transform 1 0 74520 0 1 1080
box 0 0 1 1
use contact_39  contact_39_60
timestamp 1643671299
transform 1 0 960 0 1 36600
box 0 0 1 1
use contact_39  contact_39_61
timestamp 1643671299
transform 1 0 960 0 1 36840
box 0 0 1 1
use contact_39  contact_39_62
timestamp 1643671299
transform 1 0 74400 0 1 36600
box 0 0 1 1
use contact_39  contact_39_63
timestamp 1643671299
transform 1 0 960 0 1 960
box 0 0 1 1
use contact_39  contact_39_64
timestamp 1643671299
transform 1 0 74400 0 1 960
box 0 0 1 1
use contact_39  contact_39_65
timestamp 1643671299
transform 1 0 840 0 1 36720
box 0 0 1 1
use contact_39  contact_39_66
timestamp 1643671299
transform 1 0 840 0 1 1080
box 0 0 1 1
use contact_39  contact_39_67
timestamp 1643671299
transform 1 0 1080 0 1 840
box 0 0 1 1
use contact_39  contact_39_68
timestamp 1643671299
transform 1 0 840 0 1 840
box 0 0 1 1
use contact_39  contact_39_69
timestamp 1643671299
transform 1 0 74520 0 1 840
box 0 0 1 1
use contact_39  contact_39_70
timestamp 1643671299
transform 1 0 74640 0 1 36720
box 0 0 1 1
use contact_39  contact_39_71
timestamp 1643671299
transform 1 0 1080 0 1 36840
box 0 0 1 1
use contact_32  contact_32_379
timestamp 1643671299
transform 1 0 12480 0 1 12120
box 0 0 1 1
use contact_32  contact_32_380
timestamp 1643671299
transform 1 0 12360 0 1 10920
box 0 0 1 1
use contact_32  contact_32_381
timestamp 1643671299
transform 1 0 48120 0 1 9240
box 0 0 1 1
use contact_32  contact_32_382
timestamp 1643671299
transform 1 0 46560 0 1 9240
box 0 0 1 1
use contact_32  contact_32_383
timestamp 1643671299
transform 1 0 45000 0 1 9360
box 0 0 1 1
use contact_32  contact_32_384
timestamp 1643671299
transform 1 0 43440 0 1 9360
box 0 0 1 1
use contact_32  contact_32_385
timestamp 1643671299
transform 1 0 41880 0 1 9360
box 0 0 1 1
use contact_32  contact_32_386
timestamp 1643671299
transform 1 0 40320 0 1 9240
box 0 0 1 1
use contact_32  contact_32_387
timestamp 1643671299
transform 1 0 38760 0 1 9240
box 0 0 1 1
use contact_32  contact_32_388
timestamp 1643671299
transform 1 0 37200 0 1 9240
box 0 0 1 1
use contact_32  contact_32_389
timestamp 1643671299
transform 1 0 35640 0 1 9240
box 0 0 1 1
use contact_32  contact_32_390
timestamp 1643671299
transform 1 0 34080 0 1 9240
box 0 0 1 1
use contact_32  contact_32_391
timestamp 1643671299
transform 1 0 32520 0 1 9240
box 0 0 1 1
use contact_32  contact_32_392
timestamp 1643671299
transform 1 0 30960 0 1 9240
box 0 0 1 1
use contact_32  contact_32_393
timestamp 1643671299
transform 1 0 29400 0 1 9240
box 0 0 1 1
use contact_32  contact_32_394
timestamp 1643671299
transform 1 0 27840 0 1 9240
box 0 0 1 1
use contact_32  contact_32_395
timestamp 1643671299
transform 1 0 26280 0 1 9240
box 0 0 1 1
use contact_32  contact_32_396
timestamp 1643671299
transform 1 0 24840 0 1 9360
box 0 0 1 1
use contact_32  contact_32_397
timestamp 1643671299
transform 1 0 6000 0 1 5760
box 0 0 1 1
use contact_32  contact_32_398
timestamp 1643671299
transform 1 0 15240 0 1 2520
box 0 0 1 1
use contact_32  contact_32_399
timestamp 1643671299
transform 1 0 39120 0 1 2520
box 0 0 1 1
use contact_32  contact_32_400
timestamp 1643671299
transform 1 0 37680 0 1 2520
box 0 0 1 1
use contact_32  contact_32_401
timestamp 1643671299
transform 1 0 36000 0 1 2520
box 0 0 1 1
use contact_32  contact_32_402
timestamp 1643671299
transform 1 0 34560 0 1 2520
box 0 0 1 1
use contact_32  contact_32_403
timestamp 1643671299
transform 1 0 33120 0 1 2520
box 0 0 1 1
use contact_32  contact_32_404
timestamp 1643671299
transform 1 0 31680 0 1 2520
box 0 0 1 1
use contact_32  contact_32_405
timestamp 1643671299
transform 1 0 30240 0 1 2520
box 0 0 1 1
use contact_32  contact_32_406
timestamp 1643671299
transform 1 0 28800 0 1 2520
box 0 0 1 1
use contact_32  contact_32_407
timestamp 1643671299
transform 1 0 27240 0 1 2520
box 0 0 1 1
use contact_32  contact_32_408
timestamp 1643671299
transform 1 0 25800 0 1 2520
box 0 0 1 1
use contact_32  contact_32_409
timestamp 1643671299
transform 1 0 24360 0 1 2520
box 0 0 1 1
use contact_32  contact_32_410
timestamp 1643671299
transform 1 0 22800 0 1 2520
box 0 0 1 1
use contact_32  contact_32_411
timestamp 1643671299
transform 1 0 21360 0 1 2520
box 0 0 1 1
use contact_32  contact_32_412
timestamp 1643671299
transform 1 0 19680 0 1 2520
box 0 0 1 1
use contact_32  contact_32_413
timestamp 1643671299
transform 1 0 18240 0 1 2520
box 0 0 1 1
use contact_32  contact_32_414
timestamp 1643671299
transform 1 0 16920 0 1 2520
box 0 0 1 1
use contact_37  contact_37_0
timestamp 1643671299
transform 1 0 1507 0 1 36097
box -11 -11 233 233
use contact_37  contact_37_1
timestamp 1643671299
transform 1 0 73855 0 1 36097
box -11 -11 233 233
use contact_37  contact_37_2
timestamp 1643671299
transform 1 0 73855 0 1 1453
box -11 -11 233 233
use contact_37  contact_37_3
timestamp 1643671299
transform 1 0 1507 0 1 1453
box -11 -11 233 233
use contact_17  contact_17_0
timestamp 1643671299
transform 1 0 73951 0 1 35821
box 0 0 1 1
use contact_13  contact_13_0
timestamp 1643671299
transform 1 0 73937 0 1 35813
box 0 0 1 1
use contact_21  contact_21_0
timestamp 1643671299
transform 1 0 73941 0 1 35795
box 0 0 1 1
use contact_18  contact_18_0
timestamp 1643671299
transform 1 0 73936 0 1 35470
box 0 0 1 1
use contact_17  contact_17_1
timestamp 1643671299
transform 1 0 73951 0 1 35485
box 0 0 1 1
use contact_13  contact_13_1
timestamp 1643671299
transform 1 0 73937 0 1 35477
box 0 0 1 1
use contact_21  contact_21_1
timestamp 1643671299
transform 1 0 73941 0 1 35459
box 0 0 1 1
use contact_17  contact_17_2
timestamp 1643671299
transform 1 0 73951 0 1 35149
box 0 0 1 1
use contact_13  contact_13_2
timestamp 1643671299
transform 1 0 73937 0 1 35141
box 0 0 1 1
use contact_21  contact_21_2
timestamp 1643671299
transform 1 0 73941 0 1 35123
box 0 0 1 1
use contact_17  contact_17_3
timestamp 1643671299
transform 1 0 73951 0 1 34813
box 0 0 1 1
use contact_13  contact_13_3
timestamp 1643671299
transform 1 0 73937 0 1 34805
box 0 0 1 1
use contact_21  contact_21_3
timestamp 1643671299
transform 1 0 73941 0 1 34787
box 0 0 1 1
use contact_17  contact_17_4
timestamp 1643671299
transform 1 0 73951 0 1 34477
box 0 0 1 1
use contact_13  contact_13_4
timestamp 1643671299
transform 1 0 73937 0 1 34469
box 0 0 1 1
use contact_21  contact_21_4
timestamp 1643671299
transform 1 0 73941 0 1 34451
box 0 0 1 1
use contact_17  contact_17_5
timestamp 1643671299
transform 1 0 73951 0 1 34141
box 0 0 1 1
use contact_13  contact_13_5
timestamp 1643671299
transform 1 0 73937 0 1 34133
box 0 0 1 1
use contact_21  contact_21_5
timestamp 1643671299
transform 1 0 73941 0 1 34115
box 0 0 1 1
use contact_18  contact_18_1
timestamp 1643671299
transform 1 0 73936 0 1 33790
box 0 0 1 1
use contact_17  contact_17_6
timestamp 1643671299
transform 1 0 73951 0 1 33805
box 0 0 1 1
use contact_13  contact_13_6
timestamp 1643671299
transform 1 0 73937 0 1 33797
box 0 0 1 1
use contact_21  contact_21_6
timestamp 1643671299
transform 1 0 73941 0 1 33779
box 0 0 1 1
use contact_17  contact_17_7
timestamp 1643671299
transform 1 0 73951 0 1 33469
box 0 0 1 1
use contact_13  contact_13_7
timestamp 1643671299
transform 1 0 73937 0 1 33461
box 0 0 1 1
use contact_21  contact_21_7
timestamp 1643671299
transform 1 0 73941 0 1 33443
box 0 0 1 1
use contact_17  contact_17_8
timestamp 1643671299
transform 1 0 73951 0 1 33133
box 0 0 1 1
use contact_13  contact_13_8
timestamp 1643671299
transform 1 0 73937 0 1 33125
box 0 0 1 1
use contact_21  contact_21_8
timestamp 1643671299
transform 1 0 73941 0 1 33107
box 0 0 1 1
use contact_17  contact_17_9
timestamp 1643671299
transform 1 0 73951 0 1 32797
box 0 0 1 1
use contact_13  contact_13_9
timestamp 1643671299
transform 1 0 73937 0 1 32789
box 0 0 1 1
use contact_21  contact_21_9
timestamp 1643671299
transform 1 0 73941 0 1 32771
box 0 0 1 1
use contact_17  contact_17_10
timestamp 1643671299
transform 1 0 73951 0 1 32461
box 0 0 1 1
use contact_13  contact_13_10
timestamp 1643671299
transform 1 0 73937 0 1 32453
box 0 0 1 1
use contact_21  contact_21_10
timestamp 1643671299
transform 1 0 73941 0 1 32435
box 0 0 1 1
use contact_18  contact_18_2
timestamp 1643671299
transform 1 0 73936 0 1 32110
box 0 0 1 1
use contact_17  contact_17_11
timestamp 1643671299
transform 1 0 73951 0 1 32125
box 0 0 1 1
use contact_13  contact_13_11
timestamp 1643671299
transform 1 0 73937 0 1 32117
box 0 0 1 1
use contact_21  contact_21_11
timestamp 1643671299
transform 1 0 73941 0 1 32099
box 0 0 1 1
use contact_17  contact_17_12
timestamp 1643671299
transform 1 0 73951 0 1 31789
box 0 0 1 1
use contact_13  contact_13_12
timestamp 1643671299
transform 1 0 73937 0 1 31781
box 0 0 1 1
use contact_21  contact_21_12
timestamp 1643671299
transform 1 0 73941 0 1 31763
box 0 0 1 1
use contact_17  contact_17_13
timestamp 1643671299
transform 1 0 73951 0 1 31453
box 0 0 1 1
use contact_13  contact_13_13
timestamp 1643671299
transform 1 0 73937 0 1 31445
box 0 0 1 1
use contact_21  contact_21_13
timestamp 1643671299
transform 1 0 73941 0 1 31427
box 0 0 1 1
use contact_17  contact_17_14
timestamp 1643671299
transform 1 0 73951 0 1 31117
box 0 0 1 1
use contact_13  contact_13_14
timestamp 1643671299
transform 1 0 73937 0 1 31109
box 0 0 1 1
use contact_21  contact_21_14
timestamp 1643671299
transform 1 0 73941 0 1 31091
box 0 0 1 1
use contact_17  contact_17_15
timestamp 1643671299
transform 1 0 73951 0 1 30781
box 0 0 1 1
use contact_13  contact_13_15
timestamp 1643671299
transform 1 0 73937 0 1 30773
box 0 0 1 1
use contact_21  contact_21_15
timestamp 1643671299
transform 1 0 73941 0 1 30755
box 0 0 1 1
use contact_18  contact_18_3
timestamp 1643671299
transform 1 0 73936 0 1 30430
box 0 0 1 1
use contact_17  contact_17_16
timestamp 1643671299
transform 1 0 73951 0 1 30445
box 0 0 1 1
use contact_13  contact_13_16
timestamp 1643671299
transform 1 0 73937 0 1 30437
box 0 0 1 1
use contact_21  contact_21_16
timestamp 1643671299
transform 1 0 73941 0 1 30419
box 0 0 1 1
use contact_17  contact_17_17
timestamp 1643671299
transform 1 0 73951 0 1 30109
box 0 0 1 1
use contact_13  contact_13_17
timestamp 1643671299
transform 1 0 73937 0 1 30101
box 0 0 1 1
use contact_21  contact_21_17
timestamp 1643671299
transform 1 0 73941 0 1 30083
box 0 0 1 1
use contact_17  contact_17_18
timestamp 1643671299
transform 1 0 73951 0 1 29773
box 0 0 1 1
use contact_13  contact_13_18
timestamp 1643671299
transform 1 0 73937 0 1 29765
box 0 0 1 1
use contact_21  contact_21_18
timestamp 1643671299
transform 1 0 73941 0 1 29747
box 0 0 1 1
use contact_17  contact_17_19
timestamp 1643671299
transform 1 0 73951 0 1 29437
box 0 0 1 1
use contact_13  contact_13_19
timestamp 1643671299
transform 1 0 73937 0 1 29429
box 0 0 1 1
use contact_21  contact_21_19
timestamp 1643671299
transform 1 0 73941 0 1 29411
box 0 0 1 1
use contact_17  contact_17_20
timestamp 1643671299
transform 1 0 73951 0 1 29101
box 0 0 1 1
use contact_13  contact_13_20
timestamp 1643671299
transform 1 0 73937 0 1 29093
box 0 0 1 1
use contact_21  contact_21_20
timestamp 1643671299
transform 1 0 73941 0 1 29075
box 0 0 1 1
use contact_18  contact_18_4
timestamp 1643671299
transform 1 0 73936 0 1 28750
box 0 0 1 1
use contact_17  contact_17_21
timestamp 1643671299
transform 1 0 73951 0 1 28765
box 0 0 1 1
use contact_13  contact_13_21
timestamp 1643671299
transform 1 0 73937 0 1 28757
box 0 0 1 1
use contact_21  contact_21_21
timestamp 1643671299
transform 1 0 73941 0 1 28739
box 0 0 1 1
use contact_17  contact_17_22
timestamp 1643671299
transform 1 0 73951 0 1 28429
box 0 0 1 1
use contact_13  contact_13_22
timestamp 1643671299
transform 1 0 73937 0 1 28421
box 0 0 1 1
use contact_21  contact_21_22
timestamp 1643671299
transform 1 0 73941 0 1 28403
box 0 0 1 1
use contact_17  contact_17_23
timestamp 1643671299
transform 1 0 73951 0 1 28093
box 0 0 1 1
use contact_13  contact_13_23
timestamp 1643671299
transform 1 0 73937 0 1 28085
box 0 0 1 1
use contact_21  contact_21_23
timestamp 1643671299
transform 1 0 73941 0 1 28067
box 0 0 1 1
use contact_17  contact_17_24
timestamp 1643671299
transform 1 0 73951 0 1 27757
box 0 0 1 1
use contact_13  contact_13_24
timestamp 1643671299
transform 1 0 73937 0 1 27749
box 0 0 1 1
use contact_21  contact_21_24
timestamp 1643671299
transform 1 0 73941 0 1 27731
box 0 0 1 1
use contact_17  contact_17_25
timestamp 1643671299
transform 1 0 73951 0 1 27421
box 0 0 1 1
use contact_13  contact_13_25
timestamp 1643671299
transform 1 0 73937 0 1 27413
box 0 0 1 1
use contact_21  contact_21_25
timestamp 1643671299
transform 1 0 73941 0 1 27395
box 0 0 1 1
use contact_18  contact_18_5
timestamp 1643671299
transform 1 0 73936 0 1 27070
box 0 0 1 1
use contact_17  contact_17_26
timestamp 1643671299
transform 1 0 73951 0 1 27085
box 0 0 1 1
use contact_13  contact_13_26
timestamp 1643671299
transform 1 0 73937 0 1 27077
box 0 0 1 1
use contact_21  contact_21_26
timestamp 1643671299
transform 1 0 73941 0 1 27059
box 0 0 1 1
use contact_17  contact_17_27
timestamp 1643671299
transform 1 0 73951 0 1 26749
box 0 0 1 1
use contact_13  contact_13_27
timestamp 1643671299
transform 1 0 73937 0 1 26741
box 0 0 1 1
use contact_21  contact_21_27
timestamp 1643671299
transform 1 0 73941 0 1 26723
box 0 0 1 1
use contact_17  contact_17_28
timestamp 1643671299
transform 1 0 73951 0 1 26413
box 0 0 1 1
use contact_13  contact_13_28
timestamp 1643671299
transform 1 0 73937 0 1 26405
box 0 0 1 1
use contact_21  contact_21_28
timestamp 1643671299
transform 1 0 73941 0 1 26387
box 0 0 1 1
use contact_17  contact_17_29
timestamp 1643671299
transform 1 0 73951 0 1 26077
box 0 0 1 1
use contact_13  contact_13_29
timestamp 1643671299
transform 1 0 73937 0 1 26069
box 0 0 1 1
use contact_21  contact_21_29
timestamp 1643671299
transform 1 0 73941 0 1 26051
box 0 0 1 1
use contact_17  contact_17_30
timestamp 1643671299
transform 1 0 73951 0 1 25741
box 0 0 1 1
use contact_13  contact_13_30
timestamp 1643671299
transform 1 0 73937 0 1 25733
box 0 0 1 1
use contact_21  contact_21_30
timestamp 1643671299
transform 1 0 73941 0 1 25715
box 0 0 1 1
use contact_18  contact_18_6
timestamp 1643671299
transform 1 0 73936 0 1 25390
box 0 0 1 1
use contact_17  contact_17_31
timestamp 1643671299
transform 1 0 73951 0 1 25405
box 0 0 1 1
use contact_13  contact_13_31
timestamp 1643671299
transform 1 0 73937 0 1 25397
box 0 0 1 1
use contact_21  contact_21_31
timestamp 1643671299
transform 1 0 73941 0 1 25379
box 0 0 1 1
use contact_17  contact_17_32
timestamp 1643671299
transform 1 0 73951 0 1 25069
box 0 0 1 1
use contact_13  contact_13_32
timestamp 1643671299
transform 1 0 73937 0 1 25061
box 0 0 1 1
use contact_21  contact_21_32
timestamp 1643671299
transform 1 0 73941 0 1 25043
box 0 0 1 1
use contact_17  contact_17_33
timestamp 1643671299
transform 1 0 73951 0 1 24733
box 0 0 1 1
use contact_13  contact_13_33
timestamp 1643671299
transform 1 0 73937 0 1 24725
box 0 0 1 1
use contact_21  contact_21_33
timestamp 1643671299
transform 1 0 73941 0 1 24707
box 0 0 1 1
use contact_17  contact_17_34
timestamp 1643671299
transform 1 0 73951 0 1 24397
box 0 0 1 1
use contact_13  contact_13_34
timestamp 1643671299
transform 1 0 73937 0 1 24389
box 0 0 1 1
use contact_21  contact_21_34
timestamp 1643671299
transform 1 0 73941 0 1 24371
box 0 0 1 1
use contact_17  contact_17_35
timestamp 1643671299
transform 1 0 73951 0 1 24061
box 0 0 1 1
use contact_13  contact_13_35
timestamp 1643671299
transform 1 0 73937 0 1 24053
box 0 0 1 1
use contact_21  contact_21_35
timestamp 1643671299
transform 1 0 73941 0 1 24035
box 0 0 1 1
use contact_18  contact_18_7
timestamp 1643671299
transform 1 0 73936 0 1 23710
box 0 0 1 1
use contact_17  contact_17_36
timestamp 1643671299
transform 1 0 73951 0 1 23725
box 0 0 1 1
use contact_13  contact_13_36
timestamp 1643671299
transform 1 0 73937 0 1 23717
box 0 0 1 1
use contact_21  contact_21_36
timestamp 1643671299
transform 1 0 73941 0 1 23699
box 0 0 1 1
use contact_17  contact_17_37
timestamp 1643671299
transform 1 0 73951 0 1 23389
box 0 0 1 1
use contact_13  contact_13_37
timestamp 1643671299
transform 1 0 73937 0 1 23381
box 0 0 1 1
use contact_21  contact_21_37
timestamp 1643671299
transform 1 0 73941 0 1 23363
box 0 0 1 1
use contact_17  contact_17_38
timestamp 1643671299
transform 1 0 73951 0 1 23053
box 0 0 1 1
use contact_13  contact_13_38
timestamp 1643671299
transform 1 0 73937 0 1 23045
box 0 0 1 1
use contact_21  contact_21_38
timestamp 1643671299
transform 1 0 73941 0 1 23027
box 0 0 1 1
use contact_17  contact_17_39
timestamp 1643671299
transform 1 0 73951 0 1 22717
box 0 0 1 1
use contact_13  contact_13_39
timestamp 1643671299
transform 1 0 73937 0 1 22709
box 0 0 1 1
use contact_21  contact_21_39
timestamp 1643671299
transform 1 0 73941 0 1 22691
box 0 0 1 1
use contact_17  contact_17_40
timestamp 1643671299
transform 1 0 73951 0 1 22381
box 0 0 1 1
use contact_13  contact_13_40
timestamp 1643671299
transform 1 0 73937 0 1 22373
box 0 0 1 1
use contact_21  contact_21_40
timestamp 1643671299
transform 1 0 73941 0 1 22355
box 0 0 1 1
use contact_18  contact_18_8
timestamp 1643671299
transform 1 0 73936 0 1 22030
box 0 0 1 1
use contact_17  contact_17_41
timestamp 1643671299
transform 1 0 73951 0 1 22045
box 0 0 1 1
use contact_13  contact_13_41
timestamp 1643671299
transform 1 0 73937 0 1 22037
box 0 0 1 1
use contact_21  contact_21_41
timestamp 1643671299
transform 1 0 73941 0 1 22019
box 0 0 1 1
use contact_17  contact_17_42
timestamp 1643671299
transform 1 0 73951 0 1 21709
box 0 0 1 1
use contact_13  contact_13_42
timestamp 1643671299
transform 1 0 73937 0 1 21701
box 0 0 1 1
use contact_21  contact_21_42
timestamp 1643671299
transform 1 0 73941 0 1 21683
box 0 0 1 1
use contact_17  contact_17_43
timestamp 1643671299
transform 1 0 73951 0 1 21373
box 0 0 1 1
use contact_13  contact_13_43
timestamp 1643671299
transform 1 0 73937 0 1 21365
box 0 0 1 1
use contact_21  contact_21_43
timestamp 1643671299
transform 1 0 73941 0 1 21347
box 0 0 1 1
use contact_17  contact_17_44
timestamp 1643671299
transform 1 0 73951 0 1 21037
box 0 0 1 1
use contact_13  contact_13_44
timestamp 1643671299
transform 1 0 73937 0 1 21029
box 0 0 1 1
use contact_21  contact_21_44
timestamp 1643671299
transform 1 0 73941 0 1 21011
box 0 0 1 1
use contact_17  contact_17_45
timestamp 1643671299
transform 1 0 73951 0 1 20701
box 0 0 1 1
use contact_13  contact_13_45
timestamp 1643671299
transform 1 0 73937 0 1 20693
box 0 0 1 1
use contact_21  contact_21_45
timestamp 1643671299
transform 1 0 73941 0 1 20675
box 0 0 1 1
use contact_18  contact_18_9
timestamp 1643671299
transform 1 0 73936 0 1 20350
box 0 0 1 1
use contact_17  contact_17_46
timestamp 1643671299
transform 1 0 73951 0 1 20365
box 0 0 1 1
use contact_13  contact_13_46
timestamp 1643671299
transform 1 0 73937 0 1 20357
box 0 0 1 1
use contact_21  contact_21_46
timestamp 1643671299
transform 1 0 73941 0 1 20339
box 0 0 1 1
use contact_17  contact_17_47
timestamp 1643671299
transform 1 0 73951 0 1 20029
box 0 0 1 1
use contact_13  contact_13_47
timestamp 1643671299
transform 1 0 73937 0 1 20021
box 0 0 1 1
use contact_21  contact_21_47
timestamp 1643671299
transform 1 0 73941 0 1 20003
box 0 0 1 1
use contact_17  contact_17_48
timestamp 1643671299
transform 1 0 73951 0 1 19693
box 0 0 1 1
use contact_13  contact_13_48
timestamp 1643671299
transform 1 0 73937 0 1 19685
box 0 0 1 1
use contact_21  contact_21_48
timestamp 1643671299
transform 1 0 73941 0 1 19667
box 0 0 1 1
use contact_17  contact_17_49
timestamp 1643671299
transform 1 0 73951 0 1 19357
box 0 0 1 1
use contact_13  contact_13_49
timestamp 1643671299
transform 1 0 73937 0 1 19349
box 0 0 1 1
use contact_21  contact_21_49
timestamp 1643671299
transform 1 0 73941 0 1 19331
box 0 0 1 1
use contact_17  contact_17_50
timestamp 1643671299
transform 1 0 73951 0 1 19021
box 0 0 1 1
use contact_13  contact_13_50
timestamp 1643671299
transform 1 0 73937 0 1 19013
box 0 0 1 1
use contact_21  contact_21_50
timestamp 1643671299
transform 1 0 73941 0 1 18995
box 0 0 1 1
use contact_18  contact_18_10
timestamp 1643671299
transform 1 0 73936 0 1 18670
box 0 0 1 1
use contact_17  contact_17_51
timestamp 1643671299
transform 1 0 73951 0 1 18685
box 0 0 1 1
use contact_13  contact_13_51
timestamp 1643671299
transform 1 0 73937 0 1 18677
box 0 0 1 1
use contact_21  contact_21_51
timestamp 1643671299
transform 1 0 73941 0 1 18659
box 0 0 1 1
use contact_17  contact_17_52
timestamp 1643671299
transform 1 0 73951 0 1 18349
box 0 0 1 1
use contact_13  contact_13_52
timestamp 1643671299
transform 1 0 73937 0 1 18341
box 0 0 1 1
use contact_21  contact_21_52
timestamp 1643671299
transform 1 0 73941 0 1 18323
box 0 0 1 1
use contact_17  contact_17_53
timestamp 1643671299
transform 1 0 73951 0 1 18013
box 0 0 1 1
use contact_13  contact_13_53
timestamp 1643671299
transform 1 0 73937 0 1 18005
box 0 0 1 1
use contact_21  contact_21_53
timestamp 1643671299
transform 1 0 73941 0 1 17987
box 0 0 1 1
use contact_17  contact_17_54
timestamp 1643671299
transform 1 0 73951 0 1 17677
box 0 0 1 1
use contact_13  contact_13_54
timestamp 1643671299
transform 1 0 73937 0 1 17669
box 0 0 1 1
use contact_21  contact_21_54
timestamp 1643671299
transform 1 0 73941 0 1 17651
box 0 0 1 1
use contact_17  contact_17_55
timestamp 1643671299
transform 1 0 73951 0 1 17341
box 0 0 1 1
use contact_13  contact_13_55
timestamp 1643671299
transform 1 0 73937 0 1 17333
box 0 0 1 1
use contact_21  contact_21_55
timestamp 1643671299
transform 1 0 73941 0 1 17315
box 0 0 1 1
use contact_18  contact_18_11
timestamp 1643671299
transform 1 0 73936 0 1 16990
box 0 0 1 1
use contact_17  contact_17_56
timestamp 1643671299
transform 1 0 73951 0 1 17005
box 0 0 1 1
use contact_13  contact_13_56
timestamp 1643671299
transform 1 0 73937 0 1 16997
box 0 0 1 1
use contact_21  contact_21_56
timestamp 1643671299
transform 1 0 73941 0 1 16979
box 0 0 1 1
use contact_17  contact_17_57
timestamp 1643671299
transform 1 0 73951 0 1 16669
box 0 0 1 1
use contact_13  contact_13_57
timestamp 1643671299
transform 1 0 73937 0 1 16661
box 0 0 1 1
use contact_21  contact_21_57
timestamp 1643671299
transform 1 0 73941 0 1 16643
box 0 0 1 1
use contact_17  contact_17_58
timestamp 1643671299
transform 1 0 73951 0 1 16333
box 0 0 1 1
use contact_13  contact_13_58
timestamp 1643671299
transform 1 0 73937 0 1 16325
box 0 0 1 1
use contact_21  contact_21_58
timestamp 1643671299
transform 1 0 73941 0 1 16307
box 0 0 1 1
use contact_17  contact_17_59
timestamp 1643671299
transform 1 0 73951 0 1 15997
box 0 0 1 1
use contact_13  contact_13_59
timestamp 1643671299
transform 1 0 73937 0 1 15989
box 0 0 1 1
use contact_21  contact_21_59
timestamp 1643671299
transform 1 0 73941 0 1 15971
box 0 0 1 1
use contact_17  contact_17_60
timestamp 1643671299
transform 1 0 73951 0 1 15661
box 0 0 1 1
use contact_13  contact_13_60
timestamp 1643671299
transform 1 0 73937 0 1 15653
box 0 0 1 1
use contact_21  contact_21_60
timestamp 1643671299
transform 1 0 73941 0 1 15635
box 0 0 1 1
use contact_18  contact_18_12
timestamp 1643671299
transform 1 0 73936 0 1 15310
box 0 0 1 1
use contact_17  contact_17_61
timestamp 1643671299
transform 1 0 73951 0 1 15325
box 0 0 1 1
use contact_13  contact_13_61
timestamp 1643671299
transform 1 0 73937 0 1 15317
box 0 0 1 1
use contact_21  contact_21_61
timestamp 1643671299
transform 1 0 73941 0 1 15299
box 0 0 1 1
use contact_17  contact_17_62
timestamp 1643671299
transform 1 0 73951 0 1 14989
box 0 0 1 1
use contact_13  contact_13_62
timestamp 1643671299
transform 1 0 73937 0 1 14981
box 0 0 1 1
use contact_21  contact_21_62
timestamp 1643671299
transform 1 0 73941 0 1 14963
box 0 0 1 1
use contact_17  contact_17_63
timestamp 1643671299
transform 1 0 73951 0 1 14653
box 0 0 1 1
use contact_13  contact_13_63
timestamp 1643671299
transform 1 0 73937 0 1 14645
box 0 0 1 1
use contact_21  contact_21_63
timestamp 1643671299
transform 1 0 73941 0 1 14627
box 0 0 1 1
use contact_17  contact_17_64
timestamp 1643671299
transform 1 0 73951 0 1 14317
box 0 0 1 1
use contact_13  contact_13_64
timestamp 1643671299
transform 1 0 73937 0 1 14309
box 0 0 1 1
use contact_21  contact_21_64
timestamp 1643671299
transform 1 0 73941 0 1 14291
box 0 0 1 1
use contact_17  contact_17_65
timestamp 1643671299
transform 1 0 73951 0 1 13981
box 0 0 1 1
use contact_13  contact_13_65
timestamp 1643671299
transform 1 0 73937 0 1 13973
box 0 0 1 1
use contact_21  contact_21_65
timestamp 1643671299
transform 1 0 73941 0 1 13955
box 0 0 1 1
use contact_18  contact_18_13
timestamp 1643671299
transform 1 0 73936 0 1 13630
box 0 0 1 1
use contact_17  contact_17_66
timestamp 1643671299
transform 1 0 73951 0 1 13645
box 0 0 1 1
use contact_13  contact_13_66
timestamp 1643671299
transform 1 0 73937 0 1 13637
box 0 0 1 1
use contact_21  contact_21_66
timestamp 1643671299
transform 1 0 73941 0 1 13619
box 0 0 1 1
use contact_17  contact_17_67
timestamp 1643671299
transform 1 0 73951 0 1 13309
box 0 0 1 1
use contact_13  contact_13_67
timestamp 1643671299
transform 1 0 73937 0 1 13301
box 0 0 1 1
use contact_21  contact_21_67
timestamp 1643671299
transform 1 0 73941 0 1 13283
box 0 0 1 1
use contact_17  contact_17_68
timestamp 1643671299
transform 1 0 73951 0 1 12973
box 0 0 1 1
use contact_13  contact_13_68
timestamp 1643671299
transform 1 0 73937 0 1 12965
box 0 0 1 1
use contact_21  contact_21_68
timestamp 1643671299
transform 1 0 73941 0 1 12947
box 0 0 1 1
use contact_17  contact_17_69
timestamp 1643671299
transform 1 0 73951 0 1 12637
box 0 0 1 1
use contact_13  contact_13_69
timestamp 1643671299
transform 1 0 73937 0 1 12629
box 0 0 1 1
use contact_21  contact_21_69
timestamp 1643671299
transform 1 0 73941 0 1 12611
box 0 0 1 1
use contact_17  contact_17_70
timestamp 1643671299
transform 1 0 73951 0 1 12301
box 0 0 1 1
use contact_13  contact_13_70
timestamp 1643671299
transform 1 0 73937 0 1 12293
box 0 0 1 1
use contact_21  contact_21_70
timestamp 1643671299
transform 1 0 73941 0 1 12275
box 0 0 1 1
use contact_18  contact_18_14
timestamp 1643671299
transform 1 0 73936 0 1 11950
box 0 0 1 1
use contact_17  contact_17_71
timestamp 1643671299
transform 1 0 73951 0 1 11965
box 0 0 1 1
use contact_13  contact_13_71
timestamp 1643671299
transform 1 0 73937 0 1 11957
box 0 0 1 1
use contact_21  contact_21_71
timestamp 1643671299
transform 1 0 73941 0 1 11939
box 0 0 1 1
use contact_17  contact_17_72
timestamp 1643671299
transform 1 0 73951 0 1 11629
box 0 0 1 1
use contact_13  contact_13_72
timestamp 1643671299
transform 1 0 73937 0 1 11621
box 0 0 1 1
use contact_21  contact_21_72
timestamp 1643671299
transform 1 0 73941 0 1 11603
box 0 0 1 1
use contact_17  contact_17_73
timestamp 1643671299
transform 1 0 73951 0 1 11293
box 0 0 1 1
use contact_13  contact_13_73
timestamp 1643671299
transform 1 0 73937 0 1 11285
box 0 0 1 1
use contact_21  contact_21_73
timestamp 1643671299
transform 1 0 73941 0 1 11267
box 0 0 1 1
use contact_17  contact_17_74
timestamp 1643671299
transform 1 0 73951 0 1 10957
box 0 0 1 1
use contact_13  contact_13_74
timestamp 1643671299
transform 1 0 73937 0 1 10949
box 0 0 1 1
use contact_21  contact_21_74
timestamp 1643671299
transform 1 0 73941 0 1 10931
box 0 0 1 1
use contact_17  contact_17_75
timestamp 1643671299
transform 1 0 73951 0 1 10621
box 0 0 1 1
use contact_13  contact_13_75
timestamp 1643671299
transform 1 0 73937 0 1 10613
box 0 0 1 1
use contact_21  contact_21_75
timestamp 1643671299
transform 1 0 73941 0 1 10595
box 0 0 1 1
use contact_18  contact_18_15
timestamp 1643671299
transform 1 0 73936 0 1 10270
box 0 0 1 1
use contact_17  contact_17_76
timestamp 1643671299
transform 1 0 73951 0 1 10285
box 0 0 1 1
use contact_13  contact_13_76
timestamp 1643671299
transform 1 0 73937 0 1 10277
box 0 0 1 1
use contact_21  contact_21_76
timestamp 1643671299
transform 1 0 73941 0 1 10259
box 0 0 1 1
use contact_17  contact_17_77
timestamp 1643671299
transform 1 0 73951 0 1 9949
box 0 0 1 1
use contact_13  contact_13_77
timestamp 1643671299
transform 1 0 73937 0 1 9941
box 0 0 1 1
use contact_21  contact_21_77
timestamp 1643671299
transform 1 0 73941 0 1 9923
box 0 0 1 1
use contact_17  contact_17_78
timestamp 1643671299
transform 1 0 73951 0 1 9613
box 0 0 1 1
use contact_13  contact_13_78
timestamp 1643671299
transform 1 0 73937 0 1 9605
box 0 0 1 1
use contact_21  contact_21_78
timestamp 1643671299
transform 1 0 73941 0 1 9587
box 0 0 1 1
use contact_17  contact_17_79
timestamp 1643671299
transform 1 0 73951 0 1 9277
box 0 0 1 1
use contact_13  contact_13_79
timestamp 1643671299
transform 1 0 73937 0 1 9269
box 0 0 1 1
use contact_21  contact_21_79
timestamp 1643671299
transform 1 0 73941 0 1 9251
box 0 0 1 1
use contact_17  contact_17_80
timestamp 1643671299
transform 1 0 73951 0 1 8941
box 0 0 1 1
use contact_13  contact_13_80
timestamp 1643671299
transform 1 0 73937 0 1 8933
box 0 0 1 1
use contact_21  contact_21_80
timestamp 1643671299
transform 1 0 73941 0 1 8915
box 0 0 1 1
use contact_18  contact_18_16
timestamp 1643671299
transform 1 0 73936 0 1 8590
box 0 0 1 1
use contact_17  contact_17_81
timestamp 1643671299
transform 1 0 73951 0 1 8605
box 0 0 1 1
use contact_13  contact_13_81
timestamp 1643671299
transform 1 0 73937 0 1 8597
box 0 0 1 1
use contact_21  contact_21_81
timestamp 1643671299
transform 1 0 73941 0 1 8579
box 0 0 1 1
use contact_17  contact_17_82
timestamp 1643671299
transform 1 0 73951 0 1 8269
box 0 0 1 1
use contact_13  contact_13_82
timestamp 1643671299
transform 1 0 73937 0 1 8261
box 0 0 1 1
use contact_21  contact_21_82
timestamp 1643671299
transform 1 0 73941 0 1 8243
box 0 0 1 1
use contact_17  contact_17_83
timestamp 1643671299
transform 1 0 73951 0 1 7933
box 0 0 1 1
use contact_13  contact_13_83
timestamp 1643671299
transform 1 0 73937 0 1 7925
box 0 0 1 1
use contact_21  contact_21_83
timestamp 1643671299
transform 1 0 73941 0 1 7907
box 0 0 1 1
use contact_17  contact_17_84
timestamp 1643671299
transform 1 0 73951 0 1 7597
box 0 0 1 1
use contact_13  contact_13_84
timestamp 1643671299
transform 1 0 73937 0 1 7589
box 0 0 1 1
use contact_21  contact_21_84
timestamp 1643671299
transform 1 0 73941 0 1 7571
box 0 0 1 1
use contact_17  contact_17_85
timestamp 1643671299
transform 1 0 73951 0 1 7261
box 0 0 1 1
use contact_13  contact_13_85
timestamp 1643671299
transform 1 0 73937 0 1 7253
box 0 0 1 1
use contact_21  contact_21_85
timestamp 1643671299
transform 1 0 73941 0 1 7235
box 0 0 1 1
use contact_18  contact_18_17
timestamp 1643671299
transform 1 0 73936 0 1 6910
box 0 0 1 1
use contact_17  contact_17_86
timestamp 1643671299
transform 1 0 73951 0 1 6925
box 0 0 1 1
use contact_13  contact_13_86
timestamp 1643671299
transform 1 0 73937 0 1 6917
box 0 0 1 1
use contact_21  contact_21_86
timestamp 1643671299
transform 1 0 73941 0 1 6899
box 0 0 1 1
use contact_17  contact_17_87
timestamp 1643671299
transform 1 0 73951 0 1 6589
box 0 0 1 1
use contact_13  contact_13_87
timestamp 1643671299
transform 1 0 73937 0 1 6581
box 0 0 1 1
use contact_21  contact_21_87
timestamp 1643671299
transform 1 0 73941 0 1 6563
box 0 0 1 1
use contact_17  contact_17_88
timestamp 1643671299
transform 1 0 73951 0 1 6253
box 0 0 1 1
use contact_13  contact_13_88
timestamp 1643671299
transform 1 0 73937 0 1 6245
box 0 0 1 1
use contact_21  contact_21_88
timestamp 1643671299
transform 1 0 73941 0 1 6227
box 0 0 1 1
use contact_17  contact_17_89
timestamp 1643671299
transform 1 0 73951 0 1 5917
box 0 0 1 1
use contact_13  contact_13_89
timestamp 1643671299
transform 1 0 73937 0 1 5909
box 0 0 1 1
use contact_21  contact_21_89
timestamp 1643671299
transform 1 0 73941 0 1 5891
box 0 0 1 1
use contact_17  contact_17_90
timestamp 1643671299
transform 1 0 73951 0 1 5581
box 0 0 1 1
use contact_13  contact_13_90
timestamp 1643671299
transform 1 0 73937 0 1 5573
box 0 0 1 1
use contact_21  contact_21_90
timestamp 1643671299
transform 1 0 73941 0 1 5555
box 0 0 1 1
use contact_18  contact_18_18
timestamp 1643671299
transform 1 0 73936 0 1 5230
box 0 0 1 1
use contact_17  contact_17_91
timestamp 1643671299
transform 1 0 73951 0 1 5245
box 0 0 1 1
use contact_13  contact_13_91
timestamp 1643671299
transform 1 0 73937 0 1 5237
box 0 0 1 1
use contact_21  contact_21_91
timestamp 1643671299
transform 1 0 73941 0 1 5219
box 0 0 1 1
use contact_17  contact_17_92
timestamp 1643671299
transform 1 0 73951 0 1 4909
box 0 0 1 1
use contact_13  contact_13_92
timestamp 1643671299
transform 1 0 73937 0 1 4901
box 0 0 1 1
use contact_21  contact_21_92
timestamp 1643671299
transform 1 0 73941 0 1 4883
box 0 0 1 1
use contact_17  contact_17_93
timestamp 1643671299
transform 1 0 73951 0 1 4573
box 0 0 1 1
use contact_13  contact_13_93
timestamp 1643671299
transform 1 0 73937 0 1 4565
box 0 0 1 1
use contact_21  contact_21_93
timestamp 1643671299
transform 1 0 73941 0 1 4547
box 0 0 1 1
use contact_17  contact_17_94
timestamp 1643671299
transform 1 0 73951 0 1 4237
box 0 0 1 1
use contact_13  contact_13_94
timestamp 1643671299
transform 1 0 73937 0 1 4229
box 0 0 1 1
use contact_21  contact_21_94
timestamp 1643671299
transform 1 0 73941 0 1 4211
box 0 0 1 1
use contact_17  contact_17_95
timestamp 1643671299
transform 1 0 73951 0 1 3901
box 0 0 1 1
use contact_13  contact_13_95
timestamp 1643671299
transform 1 0 73937 0 1 3893
box 0 0 1 1
use contact_21  contact_21_95
timestamp 1643671299
transform 1 0 73941 0 1 3875
box 0 0 1 1
use contact_18  contact_18_19
timestamp 1643671299
transform 1 0 73936 0 1 3550
box 0 0 1 1
use contact_17  contact_17_96
timestamp 1643671299
transform 1 0 73951 0 1 3565
box 0 0 1 1
use contact_13  contact_13_96
timestamp 1643671299
transform 1 0 73937 0 1 3557
box 0 0 1 1
use contact_21  contact_21_96
timestamp 1643671299
transform 1 0 73941 0 1 3539
box 0 0 1 1
use contact_17  contact_17_97
timestamp 1643671299
transform 1 0 73951 0 1 3229
box 0 0 1 1
use contact_13  contact_13_97
timestamp 1643671299
transform 1 0 73937 0 1 3221
box 0 0 1 1
use contact_21  contact_21_97
timestamp 1643671299
transform 1 0 73941 0 1 3203
box 0 0 1 1
use contact_17  contact_17_98
timestamp 1643671299
transform 1 0 73951 0 1 2893
box 0 0 1 1
use contact_13  contact_13_98
timestamp 1643671299
transform 1 0 73937 0 1 2885
box 0 0 1 1
use contact_21  contact_21_98
timestamp 1643671299
transform 1 0 73941 0 1 2867
box 0 0 1 1
use contact_17  contact_17_99
timestamp 1643671299
transform 1 0 73951 0 1 2557
box 0 0 1 1
use contact_13  contact_13_99
timestamp 1643671299
transform 1 0 73937 0 1 2549
box 0 0 1 1
use contact_21  contact_21_99
timestamp 1643671299
transform 1 0 73941 0 1 2531
box 0 0 1 1
use contact_17  contact_17_100
timestamp 1643671299
transform 1 0 73951 0 1 2221
box 0 0 1 1
use contact_13  contact_13_100
timestamp 1643671299
transform 1 0 73937 0 1 2213
box 0 0 1 1
use contact_21  contact_21_100
timestamp 1643671299
transform 1 0 73941 0 1 2195
box 0 0 1 1
use contact_18  contact_18_20
timestamp 1643671299
transform 1 0 73936 0 1 1870
box 0 0 1 1
use contact_17  contact_17_101
timestamp 1643671299
transform 1 0 73951 0 1 1885
box 0 0 1 1
use contact_13  contact_13_101
timestamp 1643671299
transform 1 0 73937 0 1 1877
box 0 0 1 1
use contact_21  contact_21_101
timestamp 1643671299
transform 1 0 73941 0 1 1859
box 0 0 1 1
use contact_17  contact_17_102
timestamp 1643671299
transform 1 0 1603 0 1 35821
box 0 0 1 1
use contact_13  contact_13_102
timestamp 1643671299
transform 1 0 1589 0 1 35813
box 0 0 1 1
use contact_21  contact_21_102
timestamp 1643671299
transform 1 0 1593 0 1 35795
box 0 0 1 1
use contact_18  contact_18_21
timestamp 1643671299
transform 1 0 1588 0 1 35470
box 0 0 1 1
use contact_17  contact_17_103
timestamp 1643671299
transform 1 0 1603 0 1 35485
box 0 0 1 1
use contact_13  contact_13_103
timestamp 1643671299
transform 1 0 1589 0 1 35477
box 0 0 1 1
use contact_21  contact_21_103
timestamp 1643671299
transform 1 0 1593 0 1 35459
box 0 0 1 1
use contact_17  contact_17_104
timestamp 1643671299
transform 1 0 1603 0 1 35149
box 0 0 1 1
use contact_13  contact_13_104
timestamp 1643671299
transform 1 0 1589 0 1 35141
box 0 0 1 1
use contact_21  contact_21_104
timestamp 1643671299
transform 1 0 1593 0 1 35123
box 0 0 1 1
use contact_17  contact_17_105
timestamp 1643671299
transform 1 0 1603 0 1 34813
box 0 0 1 1
use contact_13  contact_13_105
timestamp 1643671299
transform 1 0 1589 0 1 34805
box 0 0 1 1
use contact_21  contact_21_105
timestamp 1643671299
transform 1 0 1593 0 1 34787
box 0 0 1 1
use contact_17  contact_17_106
timestamp 1643671299
transform 1 0 1603 0 1 34477
box 0 0 1 1
use contact_13  contact_13_106
timestamp 1643671299
transform 1 0 1589 0 1 34469
box 0 0 1 1
use contact_21  contact_21_106
timestamp 1643671299
transform 1 0 1593 0 1 34451
box 0 0 1 1
use contact_17  contact_17_107
timestamp 1643671299
transform 1 0 1603 0 1 34141
box 0 0 1 1
use contact_13  contact_13_107
timestamp 1643671299
transform 1 0 1589 0 1 34133
box 0 0 1 1
use contact_21  contact_21_107
timestamp 1643671299
transform 1 0 1593 0 1 34115
box 0 0 1 1
use contact_18  contact_18_22
timestamp 1643671299
transform 1 0 1588 0 1 33790
box 0 0 1 1
use contact_17  contact_17_108
timestamp 1643671299
transform 1 0 1603 0 1 33805
box 0 0 1 1
use contact_13  contact_13_108
timestamp 1643671299
transform 1 0 1589 0 1 33797
box 0 0 1 1
use contact_21  contact_21_108
timestamp 1643671299
transform 1 0 1593 0 1 33779
box 0 0 1 1
use contact_17  contact_17_109
timestamp 1643671299
transform 1 0 1603 0 1 33469
box 0 0 1 1
use contact_13  contact_13_109
timestamp 1643671299
transform 1 0 1589 0 1 33461
box 0 0 1 1
use contact_21  contact_21_109
timestamp 1643671299
transform 1 0 1593 0 1 33443
box 0 0 1 1
use contact_17  contact_17_110
timestamp 1643671299
transform 1 0 1603 0 1 33133
box 0 0 1 1
use contact_13  contact_13_110
timestamp 1643671299
transform 1 0 1589 0 1 33125
box 0 0 1 1
use contact_21  contact_21_110
timestamp 1643671299
transform 1 0 1593 0 1 33107
box 0 0 1 1
use contact_17  contact_17_111
timestamp 1643671299
transform 1 0 1603 0 1 32797
box 0 0 1 1
use contact_13  contact_13_111
timestamp 1643671299
transform 1 0 1589 0 1 32789
box 0 0 1 1
use contact_21  contact_21_111
timestamp 1643671299
transform 1 0 1593 0 1 32771
box 0 0 1 1
use contact_17  contact_17_112
timestamp 1643671299
transform 1 0 1603 0 1 32461
box 0 0 1 1
use contact_13  contact_13_112
timestamp 1643671299
transform 1 0 1589 0 1 32453
box 0 0 1 1
use contact_21  contact_21_112
timestamp 1643671299
transform 1 0 1593 0 1 32435
box 0 0 1 1
use contact_18  contact_18_23
timestamp 1643671299
transform 1 0 1588 0 1 32110
box 0 0 1 1
use contact_17  contact_17_113
timestamp 1643671299
transform 1 0 1603 0 1 32125
box 0 0 1 1
use contact_13  contact_13_113
timestamp 1643671299
transform 1 0 1589 0 1 32117
box 0 0 1 1
use contact_21  contact_21_113
timestamp 1643671299
transform 1 0 1593 0 1 32099
box 0 0 1 1
use contact_17  contact_17_114
timestamp 1643671299
transform 1 0 1603 0 1 31789
box 0 0 1 1
use contact_13  contact_13_114
timestamp 1643671299
transform 1 0 1589 0 1 31781
box 0 0 1 1
use contact_21  contact_21_114
timestamp 1643671299
transform 1 0 1593 0 1 31763
box 0 0 1 1
use contact_17  contact_17_115
timestamp 1643671299
transform 1 0 1603 0 1 31453
box 0 0 1 1
use contact_13  contact_13_115
timestamp 1643671299
transform 1 0 1589 0 1 31445
box 0 0 1 1
use contact_21  contact_21_115
timestamp 1643671299
transform 1 0 1593 0 1 31427
box 0 0 1 1
use contact_17  contact_17_116
timestamp 1643671299
transform 1 0 1603 0 1 31117
box 0 0 1 1
use contact_13  contact_13_116
timestamp 1643671299
transform 1 0 1589 0 1 31109
box 0 0 1 1
use contact_21  contact_21_116
timestamp 1643671299
transform 1 0 1593 0 1 31091
box 0 0 1 1
use contact_17  contact_17_117
timestamp 1643671299
transform 1 0 1603 0 1 30781
box 0 0 1 1
use contact_13  contact_13_117
timestamp 1643671299
transform 1 0 1589 0 1 30773
box 0 0 1 1
use contact_21  contact_21_117
timestamp 1643671299
transform 1 0 1593 0 1 30755
box 0 0 1 1
use contact_18  contact_18_24
timestamp 1643671299
transform 1 0 1588 0 1 30430
box 0 0 1 1
use contact_17  contact_17_118
timestamp 1643671299
transform 1 0 1603 0 1 30445
box 0 0 1 1
use contact_13  contact_13_118
timestamp 1643671299
transform 1 0 1589 0 1 30437
box 0 0 1 1
use contact_21  contact_21_118
timestamp 1643671299
transform 1 0 1593 0 1 30419
box 0 0 1 1
use contact_17  contact_17_119
timestamp 1643671299
transform 1 0 1603 0 1 30109
box 0 0 1 1
use contact_13  contact_13_119
timestamp 1643671299
transform 1 0 1589 0 1 30101
box 0 0 1 1
use contact_21  contact_21_119
timestamp 1643671299
transform 1 0 1593 0 1 30083
box 0 0 1 1
use contact_17  contact_17_120
timestamp 1643671299
transform 1 0 1603 0 1 29773
box 0 0 1 1
use contact_13  contact_13_120
timestamp 1643671299
transform 1 0 1589 0 1 29765
box 0 0 1 1
use contact_21  contact_21_120
timestamp 1643671299
transform 1 0 1593 0 1 29747
box 0 0 1 1
use contact_17  contact_17_121
timestamp 1643671299
transform 1 0 1603 0 1 29437
box 0 0 1 1
use contact_13  contact_13_121
timestamp 1643671299
transform 1 0 1589 0 1 29429
box 0 0 1 1
use contact_21  contact_21_121
timestamp 1643671299
transform 1 0 1593 0 1 29411
box 0 0 1 1
use contact_17  contact_17_122
timestamp 1643671299
transform 1 0 1603 0 1 29101
box 0 0 1 1
use contact_13  contact_13_122
timestamp 1643671299
transform 1 0 1589 0 1 29093
box 0 0 1 1
use contact_21  contact_21_122
timestamp 1643671299
transform 1 0 1593 0 1 29075
box 0 0 1 1
use contact_18  contact_18_25
timestamp 1643671299
transform 1 0 1588 0 1 28750
box 0 0 1 1
use contact_17  contact_17_123
timestamp 1643671299
transform 1 0 1603 0 1 28765
box 0 0 1 1
use contact_13  contact_13_123
timestamp 1643671299
transform 1 0 1589 0 1 28757
box 0 0 1 1
use contact_21  contact_21_123
timestamp 1643671299
transform 1 0 1593 0 1 28739
box 0 0 1 1
use contact_17  contact_17_124
timestamp 1643671299
transform 1 0 1603 0 1 28429
box 0 0 1 1
use contact_13  contact_13_124
timestamp 1643671299
transform 1 0 1589 0 1 28421
box 0 0 1 1
use contact_21  contact_21_124
timestamp 1643671299
transform 1 0 1593 0 1 28403
box 0 0 1 1
use contact_17  contact_17_125
timestamp 1643671299
transform 1 0 1603 0 1 28093
box 0 0 1 1
use contact_13  contact_13_125
timestamp 1643671299
transform 1 0 1589 0 1 28085
box 0 0 1 1
use contact_21  contact_21_125
timestamp 1643671299
transform 1 0 1593 0 1 28067
box 0 0 1 1
use contact_17  contact_17_126
timestamp 1643671299
transform 1 0 1603 0 1 27757
box 0 0 1 1
use contact_13  contact_13_126
timestamp 1643671299
transform 1 0 1589 0 1 27749
box 0 0 1 1
use contact_21  contact_21_126
timestamp 1643671299
transform 1 0 1593 0 1 27731
box 0 0 1 1
use contact_17  contact_17_127
timestamp 1643671299
transform 1 0 1603 0 1 27421
box 0 0 1 1
use contact_13  contact_13_127
timestamp 1643671299
transform 1 0 1589 0 1 27413
box 0 0 1 1
use contact_21  contact_21_127
timestamp 1643671299
transform 1 0 1593 0 1 27395
box 0 0 1 1
use contact_18  contact_18_26
timestamp 1643671299
transform 1 0 1588 0 1 27070
box 0 0 1 1
use contact_17  contact_17_128
timestamp 1643671299
transform 1 0 1603 0 1 27085
box 0 0 1 1
use contact_13  contact_13_128
timestamp 1643671299
transform 1 0 1589 0 1 27077
box 0 0 1 1
use contact_21  contact_21_128
timestamp 1643671299
transform 1 0 1593 0 1 27059
box 0 0 1 1
use contact_17  contact_17_129
timestamp 1643671299
transform 1 0 1603 0 1 26749
box 0 0 1 1
use contact_13  contact_13_129
timestamp 1643671299
transform 1 0 1589 0 1 26741
box 0 0 1 1
use contact_21  contact_21_129
timestamp 1643671299
transform 1 0 1593 0 1 26723
box 0 0 1 1
use contact_17  contact_17_130
timestamp 1643671299
transform 1 0 1603 0 1 26413
box 0 0 1 1
use contact_13  contact_13_130
timestamp 1643671299
transform 1 0 1589 0 1 26405
box 0 0 1 1
use contact_21  contact_21_130
timestamp 1643671299
transform 1 0 1593 0 1 26387
box 0 0 1 1
use contact_17  contact_17_131
timestamp 1643671299
transform 1 0 1603 0 1 26077
box 0 0 1 1
use contact_13  contact_13_131
timestamp 1643671299
transform 1 0 1589 0 1 26069
box 0 0 1 1
use contact_21  contact_21_131
timestamp 1643671299
transform 1 0 1593 0 1 26051
box 0 0 1 1
use contact_17  contact_17_132
timestamp 1643671299
transform 1 0 1603 0 1 25741
box 0 0 1 1
use contact_13  contact_13_132
timestamp 1643671299
transform 1 0 1589 0 1 25733
box 0 0 1 1
use contact_21  contact_21_132
timestamp 1643671299
transform 1 0 1593 0 1 25715
box 0 0 1 1
use contact_18  contact_18_27
timestamp 1643671299
transform 1 0 1588 0 1 25390
box 0 0 1 1
use contact_17  contact_17_133
timestamp 1643671299
transform 1 0 1603 0 1 25405
box 0 0 1 1
use contact_13  contact_13_133
timestamp 1643671299
transform 1 0 1589 0 1 25397
box 0 0 1 1
use contact_21  contact_21_133
timestamp 1643671299
transform 1 0 1593 0 1 25379
box 0 0 1 1
use contact_17  contact_17_134
timestamp 1643671299
transform 1 0 1603 0 1 25069
box 0 0 1 1
use contact_13  contact_13_134
timestamp 1643671299
transform 1 0 1589 0 1 25061
box 0 0 1 1
use contact_21  contact_21_134
timestamp 1643671299
transform 1 0 1593 0 1 25043
box 0 0 1 1
use contact_17  contact_17_135
timestamp 1643671299
transform 1 0 1603 0 1 24733
box 0 0 1 1
use contact_13  contact_13_135
timestamp 1643671299
transform 1 0 1589 0 1 24725
box 0 0 1 1
use contact_21  contact_21_135
timestamp 1643671299
transform 1 0 1593 0 1 24707
box 0 0 1 1
use contact_17  contact_17_136
timestamp 1643671299
transform 1 0 1603 0 1 24397
box 0 0 1 1
use contact_13  contact_13_136
timestamp 1643671299
transform 1 0 1589 0 1 24389
box 0 0 1 1
use contact_21  contact_21_136
timestamp 1643671299
transform 1 0 1593 0 1 24371
box 0 0 1 1
use contact_17  contact_17_137
timestamp 1643671299
transform 1 0 1603 0 1 24061
box 0 0 1 1
use contact_13  contact_13_137
timestamp 1643671299
transform 1 0 1589 0 1 24053
box 0 0 1 1
use contact_21  contact_21_137
timestamp 1643671299
transform 1 0 1593 0 1 24035
box 0 0 1 1
use contact_18  contact_18_28
timestamp 1643671299
transform 1 0 1588 0 1 23710
box 0 0 1 1
use contact_17  contact_17_138
timestamp 1643671299
transform 1 0 1603 0 1 23725
box 0 0 1 1
use contact_13  contact_13_138
timestamp 1643671299
transform 1 0 1589 0 1 23717
box 0 0 1 1
use contact_21  contact_21_138
timestamp 1643671299
transform 1 0 1593 0 1 23699
box 0 0 1 1
use contact_17  contact_17_139
timestamp 1643671299
transform 1 0 1603 0 1 23389
box 0 0 1 1
use contact_13  contact_13_139
timestamp 1643671299
transform 1 0 1589 0 1 23381
box 0 0 1 1
use contact_21  contact_21_139
timestamp 1643671299
transform 1 0 1593 0 1 23363
box 0 0 1 1
use contact_17  contact_17_140
timestamp 1643671299
transform 1 0 1603 0 1 23053
box 0 0 1 1
use contact_13  contact_13_140
timestamp 1643671299
transform 1 0 1589 0 1 23045
box 0 0 1 1
use contact_21  contact_21_140
timestamp 1643671299
transform 1 0 1593 0 1 23027
box 0 0 1 1
use contact_17  contact_17_141
timestamp 1643671299
transform 1 0 1603 0 1 22717
box 0 0 1 1
use contact_13  contact_13_141
timestamp 1643671299
transform 1 0 1589 0 1 22709
box 0 0 1 1
use contact_21  contact_21_141
timestamp 1643671299
transform 1 0 1593 0 1 22691
box 0 0 1 1
use contact_17  contact_17_142
timestamp 1643671299
transform 1 0 1603 0 1 22381
box 0 0 1 1
use contact_13  contact_13_142
timestamp 1643671299
transform 1 0 1589 0 1 22373
box 0 0 1 1
use contact_21  contact_21_142
timestamp 1643671299
transform 1 0 1593 0 1 22355
box 0 0 1 1
use contact_18  contact_18_29
timestamp 1643671299
transform 1 0 1588 0 1 22030
box 0 0 1 1
use contact_17  contact_17_143
timestamp 1643671299
transform 1 0 1603 0 1 22045
box 0 0 1 1
use contact_13  contact_13_143
timestamp 1643671299
transform 1 0 1589 0 1 22037
box 0 0 1 1
use contact_21  contact_21_143
timestamp 1643671299
transform 1 0 1593 0 1 22019
box 0 0 1 1
use contact_17  contact_17_144
timestamp 1643671299
transform 1 0 1603 0 1 21709
box 0 0 1 1
use contact_13  contact_13_144
timestamp 1643671299
transform 1 0 1589 0 1 21701
box 0 0 1 1
use contact_21  contact_21_144
timestamp 1643671299
transform 1 0 1593 0 1 21683
box 0 0 1 1
use contact_17  contact_17_145
timestamp 1643671299
transform 1 0 1603 0 1 21373
box 0 0 1 1
use contact_13  contact_13_145
timestamp 1643671299
transform 1 0 1589 0 1 21365
box 0 0 1 1
use contact_21  contact_21_145
timestamp 1643671299
transform 1 0 1593 0 1 21347
box 0 0 1 1
use contact_17  contact_17_146
timestamp 1643671299
transform 1 0 1603 0 1 21037
box 0 0 1 1
use contact_13  contact_13_146
timestamp 1643671299
transform 1 0 1589 0 1 21029
box 0 0 1 1
use contact_21  contact_21_146
timestamp 1643671299
transform 1 0 1593 0 1 21011
box 0 0 1 1
use contact_17  contact_17_147
timestamp 1643671299
transform 1 0 1603 0 1 20701
box 0 0 1 1
use contact_13  contact_13_147
timestamp 1643671299
transform 1 0 1589 0 1 20693
box 0 0 1 1
use contact_21  contact_21_147
timestamp 1643671299
transform 1 0 1593 0 1 20675
box 0 0 1 1
use contact_18  contact_18_30
timestamp 1643671299
transform 1 0 1588 0 1 20350
box 0 0 1 1
use contact_17  contact_17_148
timestamp 1643671299
transform 1 0 1603 0 1 20365
box 0 0 1 1
use contact_13  contact_13_148
timestamp 1643671299
transform 1 0 1589 0 1 20357
box 0 0 1 1
use contact_21  contact_21_148
timestamp 1643671299
transform 1 0 1593 0 1 20339
box 0 0 1 1
use contact_17  contact_17_149
timestamp 1643671299
transform 1 0 1603 0 1 20029
box 0 0 1 1
use contact_13  contact_13_149
timestamp 1643671299
transform 1 0 1589 0 1 20021
box 0 0 1 1
use contact_21  contact_21_149
timestamp 1643671299
transform 1 0 1593 0 1 20003
box 0 0 1 1
use contact_17  contact_17_150
timestamp 1643671299
transform 1 0 1603 0 1 19693
box 0 0 1 1
use contact_13  contact_13_150
timestamp 1643671299
transform 1 0 1589 0 1 19685
box 0 0 1 1
use contact_21  contact_21_150
timestamp 1643671299
transform 1 0 1593 0 1 19667
box 0 0 1 1
use contact_17  contact_17_151
timestamp 1643671299
transform 1 0 1603 0 1 19357
box 0 0 1 1
use contact_13  contact_13_151
timestamp 1643671299
transform 1 0 1589 0 1 19349
box 0 0 1 1
use contact_21  contact_21_151
timestamp 1643671299
transform 1 0 1593 0 1 19331
box 0 0 1 1
use contact_17  contact_17_152
timestamp 1643671299
transform 1 0 1603 0 1 19021
box 0 0 1 1
use contact_13  contact_13_152
timestamp 1643671299
transform 1 0 1589 0 1 19013
box 0 0 1 1
use contact_21  contact_21_152
timestamp 1643671299
transform 1 0 1593 0 1 18995
box 0 0 1 1
use contact_18  contact_18_31
timestamp 1643671299
transform 1 0 1588 0 1 18670
box 0 0 1 1
use contact_17  contact_17_153
timestamp 1643671299
transform 1 0 1603 0 1 18685
box 0 0 1 1
use contact_13  contact_13_153
timestamp 1643671299
transform 1 0 1589 0 1 18677
box 0 0 1 1
use contact_21  contact_21_153
timestamp 1643671299
transform 1 0 1593 0 1 18659
box 0 0 1 1
use contact_17  contact_17_154
timestamp 1643671299
transform 1 0 1603 0 1 18349
box 0 0 1 1
use contact_13  contact_13_154
timestamp 1643671299
transform 1 0 1589 0 1 18341
box 0 0 1 1
use contact_21  contact_21_154
timestamp 1643671299
transform 1 0 1593 0 1 18323
box 0 0 1 1
use contact_17  contact_17_155
timestamp 1643671299
transform 1 0 1603 0 1 18013
box 0 0 1 1
use contact_13  contact_13_155
timestamp 1643671299
transform 1 0 1589 0 1 18005
box 0 0 1 1
use contact_21  contact_21_155
timestamp 1643671299
transform 1 0 1593 0 1 17987
box 0 0 1 1
use contact_17  contact_17_156
timestamp 1643671299
transform 1 0 1603 0 1 17677
box 0 0 1 1
use contact_13  contact_13_156
timestamp 1643671299
transform 1 0 1589 0 1 17669
box 0 0 1 1
use contact_21  contact_21_156
timestamp 1643671299
transform 1 0 1593 0 1 17651
box 0 0 1 1
use contact_17  contact_17_157
timestamp 1643671299
transform 1 0 1603 0 1 17341
box 0 0 1 1
use contact_13  contact_13_157
timestamp 1643671299
transform 1 0 1589 0 1 17333
box 0 0 1 1
use contact_21  contact_21_157
timestamp 1643671299
transform 1 0 1593 0 1 17315
box 0 0 1 1
use contact_18  contact_18_32
timestamp 1643671299
transform 1 0 1588 0 1 16990
box 0 0 1 1
use contact_17  contact_17_158
timestamp 1643671299
transform 1 0 1603 0 1 17005
box 0 0 1 1
use contact_13  contact_13_158
timestamp 1643671299
transform 1 0 1589 0 1 16997
box 0 0 1 1
use contact_21  contact_21_158
timestamp 1643671299
transform 1 0 1593 0 1 16979
box 0 0 1 1
use contact_17  contact_17_159
timestamp 1643671299
transform 1 0 1603 0 1 16669
box 0 0 1 1
use contact_13  contact_13_159
timestamp 1643671299
transform 1 0 1589 0 1 16661
box 0 0 1 1
use contact_21  contact_21_159
timestamp 1643671299
transform 1 0 1593 0 1 16643
box 0 0 1 1
use contact_17  contact_17_160
timestamp 1643671299
transform 1 0 1603 0 1 16333
box 0 0 1 1
use contact_13  contact_13_160
timestamp 1643671299
transform 1 0 1589 0 1 16325
box 0 0 1 1
use contact_21  contact_21_160
timestamp 1643671299
transform 1 0 1593 0 1 16307
box 0 0 1 1
use contact_17  contact_17_161
timestamp 1643671299
transform 1 0 1603 0 1 15997
box 0 0 1 1
use contact_13  contact_13_161
timestamp 1643671299
transform 1 0 1589 0 1 15989
box 0 0 1 1
use contact_21  contact_21_161
timestamp 1643671299
transform 1 0 1593 0 1 15971
box 0 0 1 1
use contact_17  contact_17_162
timestamp 1643671299
transform 1 0 1603 0 1 15661
box 0 0 1 1
use contact_13  contact_13_162
timestamp 1643671299
transform 1 0 1589 0 1 15653
box 0 0 1 1
use contact_21  contact_21_162
timestamp 1643671299
transform 1 0 1593 0 1 15635
box 0 0 1 1
use contact_18  contact_18_33
timestamp 1643671299
transform 1 0 1588 0 1 15310
box 0 0 1 1
use contact_17  contact_17_163
timestamp 1643671299
transform 1 0 1603 0 1 15325
box 0 0 1 1
use contact_13  contact_13_163
timestamp 1643671299
transform 1 0 1589 0 1 15317
box 0 0 1 1
use contact_21  contact_21_163
timestamp 1643671299
transform 1 0 1593 0 1 15299
box 0 0 1 1
use contact_17  contact_17_164
timestamp 1643671299
transform 1 0 1603 0 1 14989
box 0 0 1 1
use contact_13  contact_13_164
timestamp 1643671299
transform 1 0 1589 0 1 14981
box 0 0 1 1
use contact_21  contact_21_164
timestamp 1643671299
transform 1 0 1593 0 1 14963
box 0 0 1 1
use contact_17  contact_17_165
timestamp 1643671299
transform 1 0 1603 0 1 14653
box 0 0 1 1
use contact_13  contact_13_165
timestamp 1643671299
transform 1 0 1589 0 1 14645
box 0 0 1 1
use contact_21  contact_21_165
timestamp 1643671299
transform 1 0 1593 0 1 14627
box 0 0 1 1
use contact_17  contact_17_166
timestamp 1643671299
transform 1 0 1603 0 1 14317
box 0 0 1 1
use contact_13  contact_13_166
timestamp 1643671299
transform 1 0 1589 0 1 14309
box 0 0 1 1
use contact_21  contact_21_166
timestamp 1643671299
transform 1 0 1593 0 1 14291
box 0 0 1 1
use contact_17  contact_17_167
timestamp 1643671299
transform 1 0 1603 0 1 13981
box 0 0 1 1
use contact_13  contact_13_167
timestamp 1643671299
transform 1 0 1589 0 1 13973
box 0 0 1 1
use contact_21  contact_21_167
timestamp 1643671299
transform 1 0 1593 0 1 13955
box 0 0 1 1
use contact_18  contact_18_34
timestamp 1643671299
transform 1 0 1588 0 1 13630
box 0 0 1 1
use contact_17  contact_17_168
timestamp 1643671299
transform 1 0 1603 0 1 13645
box 0 0 1 1
use contact_13  contact_13_168
timestamp 1643671299
transform 1 0 1589 0 1 13637
box 0 0 1 1
use contact_21  contact_21_168
timestamp 1643671299
transform 1 0 1593 0 1 13619
box 0 0 1 1
use contact_17  contact_17_169
timestamp 1643671299
transform 1 0 1603 0 1 13309
box 0 0 1 1
use contact_13  contact_13_169
timestamp 1643671299
transform 1 0 1589 0 1 13301
box 0 0 1 1
use contact_21  contact_21_169
timestamp 1643671299
transform 1 0 1593 0 1 13283
box 0 0 1 1
use contact_17  contact_17_170
timestamp 1643671299
transform 1 0 1603 0 1 12973
box 0 0 1 1
use contact_13  contact_13_170
timestamp 1643671299
transform 1 0 1589 0 1 12965
box 0 0 1 1
use contact_21  contact_21_170
timestamp 1643671299
transform 1 0 1593 0 1 12947
box 0 0 1 1
use contact_17  contact_17_171
timestamp 1643671299
transform 1 0 1603 0 1 12637
box 0 0 1 1
use contact_13  contact_13_171
timestamp 1643671299
transform 1 0 1589 0 1 12629
box 0 0 1 1
use contact_21  contact_21_171
timestamp 1643671299
transform 1 0 1593 0 1 12611
box 0 0 1 1
use contact_17  contact_17_172
timestamp 1643671299
transform 1 0 1603 0 1 12301
box 0 0 1 1
use contact_13  contact_13_172
timestamp 1643671299
transform 1 0 1589 0 1 12293
box 0 0 1 1
use contact_21  contact_21_172
timestamp 1643671299
transform 1 0 1593 0 1 12275
box 0 0 1 1
use contact_18  contact_18_35
timestamp 1643671299
transform 1 0 1588 0 1 11950
box 0 0 1 1
use contact_17  contact_17_173
timestamp 1643671299
transform 1 0 1603 0 1 11965
box 0 0 1 1
use contact_13  contact_13_173
timestamp 1643671299
transform 1 0 1589 0 1 11957
box 0 0 1 1
use contact_21  contact_21_173
timestamp 1643671299
transform 1 0 1593 0 1 11939
box 0 0 1 1
use contact_17  contact_17_174
timestamp 1643671299
transform 1 0 1603 0 1 11629
box 0 0 1 1
use contact_13  contact_13_174
timestamp 1643671299
transform 1 0 1589 0 1 11621
box 0 0 1 1
use contact_21  contact_21_174
timestamp 1643671299
transform 1 0 1593 0 1 11603
box 0 0 1 1
use contact_17  contact_17_175
timestamp 1643671299
transform 1 0 1603 0 1 11293
box 0 0 1 1
use contact_13  contact_13_175
timestamp 1643671299
transform 1 0 1589 0 1 11285
box 0 0 1 1
use contact_21  contact_21_175
timestamp 1643671299
transform 1 0 1593 0 1 11267
box 0 0 1 1
use contact_17  contact_17_176
timestamp 1643671299
transform 1 0 1603 0 1 10957
box 0 0 1 1
use contact_13  contact_13_176
timestamp 1643671299
transform 1 0 1589 0 1 10949
box 0 0 1 1
use contact_21  contact_21_176
timestamp 1643671299
transform 1 0 1593 0 1 10931
box 0 0 1 1
use contact_17  contact_17_177
timestamp 1643671299
transform 1 0 1603 0 1 10621
box 0 0 1 1
use contact_13  contact_13_177
timestamp 1643671299
transform 1 0 1589 0 1 10613
box 0 0 1 1
use contact_21  contact_21_177
timestamp 1643671299
transform 1 0 1593 0 1 10595
box 0 0 1 1
use contact_18  contact_18_36
timestamp 1643671299
transform 1 0 1588 0 1 10270
box 0 0 1 1
use contact_17  contact_17_178
timestamp 1643671299
transform 1 0 1603 0 1 10285
box 0 0 1 1
use contact_13  contact_13_178
timestamp 1643671299
transform 1 0 1589 0 1 10277
box 0 0 1 1
use contact_21  contact_21_178
timestamp 1643671299
transform 1 0 1593 0 1 10259
box 0 0 1 1
use contact_17  contact_17_179
timestamp 1643671299
transform 1 0 1603 0 1 9949
box 0 0 1 1
use contact_13  contact_13_179
timestamp 1643671299
transform 1 0 1589 0 1 9941
box 0 0 1 1
use contact_21  contact_21_179
timestamp 1643671299
transform 1 0 1593 0 1 9923
box 0 0 1 1
use contact_17  contact_17_180
timestamp 1643671299
transform 1 0 1603 0 1 9613
box 0 0 1 1
use contact_13  contact_13_180
timestamp 1643671299
transform 1 0 1589 0 1 9605
box 0 0 1 1
use contact_21  contact_21_180
timestamp 1643671299
transform 1 0 1593 0 1 9587
box 0 0 1 1
use contact_17  contact_17_181
timestamp 1643671299
transform 1 0 1603 0 1 9277
box 0 0 1 1
use contact_13  contact_13_181
timestamp 1643671299
transform 1 0 1589 0 1 9269
box 0 0 1 1
use contact_21  contact_21_181
timestamp 1643671299
transform 1 0 1593 0 1 9251
box 0 0 1 1
use contact_17  contact_17_182
timestamp 1643671299
transform 1 0 1603 0 1 8941
box 0 0 1 1
use contact_13  contact_13_182
timestamp 1643671299
transform 1 0 1589 0 1 8933
box 0 0 1 1
use contact_21  contact_21_182
timestamp 1643671299
transform 1 0 1593 0 1 8915
box 0 0 1 1
use contact_18  contact_18_37
timestamp 1643671299
transform 1 0 1588 0 1 8590
box 0 0 1 1
use contact_17  contact_17_183
timestamp 1643671299
transform 1 0 1603 0 1 8605
box 0 0 1 1
use contact_13  contact_13_183
timestamp 1643671299
transform 1 0 1589 0 1 8597
box 0 0 1 1
use contact_21  contact_21_183
timestamp 1643671299
transform 1 0 1593 0 1 8579
box 0 0 1 1
use contact_17  contact_17_184
timestamp 1643671299
transform 1 0 1603 0 1 8269
box 0 0 1 1
use contact_13  contact_13_184
timestamp 1643671299
transform 1 0 1589 0 1 8261
box 0 0 1 1
use contact_21  contact_21_184
timestamp 1643671299
transform 1 0 1593 0 1 8243
box 0 0 1 1
use contact_17  contact_17_185
timestamp 1643671299
transform 1 0 1603 0 1 7933
box 0 0 1 1
use contact_13  contact_13_185
timestamp 1643671299
transform 1 0 1589 0 1 7925
box 0 0 1 1
use contact_21  contact_21_185
timestamp 1643671299
transform 1 0 1593 0 1 7907
box 0 0 1 1
use contact_17  contact_17_186
timestamp 1643671299
transform 1 0 1603 0 1 7597
box 0 0 1 1
use contact_13  contact_13_186
timestamp 1643671299
transform 1 0 1589 0 1 7589
box 0 0 1 1
use contact_21  contact_21_186
timestamp 1643671299
transform 1 0 1593 0 1 7571
box 0 0 1 1
use contact_17  contact_17_187
timestamp 1643671299
transform 1 0 1603 0 1 7261
box 0 0 1 1
use contact_13  contact_13_187
timestamp 1643671299
transform 1 0 1589 0 1 7253
box 0 0 1 1
use contact_21  contact_21_187
timestamp 1643671299
transform 1 0 1593 0 1 7235
box 0 0 1 1
use contact_18  contact_18_38
timestamp 1643671299
transform 1 0 1588 0 1 6910
box 0 0 1 1
use contact_17  contact_17_188
timestamp 1643671299
transform 1 0 1603 0 1 6925
box 0 0 1 1
use contact_13  contact_13_188
timestamp 1643671299
transform 1 0 1589 0 1 6917
box 0 0 1 1
use contact_21  contact_21_188
timestamp 1643671299
transform 1 0 1593 0 1 6899
box 0 0 1 1
use contact_17  contact_17_189
timestamp 1643671299
transform 1 0 1603 0 1 6589
box 0 0 1 1
use contact_13  contact_13_189
timestamp 1643671299
transform 1 0 1589 0 1 6581
box 0 0 1 1
use contact_21  contact_21_189
timestamp 1643671299
transform 1 0 1593 0 1 6563
box 0 0 1 1
use contact_17  contact_17_190
timestamp 1643671299
transform 1 0 1603 0 1 6253
box 0 0 1 1
use contact_13  contact_13_190
timestamp 1643671299
transform 1 0 1589 0 1 6245
box 0 0 1 1
use contact_21  contact_21_190
timestamp 1643671299
transform 1 0 1593 0 1 6227
box 0 0 1 1
use contact_17  contact_17_191
timestamp 1643671299
transform 1 0 1603 0 1 5917
box 0 0 1 1
use contact_13  contact_13_191
timestamp 1643671299
transform 1 0 1589 0 1 5909
box 0 0 1 1
use contact_21  contact_21_191
timestamp 1643671299
transform 1 0 1593 0 1 5891
box 0 0 1 1
use contact_17  contact_17_192
timestamp 1643671299
transform 1 0 1603 0 1 5581
box 0 0 1 1
use contact_13  contact_13_192
timestamp 1643671299
transform 1 0 1589 0 1 5573
box 0 0 1 1
use contact_21  contact_21_192
timestamp 1643671299
transform 1 0 1593 0 1 5555
box 0 0 1 1
use contact_18  contact_18_39
timestamp 1643671299
transform 1 0 1588 0 1 5230
box 0 0 1 1
use contact_17  contact_17_193
timestamp 1643671299
transform 1 0 1603 0 1 5245
box 0 0 1 1
use contact_13  contact_13_193
timestamp 1643671299
transform 1 0 1589 0 1 5237
box 0 0 1 1
use contact_21  contact_21_193
timestamp 1643671299
transform 1 0 1593 0 1 5219
box 0 0 1 1
use contact_17  contact_17_194
timestamp 1643671299
transform 1 0 1603 0 1 4909
box 0 0 1 1
use contact_13  contact_13_194
timestamp 1643671299
transform 1 0 1589 0 1 4901
box 0 0 1 1
use contact_21  contact_21_194
timestamp 1643671299
transform 1 0 1593 0 1 4883
box 0 0 1 1
use contact_17  contact_17_195
timestamp 1643671299
transform 1 0 1603 0 1 4573
box 0 0 1 1
use contact_13  contact_13_195
timestamp 1643671299
transform 1 0 1589 0 1 4565
box 0 0 1 1
use contact_21  contact_21_195
timestamp 1643671299
transform 1 0 1593 0 1 4547
box 0 0 1 1
use contact_17  contact_17_196
timestamp 1643671299
transform 1 0 1603 0 1 4237
box 0 0 1 1
use contact_13  contact_13_196
timestamp 1643671299
transform 1 0 1589 0 1 4229
box 0 0 1 1
use contact_21  contact_21_196
timestamp 1643671299
transform 1 0 1593 0 1 4211
box 0 0 1 1
use contact_17  contact_17_197
timestamp 1643671299
transform 1 0 1603 0 1 3901
box 0 0 1 1
use contact_13  contact_13_197
timestamp 1643671299
transform 1 0 1589 0 1 3893
box 0 0 1 1
use contact_21  contact_21_197
timestamp 1643671299
transform 1 0 1593 0 1 3875
box 0 0 1 1
use contact_18  contact_18_40
timestamp 1643671299
transform 1 0 1588 0 1 3550
box 0 0 1 1
use contact_17  contact_17_198
timestamp 1643671299
transform 1 0 1603 0 1 3565
box 0 0 1 1
use contact_13  contact_13_198
timestamp 1643671299
transform 1 0 1589 0 1 3557
box 0 0 1 1
use contact_21  contact_21_198
timestamp 1643671299
transform 1 0 1593 0 1 3539
box 0 0 1 1
use contact_17  contact_17_199
timestamp 1643671299
transform 1 0 1603 0 1 3229
box 0 0 1 1
use contact_13  contact_13_199
timestamp 1643671299
transform 1 0 1589 0 1 3221
box 0 0 1 1
use contact_21  contact_21_199
timestamp 1643671299
transform 1 0 1593 0 1 3203
box 0 0 1 1
use contact_17  contact_17_200
timestamp 1643671299
transform 1 0 1603 0 1 2893
box 0 0 1 1
use contact_13  contact_13_200
timestamp 1643671299
transform 1 0 1589 0 1 2885
box 0 0 1 1
use contact_21  contact_21_200
timestamp 1643671299
transform 1 0 1593 0 1 2867
box 0 0 1 1
use contact_17  contact_17_201
timestamp 1643671299
transform 1 0 1603 0 1 2557
box 0 0 1 1
use contact_13  contact_13_201
timestamp 1643671299
transform 1 0 1589 0 1 2549
box 0 0 1 1
use contact_21  contact_21_201
timestamp 1643671299
transform 1 0 1593 0 1 2531
box 0 0 1 1
use contact_17  contact_17_202
timestamp 1643671299
transform 1 0 1603 0 1 2221
box 0 0 1 1
use contact_13  contact_13_202
timestamp 1643671299
transform 1 0 1589 0 1 2213
box 0 0 1 1
use contact_21  contact_21_202
timestamp 1643671299
transform 1 0 1593 0 1 2195
box 0 0 1 1
use contact_18  contact_18_41
timestamp 1643671299
transform 1 0 1588 0 1 1870
box 0 0 1 1
use contact_17  contact_17_203
timestamp 1643671299
transform 1 0 1603 0 1 1885
box 0 0 1 1
use contact_13  contact_13_203
timestamp 1643671299
transform 1 0 1589 0 1 1877
box 0 0 1 1
use contact_21  contact_21_203
timestamp 1643671299
transform 1 0 1593 0 1 1859
box 0 0 1 1
use contact_13  contact_13_204
timestamp 1643671299
transform 1 0 73493 0 1 36185
box 0 0 1 1
use contact_21  contact_21_204
timestamp 1643671299
transform 1 0 73497 0 1 36167
box 0 0 1 1
use contact_13  contact_13_205
timestamp 1643671299
transform 1 0 73157 0 1 36185
box 0 0 1 1
use contact_21  contact_21_205
timestamp 1643671299
transform 1 0 73161 0 1 36167
box 0 0 1 1
use contact_13  contact_13_206
timestamp 1643671299
transform 1 0 72821 0 1 36185
box 0 0 1 1
use contact_21  contact_21_206
timestamp 1643671299
transform 1 0 72825 0 1 36167
box 0 0 1 1
use contact_18  contact_18_42
timestamp 1643671299
transform 1 0 72484 0 1 36178
box 0 0 1 1
use contact_17  contact_17_204
timestamp 1643671299
transform 1 0 72499 0 1 36193
box 0 0 1 1
use contact_13  contact_13_207
timestamp 1643671299
transform 1 0 72485 0 1 36185
box 0 0 1 1
use contact_21  contact_21_207
timestamp 1643671299
transform 1 0 72489 0 1 36167
box 0 0 1 1
use contact_13  contact_13_208
timestamp 1643671299
transform 1 0 72149 0 1 36185
box 0 0 1 1
use contact_21  contact_21_208
timestamp 1643671299
transform 1 0 72153 0 1 36167
box 0 0 1 1
use contact_13  contact_13_209
timestamp 1643671299
transform 1 0 71813 0 1 36185
box 0 0 1 1
use contact_21  contact_21_209
timestamp 1643671299
transform 1 0 71817 0 1 36167
box 0 0 1 1
use contact_13  contact_13_210
timestamp 1643671299
transform 1 0 71477 0 1 36185
box 0 0 1 1
use contact_21  contact_21_210
timestamp 1643671299
transform 1 0 71481 0 1 36167
box 0 0 1 1
use contact_13  contact_13_211
timestamp 1643671299
transform 1 0 71141 0 1 36185
box 0 0 1 1
use contact_21  contact_21_211
timestamp 1643671299
transform 1 0 71145 0 1 36167
box 0 0 1 1
use contact_18  contact_18_43
timestamp 1643671299
transform 1 0 70804 0 1 36178
box 0 0 1 1
use contact_17  contact_17_205
timestamp 1643671299
transform 1 0 70819 0 1 36193
box 0 0 1 1
use contact_13  contact_13_212
timestamp 1643671299
transform 1 0 70805 0 1 36185
box 0 0 1 1
use contact_21  contact_21_212
timestamp 1643671299
transform 1 0 70809 0 1 36167
box 0 0 1 1
use contact_13  contact_13_213
timestamp 1643671299
transform 1 0 70469 0 1 36185
box 0 0 1 1
use contact_21  contact_21_213
timestamp 1643671299
transform 1 0 70473 0 1 36167
box 0 0 1 1
use contact_13  contact_13_214
timestamp 1643671299
transform 1 0 70133 0 1 36185
box 0 0 1 1
use contact_21  contact_21_214
timestamp 1643671299
transform 1 0 70137 0 1 36167
box 0 0 1 1
use contact_13  contact_13_215
timestamp 1643671299
transform 1 0 69797 0 1 36185
box 0 0 1 1
use contact_21  contact_21_215
timestamp 1643671299
transform 1 0 69801 0 1 36167
box 0 0 1 1
use contact_13  contact_13_216
timestamp 1643671299
transform 1 0 69461 0 1 36185
box 0 0 1 1
use contact_21  contact_21_216
timestamp 1643671299
transform 1 0 69465 0 1 36167
box 0 0 1 1
use contact_18  contact_18_44
timestamp 1643671299
transform 1 0 69124 0 1 36178
box 0 0 1 1
use contact_17  contact_17_206
timestamp 1643671299
transform 1 0 69139 0 1 36193
box 0 0 1 1
use contact_13  contact_13_217
timestamp 1643671299
transform 1 0 69125 0 1 36185
box 0 0 1 1
use contact_21  contact_21_217
timestamp 1643671299
transform 1 0 69129 0 1 36167
box 0 0 1 1
use contact_13  contact_13_218
timestamp 1643671299
transform 1 0 68789 0 1 36185
box 0 0 1 1
use contact_21  contact_21_218
timestamp 1643671299
transform 1 0 68793 0 1 36167
box 0 0 1 1
use contact_13  contact_13_219
timestamp 1643671299
transform 1 0 68453 0 1 36185
box 0 0 1 1
use contact_21  contact_21_219
timestamp 1643671299
transform 1 0 68457 0 1 36167
box 0 0 1 1
use contact_13  contact_13_220
timestamp 1643671299
transform 1 0 68117 0 1 36185
box 0 0 1 1
use contact_21  contact_21_220
timestamp 1643671299
transform 1 0 68121 0 1 36167
box 0 0 1 1
use contact_13  contact_13_221
timestamp 1643671299
transform 1 0 67781 0 1 36185
box 0 0 1 1
use contact_21  contact_21_221
timestamp 1643671299
transform 1 0 67785 0 1 36167
box 0 0 1 1
use contact_18  contact_18_45
timestamp 1643671299
transform 1 0 67444 0 1 36178
box 0 0 1 1
use contact_17  contact_17_207
timestamp 1643671299
transform 1 0 67459 0 1 36193
box 0 0 1 1
use contact_13  contact_13_222
timestamp 1643671299
transform 1 0 67445 0 1 36185
box 0 0 1 1
use contact_21  contact_21_222
timestamp 1643671299
transform 1 0 67449 0 1 36167
box 0 0 1 1
use contact_13  contact_13_223
timestamp 1643671299
transform 1 0 67109 0 1 36185
box 0 0 1 1
use contact_21  contact_21_223
timestamp 1643671299
transform 1 0 67113 0 1 36167
box 0 0 1 1
use contact_13  contact_13_224
timestamp 1643671299
transform 1 0 66773 0 1 36185
box 0 0 1 1
use contact_21  contact_21_224
timestamp 1643671299
transform 1 0 66777 0 1 36167
box 0 0 1 1
use contact_13  contact_13_225
timestamp 1643671299
transform 1 0 66437 0 1 36185
box 0 0 1 1
use contact_21  contact_21_225
timestamp 1643671299
transform 1 0 66441 0 1 36167
box 0 0 1 1
use contact_13  contact_13_226
timestamp 1643671299
transform 1 0 66101 0 1 36185
box 0 0 1 1
use contact_21  contact_21_226
timestamp 1643671299
transform 1 0 66105 0 1 36167
box 0 0 1 1
use contact_18  contact_18_46
timestamp 1643671299
transform 1 0 65764 0 1 36178
box 0 0 1 1
use contact_17  contact_17_208
timestamp 1643671299
transform 1 0 65779 0 1 36193
box 0 0 1 1
use contact_13  contact_13_227
timestamp 1643671299
transform 1 0 65765 0 1 36185
box 0 0 1 1
use contact_21  contact_21_227
timestamp 1643671299
transform 1 0 65769 0 1 36167
box 0 0 1 1
use contact_13  contact_13_228
timestamp 1643671299
transform 1 0 65429 0 1 36185
box 0 0 1 1
use contact_21  contact_21_228
timestamp 1643671299
transform 1 0 65433 0 1 36167
box 0 0 1 1
use contact_13  contact_13_229
timestamp 1643671299
transform 1 0 65093 0 1 36185
box 0 0 1 1
use contact_21  contact_21_229
timestamp 1643671299
transform 1 0 65097 0 1 36167
box 0 0 1 1
use contact_13  contact_13_230
timestamp 1643671299
transform 1 0 64757 0 1 36185
box 0 0 1 1
use contact_21  contact_21_230
timestamp 1643671299
transform 1 0 64761 0 1 36167
box 0 0 1 1
use contact_13  contact_13_231
timestamp 1643671299
transform 1 0 64421 0 1 36185
box 0 0 1 1
use contact_21  contact_21_231
timestamp 1643671299
transform 1 0 64425 0 1 36167
box 0 0 1 1
use contact_18  contact_18_47
timestamp 1643671299
transform 1 0 64084 0 1 36178
box 0 0 1 1
use contact_17  contact_17_209
timestamp 1643671299
transform 1 0 64099 0 1 36193
box 0 0 1 1
use contact_13  contact_13_232
timestamp 1643671299
transform 1 0 64085 0 1 36185
box 0 0 1 1
use contact_21  contact_21_232
timestamp 1643671299
transform 1 0 64089 0 1 36167
box 0 0 1 1
use contact_13  contact_13_233
timestamp 1643671299
transform 1 0 63749 0 1 36185
box 0 0 1 1
use contact_21  contact_21_233
timestamp 1643671299
transform 1 0 63753 0 1 36167
box 0 0 1 1
use contact_13  contact_13_234
timestamp 1643671299
transform 1 0 63413 0 1 36185
box 0 0 1 1
use contact_21  contact_21_234
timestamp 1643671299
transform 1 0 63417 0 1 36167
box 0 0 1 1
use contact_13  contact_13_235
timestamp 1643671299
transform 1 0 63077 0 1 36185
box 0 0 1 1
use contact_21  contact_21_235
timestamp 1643671299
transform 1 0 63081 0 1 36167
box 0 0 1 1
use contact_13  contact_13_236
timestamp 1643671299
transform 1 0 62741 0 1 36185
box 0 0 1 1
use contact_21  contact_21_236
timestamp 1643671299
transform 1 0 62745 0 1 36167
box 0 0 1 1
use contact_18  contact_18_48
timestamp 1643671299
transform 1 0 62404 0 1 36178
box 0 0 1 1
use contact_17  contact_17_210
timestamp 1643671299
transform 1 0 62419 0 1 36193
box 0 0 1 1
use contact_13  contact_13_237
timestamp 1643671299
transform 1 0 62405 0 1 36185
box 0 0 1 1
use contact_21  contact_21_237
timestamp 1643671299
transform 1 0 62409 0 1 36167
box 0 0 1 1
use contact_13  contact_13_238
timestamp 1643671299
transform 1 0 62069 0 1 36185
box 0 0 1 1
use contact_21  contact_21_238
timestamp 1643671299
transform 1 0 62073 0 1 36167
box 0 0 1 1
use contact_13  contact_13_239
timestamp 1643671299
transform 1 0 61733 0 1 36185
box 0 0 1 1
use contact_21  contact_21_239
timestamp 1643671299
transform 1 0 61737 0 1 36167
box 0 0 1 1
use contact_13  contact_13_240
timestamp 1643671299
transform 1 0 61397 0 1 36185
box 0 0 1 1
use contact_21  contact_21_240
timestamp 1643671299
transform 1 0 61401 0 1 36167
box 0 0 1 1
use contact_13  contact_13_241
timestamp 1643671299
transform 1 0 61061 0 1 36185
box 0 0 1 1
use contact_21  contact_21_241
timestamp 1643671299
transform 1 0 61065 0 1 36167
box 0 0 1 1
use contact_18  contact_18_49
timestamp 1643671299
transform 1 0 60724 0 1 36178
box 0 0 1 1
use contact_17  contact_17_211
timestamp 1643671299
transform 1 0 60739 0 1 36193
box 0 0 1 1
use contact_13  contact_13_242
timestamp 1643671299
transform 1 0 60725 0 1 36185
box 0 0 1 1
use contact_21  contact_21_242
timestamp 1643671299
transform 1 0 60729 0 1 36167
box 0 0 1 1
use contact_13  contact_13_243
timestamp 1643671299
transform 1 0 60389 0 1 36185
box 0 0 1 1
use contact_21  contact_21_243
timestamp 1643671299
transform 1 0 60393 0 1 36167
box 0 0 1 1
use contact_13  contact_13_244
timestamp 1643671299
transform 1 0 60053 0 1 36185
box 0 0 1 1
use contact_21  contact_21_244
timestamp 1643671299
transform 1 0 60057 0 1 36167
box 0 0 1 1
use contact_13  contact_13_245
timestamp 1643671299
transform 1 0 59717 0 1 36185
box 0 0 1 1
use contact_21  contact_21_245
timestamp 1643671299
transform 1 0 59721 0 1 36167
box 0 0 1 1
use contact_13  contact_13_246
timestamp 1643671299
transform 1 0 59381 0 1 36185
box 0 0 1 1
use contact_21  contact_21_246
timestamp 1643671299
transform 1 0 59385 0 1 36167
box 0 0 1 1
use contact_18  contact_18_50
timestamp 1643671299
transform 1 0 59044 0 1 36178
box 0 0 1 1
use contact_17  contact_17_212
timestamp 1643671299
transform 1 0 59059 0 1 36193
box 0 0 1 1
use contact_13  contact_13_247
timestamp 1643671299
transform 1 0 59045 0 1 36185
box 0 0 1 1
use contact_21  contact_21_247
timestamp 1643671299
transform 1 0 59049 0 1 36167
box 0 0 1 1
use contact_13  contact_13_248
timestamp 1643671299
transform 1 0 58709 0 1 36185
box 0 0 1 1
use contact_21  contact_21_248
timestamp 1643671299
transform 1 0 58713 0 1 36167
box 0 0 1 1
use contact_13  contact_13_249
timestamp 1643671299
transform 1 0 58373 0 1 36185
box 0 0 1 1
use contact_21  contact_21_249
timestamp 1643671299
transform 1 0 58377 0 1 36167
box 0 0 1 1
use contact_13  contact_13_250
timestamp 1643671299
transform 1 0 58037 0 1 36185
box 0 0 1 1
use contact_21  contact_21_250
timestamp 1643671299
transform 1 0 58041 0 1 36167
box 0 0 1 1
use contact_13  contact_13_251
timestamp 1643671299
transform 1 0 57701 0 1 36185
box 0 0 1 1
use contact_21  contact_21_251
timestamp 1643671299
transform 1 0 57705 0 1 36167
box 0 0 1 1
use contact_18  contact_18_51
timestamp 1643671299
transform 1 0 57364 0 1 36178
box 0 0 1 1
use contact_17  contact_17_213
timestamp 1643671299
transform 1 0 57379 0 1 36193
box 0 0 1 1
use contact_13  contact_13_252
timestamp 1643671299
transform 1 0 57365 0 1 36185
box 0 0 1 1
use contact_21  contact_21_252
timestamp 1643671299
transform 1 0 57369 0 1 36167
box 0 0 1 1
use contact_13  contact_13_253
timestamp 1643671299
transform 1 0 57029 0 1 36185
box 0 0 1 1
use contact_21  contact_21_253
timestamp 1643671299
transform 1 0 57033 0 1 36167
box 0 0 1 1
use contact_13  contact_13_254
timestamp 1643671299
transform 1 0 56693 0 1 36185
box 0 0 1 1
use contact_21  contact_21_254
timestamp 1643671299
transform 1 0 56697 0 1 36167
box 0 0 1 1
use contact_13  contact_13_255
timestamp 1643671299
transform 1 0 56357 0 1 36185
box 0 0 1 1
use contact_21  contact_21_255
timestamp 1643671299
transform 1 0 56361 0 1 36167
box 0 0 1 1
use contact_13  contact_13_256
timestamp 1643671299
transform 1 0 56021 0 1 36185
box 0 0 1 1
use contact_21  contact_21_256
timestamp 1643671299
transform 1 0 56025 0 1 36167
box 0 0 1 1
use contact_18  contact_18_52
timestamp 1643671299
transform 1 0 55684 0 1 36178
box 0 0 1 1
use contact_17  contact_17_214
timestamp 1643671299
transform 1 0 55699 0 1 36193
box 0 0 1 1
use contact_13  contact_13_257
timestamp 1643671299
transform 1 0 55685 0 1 36185
box 0 0 1 1
use contact_21  contact_21_257
timestamp 1643671299
transform 1 0 55689 0 1 36167
box 0 0 1 1
use contact_13  contact_13_258
timestamp 1643671299
transform 1 0 55349 0 1 36185
box 0 0 1 1
use contact_21  contact_21_258
timestamp 1643671299
transform 1 0 55353 0 1 36167
box 0 0 1 1
use contact_13  contact_13_259
timestamp 1643671299
transform 1 0 55013 0 1 36185
box 0 0 1 1
use contact_21  contact_21_259
timestamp 1643671299
transform 1 0 55017 0 1 36167
box 0 0 1 1
use contact_13  contact_13_260
timestamp 1643671299
transform 1 0 54677 0 1 36185
box 0 0 1 1
use contact_21  contact_21_260
timestamp 1643671299
transform 1 0 54681 0 1 36167
box 0 0 1 1
use contact_13  contact_13_261
timestamp 1643671299
transform 1 0 54341 0 1 36185
box 0 0 1 1
use contact_21  contact_21_261
timestamp 1643671299
transform 1 0 54345 0 1 36167
box 0 0 1 1
use contact_18  contact_18_53
timestamp 1643671299
transform 1 0 54004 0 1 36178
box 0 0 1 1
use contact_17  contact_17_215
timestamp 1643671299
transform 1 0 54019 0 1 36193
box 0 0 1 1
use contact_13  contact_13_262
timestamp 1643671299
transform 1 0 54005 0 1 36185
box 0 0 1 1
use contact_21  contact_21_262
timestamp 1643671299
transform 1 0 54009 0 1 36167
box 0 0 1 1
use contact_13  contact_13_263
timestamp 1643671299
transform 1 0 53669 0 1 36185
box 0 0 1 1
use contact_21  contact_21_263
timestamp 1643671299
transform 1 0 53673 0 1 36167
box 0 0 1 1
use contact_13  contact_13_264
timestamp 1643671299
transform 1 0 53333 0 1 36185
box 0 0 1 1
use contact_21  contact_21_264
timestamp 1643671299
transform 1 0 53337 0 1 36167
box 0 0 1 1
use contact_13  contact_13_265
timestamp 1643671299
transform 1 0 52997 0 1 36185
box 0 0 1 1
use contact_21  contact_21_265
timestamp 1643671299
transform 1 0 53001 0 1 36167
box 0 0 1 1
use contact_13  contact_13_266
timestamp 1643671299
transform 1 0 52661 0 1 36185
box 0 0 1 1
use contact_21  contact_21_266
timestamp 1643671299
transform 1 0 52665 0 1 36167
box 0 0 1 1
use contact_18  contact_18_54
timestamp 1643671299
transform 1 0 52324 0 1 36178
box 0 0 1 1
use contact_17  contact_17_216
timestamp 1643671299
transform 1 0 52339 0 1 36193
box 0 0 1 1
use contact_13  contact_13_267
timestamp 1643671299
transform 1 0 52325 0 1 36185
box 0 0 1 1
use contact_21  contact_21_267
timestamp 1643671299
transform 1 0 52329 0 1 36167
box 0 0 1 1
use contact_13  contact_13_268
timestamp 1643671299
transform 1 0 51989 0 1 36185
box 0 0 1 1
use contact_21  contact_21_268
timestamp 1643671299
transform 1 0 51993 0 1 36167
box 0 0 1 1
use contact_13  contact_13_269
timestamp 1643671299
transform 1 0 51653 0 1 36185
box 0 0 1 1
use contact_21  contact_21_269
timestamp 1643671299
transform 1 0 51657 0 1 36167
box 0 0 1 1
use contact_13  contact_13_270
timestamp 1643671299
transform 1 0 51317 0 1 36185
box 0 0 1 1
use contact_21  contact_21_270
timestamp 1643671299
transform 1 0 51321 0 1 36167
box 0 0 1 1
use contact_13  contact_13_271
timestamp 1643671299
transform 1 0 50981 0 1 36185
box 0 0 1 1
use contact_21  contact_21_271
timestamp 1643671299
transform 1 0 50985 0 1 36167
box 0 0 1 1
use contact_18  contact_18_55
timestamp 1643671299
transform 1 0 50644 0 1 36178
box 0 0 1 1
use contact_17  contact_17_217
timestamp 1643671299
transform 1 0 50659 0 1 36193
box 0 0 1 1
use contact_13  contact_13_272
timestamp 1643671299
transform 1 0 50645 0 1 36185
box 0 0 1 1
use contact_21  contact_21_272
timestamp 1643671299
transform 1 0 50649 0 1 36167
box 0 0 1 1
use contact_13  contact_13_273
timestamp 1643671299
transform 1 0 50309 0 1 36185
box 0 0 1 1
use contact_21  contact_21_273
timestamp 1643671299
transform 1 0 50313 0 1 36167
box 0 0 1 1
use contact_13  contact_13_274
timestamp 1643671299
transform 1 0 49973 0 1 36185
box 0 0 1 1
use contact_21  contact_21_274
timestamp 1643671299
transform 1 0 49977 0 1 36167
box 0 0 1 1
use contact_13  contact_13_275
timestamp 1643671299
transform 1 0 49637 0 1 36185
box 0 0 1 1
use contact_21  contact_21_275
timestamp 1643671299
transform 1 0 49641 0 1 36167
box 0 0 1 1
use contact_13  contact_13_276
timestamp 1643671299
transform 1 0 49301 0 1 36185
box 0 0 1 1
use contact_21  contact_21_276
timestamp 1643671299
transform 1 0 49305 0 1 36167
box 0 0 1 1
use contact_18  contact_18_56
timestamp 1643671299
transform 1 0 48964 0 1 36178
box 0 0 1 1
use contact_17  contact_17_218
timestamp 1643671299
transform 1 0 48979 0 1 36193
box 0 0 1 1
use contact_13  contact_13_277
timestamp 1643671299
transform 1 0 48965 0 1 36185
box 0 0 1 1
use contact_21  contact_21_277
timestamp 1643671299
transform 1 0 48969 0 1 36167
box 0 0 1 1
use contact_13  contact_13_278
timestamp 1643671299
transform 1 0 48629 0 1 36185
box 0 0 1 1
use contact_21  contact_21_278
timestamp 1643671299
transform 1 0 48633 0 1 36167
box 0 0 1 1
use contact_13  contact_13_279
timestamp 1643671299
transform 1 0 48293 0 1 36185
box 0 0 1 1
use contact_21  contact_21_279
timestamp 1643671299
transform 1 0 48297 0 1 36167
box 0 0 1 1
use contact_13  contact_13_280
timestamp 1643671299
transform 1 0 47957 0 1 36185
box 0 0 1 1
use contact_21  contact_21_280
timestamp 1643671299
transform 1 0 47961 0 1 36167
box 0 0 1 1
use contact_13  contact_13_281
timestamp 1643671299
transform 1 0 47621 0 1 36185
box 0 0 1 1
use contact_21  contact_21_281
timestamp 1643671299
transform 1 0 47625 0 1 36167
box 0 0 1 1
use contact_18  contact_18_57
timestamp 1643671299
transform 1 0 47284 0 1 36178
box 0 0 1 1
use contact_17  contact_17_219
timestamp 1643671299
transform 1 0 47299 0 1 36193
box 0 0 1 1
use contact_13  contact_13_282
timestamp 1643671299
transform 1 0 47285 0 1 36185
box 0 0 1 1
use contact_21  contact_21_282
timestamp 1643671299
transform 1 0 47289 0 1 36167
box 0 0 1 1
use contact_13  contact_13_283
timestamp 1643671299
transform 1 0 46949 0 1 36185
box 0 0 1 1
use contact_21  contact_21_283
timestamp 1643671299
transform 1 0 46953 0 1 36167
box 0 0 1 1
use contact_13  contact_13_284
timestamp 1643671299
transform 1 0 46613 0 1 36185
box 0 0 1 1
use contact_21  contact_21_284
timestamp 1643671299
transform 1 0 46617 0 1 36167
box 0 0 1 1
use contact_13  contact_13_285
timestamp 1643671299
transform 1 0 46277 0 1 36185
box 0 0 1 1
use contact_21  contact_21_285
timestamp 1643671299
transform 1 0 46281 0 1 36167
box 0 0 1 1
use contact_13  contact_13_286
timestamp 1643671299
transform 1 0 45941 0 1 36185
box 0 0 1 1
use contact_21  contact_21_286
timestamp 1643671299
transform 1 0 45945 0 1 36167
box 0 0 1 1
use contact_18  contact_18_58
timestamp 1643671299
transform 1 0 45604 0 1 36178
box 0 0 1 1
use contact_17  contact_17_220
timestamp 1643671299
transform 1 0 45619 0 1 36193
box 0 0 1 1
use contact_13  contact_13_287
timestamp 1643671299
transform 1 0 45605 0 1 36185
box 0 0 1 1
use contact_21  contact_21_287
timestamp 1643671299
transform 1 0 45609 0 1 36167
box 0 0 1 1
use contact_13  contact_13_288
timestamp 1643671299
transform 1 0 45269 0 1 36185
box 0 0 1 1
use contact_21  contact_21_288
timestamp 1643671299
transform 1 0 45273 0 1 36167
box 0 0 1 1
use contact_13  contact_13_289
timestamp 1643671299
transform 1 0 44933 0 1 36185
box 0 0 1 1
use contact_21  contact_21_289
timestamp 1643671299
transform 1 0 44937 0 1 36167
box 0 0 1 1
use contact_13  contact_13_290
timestamp 1643671299
transform 1 0 44597 0 1 36185
box 0 0 1 1
use contact_21  contact_21_290
timestamp 1643671299
transform 1 0 44601 0 1 36167
box 0 0 1 1
use contact_13  contact_13_291
timestamp 1643671299
transform 1 0 44261 0 1 36185
box 0 0 1 1
use contact_21  contact_21_291
timestamp 1643671299
transform 1 0 44265 0 1 36167
box 0 0 1 1
use contact_18  contact_18_59
timestamp 1643671299
transform 1 0 43924 0 1 36178
box 0 0 1 1
use contact_17  contact_17_221
timestamp 1643671299
transform 1 0 43939 0 1 36193
box 0 0 1 1
use contact_13  contact_13_292
timestamp 1643671299
transform 1 0 43925 0 1 36185
box 0 0 1 1
use contact_21  contact_21_292
timestamp 1643671299
transform 1 0 43929 0 1 36167
box 0 0 1 1
use contact_13  contact_13_293
timestamp 1643671299
transform 1 0 43589 0 1 36185
box 0 0 1 1
use contact_21  contact_21_293
timestamp 1643671299
transform 1 0 43593 0 1 36167
box 0 0 1 1
use contact_13  contact_13_294
timestamp 1643671299
transform 1 0 43253 0 1 36185
box 0 0 1 1
use contact_21  contact_21_294
timestamp 1643671299
transform 1 0 43257 0 1 36167
box 0 0 1 1
use contact_13  contact_13_295
timestamp 1643671299
transform 1 0 42917 0 1 36185
box 0 0 1 1
use contact_21  contact_21_295
timestamp 1643671299
transform 1 0 42921 0 1 36167
box 0 0 1 1
use contact_13  contact_13_296
timestamp 1643671299
transform 1 0 42581 0 1 36185
box 0 0 1 1
use contact_21  contact_21_296
timestamp 1643671299
transform 1 0 42585 0 1 36167
box 0 0 1 1
use contact_18  contact_18_60
timestamp 1643671299
transform 1 0 42244 0 1 36178
box 0 0 1 1
use contact_17  contact_17_222
timestamp 1643671299
transform 1 0 42259 0 1 36193
box 0 0 1 1
use contact_13  contact_13_297
timestamp 1643671299
transform 1 0 42245 0 1 36185
box 0 0 1 1
use contact_21  contact_21_297
timestamp 1643671299
transform 1 0 42249 0 1 36167
box 0 0 1 1
use contact_13  contact_13_298
timestamp 1643671299
transform 1 0 41909 0 1 36185
box 0 0 1 1
use contact_21  contact_21_298
timestamp 1643671299
transform 1 0 41913 0 1 36167
box 0 0 1 1
use contact_13  contact_13_299
timestamp 1643671299
transform 1 0 41573 0 1 36185
box 0 0 1 1
use contact_21  contact_21_299
timestamp 1643671299
transform 1 0 41577 0 1 36167
box 0 0 1 1
use contact_13  contact_13_300
timestamp 1643671299
transform 1 0 41237 0 1 36185
box 0 0 1 1
use contact_21  contact_21_300
timestamp 1643671299
transform 1 0 41241 0 1 36167
box 0 0 1 1
use contact_13  contact_13_301
timestamp 1643671299
transform 1 0 40901 0 1 36185
box 0 0 1 1
use contact_21  contact_21_301
timestamp 1643671299
transform 1 0 40905 0 1 36167
box 0 0 1 1
use contact_18  contact_18_61
timestamp 1643671299
transform 1 0 40564 0 1 36178
box 0 0 1 1
use contact_17  contact_17_223
timestamp 1643671299
transform 1 0 40579 0 1 36193
box 0 0 1 1
use contact_13  contact_13_302
timestamp 1643671299
transform 1 0 40565 0 1 36185
box 0 0 1 1
use contact_21  contact_21_302
timestamp 1643671299
transform 1 0 40569 0 1 36167
box 0 0 1 1
use contact_13  contact_13_303
timestamp 1643671299
transform 1 0 40229 0 1 36185
box 0 0 1 1
use contact_21  contact_21_303
timestamp 1643671299
transform 1 0 40233 0 1 36167
box 0 0 1 1
use contact_13  contact_13_304
timestamp 1643671299
transform 1 0 39893 0 1 36185
box 0 0 1 1
use contact_21  contact_21_304
timestamp 1643671299
transform 1 0 39897 0 1 36167
box 0 0 1 1
use contact_13  contact_13_305
timestamp 1643671299
transform 1 0 39557 0 1 36185
box 0 0 1 1
use contact_21  contact_21_305
timestamp 1643671299
transform 1 0 39561 0 1 36167
box 0 0 1 1
use contact_13  contact_13_306
timestamp 1643671299
transform 1 0 39221 0 1 36185
box 0 0 1 1
use contact_21  contact_21_306
timestamp 1643671299
transform 1 0 39225 0 1 36167
box 0 0 1 1
use contact_18  contact_18_62
timestamp 1643671299
transform 1 0 38884 0 1 36178
box 0 0 1 1
use contact_17  contact_17_224
timestamp 1643671299
transform 1 0 38899 0 1 36193
box 0 0 1 1
use contact_13  contact_13_307
timestamp 1643671299
transform 1 0 38885 0 1 36185
box 0 0 1 1
use contact_21  contact_21_307
timestamp 1643671299
transform 1 0 38889 0 1 36167
box 0 0 1 1
use contact_13  contact_13_308
timestamp 1643671299
transform 1 0 38549 0 1 36185
box 0 0 1 1
use contact_21  contact_21_308
timestamp 1643671299
transform 1 0 38553 0 1 36167
box 0 0 1 1
use contact_13  contact_13_309
timestamp 1643671299
transform 1 0 38213 0 1 36185
box 0 0 1 1
use contact_21  contact_21_309
timestamp 1643671299
transform 1 0 38217 0 1 36167
box 0 0 1 1
use contact_13  contact_13_310
timestamp 1643671299
transform 1 0 37877 0 1 36185
box 0 0 1 1
use contact_21  contact_21_310
timestamp 1643671299
transform 1 0 37881 0 1 36167
box 0 0 1 1
use contact_13  contact_13_311
timestamp 1643671299
transform 1 0 37541 0 1 36185
box 0 0 1 1
use contact_21  contact_21_311
timestamp 1643671299
transform 1 0 37545 0 1 36167
box 0 0 1 1
use contact_18  contact_18_63
timestamp 1643671299
transform 1 0 37204 0 1 36178
box 0 0 1 1
use contact_17  contact_17_225
timestamp 1643671299
transform 1 0 37219 0 1 36193
box 0 0 1 1
use contact_13  contact_13_312
timestamp 1643671299
transform 1 0 37205 0 1 36185
box 0 0 1 1
use contact_21  contact_21_312
timestamp 1643671299
transform 1 0 37209 0 1 36167
box 0 0 1 1
use contact_13  contact_13_313
timestamp 1643671299
transform 1 0 36869 0 1 36185
box 0 0 1 1
use contact_21  contact_21_313
timestamp 1643671299
transform 1 0 36873 0 1 36167
box 0 0 1 1
use contact_13  contact_13_314
timestamp 1643671299
transform 1 0 36533 0 1 36185
box 0 0 1 1
use contact_21  contact_21_314
timestamp 1643671299
transform 1 0 36537 0 1 36167
box 0 0 1 1
use contact_13  contact_13_315
timestamp 1643671299
transform 1 0 36197 0 1 36185
box 0 0 1 1
use contact_21  contact_21_315
timestamp 1643671299
transform 1 0 36201 0 1 36167
box 0 0 1 1
use contact_13  contact_13_316
timestamp 1643671299
transform 1 0 35861 0 1 36185
box 0 0 1 1
use contact_21  contact_21_316
timestamp 1643671299
transform 1 0 35865 0 1 36167
box 0 0 1 1
use contact_18  contact_18_64
timestamp 1643671299
transform 1 0 35524 0 1 36178
box 0 0 1 1
use contact_17  contact_17_226
timestamp 1643671299
transform 1 0 35539 0 1 36193
box 0 0 1 1
use contact_13  contact_13_317
timestamp 1643671299
transform 1 0 35525 0 1 36185
box 0 0 1 1
use contact_21  contact_21_317
timestamp 1643671299
transform 1 0 35529 0 1 36167
box 0 0 1 1
use contact_13  contact_13_318
timestamp 1643671299
transform 1 0 35189 0 1 36185
box 0 0 1 1
use contact_21  contact_21_318
timestamp 1643671299
transform 1 0 35193 0 1 36167
box 0 0 1 1
use contact_13  contact_13_319
timestamp 1643671299
transform 1 0 34853 0 1 36185
box 0 0 1 1
use contact_21  contact_21_319
timestamp 1643671299
transform 1 0 34857 0 1 36167
box 0 0 1 1
use contact_13  contact_13_320
timestamp 1643671299
transform 1 0 34517 0 1 36185
box 0 0 1 1
use contact_21  contact_21_320
timestamp 1643671299
transform 1 0 34521 0 1 36167
box 0 0 1 1
use contact_13  contact_13_321
timestamp 1643671299
transform 1 0 34181 0 1 36185
box 0 0 1 1
use contact_21  contact_21_321
timestamp 1643671299
transform 1 0 34185 0 1 36167
box 0 0 1 1
use contact_18  contact_18_65
timestamp 1643671299
transform 1 0 33844 0 1 36178
box 0 0 1 1
use contact_17  contact_17_227
timestamp 1643671299
transform 1 0 33859 0 1 36193
box 0 0 1 1
use contact_13  contact_13_322
timestamp 1643671299
transform 1 0 33845 0 1 36185
box 0 0 1 1
use contact_21  contact_21_322
timestamp 1643671299
transform 1 0 33849 0 1 36167
box 0 0 1 1
use contact_13  contact_13_323
timestamp 1643671299
transform 1 0 33509 0 1 36185
box 0 0 1 1
use contact_21  contact_21_323
timestamp 1643671299
transform 1 0 33513 0 1 36167
box 0 0 1 1
use contact_13  contact_13_324
timestamp 1643671299
transform 1 0 33173 0 1 36185
box 0 0 1 1
use contact_21  contact_21_324
timestamp 1643671299
transform 1 0 33177 0 1 36167
box 0 0 1 1
use contact_13  contact_13_325
timestamp 1643671299
transform 1 0 32837 0 1 36185
box 0 0 1 1
use contact_21  contact_21_325
timestamp 1643671299
transform 1 0 32841 0 1 36167
box 0 0 1 1
use contact_13  contact_13_326
timestamp 1643671299
transform 1 0 32501 0 1 36185
box 0 0 1 1
use contact_21  contact_21_326
timestamp 1643671299
transform 1 0 32505 0 1 36167
box 0 0 1 1
use contact_18  contact_18_66
timestamp 1643671299
transform 1 0 32164 0 1 36178
box 0 0 1 1
use contact_17  contact_17_228
timestamp 1643671299
transform 1 0 32179 0 1 36193
box 0 0 1 1
use contact_13  contact_13_327
timestamp 1643671299
transform 1 0 32165 0 1 36185
box 0 0 1 1
use contact_21  contact_21_327
timestamp 1643671299
transform 1 0 32169 0 1 36167
box 0 0 1 1
use contact_13  contact_13_328
timestamp 1643671299
transform 1 0 31829 0 1 36185
box 0 0 1 1
use contact_21  contact_21_328
timestamp 1643671299
transform 1 0 31833 0 1 36167
box 0 0 1 1
use contact_13  contact_13_329
timestamp 1643671299
transform 1 0 31493 0 1 36185
box 0 0 1 1
use contact_21  contact_21_329
timestamp 1643671299
transform 1 0 31497 0 1 36167
box 0 0 1 1
use contact_13  contact_13_330
timestamp 1643671299
transform 1 0 31157 0 1 36185
box 0 0 1 1
use contact_21  contact_21_330
timestamp 1643671299
transform 1 0 31161 0 1 36167
box 0 0 1 1
use contact_13  contact_13_331
timestamp 1643671299
transform 1 0 30821 0 1 36185
box 0 0 1 1
use contact_21  contact_21_331
timestamp 1643671299
transform 1 0 30825 0 1 36167
box 0 0 1 1
use contact_18  contact_18_67
timestamp 1643671299
transform 1 0 30484 0 1 36178
box 0 0 1 1
use contact_17  contact_17_229
timestamp 1643671299
transform 1 0 30499 0 1 36193
box 0 0 1 1
use contact_13  contact_13_332
timestamp 1643671299
transform 1 0 30485 0 1 36185
box 0 0 1 1
use contact_21  contact_21_332
timestamp 1643671299
transform 1 0 30489 0 1 36167
box 0 0 1 1
use contact_13  contact_13_333
timestamp 1643671299
transform 1 0 30149 0 1 36185
box 0 0 1 1
use contact_21  contact_21_333
timestamp 1643671299
transform 1 0 30153 0 1 36167
box 0 0 1 1
use contact_13  contact_13_334
timestamp 1643671299
transform 1 0 29813 0 1 36185
box 0 0 1 1
use contact_21  contact_21_334
timestamp 1643671299
transform 1 0 29817 0 1 36167
box 0 0 1 1
use contact_13  contact_13_335
timestamp 1643671299
transform 1 0 29477 0 1 36185
box 0 0 1 1
use contact_21  contact_21_335
timestamp 1643671299
transform 1 0 29481 0 1 36167
box 0 0 1 1
use contact_13  contact_13_336
timestamp 1643671299
transform 1 0 29141 0 1 36185
box 0 0 1 1
use contact_21  contact_21_336
timestamp 1643671299
transform 1 0 29145 0 1 36167
box 0 0 1 1
use contact_18  contact_18_68
timestamp 1643671299
transform 1 0 28804 0 1 36178
box 0 0 1 1
use contact_17  contact_17_230
timestamp 1643671299
transform 1 0 28819 0 1 36193
box 0 0 1 1
use contact_13  contact_13_337
timestamp 1643671299
transform 1 0 28805 0 1 36185
box 0 0 1 1
use contact_21  contact_21_337
timestamp 1643671299
transform 1 0 28809 0 1 36167
box 0 0 1 1
use contact_13  contact_13_338
timestamp 1643671299
transform 1 0 28469 0 1 36185
box 0 0 1 1
use contact_21  contact_21_338
timestamp 1643671299
transform 1 0 28473 0 1 36167
box 0 0 1 1
use contact_13  contact_13_339
timestamp 1643671299
transform 1 0 28133 0 1 36185
box 0 0 1 1
use contact_21  contact_21_339
timestamp 1643671299
transform 1 0 28137 0 1 36167
box 0 0 1 1
use contact_13  contact_13_340
timestamp 1643671299
transform 1 0 27797 0 1 36185
box 0 0 1 1
use contact_21  contact_21_340
timestamp 1643671299
transform 1 0 27801 0 1 36167
box 0 0 1 1
use contact_13  contact_13_341
timestamp 1643671299
transform 1 0 27461 0 1 36185
box 0 0 1 1
use contact_21  contact_21_341
timestamp 1643671299
transform 1 0 27465 0 1 36167
box 0 0 1 1
use contact_18  contact_18_69
timestamp 1643671299
transform 1 0 27124 0 1 36178
box 0 0 1 1
use contact_17  contact_17_231
timestamp 1643671299
transform 1 0 27139 0 1 36193
box 0 0 1 1
use contact_13  contact_13_342
timestamp 1643671299
transform 1 0 27125 0 1 36185
box 0 0 1 1
use contact_21  contact_21_342
timestamp 1643671299
transform 1 0 27129 0 1 36167
box 0 0 1 1
use contact_13  contact_13_343
timestamp 1643671299
transform 1 0 26789 0 1 36185
box 0 0 1 1
use contact_21  contact_21_343
timestamp 1643671299
transform 1 0 26793 0 1 36167
box 0 0 1 1
use contact_13  contact_13_344
timestamp 1643671299
transform 1 0 26453 0 1 36185
box 0 0 1 1
use contact_21  contact_21_344
timestamp 1643671299
transform 1 0 26457 0 1 36167
box 0 0 1 1
use contact_13  contact_13_345
timestamp 1643671299
transform 1 0 26117 0 1 36185
box 0 0 1 1
use contact_21  contact_21_345
timestamp 1643671299
transform 1 0 26121 0 1 36167
box 0 0 1 1
use contact_13  contact_13_346
timestamp 1643671299
transform 1 0 25781 0 1 36185
box 0 0 1 1
use contact_21  contact_21_346
timestamp 1643671299
transform 1 0 25785 0 1 36167
box 0 0 1 1
use contact_18  contact_18_70
timestamp 1643671299
transform 1 0 25444 0 1 36178
box 0 0 1 1
use contact_17  contact_17_232
timestamp 1643671299
transform 1 0 25459 0 1 36193
box 0 0 1 1
use contact_13  contact_13_347
timestamp 1643671299
transform 1 0 25445 0 1 36185
box 0 0 1 1
use contact_21  contact_21_347
timestamp 1643671299
transform 1 0 25449 0 1 36167
box 0 0 1 1
use contact_13  contact_13_348
timestamp 1643671299
transform 1 0 25109 0 1 36185
box 0 0 1 1
use contact_21  contact_21_348
timestamp 1643671299
transform 1 0 25113 0 1 36167
box 0 0 1 1
use contact_13  contact_13_349
timestamp 1643671299
transform 1 0 24773 0 1 36185
box 0 0 1 1
use contact_21  contact_21_349
timestamp 1643671299
transform 1 0 24777 0 1 36167
box 0 0 1 1
use contact_13  contact_13_350
timestamp 1643671299
transform 1 0 24437 0 1 36185
box 0 0 1 1
use contact_21  contact_21_350
timestamp 1643671299
transform 1 0 24441 0 1 36167
box 0 0 1 1
use contact_13  contact_13_351
timestamp 1643671299
transform 1 0 24101 0 1 36185
box 0 0 1 1
use contact_21  contact_21_351
timestamp 1643671299
transform 1 0 24105 0 1 36167
box 0 0 1 1
use contact_18  contact_18_71
timestamp 1643671299
transform 1 0 23764 0 1 36178
box 0 0 1 1
use contact_17  contact_17_233
timestamp 1643671299
transform 1 0 23779 0 1 36193
box 0 0 1 1
use contact_13  contact_13_352
timestamp 1643671299
transform 1 0 23765 0 1 36185
box 0 0 1 1
use contact_21  contact_21_352
timestamp 1643671299
transform 1 0 23769 0 1 36167
box 0 0 1 1
use contact_13  contact_13_353
timestamp 1643671299
transform 1 0 23429 0 1 36185
box 0 0 1 1
use contact_21  contact_21_353
timestamp 1643671299
transform 1 0 23433 0 1 36167
box 0 0 1 1
use contact_13  contact_13_354
timestamp 1643671299
transform 1 0 23093 0 1 36185
box 0 0 1 1
use contact_21  contact_21_354
timestamp 1643671299
transform 1 0 23097 0 1 36167
box 0 0 1 1
use contact_13  contact_13_355
timestamp 1643671299
transform 1 0 22757 0 1 36185
box 0 0 1 1
use contact_21  contact_21_355
timestamp 1643671299
transform 1 0 22761 0 1 36167
box 0 0 1 1
use contact_13  contact_13_356
timestamp 1643671299
transform 1 0 22421 0 1 36185
box 0 0 1 1
use contact_21  contact_21_356
timestamp 1643671299
transform 1 0 22425 0 1 36167
box 0 0 1 1
use contact_18  contact_18_72
timestamp 1643671299
transform 1 0 22084 0 1 36178
box 0 0 1 1
use contact_17  contact_17_234
timestamp 1643671299
transform 1 0 22099 0 1 36193
box 0 0 1 1
use contact_13  contact_13_357
timestamp 1643671299
transform 1 0 22085 0 1 36185
box 0 0 1 1
use contact_21  contact_21_357
timestamp 1643671299
transform 1 0 22089 0 1 36167
box 0 0 1 1
use contact_13  contact_13_358
timestamp 1643671299
transform 1 0 21749 0 1 36185
box 0 0 1 1
use contact_21  contact_21_358
timestamp 1643671299
transform 1 0 21753 0 1 36167
box 0 0 1 1
use contact_13  contact_13_359
timestamp 1643671299
transform 1 0 21413 0 1 36185
box 0 0 1 1
use contact_21  contact_21_359
timestamp 1643671299
transform 1 0 21417 0 1 36167
box 0 0 1 1
use contact_13  contact_13_360
timestamp 1643671299
transform 1 0 21077 0 1 36185
box 0 0 1 1
use contact_21  contact_21_360
timestamp 1643671299
transform 1 0 21081 0 1 36167
box 0 0 1 1
use contact_13  contact_13_361
timestamp 1643671299
transform 1 0 20741 0 1 36185
box 0 0 1 1
use contact_21  contact_21_361
timestamp 1643671299
transform 1 0 20745 0 1 36167
box 0 0 1 1
use contact_18  contact_18_73
timestamp 1643671299
transform 1 0 20404 0 1 36178
box 0 0 1 1
use contact_17  contact_17_235
timestamp 1643671299
transform 1 0 20419 0 1 36193
box 0 0 1 1
use contact_13  contact_13_362
timestamp 1643671299
transform 1 0 20405 0 1 36185
box 0 0 1 1
use contact_21  contact_21_362
timestamp 1643671299
transform 1 0 20409 0 1 36167
box 0 0 1 1
use contact_13  contact_13_363
timestamp 1643671299
transform 1 0 20069 0 1 36185
box 0 0 1 1
use contact_21  contact_21_363
timestamp 1643671299
transform 1 0 20073 0 1 36167
box 0 0 1 1
use contact_13  contact_13_364
timestamp 1643671299
transform 1 0 19733 0 1 36185
box 0 0 1 1
use contact_21  contact_21_364
timestamp 1643671299
transform 1 0 19737 0 1 36167
box 0 0 1 1
use contact_13  contact_13_365
timestamp 1643671299
transform 1 0 19397 0 1 36185
box 0 0 1 1
use contact_21  contact_21_365
timestamp 1643671299
transform 1 0 19401 0 1 36167
box 0 0 1 1
use contact_13  contact_13_366
timestamp 1643671299
transform 1 0 19061 0 1 36185
box 0 0 1 1
use contact_21  contact_21_366
timestamp 1643671299
transform 1 0 19065 0 1 36167
box 0 0 1 1
use contact_18  contact_18_74
timestamp 1643671299
transform 1 0 18724 0 1 36178
box 0 0 1 1
use contact_17  contact_17_236
timestamp 1643671299
transform 1 0 18739 0 1 36193
box 0 0 1 1
use contact_13  contact_13_367
timestamp 1643671299
transform 1 0 18725 0 1 36185
box 0 0 1 1
use contact_21  contact_21_367
timestamp 1643671299
transform 1 0 18729 0 1 36167
box 0 0 1 1
use contact_13  contact_13_368
timestamp 1643671299
transform 1 0 18389 0 1 36185
box 0 0 1 1
use contact_21  contact_21_368
timestamp 1643671299
transform 1 0 18393 0 1 36167
box 0 0 1 1
use contact_13  contact_13_369
timestamp 1643671299
transform 1 0 18053 0 1 36185
box 0 0 1 1
use contact_21  contact_21_369
timestamp 1643671299
transform 1 0 18057 0 1 36167
box 0 0 1 1
use contact_13  contact_13_370
timestamp 1643671299
transform 1 0 17717 0 1 36185
box 0 0 1 1
use contact_21  contact_21_370
timestamp 1643671299
transform 1 0 17721 0 1 36167
box 0 0 1 1
use contact_13  contact_13_371
timestamp 1643671299
transform 1 0 17381 0 1 36185
box 0 0 1 1
use contact_21  contact_21_371
timestamp 1643671299
transform 1 0 17385 0 1 36167
box 0 0 1 1
use contact_18  contact_18_75
timestamp 1643671299
transform 1 0 17044 0 1 36178
box 0 0 1 1
use contact_17  contact_17_237
timestamp 1643671299
transform 1 0 17059 0 1 36193
box 0 0 1 1
use contact_13  contact_13_372
timestamp 1643671299
transform 1 0 17045 0 1 36185
box 0 0 1 1
use contact_21  contact_21_372
timestamp 1643671299
transform 1 0 17049 0 1 36167
box 0 0 1 1
use contact_13  contact_13_373
timestamp 1643671299
transform 1 0 16709 0 1 36185
box 0 0 1 1
use contact_21  contact_21_373
timestamp 1643671299
transform 1 0 16713 0 1 36167
box 0 0 1 1
use contact_13  contact_13_374
timestamp 1643671299
transform 1 0 16373 0 1 36185
box 0 0 1 1
use contact_21  contact_21_374
timestamp 1643671299
transform 1 0 16377 0 1 36167
box 0 0 1 1
use contact_13  contact_13_375
timestamp 1643671299
transform 1 0 16037 0 1 36185
box 0 0 1 1
use contact_21  contact_21_375
timestamp 1643671299
transform 1 0 16041 0 1 36167
box 0 0 1 1
use contact_13  contact_13_376
timestamp 1643671299
transform 1 0 15701 0 1 36185
box 0 0 1 1
use contact_21  contact_21_376
timestamp 1643671299
transform 1 0 15705 0 1 36167
box 0 0 1 1
use contact_18  contact_18_76
timestamp 1643671299
transform 1 0 15364 0 1 36178
box 0 0 1 1
use contact_17  contact_17_238
timestamp 1643671299
transform 1 0 15379 0 1 36193
box 0 0 1 1
use contact_13  contact_13_377
timestamp 1643671299
transform 1 0 15365 0 1 36185
box 0 0 1 1
use contact_21  contact_21_377
timestamp 1643671299
transform 1 0 15369 0 1 36167
box 0 0 1 1
use contact_13  contact_13_378
timestamp 1643671299
transform 1 0 15029 0 1 36185
box 0 0 1 1
use contact_21  contact_21_378
timestamp 1643671299
transform 1 0 15033 0 1 36167
box 0 0 1 1
use contact_13  contact_13_379
timestamp 1643671299
transform 1 0 14693 0 1 36185
box 0 0 1 1
use contact_21  contact_21_379
timestamp 1643671299
transform 1 0 14697 0 1 36167
box 0 0 1 1
use contact_13  contact_13_380
timestamp 1643671299
transform 1 0 14357 0 1 36185
box 0 0 1 1
use contact_21  contact_21_380
timestamp 1643671299
transform 1 0 14361 0 1 36167
box 0 0 1 1
use contact_13  contact_13_381
timestamp 1643671299
transform 1 0 14021 0 1 36185
box 0 0 1 1
use contact_21  contact_21_381
timestamp 1643671299
transform 1 0 14025 0 1 36167
box 0 0 1 1
use contact_18  contact_18_77
timestamp 1643671299
transform 1 0 13684 0 1 36178
box 0 0 1 1
use contact_17  contact_17_239
timestamp 1643671299
transform 1 0 13699 0 1 36193
box 0 0 1 1
use contact_13  contact_13_382
timestamp 1643671299
transform 1 0 13685 0 1 36185
box 0 0 1 1
use contact_21  contact_21_382
timestamp 1643671299
transform 1 0 13689 0 1 36167
box 0 0 1 1
use contact_13  contact_13_383
timestamp 1643671299
transform 1 0 13349 0 1 36185
box 0 0 1 1
use contact_21  contact_21_383
timestamp 1643671299
transform 1 0 13353 0 1 36167
box 0 0 1 1
use contact_13  contact_13_384
timestamp 1643671299
transform 1 0 13013 0 1 36185
box 0 0 1 1
use contact_21  contact_21_384
timestamp 1643671299
transform 1 0 13017 0 1 36167
box 0 0 1 1
use contact_13  contact_13_385
timestamp 1643671299
transform 1 0 12677 0 1 36185
box 0 0 1 1
use contact_21  contact_21_385
timestamp 1643671299
transform 1 0 12681 0 1 36167
box 0 0 1 1
use contact_13  contact_13_386
timestamp 1643671299
transform 1 0 12341 0 1 36185
box 0 0 1 1
use contact_21  contact_21_386
timestamp 1643671299
transform 1 0 12345 0 1 36167
box 0 0 1 1
use contact_18  contact_18_78
timestamp 1643671299
transform 1 0 12004 0 1 36178
box 0 0 1 1
use contact_17  contact_17_240
timestamp 1643671299
transform 1 0 12019 0 1 36193
box 0 0 1 1
use contact_13  contact_13_387
timestamp 1643671299
transform 1 0 12005 0 1 36185
box 0 0 1 1
use contact_21  contact_21_387
timestamp 1643671299
transform 1 0 12009 0 1 36167
box 0 0 1 1
use contact_13  contact_13_388
timestamp 1643671299
transform 1 0 11669 0 1 36185
box 0 0 1 1
use contact_21  contact_21_388
timestamp 1643671299
transform 1 0 11673 0 1 36167
box 0 0 1 1
use contact_13  contact_13_389
timestamp 1643671299
transform 1 0 11333 0 1 36185
box 0 0 1 1
use contact_21  contact_21_389
timestamp 1643671299
transform 1 0 11337 0 1 36167
box 0 0 1 1
use contact_13  contact_13_390
timestamp 1643671299
transform 1 0 10997 0 1 36185
box 0 0 1 1
use contact_21  contact_21_390
timestamp 1643671299
transform 1 0 11001 0 1 36167
box 0 0 1 1
use contact_13  contact_13_391
timestamp 1643671299
transform 1 0 10661 0 1 36185
box 0 0 1 1
use contact_21  contact_21_391
timestamp 1643671299
transform 1 0 10665 0 1 36167
box 0 0 1 1
use contact_18  contact_18_79
timestamp 1643671299
transform 1 0 10324 0 1 36178
box 0 0 1 1
use contact_17  contact_17_241
timestamp 1643671299
transform 1 0 10339 0 1 36193
box 0 0 1 1
use contact_13  contact_13_392
timestamp 1643671299
transform 1 0 10325 0 1 36185
box 0 0 1 1
use contact_21  contact_21_392
timestamp 1643671299
transform 1 0 10329 0 1 36167
box 0 0 1 1
use contact_13  contact_13_393
timestamp 1643671299
transform 1 0 9989 0 1 36185
box 0 0 1 1
use contact_21  contact_21_393
timestamp 1643671299
transform 1 0 9993 0 1 36167
box 0 0 1 1
use contact_13  contact_13_394
timestamp 1643671299
transform 1 0 9653 0 1 36185
box 0 0 1 1
use contact_21  contact_21_394
timestamp 1643671299
transform 1 0 9657 0 1 36167
box 0 0 1 1
use contact_13  contact_13_395
timestamp 1643671299
transform 1 0 9317 0 1 36185
box 0 0 1 1
use contact_21  contact_21_395
timestamp 1643671299
transform 1 0 9321 0 1 36167
box 0 0 1 1
use contact_13  contact_13_396
timestamp 1643671299
transform 1 0 8981 0 1 36185
box 0 0 1 1
use contact_21  contact_21_396
timestamp 1643671299
transform 1 0 8985 0 1 36167
box 0 0 1 1
use contact_18  contact_18_80
timestamp 1643671299
transform 1 0 8644 0 1 36178
box 0 0 1 1
use contact_17  contact_17_242
timestamp 1643671299
transform 1 0 8659 0 1 36193
box 0 0 1 1
use contact_13  contact_13_397
timestamp 1643671299
transform 1 0 8645 0 1 36185
box 0 0 1 1
use contact_21  contact_21_397
timestamp 1643671299
transform 1 0 8649 0 1 36167
box 0 0 1 1
use contact_13  contact_13_398
timestamp 1643671299
transform 1 0 8309 0 1 36185
box 0 0 1 1
use contact_21  contact_21_398
timestamp 1643671299
transform 1 0 8313 0 1 36167
box 0 0 1 1
use contact_13  contact_13_399
timestamp 1643671299
transform 1 0 7973 0 1 36185
box 0 0 1 1
use contact_21  contact_21_399
timestamp 1643671299
transform 1 0 7977 0 1 36167
box 0 0 1 1
use contact_13  contact_13_400
timestamp 1643671299
transform 1 0 7637 0 1 36185
box 0 0 1 1
use contact_21  contact_21_400
timestamp 1643671299
transform 1 0 7641 0 1 36167
box 0 0 1 1
use contact_13  contact_13_401
timestamp 1643671299
transform 1 0 7301 0 1 36185
box 0 0 1 1
use contact_21  contact_21_401
timestamp 1643671299
transform 1 0 7305 0 1 36167
box 0 0 1 1
use contact_18  contact_18_81
timestamp 1643671299
transform 1 0 6964 0 1 36178
box 0 0 1 1
use contact_17  contact_17_243
timestamp 1643671299
transform 1 0 6979 0 1 36193
box 0 0 1 1
use contact_13  contact_13_402
timestamp 1643671299
transform 1 0 6965 0 1 36185
box 0 0 1 1
use contact_21  contact_21_402
timestamp 1643671299
transform 1 0 6969 0 1 36167
box 0 0 1 1
use contact_13  contact_13_403
timestamp 1643671299
transform 1 0 6629 0 1 36185
box 0 0 1 1
use contact_21  contact_21_403
timestamp 1643671299
transform 1 0 6633 0 1 36167
box 0 0 1 1
use contact_13  contact_13_404
timestamp 1643671299
transform 1 0 6293 0 1 36185
box 0 0 1 1
use contact_21  contact_21_404
timestamp 1643671299
transform 1 0 6297 0 1 36167
box 0 0 1 1
use contact_13  contact_13_405
timestamp 1643671299
transform 1 0 5957 0 1 36185
box 0 0 1 1
use contact_21  contact_21_405
timestamp 1643671299
transform 1 0 5961 0 1 36167
box 0 0 1 1
use contact_13  contact_13_406
timestamp 1643671299
transform 1 0 5621 0 1 36185
box 0 0 1 1
use contact_21  contact_21_406
timestamp 1643671299
transform 1 0 5625 0 1 36167
box 0 0 1 1
use contact_18  contact_18_82
timestamp 1643671299
transform 1 0 5284 0 1 36178
box 0 0 1 1
use contact_17  contact_17_244
timestamp 1643671299
transform 1 0 5299 0 1 36193
box 0 0 1 1
use contact_13  contact_13_407
timestamp 1643671299
transform 1 0 5285 0 1 36185
box 0 0 1 1
use contact_21  contact_21_407
timestamp 1643671299
transform 1 0 5289 0 1 36167
box 0 0 1 1
use contact_13  contact_13_408
timestamp 1643671299
transform 1 0 4949 0 1 36185
box 0 0 1 1
use contact_21  contact_21_408
timestamp 1643671299
transform 1 0 4953 0 1 36167
box 0 0 1 1
use contact_13  contact_13_409
timestamp 1643671299
transform 1 0 4613 0 1 36185
box 0 0 1 1
use contact_21  contact_21_409
timestamp 1643671299
transform 1 0 4617 0 1 36167
box 0 0 1 1
use contact_13  contact_13_410
timestamp 1643671299
transform 1 0 4277 0 1 36185
box 0 0 1 1
use contact_21  contact_21_410
timestamp 1643671299
transform 1 0 4281 0 1 36167
box 0 0 1 1
use contact_13  contact_13_411
timestamp 1643671299
transform 1 0 3941 0 1 36185
box 0 0 1 1
use contact_21  contact_21_411
timestamp 1643671299
transform 1 0 3945 0 1 36167
box 0 0 1 1
use contact_18  contact_18_83
timestamp 1643671299
transform 1 0 3604 0 1 36178
box 0 0 1 1
use contact_17  contact_17_245
timestamp 1643671299
transform 1 0 3619 0 1 36193
box 0 0 1 1
use contact_13  contact_13_412
timestamp 1643671299
transform 1 0 3605 0 1 36185
box 0 0 1 1
use contact_21  contact_21_412
timestamp 1643671299
transform 1 0 3609 0 1 36167
box 0 0 1 1
use contact_13  contact_13_413
timestamp 1643671299
transform 1 0 3269 0 1 36185
box 0 0 1 1
use contact_21  contact_21_413
timestamp 1643671299
transform 1 0 3273 0 1 36167
box 0 0 1 1
use contact_13  contact_13_414
timestamp 1643671299
transform 1 0 2933 0 1 36185
box 0 0 1 1
use contact_21  contact_21_414
timestamp 1643671299
transform 1 0 2937 0 1 36167
box 0 0 1 1
use contact_13  contact_13_415
timestamp 1643671299
transform 1 0 2597 0 1 36185
box 0 0 1 1
use contact_21  contact_21_415
timestamp 1643671299
transform 1 0 2601 0 1 36167
box 0 0 1 1
use contact_13  contact_13_416
timestamp 1643671299
transform 1 0 2261 0 1 36185
box 0 0 1 1
use contact_21  contact_21_416
timestamp 1643671299
transform 1 0 2265 0 1 36167
box 0 0 1 1
use contact_18  contact_18_84
timestamp 1643671299
transform 1 0 1924 0 1 36178
box 0 0 1 1
use contact_17  contact_17_246
timestamp 1643671299
transform 1 0 1939 0 1 36193
box 0 0 1 1
use contact_13  contact_13_417
timestamp 1643671299
transform 1 0 1925 0 1 36185
box 0 0 1 1
use contact_21  contact_21_417
timestamp 1643671299
transform 1 0 1929 0 1 36167
box 0 0 1 1
use contact_13  contact_13_418
timestamp 1643671299
transform 1 0 73493 0 1 1541
box 0 0 1 1
use contact_21  contact_21_418
timestamp 1643671299
transform 1 0 73497 0 1 1523
box 0 0 1 1
use contact_13  contact_13_419
timestamp 1643671299
transform 1 0 73157 0 1 1541
box 0 0 1 1
use contact_21  contact_21_419
timestamp 1643671299
transform 1 0 73161 0 1 1523
box 0 0 1 1
use contact_13  contact_13_420
timestamp 1643671299
transform 1 0 72821 0 1 1541
box 0 0 1 1
use contact_21  contact_21_420
timestamp 1643671299
transform 1 0 72825 0 1 1523
box 0 0 1 1
use contact_18  contact_18_85
timestamp 1643671299
transform 1 0 72484 0 1 1534
box 0 0 1 1
use contact_17  contact_17_247
timestamp 1643671299
transform 1 0 72499 0 1 1549
box 0 0 1 1
use contact_13  contact_13_421
timestamp 1643671299
transform 1 0 72485 0 1 1541
box 0 0 1 1
use contact_21  contact_21_421
timestamp 1643671299
transform 1 0 72489 0 1 1523
box 0 0 1 1
use contact_13  contact_13_422
timestamp 1643671299
transform 1 0 72149 0 1 1541
box 0 0 1 1
use contact_21  contact_21_422
timestamp 1643671299
transform 1 0 72153 0 1 1523
box 0 0 1 1
use contact_13  contact_13_423
timestamp 1643671299
transform 1 0 71813 0 1 1541
box 0 0 1 1
use contact_21  contact_21_423
timestamp 1643671299
transform 1 0 71817 0 1 1523
box 0 0 1 1
use contact_13  contact_13_424
timestamp 1643671299
transform 1 0 71477 0 1 1541
box 0 0 1 1
use contact_21  contact_21_424
timestamp 1643671299
transform 1 0 71481 0 1 1523
box 0 0 1 1
use contact_13  contact_13_425
timestamp 1643671299
transform 1 0 71141 0 1 1541
box 0 0 1 1
use contact_21  contact_21_425
timestamp 1643671299
transform 1 0 71145 0 1 1523
box 0 0 1 1
use contact_18  contact_18_86
timestamp 1643671299
transform 1 0 70804 0 1 1534
box 0 0 1 1
use contact_17  contact_17_248
timestamp 1643671299
transform 1 0 70819 0 1 1549
box 0 0 1 1
use contact_13  contact_13_426
timestamp 1643671299
transform 1 0 70805 0 1 1541
box 0 0 1 1
use contact_21  contact_21_426
timestamp 1643671299
transform 1 0 70809 0 1 1523
box 0 0 1 1
use contact_13  contact_13_427
timestamp 1643671299
transform 1 0 70469 0 1 1541
box 0 0 1 1
use contact_21  contact_21_427
timestamp 1643671299
transform 1 0 70473 0 1 1523
box 0 0 1 1
use contact_13  contact_13_428
timestamp 1643671299
transform 1 0 70133 0 1 1541
box 0 0 1 1
use contact_21  contact_21_428
timestamp 1643671299
transform 1 0 70137 0 1 1523
box 0 0 1 1
use contact_13  contact_13_429
timestamp 1643671299
transform 1 0 69797 0 1 1541
box 0 0 1 1
use contact_21  contact_21_429
timestamp 1643671299
transform 1 0 69801 0 1 1523
box 0 0 1 1
use contact_13  contact_13_430
timestamp 1643671299
transform 1 0 69461 0 1 1541
box 0 0 1 1
use contact_21  contact_21_430
timestamp 1643671299
transform 1 0 69465 0 1 1523
box 0 0 1 1
use contact_18  contact_18_87
timestamp 1643671299
transform 1 0 69124 0 1 1534
box 0 0 1 1
use contact_17  contact_17_249
timestamp 1643671299
transform 1 0 69139 0 1 1549
box 0 0 1 1
use contact_13  contact_13_431
timestamp 1643671299
transform 1 0 69125 0 1 1541
box 0 0 1 1
use contact_21  contact_21_431
timestamp 1643671299
transform 1 0 69129 0 1 1523
box 0 0 1 1
use contact_13  contact_13_432
timestamp 1643671299
transform 1 0 68789 0 1 1541
box 0 0 1 1
use contact_21  contact_21_432
timestamp 1643671299
transform 1 0 68793 0 1 1523
box 0 0 1 1
use contact_13  contact_13_433
timestamp 1643671299
transform 1 0 68453 0 1 1541
box 0 0 1 1
use contact_21  contact_21_433
timestamp 1643671299
transform 1 0 68457 0 1 1523
box 0 0 1 1
use contact_13  contact_13_434
timestamp 1643671299
transform 1 0 68117 0 1 1541
box 0 0 1 1
use contact_21  contact_21_434
timestamp 1643671299
transform 1 0 68121 0 1 1523
box 0 0 1 1
use contact_13  contact_13_435
timestamp 1643671299
transform 1 0 67781 0 1 1541
box 0 0 1 1
use contact_21  contact_21_435
timestamp 1643671299
transform 1 0 67785 0 1 1523
box 0 0 1 1
use contact_18  contact_18_88
timestamp 1643671299
transform 1 0 67444 0 1 1534
box 0 0 1 1
use contact_17  contact_17_250
timestamp 1643671299
transform 1 0 67459 0 1 1549
box 0 0 1 1
use contact_13  contact_13_436
timestamp 1643671299
transform 1 0 67445 0 1 1541
box 0 0 1 1
use contact_21  contact_21_436
timestamp 1643671299
transform 1 0 67449 0 1 1523
box 0 0 1 1
use contact_13  contact_13_437
timestamp 1643671299
transform 1 0 67109 0 1 1541
box 0 0 1 1
use contact_21  contact_21_437
timestamp 1643671299
transform 1 0 67113 0 1 1523
box 0 0 1 1
use contact_13  contact_13_438
timestamp 1643671299
transform 1 0 66773 0 1 1541
box 0 0 1 1
use contact_21  contact_21_438
timestamp 1643671299
transform 1 0 66777 0 1 1523
box 0 0 1 1
use contact_13  contact_13_439
timestamp 1643671299
transform 1 0 66437 0 1 1541
box 0 0 1 1
use contact_21  contact_21_439
timestamp 1643671299
transform 1 0 66441 0 1 1523
box 0 0 1 1
use contact_13  contact_13_440
timestamp 1643671299
transform 1 0 66101 0 1 1541
box 0 0 1 1
use contact_21  contact_21_440
timestamp 1643671299
transform 1 0 66105 0 1 1523
box 0 0 1 1
use contact_18  contact_18_89
timestamp 1643671299
transform 1 0 65764 0 1 1534
box 0 0 1 1
use contact_17  contact_17_251
timestamp 1643671299
transform 1 0 65779 0 1 1549
box 0 0 1 1
use contact_13  contact_13_441
timestamp 1643671299
transform 1 0 65765 0 1 1541
box 0 0 1 1
use contact_21  contact_21_441
timestamp 1643671299
transform 1 0 65769 0 1 1523
box 0 0 1 1
use contact_13  contact_13_442
timestamp 1643671299
transform 1 0 65429 0 1 1541
box 0 0 1 1
use contact_21  contact_21_442
timestamp 1643671299
transform 1 0 65433 0 1 1523
box 0 0 1 1
use contact_13  contact_13_443
timestamp 1643671299
transform 1 0 65093 0 1 1541
box 0 0 1 1
use contact_21  contact_21_443
timestamp 1643671299
transform 1 0 65097 0 1 1523
box 0 0 1 1
use contact_13  contact_13_444
timestamp 1643671299
transform 1 0 64757 0 1 1541
box 0 0 1 1
use contact_21  contact_21_444
timestamp 1643671299
transform 1 0 64761 0 1 1523
box 0 0 1 1
use contact_13  contact_13_445
timestamp 1643671299
transform 1 0 64421 0 1 1541
box 0 0 1 1
use contact_21  contact_21_445
timestamp 1643671299
transform 1 0 64425 0 1 1523
box 0 0 1 1
use contact_18  contact_18_90
timestamp 1643671299
transform 1 0 64084 0 1 1534
box 0 0 1 1
use contact_17  contact_17_252
timestamp 1643671299
transform 1 0 64099 0 1 1549
box 0 0 1 1
use contact_13  contact_13_446
timestamp 1643671299
transform 1 0 64085 0 1 1541
box 0 0 1 1
use contact_21  contact_21_446
timestamp 1643671299
transform 1 0 64089 0 1 1523
box 0 0 1 1
use contact_13  contact_13_447
timestamp 1643671299
transform 1 0 63749 0 1 1541
box 0 0 1 1
use contact_21  contact_21_447
timestamp 1643671299
transform 1 0 63753 0 1 1523
box 0 0 1 1
use contact_13  contact_13_448
timestamp 1643671299
transform 1 0 63413 0 1 1541
box 0 0 1 1
use contact_21  contact_21_448
timestamp 1643671299
transform 1 0 63417 0 1 1523
box 0 0 1 1
use contact_13  contact_13_449
timestamp 1643671299
transform 1 0 63077 0 1 1541
box 0 0 1 1
use contact_21  contact_21_449
timestamp 1643671299
transform 1 0 63081 0 1 1523
box 0 0 1 1
use contact_13  contact_13_450
timestamp 1643671299
transform 1 0 62741 0 1 1541
box 0 0 1 1
use contact_21  contact_21_450
timestamp 1643671299
transform 1 0 62745 0 1 1523
box 0 0 1 1
use contact_18  contact_18_91
timestamp 1643671299
transform 1 0 62404 0 1 1534
box 0 0 1 1
use contact_17  contact_17_253
timestamp 1643671299
transform 1 0 62419 0 1 1549
box 0 0 1 1
use contact_13  contact_13_451
timestamp 1643671299
transform 1 0 62405 0 1 1541
box 0 0 1 1
use contact_21  contact_21_451
timestamp 1643671299
transform 1 0 62409 0 1 1523
box 0 0 1 1
use contact_13  contact_13_452
timestamp 1643671299
transform 1 0 62069 0 1 1541
box 0 0 1 1
use contact_21  contact_21_452
timestamp 1643671299
transform 1 0 62073 0 1 1523
box 0 0 1 1
use contact_13  contact_13_453
timestamp 1643671299
transform 1 0 61733 0 1 1541
box 0 0 1 1
use contact_21  contact_21_453
timestamp 1643671299
transform 1 0 61737 0 1 1523
box 0 0 1 1
use contact_13  contact_13_454
timestamp 1643671299
transform 1 0 61397 0 1 1541
box 0 0 1 1
use contact_21  contact_21_454
timestamp 1643671299
transform 1 0 61401 0 1 1523
box 0 0 1 1
use contact_13  contact_13_455
timestamp 1643671299
transform 1 0 61061 0 1 1541
box 0 0 1 1
use contact_21  contact_21_455
timestamp 1643671299
transform 1 0 61065 0 1 1523
box 0 0 1 1
use contact_18  contact_18_92
timestamp 1643671299
transform 1 0 60724 0 1 1534
box 0 0 1 1
use contact_17  contact_17_254
timestamp 1643671299
transform 1 0 60739 0 1 1549
box 0 0 1 1
use contact_13  contact_13_456
timestamp 1643671299
transform 1 0 60725 0 1 1541
box 0 0 1 1
use contact_21  contact_21_456
timestamp 1643671299
transform 1 0 60729 0 1 1523
box 0 0 1 1
use contact_13  contact_13_457
timestamp 1643671299
transform 1 0 60389 0 1 1541
box 0 0 1 1
use contact_21  contact_21_457
timestamp 1643671299
transform 1 0 60393 0 1 1523
box 0 0 1 1
use contact_13  contact_13_458
timestamp 1643671299
transform 1 0 60053 0 1 1541
box 0 0 1 1
use contact_21  contact_21_458
timestamp 1643671299
transform 1 0 60057 0 1 1523
box 0 0 1 1
use contact_13  contact_13_459
timestamp 1643671299
transform 1 0 59717 0 1 1541
box 0 0 1 1
use contact_21  contact_21_459
timestamp 1643671299
transform 1 0 59721 0 1 1523
box 0 0 1 1
use contact_13  contact_13_460
timestamp 1643671299
transform 1 0 59381 0 1 1541
box 0 0 1 1
use contact_21  contact_21_460
timestamp 1643671299
transform 1 0 59385 0 1 1523
box 0 0 1 1
use contact_18  contact_18_93
timestamp 1643671299
transform 1 0 59044 0 1 1534
box 0 0 1 1
use contact_17  contact_17_255
timestamp 1643671299
transform 1 0 59059 0 1 1549
box 0 0 1 1
use contact_13  contact_13_461
timestamp 1643671299
transform 1 0 59045 0 1 1541
box 0 0 1 1
use contact_21  contact_21_461
timestamp 1643671299
transform 1 0 59049 0 1 1523
box 0 0 1 1
use contact_13  contact_13_462
timestamp 1643671299
transform 1 0 58709 0 1 1541
box 0 0 1 1
use contact_21  contact_21_462
timestamp 1643671299
transform 1 0 58713 0 1 1523
box 0 0 1 1
use contact_13  contact_13_463
timestamp 1643671299
transform 1 0 58373 0 1 1541
box 0 0 1 1
use contact_21  contact_21_463
timestamp 1643671299
transform 1 0 58377 0 1 1523
box 0 0 1 1
use contact_13  contact_13_464
timestamp 1643671299
transform 1 0 58037 0 1 1541
box 0 0 1 1
use contact_21  contact_21_464
timestamp 1643671299
transform 1 0 58041 0 1 1523
box 0 0 1 1
use contact_13  contact_13_465
timestamp 1643671299
transform 1 0 57701 0 1 1541
box 0 0 1 1
use contact_21  contact_21_465
timestamp 1643671299
transform 1 0 57705 0 1 1523
box 0 0 1 1
use contact_18  contact_18_94
timestamp 1643671299
transform 1 0 57364 0 1 1534
box 0 0 1 1
use contact_17  contact_17_256
timestamp 1643671299
transform 1 0 57379 0 1 1549
box 0 0 1 1
use contact_13  contact_13_466
timestamp 1643671299
transform 1 0 57365 0 1 1541
box 0 0 1 1
use contact_21  contact_21_466
timestamp 1643671299
transform 1 0 57369 0 1 1523
box 0 0 1 1
use contact_13  contact_13_467
timestamp 1643671299
transform 1 0 57029 0 1 1541
box 0 0 1 1
use contact_21  contact_21_467
timestamp 1643671299
transform 1 0 57033 0 1 1523
box 0 0 1 1
use contact_13  contact_13_468
timestamp 1643671299
transform 1 0 56693 0 1 1541
box 0 0 1 1
use contact_21  contact_21_468
timestamp 1643671299
transform 1 0 56697 0 1 1523
box 0 0 1 1
use contact_13  contact_13_469
timestamp 1643671299
transform 1 0 56357 0 1 1541
box 0 0 1 1
use contact_21  contact_21_469
timestamp 1643671299
transform 1 0 56361 0 1 1523
box 0 0 1 1
use contact_13  contact_13_470
timestamp 1643671299
transform 1 0 56021 0 1 1541
box 0 0 1 1
use contact_21  contact_21_470
timestamp 1643671299
transform 1 0 56025 0 1 1523
box 0 0 1 1
use contact_18  contact_18_95
timestamp 1643671299
transform 1 0 55684 0 1 1534
box 0 0 1 1
use contact_17  contact_17_257
timestamp 1643671299
transform 1 0 55699 0 1 1549
box 0 0 1 1
use contact_13  contact_13_471
timestamp 1643671299
transform 1 0 55685 0 1 1541
box 0 0 1 1
use contact_21  contact_21_471
timestamp 1643671299
transform 1 0 55689 0 1 1523
box 0 0 1 1
use contact_13  contact_13_472
timestamp 1643671299
transform 1 0 55349 0 1 1541
box 0 0 1 1
use contact_21  contact_21_472
timestamp 1643671299
transform 1 0 55353 0 1 1523
box 0 0 1 1
use contact_13  contact_13_473
timestamp 1643671299
transform 1 0 55013 0 1 1541
box 0 0 1 1
use contact_21  contact_21_473
timestamp 1643671299
transform 1 0 55017 0 1 1523
box 0 0 1 1
use contact_13  contact_13_474
timestamp 1643671299
transform 1 0 54677 0 1 1541
box 0 0 1 1
use contact_21  contact_21_474
timestamp 1643671299
transform 1 0 54681 0 1 1523
box 0 0 1 1
use contact_13  contact_13_475
timestamp 1643671299
transform 1 0 54341 0 1 1541
box 0 0 1 1
use contact_21  contact_21_475
timestamp 1643671299
transform 1 0 54345 0 1 1523
box 0 0 1 1
use contact_18  contact_18_96
timestamp 1643671299
transform 1 0 54004 0 1 1534
box 0 0 1 1
use contact_17  contact_17_258
timestamp 1643671299
transform 1 0 54019 0 1 1549
box 0 0 1 1
use contact_13  contact_13_476
timestamp 1643671299
transform 1 0 54005 0 1 1541
box 0 0 1 1
use contact_21  contact_21_476
timestamp 1643671299
transform 1 0 54009 0 1 1523
box 0 0 1 1
use contact_13  contact_13_477
timestamp 1643671299
transform 1 0 53669 0 1 1541
box 0 0 1 1
use contact_21  contact_21_477
timestamp 1643671299
transform 1 0 53673 0 1 1523
box 0 0 1 1
use contact_13  contact_13_478
timestamp 1643671299
transform 1 0 53333 0 1 1541
box 0 0 1 1
use contact_21  contact_21_478
timestamp 1643671299
transform 1 0 53337 0 1 1523
box 0 0 1 1
use contact_13  contact_13_479
timestamp 1643671299
transform 1 0 52997 0 1 1541
box 0 0 1 1
use contact_21  contact_21_479
timestamp 1643671299
transform 1 0 53001 0 1 1523
box 0 0 1 1
use contact_13  contact_13_480
timestamp 1643671299
transform 1 0 52661 0 1 1541
box 0 0 1 1
use contact_21  contact_21_480
timestamp 1643671299
transform 1 0 52665 0 1 1523
box 0 0 1 1
use contact_18  contact_18_97
timestamp 1643671299
transform 1 0 52324 0 1 1534
box 0 0 1 1
use contact_17  contact_17_259
timestamp 1643671299
transform 1 0 52339 0 1 1549
box 0 0 1 1
use contact_13  contact_13_481
timestamp 1643671299
transform 1 0 52325 0 1 1541
box 0 0 1 1
use contact_21  contact_21_481
timestamp 1643671299
transform 1 0 52329 0 1 1523
box 0 0 1 1
use contact_13  contact_13_482
timestamp 1643671299
transform 1 0 51989 0 1 1541
box 0 0 1 1
use contact_21  contact_21_482
timestamp 1643671299
transform 1 0 51993 0 1 1523
box 0 0 1 1
use contact_13  contact_13_483
timestamp 1643671299
transform 1 0 51653 0 1 1541
box 0 0 1 1
use contact_21  contact_21_483
timestamp 1643671299
transform 1 0 51657 0 1 1523
box 0 0 1 1
use contact_13  contact_13_484
timestamp 1643671299
transform 1 0 51317 0 1 1541
box 0 0 1 1
use contact_21  contact_21_484
timestamp 1643671299
transform 1 0 51321 0 1 1523
box 0 0 1 1
use contact_13  contact_13_485
timestamp 1643671299
transform 1 0 50981 0 1 1541
box 0 0 1 1
use contact_21  contact_21_485
timestamp 1643671299
transform 1 0 50985 0 1 1523
box 0 0 1 1
use contact_18  contact_18_98
timestamp 1643671299
transform 1 0 50644 0 1 1534
box 0 0 1 1
use contact_17  contact_17_260
timestamp 1643671299
transform 1 0 50659 0 1 1549
box 0 0 1 1
use contact_13  contact_13_486
timestamp 1643671299
transform 1 0 50645 0 1 1541
box 0 0 1 1
use contact_21  contact_21_486
timestamp 1643671299
transform 1 0 50649 0 1 1523
box 0 0 1 1
use contact_13  contact_13_487
timestamp 1643671299
transform 1 0 50309 0 1 1541
box 0 0 1 1
use contact_21  contact_21_487
timestamp 1643671299
transform 1 0 50313 0 1 1523
box 0 0 1 1
use contact_13  contact_13_488
timestamp 1643671299
transform 1 0 49973 0 1 1541
box 0 0 1 1
use contact_21  contact_21_488
timestamp 1643671299
transform 1 0 49977 0 1 1523
box 0 0 1 1
use contact_13  contact_13_489
timestamp 1643671299
transform 1 0 49637 0 1 1541
box 0 0 1 1
use contact_21  contact_21_489
timestamp 1643671299
transform 1 0 49641 0 1 1523
box 0 0 1 1
use contact_13  contact_13_490
timestamp 1643671299
transform 1 0 49301 0 1 1541
box 0 0 1 1
use contact_21  contact_21_490
timestamp 1643671299
transform 1 0 49305 0 1 1523
box 0 0 1 1
use contact_18  contact_18_99
timestamp 1643671299
transform 1 0 48964 0 1 1534
box 0 0 1 1
use contact_17  contact_17_261
timestamp 1643671299
transform 1 0 48979 0 1 1549
box 0 0 1 1
use contact_13  contact_13_491
timestamp 1643671299
transform 1 0 48965 0 1 1541
box 0 0 1 1
use contact_21  contact_21_491
timestamp 1643671299
transform 1 0 48969 0 1 1523
box 0 0 1 1
use contact_13  contact_13_492
timestamp 1643671299
transform 1 0 48629 0 1 1541
box 0 0 1 1
use contact_21  contact_21_492
timestamp 1643671299
transform 1 0 48633 0 1 1523
box 0 0 1 1
use contact_13  contact_13_493
timestamp 1643671299
transform 1 0 48293 0 1 1541
box 0 0 1 1
use contact_21  contact_21_493
timestamp 1643671299
transform 1 0 48297 0 1 1523
box 0 0 1 1
use contact_13  contact_13_494
timestamp 1643671299
transform 1 0 47957 0 1 1541
box 0 0 1 1
use contact_21  contact_21_494
timestamp 1643671299
transform 1 0 47961 0 1 1523
box 0 0 1 1
use contact_13  contact_13_495
timestamp 1643671299
transform 1 0 47621 0 1 1541
box 0 0 1 1
use contact_21  contact_21_495
timestamp 1643671299
transform 1 0 47625 0 1 1523
box 0 0 1 1
use contact_18  contact_18_100
timestamp 1643671299
transform 1 0 47284 0 1 1534
box 0 0 1 1
use contact_17  contact_17_262
timestamp 1643671299
transform 1 0 47299 0 1 1549
box 0 0 1 1
use contact_13  contact_13_496
timestamp 1643671299
transform 1 0 47285 0 1 1541
box 0 0 1 1
use contact_21  contact_21_496
timestamp 1643671299
transform 1 0 47289 0 1 1523
box 0 0 1 1
use contact_13  contact_13_497
timestamp 1643671299
transform 1 0 46949 0 1 1541
box 0 0 1 1
use contact_21  contact_21_497
timestamp 1643671299
transform 1 0 46953 0 1 1523
box 0 0 1 1
use contact_13  contact_13_498
timestamp 1643671299
transform 1 0 46613 0 1 1541
box 0 0 1 1
use contact_21  contact_21_498
timestamp 1643671299
transform 1 0 46617 0 1 1523
box 0 0 1 1
use contact_13  contact_13_499
timestamp 1643671299
transform 1 0 46277 0 1 1541
box 0 0 1 1
use contact_21  contact_21_499
timestamp 1643671299
transform 1 0 46281 0 1 1523
box 0 0 1 1
use contact_13  contact_13_500
timestamp 1643671299
transform 1 0 45941 0 1 1541
box 0 0 1 1
use contact_21  contact_21_500
timestamp 1643671299
transform 1 0 45945 0 1 1523
box 0 0 1 1
use contact_18  contact_18_101
timestamp 1643671299
transform 1 0 45604 0 1 1534
box 0 0 1 1
use contact_17  contact_17_263
timestamp 1643671299
transform 1 0 45619 0 1 1549
box 0 0 1 1
use contact_13  contact_13_501
timestamp 1643671299
transform 1 0 45605 0 1 1541
box 0 0 1 1
use contact_21  contact_21_501
timestamp 1643671299
transform 1 0 45609 0 1 1523
box 0 0 1 1
use contact_13  contact_13_502
timestamp 1643671299
transform 1 0 45269 0 1 1541
box 0 0 1 1
use contact_21  contact_21_502
timestamp 1643671299
transform 1 0 45273 0 1 1523
box 0 0 1 1
use contact_13  contact_13_503
timestamp 1643671299
transform 1 0 44933 0 1 1541
box 0 0 1 1
use contact_21  contact_21_503
timestamp 1643671299
transform 1 0 44937 0 1 1523
box 0 0 1 1
use contact_13  contact_13_504
timestamp 1643671299
transform 1 0 44597 0 1 1541
box 0 0 1 1
use contact_21  contact_21_504
timestamp 1643671299
transform 1 0 44601 0 1 1523
box 0 0 1 1
use contact_13  contact_13_505
timestamp 1643671299
transform 1 0 44261 0 1 1541
box 0 0 1 1
use contact_21  contact_21_505
timestamp 1643671299
transform 1 0 44265 0 1 1523
box 0 0 1 1
use contact_18  contact_18_102
timestamp 1643671299
transform 1 0 43924 0 1 1534
box 0 0 1 1
use contact_17  contact_17_264
timestamp 1643671299
transform 1 0 43939 0 1 1549
box 0 0 1 1
use contact_13  contact_13_506
timestamp 1643671299
transform 1 0 43925 0 1 1541
box 0 0 1 1
use contact_21  contact_21_506
timestamp 1643671299
transform 1 0 43929 0 1 1523
box 0 0 1 1
use contact_13  contact_13_507
timestamp 1643671299
transform 1 0 43589 0 1 1541
box 0 0 1 1
use contact_21  contact_21_507
timestamp 1643671299
transform 1 0 43593 0 1 1523
box 0 0 1 1
use contact_13  contact_13_508
timestamp 1643671299
transform 1 0 43253 0 1 1541
box 0 0 1 1
use contact_21  contact_21_508
timestamp 1643671299
transform 1 0 43257 0 1 1523
box 0 0 1 1
use contact_13  contact_13_509
timestamp 1643671299
transform 1 0 42917 0 1 1541
box 0 0 1 1
use contact_21  contact_21_509
timestamp 1643671299
transform 1 0 42921 0 1 1523
box 0 0 1 1
use contact_13  contact_13_510
timestamp 1643671299
transform 1 0 42581 0 1 1541
box 0 0 1 1
use contact_21  contact_21_510
timestamp 1643671299
transform 1 0 42585 0 1 1523
box 0 0 1 1
use contact_18  contact_18_103
timestamp 1643671299
transform 1 0 42244 0 1 1534
box 0 0 1 1
use contact_17  contact_17_265
timestamp 1643671299
transform 1 0 42259 0 1 1549
box 0 0 1 1
use contact_13  contact_13_511
timestamp 1643671299
transform 1 0 42245 0 1 1541
box 0 0 1 1
use contact_21  contact_21_511
timestamp 1643671299
transform 1 0 42249 0 1 1523
box 0 0 1 1
use contact_13  contact_13_512
timestamp 1643671299
transform 1 0 41909 0 1 1541
box 0 0 1 1
use contact_21  contact_21_512
timestamp 1643671299
transform 1 0 41913 0 1 1523
box 0 0 1 1
use contact_13  contact_13_513
timestamp 1643671299
transform 1 0 41573 0 1 1541
box 0 0 1 1
use contact_21  contact_21_513
timestamp 1643671299
transform 1 0 41577 0 1 1523
box 0 0 1 1
use contact_13  contact_13_514
timestamp 1643671299
transform 1 0 41237 0 1 1541
box 0 0 1 1
use contact_21  contact_21_514
timestamp 1643671299
transform 1 0 41241 0 1 1523
box 0 0 1 1
use contact_13  contact_13_515
timestamp 1643671299
transform 1 0 40901 0 1 1541
box 0 0 1 1
use contact_21  contact_21_515
timestamp 1643671299
transform 1 0 40905 0 1 1523
box 0 0 1 1
use contact_18  contact_18_104
timestamp 1643671299
transform 1 0 40564 0 1 1534
box 0 0 1 1
use contact_17  contact_17_266
timestamp 1643671299
transform 1 0 40579 0 1 1549
box 0 0 1 1
use contact_13  contact_13_516
timestamp 1643671299
transform 1 0 40565 0 1 1541
box 0 0 1 1
use contact_21  contact_21_516
timestamp 1643671299
transform 1 0 40569 0 1 1523
box 0 0 1 1
use contact_13  contact_13_517
timestamp 1643671299
transform 1 0 40229 0 1 1541
box 0 0 1 1
use contact_21  contact_21_517
timestamp 1643671299
transform 1 0 40233 0 1 1523
box 0 0 1 1
use contact_13  contact_13_518
timestamp 1643671299
transform 1 0 39893 0 1 1541
box 0 0 1 1
use contact_21  contact_21_518
timestamp 1643671299
transform 1 0 39897 0 1 1523
box 0 0 1 1
use contact_13  contact_13_519
timestamp 1643671299
transform 1 0 39557 0 1 1541
box 0 0 1 1
use contact_21  contact_21_519
timestamp 1643671299
transform 1 0 39561 0 1 1523
box 0 0 1 1
use contact_13  contact_13_520
timestamp 1643671299
transform 1 0 39221 0 1 1541
box 0 0 1 1
use contact_21  contact_21_520
timestamp 1643671299
transform 1 0 39225 0 1 1523
box 0 0 1 1
use contact_18  contact_18_105
timestamp 1643671299
transform 1 0 38884 0 1 1534
box 0 0 1 1
use contact_17  contact_17_267
timestamp 1643671299
transform 1 0 38899 0 1 1549
box 0 0 1 1
use contact_13  contact_13_521
timestamp 1643671299
transform 1 0 38885 0 1 1541
box 0 0 1 1
use contact_21  contact_21_521
timestamp 1643671299
transform 1 0 38889 0 1 1523
box 0 0 1 1
use contact_13  contact_13_522
timestamp 1643671299
transform 1 0 38549 0 1 1541
box 0 0 1 1
use contact_21  contact_21_522
timestamp 1643671299
transform 1 0 38553 0 1 1523
box 0 0 1 1
use contact_13  contact_13_523
timestamp 1643671299
transform 1 0 38213 0 1 1541
box 0 0 1 1
use contact_21  contact_21_523
timestamp 1643671299
transform 1 0 38217 0 1 1523
box 0 0 1 1
use contact_13  contact_13_524
timestamp 1643671299
transform 1 0 37877 0 1 1541
box 0 0 1 1
use contact_21  contact_21_524
timestamp 1643671299
transform 1 0 37881 0 1 1523
box 0 0 1 1
use contact_13  contact_13_525
timestamp 1643671299
transform 1 0 37541 0 1 1541
box 0 0 1 1
use contact_21  contact_21_525
timestamp 1643671299
transform 1 0 37545 0 1 1523
box 0 0 1 1
use contact_18  contact_18_106
timestamp 1643671299
transform 1 0 37204 0 1 1534
box 0 0 1 1
use contact_17  contact_17_268
timestamp 1643671299
transform 1 0 37219 0 1 1549
box 0 0 1 1
use contact_13  contact_13_526
timestamp 1643671299
transform 1 0 37205 0 1 1541
box 0 0 1 1
use contact_21  contact_21_526
timestamp 1643671299
transform 1 0 37209 0 1 1523
box 0 0 1 1
use contact_13  contact_13_527
timestamp 1643671299
transform 1 0 36869 0 1 1541
box 0 0 1 1
use contact_21  contact_21_527
timestamp 1643671299
transform 1 0 36873 0 1 1523
box 0 0 1 1
use contact_13  contact_13_528
timestamp 1643671299
transform 1 0 36533 0 1 1541
box 0 0 1 1
use contact_21  contact_21_528
timestamp 1643671299
transform 1 0 36537 0 1 1523
box 0 0 1 1
use contact_13  contact_13_529
timestamp 1643671299
transform 1 0 36197 0 1 1541
box 0 0 1 1
use contact_21  contact_21_529
timestamp 1643671299
transform 1 0 36201 0 1 1523
box 0 0 1 1
use contact_13  contact_13_530
timestamp 1643671299
transform 1 0 35861 0 1 1541
box 0 0 1 1
use contact_21  contact_21_530
timestamp 1643671299
transform 1 0 35865 0 1 1523
box 0 0 1 1
use contact_18  contact_18_107
timestamp 1643671299
transform 1 0 35524 0 1 1534
box 0 0 1 1
use contact_17  contact_17_269
timestamp 1643671299
transform 1 0 35539 0 1 1549
box 0 0 1 1
use contact_13  contact_13_531
timestamp 1643671299
transform 1 0 35525 0 1 1541
box 0 0 1 1
use contact_21  contact_21_531
timestamp 1643671299
transform 1 0 35529 0 1 1523
box 0 0 1 1
use contact_13  contact_13_532
timestamp 1643671299
transform 1 0 35189 0 1 1541
box 0 0 1 1
use contact_21  contact_21_532
timestamp 1643671299
transform 1 0 35193 0 1 1523
box 0 0 1 1
use contact_13  contact_13_533
timestamp 1643671299
transform 1 0 34853 0 1 1541
box 0 0 1 1
use contact_21  contact_21_533
timestamp 1643671299
transform 1 0 34857 0 1 1523
box 0 0 1 1
use contact_13  contact_13_534
timestamp 1643671299
transform 1 0 34517 0 1 1541
box 0 0 1 1
use contact_21  contact_21_534
timestamp 1643671299
transform 1 0 34521 0 1 1523
box 0 0 1 1
use contact_13  contact_13_535
timestamp 1643671299
transform 1 0 34181 0 1 1541
box 0 0 1 1
use contact_21  contact_21_535
timestamp 1643671299
transform 1 0 34185 0 1 1523
box 0 0 1 1
use contact_18  contact_18_108
timestamp 1643671299
transform 1 0 33844 0 1 1534
box 0 0 1 1
use contact_17  contact_17_270
timestamp 1643671299
transform 1 0 33859 0 1 1549
box 0 0 1 1
use contact_13  contact_13_536
timestamp 1643671299
transform 1 0 33845 0 1 1541
box 0 0 1 1
use contact_21  contact_21_536
timestamp 1643671299
transform 1 0 33849 0 1 1523
box 0 0 1 1
use contact_13  contact_13_537
timestamp 1643671299
transform 1 0 33509 0 1 1541
box 0 0 1 1
use contact_21  contact_21_537
timestamp 1643671299
transform 1 0 33513 0 1 1523
box 0 0 1 1
use contact_13  contact_13_538
timestamp 1643671299
transform 1 0 33173 0 1 1541
box 0 0 1 1
use contact_21  contact_21_538
timestamp 1643671299
transform 1 0 33177 0 1 1523
box 0 0 1 1
use contact_13  contact_13_539
timestamp 1643671299
transform 1 0 32837 0 1 1541
box 0 0 1 1
use contact_21  contact_21_539
timestamp 1643671299
transform 1 0 32841 0 1 1523
box 0 0 1 1
use contact_13  contact_13_540
timestamp 1643671299
transform 1 0 32501 0 1 1541
box 0 0 1 1
use contact_21  contact_21_540
timestamp 1643671299
transform 1 0 32505 0 1 1523
box 0 0 1 1
use contact_18  contact_18_109
timestamp 1643671299
transform 1 0 32164 0 1 1534
box 0 0 1 1
use contact_17  contact_17_271
timestamp 1643671299
transform 1 0 32179 0 1 1549
box 0 0 1 1
use contact_13  contact_13_541
timestamp 1643671299
transform 1 0 32165 0 1 1541
box 0 0 1 1
use contact_21  contact_21_541
timestamp 1643671299
transform 1 0 32169 0 1 1523
box 0 0 1 1
use contact_13  contact_13_542
timestamp 1643671299
transform 1 0 31829 0 1 1541
box 0 0 1 1
use contact_21  contact_21_542
timestamp 1643671299
transform 1 0 31833 0 1 1523
box 0 0 1 1
use contact_13  contact_13_543
timestamp 1643671299
transform 1 0 31493 0 1 1541
box 0 0 1 1
use contact_21  contact_21_543
timestamp 1643671299
transform 1 0 31497 0 1 1523
box 0 0 1 1
use contact_13  contact_13_544
timestamp 1643671299
transform 1 0 31157 0 1 1541
box 0 0 1 1
use contact_21  contact_21_544
timestamp 1643671299
transform 1 0 31161 0 1 1523
box 0 0 1 1
use contact_13  contact_13_545
timestamp 1643671299
transform 1 0 30821 0 1 1541
box 0 0 1 1
use contact_21  contact_21_545
timestamp 1643671299
transform 1 0 30825 0 1 1523
box 0 0 1 1
use contact_18  contact_18_110
timestamp 1643671299
transform 1 0 30484 0 1 1534
box 0 0 1 1
use contact_17  contact_17_272
timestamp 1643671299
transform 1 0 30499 0 1 1549
box 0 0 1 1
use contact_13  contact_13_546
timestamp 1643671299
transform 1 0 30485 0 1 1541
box 0 0 1 1
use contact_21  contact_21_546
timestamp 1643671299
transform 1 0 30489 0 1 1523
box 0 0 1 1
use contact_13  contact_13_547
timestamp 1643671299
transform 1 0 30149 0 1 1541
box 0 0 1 1
use contact_21  contact_21_547
timestamp 1643671299
transform 1 0 30153 0 1 1523
box 0 0 1 1
use contact_13  contact_13_548
timestamp 1643671299
transform 1 0 29813 0 1 1541
box 0 0 1 1
use contact_21  contact_21_548
timestamp 1643671299
transform 1 0 29817 0 1 1523
box 0 0 1 1
use contact_13  contact_13_549
timestamp 1643671299
transform 1 0 29477 0 1 1541
box 0 0 1 1
use contact_21  contact_21_549
timestamp 1643671299
transform 1 0 29481 0 1 1523
box 0 0 1 1
use contact_13  contact_13_550
timestamp 1643671299
transform 1 0 29141 0 1 1541
box 0 0 1 1
use contact_21  contact_21_550
timestamp 1643671299
transform 1 0 29145 0 1 1523
box 0 0 1 1
use contact_18  contact_18_111
timestamp 1643671299
transform 1 0 28804 0 1 1534
box 0 0 1 1
use contact_17  contact_17_273
timestamp 1643671299
transform 1 0 28819 0 1 1549
box 0 0 1 1
use contact_13  contact_13_551
timestamp 1643671299
transform 1 0 28805 0 1 1541
box 0 0 1 1
use contact_21  contact_21_551
timestamp 1643671299
transform 1 0 28809 0 1 1523
box 0 0 1 1
use contact_13  contact_13_552
timestamp 1643671299
transform 1 0 28469 0 1 1541
box 0 0 1 1
use contact_21  contact_21_552
timestamp 1643671299
transform 1 0 28473 0 1 1523
box 0 0 1 1
use contact_13  contact_13_553
timestamp 1643671299
transform 1 0 28133 0 1 1541
box 0 0 1 1
use contact_21  contact_21_553
timestamp 1643671299
transform 1 0 28137 0 1 1523
box 0 0 1 1
use contact_13  contact_13_554
timestamp 1643671299
transform 1 0 27797 0 1 1541
box 0 0 1 1
use contact_21  contact_21_554
timestamp 1643671299
transform 1 0 27801 0 1 1523
box 0 0 1 1
use contact_13  contact_13_555
timestamp 1643671299
transform 1 0 27461 0 1 1541
box 0 0 1 1
use contact_21  contact_21_555
timestamp 1643671299
transform 1 0 27465 0 1 1523
box 0 0 1 1
use contact_18  contact_18_112
timestamp 1643671299
transform 1 0 27124 0 1 1534
box 0 0 1 1
use contact_17  contact_17_274
timestamp 1643671299
transform 1 0 27139 0 1 1549
box 0 0 1 1
use contact_13  contact_13_556
timestamp 1643671299
transform 1 0 27125 0 1 1541
box 0 0 1 1
use contact_21  contact_21_556
timestamp 1643671299
transform 1 0 27129 0 1 1523
box 0 0 1 1
use contact_13  contact_13_557
timestamp 1643671299
transform 1 0 26789 0 1 1541
box 0 0 1 1
use contact_21  contact_21_557
timestamp 1643671299
transform 1 0 26793 0 1 1523
box 0 0 1 1
use contact_13  contact_13_558
timestamp 1643671299
transform 1 0 26453 0 1 1541
box 0 0 1 1
use contact_21  contact_21_558
timestamp 1643671299
transform 1 0 26457 0 1 1523
box 0 0 1 1
use contact_13  contact_13_559
timestamp 1643671299
transform 1 0 26117 0 1 1541
box 0 0 1 1
use contact_21  contact_21_559
timestamp 1643671299
transform 1 0 26121 0 1 1523
box 0 0 1 1
use contact_13  contact_13_560
timestamp 1643671299
transform 1 0 25781 0 1 1541
box 0 0 1 1
use contact_21  contact_21_560
timestamp 1643671299
transform 1 0 25785 0 1 1523
box 0 0 1 1
use contact_18  contact_18_113
timestamp 1643671299
transform 1 0 25444 0 1 1534
box 0 0 1 1
use contact_17  contact_17_275
timestamp 1643671299
transform 1 0 25459 0 1 1549
box 0 0 1 1
use contact_13  contact_13_561
timestamp 1643671299
transform 1 0 25445 0 1 1541
box 0 0 1 1
use contact_21  contact_21_561
timestamp 1643671299
transform 1 0 25449 0 1 1523
box 0 0 1 1
use contact_13  contact_13_562
timestamp 1643671299
transform 1 0 25109 0 1 1541
box 0 0 1 1
use contact_21  contact_21_562
timestamp 1643671299
transform 1 0 25113 0 1 1523
box 0 0 1 1
use contact_13  contact_13_563
timestamp 1643671299
transform 1 0 24773 0 1 1541
box 0 0 1 1
use contact_21  contact_21_563
timestamp 1643671299
transform 1 0 24777 0 1 1523
box 0 0 1 1
use contact_13  contact_13_564
timestamp 1643671299
transform 1 0 24437 0 1 1541
box 0 0 1 1
use contact_21  contact_21_564
timestamp 1643671299
transform 1 0 24441 0 1 1523
box 0 0 1 1
use contact_13  contact_13_565
timestamp 1643671299
transform 1 0 24101 0 1 1541
box 0 0 1 1
use contact_21  contact_21_565
timestamp 1643671299
transform 1 0 24105 0 1 1523
box 0 0 1 1
use contact_18  contact_18_114
timestamp 1643671299
transform 1 0 23764 0 1 1534
box 0 0 1 1
use contact_17  contact_17_276
timestamp 1643671299
transform 1 0 23779 0 1 1549
box 0 0 1 1
use contact_13  contact_13_566
timestamp 1643671299
transform 1 0 23765 0 1 1541
box 0 0 1 1
use contact_21  contact_21_566
timestamp 1643671299
transform 1 0 23769 0 1 1523
box 0 0 1 1
use contact_13  contact_13_567
timestamp 1643671299
transform 1 0 23429 0 1 1541
box 0 0 1 1
use contact_21  contact_21_567
timestamp 1643671299
transform 1 0 23433 0 1 1523
box 0 0 1 1
use contact_13  contact_13_568
timestamp 1643671299
transform 1 0 23093 0 1 1541
box 0 0 1 1
use contact_21  contact_21_568
timestamp 1643671299
transform 1 0 23097 0 1 1523
box 0 0 1 1
use contact_13  contact_13_569
timestamp 1643671299
transform 1 0 22757 0 1 1541
box 0 0 1 1
use contact_21  contact_21_569
timestamp 1643671299
transform 1 0 22761 0 1 1523
box 0 0 1 1
use contact_13  contact_13_570
timestamp 1643671299
transform 1 0 22421 0 1 1541
box 0 0 1 1
use contact_21  contact_21_570
timestamp 1643671299
transform 1 0 22425 0 1 1523
box 0 0 1 1
use contact_18  contact_18_115
timestamp 1643671299
transform 1 0 22084 0 1 1534
box 0 0 1 1
use contact_17  contact_17_277
timestamp 1643671299
transform 1 0 22099 0 1 1549
box 0 0 1 1
use contact_13  contact_13_571
timestamp 1643671299
transform 1 0 22085 0 1 1541
box 0 0 1 1
use contact_21  contact_21_571
timestamp 1643671299
transform 1 0 22089 0 1 1523
box 0 0 1 1
use contact_13  contact_13_572
timestamp 1643671299
transform 1 0 21749 0 1 1541
box 0 0 1 1
use contact_21  contact_21_572
timestamp 1643671299
transform 1 0 21753 0 1 1523
box 0 0 1 1
use contact_13  contact_13_573
timestamp 1643671299
transform 1 0 21413 0 1 1541
box 0 0 1 1
use contact_21  contact_21_573
timestamp 1643671299
transform 1 0 21417 0 1 1523
box 0 0 1 1
use contact_13  contact_13_574
timestamp 1643671299
transform 1 0 21077 0 1 1541
box 0 0 1 1
use contact_21  contact_21_574
timestamp 1643671299
transform 1 0 21081 0 1 1523
box 0 0 1 1
use contact_13  contact_13_575
timestamp 1643671299
transform 1 0 20741 0 1 1541
box 0 0 1 1
use contact_21  contact_21_575
timestamp 1643671299
transform 1 0 20745 0 1 1523
box 0 0 1 1
use contact_18  contact_18_116
timestamp 1643671299
transform 1 0 20404 0 1 1534
box 0 0 1 1
use contact_17  contact_17_278
timestamp 1643671299
transform 1 0 20419 0 1 1549
box 0 0 1 1
use contact_13  contact_13_576
timestamp 1643671299
transform 1 0 20405 0 1 1541
box 0 0 1 1
use contact_21  contact_21_576
timestamp 1643671299
transform 1 0 20409 0 1 1523
box 0 0 1 1
use contact_13  contact_13_577
timestamp 1643671299
transform 1 0 20069 0 1 1541
box 0 0 1 1
use contact_21  contact_21_577
timestamp 1643671299
transform 1 0 20073 0 1 1523
box 0 0 1 1
use contact_13  contact_13_578
timestamp 1643671299
transform 1 0 19733 0 1 1541
box 0 0 1 1
use contact_21  contact_21_578
timestamp 1643671299
transform 1 0 19737 0 1 1523
box 0 0 1 1
use contact_13  contact_13_579
timestamp 1643671299
transform 1 0 19397 0 1 1541
box 0 0 1 1
use contact_21  contact_21_579
timestamp 1643671299
transform 1 0 19401 0 1 1523
box 0 0 1 1
use contact_13  contact_13_580
timestamp 1643671299
transform 1 0 19061 0 1 1541
box 0 0 1 1
use contact_21  contact_21_580
timestamp 1643671299
transform 1 0 19065 0 1 1523
box 0 0 1 1
use contact_18  contact_18_117
timestamp 1643671299
transform 1 0 18724 0 1 1534
box 0 0 1 1
use contact_17  contact_17_279
timestamp 1643671299
transform 1 0 18739 0 1 1549
box 0 0 1 1
use contact_13  contact_13_581
timestamp 1643671299
transform 1 0 18725 0 1 1541
box 0 0 1 1
use contact_21  contact_21_581
timestamp 1643671299
transform 1 0 18729 0 1 1523
box 0 0 1 1
use contact_13  contact_13_582
timestamp 1643671299
transform 1 0 18389 0 1 1541
box 0 0 1 1
use contact_21  contact_21_582
timestamp 1643671299
transform 1 0 18393 0 1 1523
box 0 0 1 1
use contact_13  contact_13_583
timestamp 1643671299
transform 1 0 18053 0 1 1541
box 0 0 1 1
use contact_21  contact_21_583
timestamp 1643671299
transform 1 0 18057 0 1 1523
box 0 0 1 1
use contact_13  contact_13_584
timestamp 1643671299
transform 1 0 17717 0 1 1541
box 0 0 1 1
use contact_21  contact_21_584
timestamp 1643671299
transform 1 0 17721 0 1 1523
box 0 0 1 1
use contact_13  contact_13_585
timestamp 1643671299
transform 1 0 17381 0 1 1541
box 0 0 1 1
use contact_21  contact_21_585
timestamp 1643671299
transform 1 0 17385 0 1 1523
box 0 0 1 1
use contact_18  contact_18_118
timestamp 1643671299
transform 1 0 17044 0 1 1534
box 0 0 1 1
use contact_17  contact_17_280
timestamp 1643671299
transform 1 0 17059 0 1 1549
box 0 0 1 1
use contact_13  contact_13_586
timestamp 1643671299
transform 1 0 17045 0 1 1541
box 0 0 1 1
use contact_21  contact_21_586
timestamp 1643671299
transform 1 0 17049 0 1 1523
box 0 0 1 1
use contact_13  contact_13_587
timestamp 1643671299
transform 1 0 16709 0 1 1541
box 0 0 1 1
use contact_21  contact_21_587
timestamp 1643671299
transform 1 0 16713 0 1 1523
box 0 0 1 1
use contact_13  contact_13_588
timestamp 1643671299
transform 1 0 16373 0 1 1541
box 0 0 1 1
use contact_21  contact_21_588
timestamp 1643671299
transform 1 0 16377 0 1 1523
box 0 0 1 1
use contact_13  contact_13_589
timestamp 1643671299
transform 1 0 16037 0 1 1541
box 0 0 1 1
use contact_21  contact_21_589
timestamp 1643671299
transform 1 0 16041 0 1 1523
box 0 0 1 1
use contact_13  contact_13_590
timestamp 1643671299
transform 1 0 15701 0 1 1541
box 0 0 1 1
use contact_21  contact_21_590
timestamp 1643671299
transform 1 0 15705 0 1 1523
box 0 0 1 1
use contact_18  contact_18_119
timestamp 1643671299
transform 1 0 15364 0 1 1534
box 0 0 1 1
use contact_17  contact_17_281
timestamp 1643671299
transform 1 0 15379 0 1 1549
box 0 0 1 1
use contact_13  contact_13_591
timestamp 1643671299
transform 1 0 15365 0 1 1541
box 0 0 1 1
use contact_21  contact_21_591
timestamp 1643671299
transform 1 0 15369 0 1 1523
box 0 0 1 1
use contact_13  contact_13_592
timestamp 1643671299
transform 1 0 15029 0 1 1541
box 0 0 1 1
use contact_21  contact_21_592
timestamp 1643671299
transform 1 0 15033 0 1 1523
box 0 0 1 1
use contact_13  contact_13_593
timestamp 1643671299
transform 1 0 14693 0 1 1541
box 0 0 1 1
use contact_21  contact_21_593
timestamp 1643671299
transform 1 0 14697 0 1 1523
box 0 0 1 1
use contact_13  contact_13_594
timestamp 1643671299
transform 1 0 14357 0 1 1541
box 0 0 1 1
use contact_21  contact_21_594
timestamp 1643671299
transform 1 0 14361 0 1 1523
box 0 0 1 1
use contact_13  contact_13_595
timestamp 1643671299
transform 1 0 14021 0 1 1541
box 0 0 1 1
use contact_21  contact_21_595
timestamp 1643671299
transform 1 0 14025 0 1 1523
box 0 0 1 1
use contact_18  contact_18_120
timestamp 1643671299
transform 1 0 13684 0 1 1534
box 0 0 1 1
use contact_17  contact_17_282
timestamp 1643671299
transform 1 0 13699 0 1 1549
box 0 0 1 1
use contact_13  contact_13_596
timestamp 1643671299
transform 1 0 13685 0 1 1541
box 0 0 1 1
use contact_21  contact_21_596
timestamp 1643671299
transform 1 0 13689 0 1 1523
box 0 0 1 1
use contact_13  contact_13_597
timestamp 1643671299
transform 1 0 13349 0 1 1541
box 0 0 1 1
use contact_21  contact_21_597
timestamp 1643671299
transform 1 0 13353 0 1 1523
box 0 0 1 1
use contact_13  contact_13_598
timestamp 1643671299
transform 1 0 13013 0 1 1541
box 0 0 1 1
use contact_21  contact_21_598
timestamp 1643671299
transform 1 0 13017 0 1 1523
box 0 0 1 1
use contact_13  contact_13_599
timestamp 1643671299
transform 1 0 12677 0 1 1541
box 0 0 1 1
use contact_21  contact_21_599
timestamp 1643671299
transform 1 0 12681 0 1 1523
box 0 0 1 1
use contact_13  contact_13_600
timestamp 1643671299
transform 1 0 12341 0 1 1541
box 0 0 1 1
use contact_21  contact_21_600
timestamp 1643671299
transform 1 0 12345 0 1 1523
box 0 0 1 1
use contact_18  contact_18_121
timestamp 1643671299
transform 1 0 12004 0 1 1534
box 0 0 1 1
use contact_17  contact_17_283
timestamp 1643671299
transform 1 0 12019 0 1 1549
box 0 0 1 1
use contact_13  contact_13_601
timestamp 1643671299
transform 1 0 12005 0 1 1541
box 0 0 1 1
use contact_21  contact_21_601
timestamp 1643671299
transform 1 0 12009 0 1 1523
box 0 0 1 1
use contact_13  contact_13_602
timestamp 1643671299
transform 1 0 11669 0 1 1541
box 0 0 1 1
use contact_21  contact_21_602
timestamp 1643671299
transform 1 0 11673 0 1 1523
box 0 0 1 1
use contact_13  contact_13_603
timestamp 1643671299
transform 1 0 11333 0 1 1541
box 0 0 1 1
use contact_21  contact_21_603
timestamp 1643671299
transform 1 0 11337 0 1 1523
box 0 0 1 1
use contact_13  contact_13_604
timestamp 1643671299
transform 1 0 10997 0 1 1541
box 0 0 1 1
use contact_21  contact_21_604
timestamp 1643671299
transform 1 0 11001 0 1 1523
box 0 0 1 1
use contact_13  contact_13_605
timestamp 1643671299
transform 1 0 10661 0 1 1541
box 0 0 1 1
use contact_21  contact_21_605
timestamp 1643671299
transform 1 0 10665 0 1 1523
box 0 0 1 1
use contact_18  contact_18_122
timestamp 1643671299
transform 1 0 10324 0 1 1534
box 0 0 1 1
use contact_17  contact_17_284
timestamp 1643671299
transform 1 0 10339 0 1 1549
box 0 0 1 1
use contact_13  contact_13_606
timestamp 1643671299
transform 1 0 10325 0 1 1541
box 0 0 1 1
use contact_21  contact_21_606
timestamp 1643671299
transform 1 0 10329 0 1 1523
box 0 0 1 1
use contact_13  contact_13_607
timestamp 1643671299
transform 1 0 9989 0 1 1541
box 0 0 1 1
use contact_21  contact_21_607
timestamp 1643671299
transform 1 0 9993 0 1 1523
box 0 0 1 1
use contact_13  contact_13_608
timestamp 1643671299
transform 1 0 9653 0 1 1541
box 0 0 1 1
use contact_21  contact_21_608
timestamp 1643671299
transform 1 0 9657 0 1 1523
box 0 0 1 1
use contact_13  contact_13_609
timestamp 1643671299
transform 1 0 9317 0 1 1541
box 0 0 1 1
use contact_21  contact_21_609
timestamp 1643671299
transform 1 0 9321 0 1 1523
box 0 0 1 1
use contact_13  contact_13_610
timestamp 1643671299
transform 1 0 8981 0 1 1541
box 0 0 1 1
use contact_21  contact_21_610
timestamp 1643671299
transform 1 0 8985 0 1 1523
box 0 0 1 1
use contact_18  contact_18_123
timestamp 1643671299
transform 1 0 8644 0 1 1534
box 0 0 1 1
use contact_17  contact_17_285
timestamp 1643671299
transform 1 0 8659 0 1 1549
box 0 0 1 1
use contact_13  contact_13_611
timestamp 1643671299
transform 1 0 8645 0 1 1541
box 0 0 1 1
use contact_21  contact_21_611
timestamp 1643671299
transform 1 0 8649 0 1 1523
box 0 0 1 1
use contact_13  contact_13_612
timestamp 1643671299
transform 1 0 8309 0 1 1541
box 0 0 1 1
use contact_21  contact_21_612
timestamp 1643671299
transform 1 0 8313 0 1 1523
box 0 0 1 1
use contact_13  contact_13_613
timestamp 1643671299
transform 1 0 7973 0 1 1541
box 0 0 1 1
use contact_21  contact_21_613
timestamp 1643671299
transform 1 0 7977 0 1 1523
box 0 0 1 1
use contact_13  contact_13_614
timestamp 1643671299
transform 1 0 7637 0 1 1541
box 0 0 1 1
use contact_21  contact_21_614
timestamp 1643671299
transform 1 0 7641 0 1 1523
box 0 0 1 1
use contact_13  contact_13_615
timestamp 1643671299
transform 1 0 7301 0 1 1541
box 0 0 1 1
use contact_21  contact_21_615
timestamp 1643671299
transform 1 0 7305 0 1 1523
box 0 0 1 1
use contact_18  contact_18_124
timestamp 1643671299
transform 1 0 6964 0 1 1534
box 0 0 1 1
use contact_17  contact_17_286
timestamp 1643671299
transform 1 0 6979 0 1 1549
box 0 0 1 1
use contact_13  contact_13_616
timestamp 1643671299
transform 1 0 6965 0 1 1541
box 0 0 1 1
use contact_21  contact_21_616
timestamp 1643671299
transform 1 0 6969 0 1 1523
box 0 0 1 1
use contact_13  contact_13_617
timestamp 1643671299
transform 1 0 6629 0 1 1541
box 0 0 1 1
use contact_21  contact_21_617
timestamp 1643671299
transform 1 0 6633 0 1 1523
box 0 0 1 1
use contact_13  contact_13_618
timestamp 1643671299
transform 1 0 6293 0 1 1541
box 0 0 1 1
use contact_21  contact_21_618
timestamp 1643671299
transform 1 0 6297 0 1 1523
box 0 0 1 1
use contact_13  contact_13_619
timestamp 1643671299
transform 1 0 5957 0 1 1541
box 0 0 1 1
use contact_21  contact_21_619
timestamp 1643671299
transform 1 0 5961 0 1 1523
box 0 0 1 1
use contact_13  contact_13_620
timestamp 1643671299
transform 1 0 5621 0 1 1541
box 0 0 1 1
use contact_21  contact_21_620
timestamp 1643671299
transform 1 0 5625 0 1 1523
box 0 0 1 1
use contact_18  contact_18_125
timestamp 1643671299
transform 1 0 5284 0 1 1534
box 0 0 1 1
use contact_17  contact_17_287
timestamp 1643671299
transform 1 0 5299 0 1 1549
box 0 0 1 1
use contact_13  contact_13_621
timestamp 1643671299
transform 1 0 5285 0 1 1541
box 0 0 1 1
use contact_21  contact_21_621
timestamp 1643671299
transform 1 0 5289 0 1 1523
box 0 0 1 1
use contact_13  contact_13_622
timestamp 1643671299
transform 1 0 4949 0 1 1541
box 0 0 1 1
use contact_21  contact_21_622
timestamp 1643671299
transform 1 0 4953 0 1 1523
box 0 0 1 1
use contact_13  contact_13_623
timestamp 1643671299
transform 1 0 4613 0 1 1541
box 0 0 1 1
use contact_21  contact_21_623
timestamp 1643671299
transform 1 0 4617 0 1 1523
box 0 0 1 1
use contact_13  contact_13_624
timestamp 1643671299
transform 1 0 4277 0 1 1541
box 0 0 1 1
use contact_21  contact_21_624
timestamp 1643671299
transform 1 0 4281 0 1 1523
box 0 0 1 1
use contact_13  contact_13_625
timestamp 1643671299
transform 1 0 3941 0 1 1541
box 0 0 1 1
use contact_21  contact_21_625
timestamp 1643671299
transform 1 0 3945 0 1 1523
box 0 0 1 1
use contact_18  contact_18_126
timestamp 1643671299
transform 1 0 3604 0 1 1534
box 0 0 1 1
use contact_17  contact_17_288
timestamp 1643671299
transform 1 0 3619 0 1 1549
box 0 0 1 1
use contact_13  contact_13_626
timestamp 1643671299
transform 1 0 3605 0 1 1541
box 0 0 1 1
use contact_21  contact_21_626
timestamp 1643671299
transform 1 0 3609 0 1 1523
box 0 0 1 1
use contact_13  contact_13_627
timestamp 1643671299
transform 1 0 3269 0 1 1541
box 0 0 1 1
use contact_21  contact_21_627
timestamp 1643671299
transform 1 0 3273 0 1 1523
box 0 0 1 1
use contact_13  contact_13_628
timestamp 1643671299
transform 1 0 2933 0 1 1541
box 0 0 1 1
use contact_21  contact_21_628
timestamp 1643671299
transform 1 0 2937 0 1 1523
box 0 0 1 1
use contact_13  contact_13_629
timestamp 1643671299
transform 1 0 2597 0 1 1541
box 0 0 1 1
use contact_21  contact_21_629
timestamp 1643671299
transform 1 0 2601 0 1 1523
box 0 0 1 1
use contact_13  contact_13_630
timestamp 1643671299
transform 1 0 2261 0 1 1541
box 0 0 1 1
use contact_21  contact_21_630
timestamp 1643671299
transform 1 0 2265 0 1 1523
box 0 0 1 1
use contact_18  contact_18_127
timestamp 1643671299
transform 1 0 1924 0 1 1534
box 0 0 1 1
use contact_17  contact_17_289
timestamp 1643671299
transform 1 0 1939 0 1 1549
box 0 0 1 1
use contact_13  contact_13_631
timestamp 1643671299
transform 1 0 1925 0 1 1541
box 0 0 1 1
use contact_21  contact_21_631
timestamp 1643671299
transform 1 0 1929 0 1 1523
box 0 0 1 1
use contact_18  contact_18_128
timestamp 1643671299
transform 1 0 12389 0 1 15512
box 0 0 1 1
use contact_18  contact_18_129
timestamp 1643671299
transform 1 0 12389 0 1 14328
box 0 0 1 1
use contact_18  contact_18_130
timestamp 1643671299
transform 1 0 12389 0 1 13836
box 0 0 1 1
use contact_18  contact_18_131
timestamp 1643671299
transform 1 0 12389 0 1 12652
box 0 0 1 1
use contact_18  contact_18_132
timestamp 1643671299
transform 1 0 12389 0 1 12160
box 0 0 1 1
use contact_18  contact_18_133
timestamp 1643671299
transform 1 0 12389 0 1 10976
box 0 0 1 1
use contact_18  contact_18_134
timestamp 1643671299
transform 1 0 15353 0 1 2620
box 0 0 1 1
use contact_18  contact_18_135
timestamp 1643671299
transform 1 0 48060 0 1 9250
box 0 0 1 1
use contact_18  contact_18_136
timestamp 1643671299
transform 1 0 48060 0 1 9250
box 0 0 1 1
use contact_18  contact_18_137
timestamp 1643671299
transform 1 0 46504 0 1 9250
box 0 0 1 1
use contact_18  contact_18_138
timestamp 1643671299
transform 1 0 46504 0 1 9250
box 0 0 1 1
use contact_18  contact_18_139
timestamp 1643671299
transform 1 0 44948 0 1 9250
box 0 0 1 1
use contact_18  contact_18_140
timestamp 1643671299
transform 1 0 44948 0 1 9250
box 0 0 1 1
use contact_18  contact_18_141
timestamp 1643671299
transform 1 0 43392 0 1 9250
box 0 0 1 1
use contact_18  contact_18_142
timestamp 1643671299
transform 1 0 43392 0 1 9250
box 0 0 1 1
use contact_18  contact_18_143
timestamp 1643671299
transform 1 0 41836 0 1 9250
box 0 0 1 1
use contact_18  contact_18_144
timestamp 1643671299
transform 1 0 41836 0 1 9250
box 0 0 1 1
use contact_18  contact_18_145
timestamp 1643671299
transform 1 0 40280 0 1 9250
box 0 0 1 1
use contact_18  contact_18_146
timestamp 1643671299
transform 1 0 40280 0 1 9250
box 0 0 1 1
use contact_18  contact_18_147
timestamp 1643671299
transform 1 0 38724 0 1 9250
box 0 0 1 1
use contact_18  contact_18_148
timestamp 1643671299
transform 1 0 38724 0 1 9250
box 0 0 1 1
use contact_18  contact_18_149
timestamp 1643671299
transform 1 0 37168 0 1 9250
box 0 0 1 1
use contact_18  contact_18_150
timestamp 1643671299
transform 1 0 37168 0 1 9250
box 0 0 1 1
use contact_18  contact_18_151
timestamp 1643671299
transform 1 0 35612 0 1 9250
box 0 0 1 1
use contact_18  contact_18_152
timestamp 1643671299
transform 1 0 35612 0 1 9250
box 0 0 1 1
use contact_18  contact_18_153
timestamp 1643671299
transform 1 0 34056 0 1 9250
box 0 0 1 1
use contact_18  contact_18_154
timestamp 1643671299
transform 1 0 34056 0 1 9250
box 0 0 1 1
use contact_18  contact_18_155
timestamp 1643671299
transform 1 0 32500 0 1 9250
box 0 0 1 1
use contact_18  contact_18_156
timestamp 1643671299
transform 1 0 32500 0 1 9250
box 0 0 1 1
use contact_18  contact_18_157
timestamp 1643671299
transform 1 0 30944 0 1 9250
box 0 0 1 1
use contact_18  contact_18_158
timestamp 1643671299
transform 1 0 30944 0 1 9250
box 0 0 1 1
use contact_18  contact_18_159
timestamp 1643671299
transform 1 0 29388 0 1 9250
box 0 0 1 1
use contact_18  contact_18_160
timestamp 1643671299
transform 1 0 29388 0 1 9250
box 0 0 1 1
use contact_18  contact_18_161
timestamp 1643671299
transform 1 0 27832 0 1 9250
box 0 0 1 1
use contact_18  contact_18_162
timestamp 1643671299
transform 1 0 27832 0 1 9250
box 0 0 1 1
use contact_18  contact_18_163
timestamp 1643671299
transform 1 0 26276 0 1 9250
box 0 0 1 1
use contact_18  contact_18_164
timestamp 1643671299
transform 1 0 26276 0 1 9250
box 0 0 1 1
use contact_18  contact_18_165
timestamp 1643671299
transform 1 0 24720 0 1 9250
box 0 0 1 1
use contact_18  contact_18_166
timestamp 1643671299
transform 1 0 24720 0 1 9250
box 0 0 1 1
use contact_18  contact_18_167
timestamp 1643671299
transform 1 0 39065 0 1 2620
box 0 0 1 1
use contact_18  contact_18_168
timestamp 1643671299
transform 1 0 37583 0 1 2620
box 0 0 1 1
use contact_18  contact_18_169
timestamp 1643671299
transform 1 0 36101 0 1 2620
box 0 0 1 1
use contact_18  contact_18_170
timestamp 1643671299
transform 1 0 34619 0 1 2620
box 0 0 1 1
use contact_18  contact_18_171
timestamp 1643671299
transform 1 0 33137 0 1 2620
box 0 0 1 1
use contact_18  contact_18_172
timestamp 1643671299
transform 1 0 31655 0 1 2620
box 0 0 1 1
use contact_18  contact_18_173
timestamp 1643671299
transform 1 0 30173 0 1 2620
box 0 0 1 1
use contact_18  contact_18_174
timestamp 1643671299
transform 1 0 28691 0 1 2620
box 0 0 1 1
use contact_18  contact_18_175
timestamp 1643671299
transform 1 0 27209 0 1 2620
box 0 0 1 1
use contact_18  contact_18_176
timestamp 1643671299
transform 1 0 25727 0 1 2620
box 0 0 1 1
use contact_18  contact_18_177
timestamp 1643671299
transform 1 0 24245 0 1 2620
box 0 0 1 1
use contact_18  contact_18_178
timestamp 1643671299
transform 1 0 22763 0 1 2620
box 0 0 1 1
use contact_18  contact_18_179
timestamp 1643671299
transform 1 0 21281 0 1 2620
box 0 0 1 1
use contact_18  contact_18_180
timestamp 1643671299
transform 1 0 19799 0 1 2620
box 0 0 1 1
use contact_18  contact_18_181
timestamp 1643671299
transform 1 0 18317 0 1 2620
box 0 0 1 1
use contact_18  contact_18_182
timestamp 1643671299
transform 1 0 16835 0 1 2620
box 0 0 1 1
use contact_18  contact_18_183
timestamp 1643671299
transform 1 0 5995 0 1 5823
box 0 0 1 1
use contact_18  contact_18_184
timestamp 1643671299
transform 1 0 2635 0 1 6038
box 0 0 1 1
use contact_18  contact_18_185
timestamp 1643671299
transform 1 0 2635 0 1 4854
box 0 0 1 1
use contact_18  contact_18_186
timestamp 1643671299
transform 1 0 14155 0 1 15516
box 0 0 1 1
use contact_18  contact_18_187
timestamp 1643671299
transform 1 0 13469 0 1 15516
box 0 0 1 1
use contact_18  contact_18_188
timestamp 1643671299
transform 1 0 14087 0 1 14324
box 0 0 1 1
use contact_18  contact_18_189
timestamp 1643671299
transform 1 0 13469 0 1 14324
box 0 0 1 1
use contact_18  contact_18_190
timestamp 1643671299
transform 1 0 14019 0 1 13840
box 0 0 1 1
use contact_18  contact_18_191
timestamp 1643671299
transform 1 0 13469 0 1 13840
box 0 0 1 1
use contact_18  contact_18_192
timestamp 1643671299
transform 1 0 13951 0 1 12648
box 0 0 1 1
use contact_18  contact_18_193
timestamp 1643671299
transform 1 0 13469 0 1 12648
box 0 0 1 1
use contact_18  contact_18_194
timestamp 1643671299
transform 1 0 13883 0 1 12164
box 0 0 1 1
use contact_18  contact_18_195
timestamp 1643671299
transform 1 0 13469 0 1 12164
box 0 0 1 1
use contact_18  contact_18_196
timestamp 1643671299
transform 1 0 13815 0 1 10972
box 0 0 1 1
use contact_18  contact_18_197
timestamp 1643671299
transform 1 0 13469 0 1 10972
box 0 0 1 1
use contact_18  contact_18_198
timestamp 1643671299
transform 1 0 18476 0 1 10097
box 0 0 1 1
use contact_18  contact_18_199
timestamp 1643671299
transform 1 0 13664 0 1 10097
box 0 0 1 1
use contact_18  contact_18_200
timestamp 1643671299
transform 1 0 45166 0 1 9171
box 0 0 1 1
use contact_18  contact_18_201
timestamp 1643671299
transform 1 0 13664 0 1 9171
box 0 0 1 1
use contact_18  contact_18_202
timestamp 1643671299
transform 1 0 19610 0 1 8427
box 0 0 1 1
use contact_18  contact_18_203
timestamp 1643671299
transform 1 0 13664 0 1 8427
box 0 0 1 1
use contact_30  contact_30_0
timestamp 1643671299
transform 1 0 12114 0 1 2674
box 0 0 1 1
use contact_30  contact_30_1
timestamp 1643671299
transform 1 0 12114 0 1 2674
box 0 0 1 1
use contact_30  contact_30_2
timestamp 1643671299
transform 1 0 12114 0 1 11030
box 0 0 1 1
use data_dff  data_dff_0
timestamp 1643671299
transform 1 0 16658 0 1 2404
box -3 -42 23712 916
use col_addr_dff  col_addr_dff_0
timestamp 1643671299
transform 1 0 15176 0 1 2404
box -3 -42 1482 916
use row_addr_dff  row_addr_dff_0
timestamp 1643671299
transform 1 0 12212 0 1 10760
box -3 -42 1482 6746
use control_logic_multiport  control_logic_multiport_0
timestamp 1643671299
transform 1 0 2458 0 1 4638
box -30 -42 11236 5918
use bank  bank_0
timestamp 1643671299
transform 1 0 13830 0 1 4950
box -11 0 59212 30418
<< labels >>
rlabel metal3 s 2634 4854 2694 4914 4 web
rlabel metal3 s 2634 6038 2694 6098 4 csb
rlabel metal4 s 6000 0 6060 180 4 clk
rlabel metal4 s 16920 0 16980 180 4 din0[0]
rlabel metal4 s 18240 0 18300 180 4 din0[1]
rlabel metal4 s 19680 0 19740 180 4 din0[2]
rlabel metal4 s 21360 0 21420 180 4 din0[3]
rlabel metal4 s 22800 0 22860 180 4 din0[4]
rlabel metal4 s 24360 0 24420 180 4 din0[5]
rlabel metal4 s 25800 0 25860 180 4 din0[6]
rlabel metal4 s 27240 0 27300 180 4 din0[7]
rlabel metal4 s 28800 0 28860 180 4 din0[8]
rlabel metal4 s 30240 0 30300 180 4 din0[9]
rlabel metal4 s 31680 0 31740 180 4 din0[10]
rlabel metal4 s 33120 0 33180 180 4 din0[11]
rlabel metal4 s 34560 0 34620 180 4 din0[12]
rlabel metal4 s 36000 0 36060 180 4 din0[13]
rlabel metal4 s 37680 0 37740 180 4 din0[14]
rlabel metal4 s 39120 0 39180 180 4 din0[15]
rlabel metal4 s 24840 0 24900 180 4 dout0[0]
rlabel metal3 s 24720 9250 24780 9310 4 dout1[0]
rlabel metal4 s 26280 0 26340 180 4 dout0[1]
rlabel metal3 s 26276 9250 26336 9310 4 dout1[1]
rlabel metal4 s 27840 0 27900 180 4 dout0[2]
rlabel metal3 s 27832 9250 27892 9310 4 dout1[2]
rlabel metal4 s 29400 0 29460 180 4 dout0[3]
rlabel metal3 s 29388 9250 29448 9310 4 dout1[3]
rlabel metal4 s 30960 0 31020 180 4 dout0[4]
rlabel metal3 s 30944 9250 31004 9310 4 dout1[4]
rlabel metal4 s 32520 0 32580 180 4 dout0[5]
rlabel metal3 s 32500 9250 32560 9310 4 dout1[5]
rlabel metal4 s 34080 0 34140 180 4 dout0[6]
rlabel metal3 s 34056 9250 34116 9310 4 dout1[6]
rlabel metal4 s 35640 0 35700 180 4 dout0[7]
rlabel metal3 s 35612 9250 35672 9310 4 dout1[7]
rlabel metal4 s 37200 0 37260 180 4 dout0[8]
rlabel metal3 s 37168 9250 37228 9310 4 dout1[8]
rlabel metal4 s 38760 0 38820 180 4 dout0[9]
rlabel metal3 s 38724 9250 38784 9310 4 dout1[9]
rlabel metal4 s 40320 0 40380 180 4 dout0[10]
rlabel metal3 s 40280 9250 40340 9310 4 dout1[10]
rlabel metal4 s 41880 0 41940 180 4 dout0[11]
rlabel metal3 s 41836 9250 41896 9310 4 dout1[11]
rlabel metal4 s 43440 0 43500 180 4 dout0[12]
rlabel metal3 s 43392 9250 43452 9310 4 dout1[12]
rlabel metal4 s 45000 0 45060 180 4 dout0[13]
rlabel metal3 s 44948 9250 45008 9310 4 dout1[13]
rlabel metal4 s 46560 0 46620 180 4 dout0[14]
rlabel metal3 s 46504 9250 46564 9310 4 dout1[14]
rlabel metal4 s 48120 0 48180 180 4 dout0[15]
rlabel metal3 s 48060 9250 48120 9310 4 dout1[15]
rlabel metal4 s 15240 0 15300 180 4 addr0
rlabel metal4 s 12360 0 12420 180 4 addr1[1]
rlabel metal4 s 12480 0 12540 180 4 addr1[2]
rlabel metal3 s 0 12600 180 12660 4 addr1[3]
rlabel metal3 s 0 13800 180 13860 4 addr1[4]
rlabel metal3 s 0 14280 180 14340 4 addr1[5]
rlabel metal3 s 0 15480 180 15540 4 addr1[6]
rlabel metal4 s 74400 840 74700 36900 4 vdd
rlabel metal3 s 840 840 74700 1140 4 vdd
rlabel metal4 s 840 840 1140 36900 4 vdd
rlabel metal3 s 840 36600 74700 36900 4 vdd
rlabel metal4 s 240 240 540 37500 4 gnd
rlabel metal4 s 75000 240 75300 37500 4 gnd
rlabel metal3 s 240 37200 75300 37500 4 gnd
rlabel metal3 s 240 240 75300 540 4 gnd
<< properties >>
string FIXED_BBOX 0 0 75300 37500
string GDS_FILE sram_0rw2r1w_16_32_sky130A.gds
string GDS_END 318874
string GDS_START 126
<< end >>
