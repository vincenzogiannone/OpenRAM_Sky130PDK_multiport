magic
tech sky130A
magscale 1 2
timestamp 1644969367
<< checkpaint >>
rect -1296 -1277 5228 2155
<< nwell >>
rect -36 402 3968 895
<< locali >>
rect 0 821 3932 855
rect 48 336 114 402
rect 1911 352 1945 386
rect 0 -17 3932 17
use pinv_14  pinv_14_0
timestamp 1644969367
transform 1 0 0 0 1 0
box -36 -17 3968 895
<< labels >>
rlabel locali s 1928 369 1928 369 4 Z
rlabel locali s 81 369 81 369 4 A
rlabel locali s 1966 0 1966 0 4 gnd
rlabel locali s 1966 838 1966 838 4 vdd
<< properties >>
string FIXED_BBOX 0 0 3932 838
string GDS_FILE sram_0rw2r1w_32_128_sky130A.gds
string GDS_END 3394646
string GDS_START 3393800
<< end >>
