magic
tech sky130A
magscale 1 2
timestamp 1643671299
<< checkpaint >>
rect -1319 -1316 3629 1602
<< nwell >>
rect -54 228 2364 342
rect -59 60 2369 228
rect -54 -54 2364 60
<< scpmos >>
rect 60 0 90 288
rect 168 0 198 288
rect 276 0 306 288
rect 384 0 414 288
rect 492 0 522 288
rect 600 0 630 288
rect 708 0 738 288
rect 816 0 846 288
rect 924 0 954 288
rect 1032 0 1062 288
rect 1140 0 1170 288
rect 1248 0 1278 288
rect 1356 0 1386 288
rect 1464 0 1494 288
rect 1572 0 1602 288
rect 1680 0 1710 288
rect 1788 0 1818 288
rect 1896 0 1926 288
rect 2004 0 2034 288
rect 2112 0 2142 288
rect 2220 0 2250 288
<< pdiff >>
rect 0 161 60 288
rect 0 127 8 161
rect 42 127 60 161
rect 0 0 60 127
rect 90 161 168 288
rect 90 127 112 161
rect 146 127 168 161
rect 90 0 168 127
rect 198 161 276 288
rect 198 127 220 161
rect 254 127 276 161
rect 198 0 276 127
rect 306 161 384 288
rect 306 127 328 161
rect 362 127 384 161
rect 306 0 384 127
rect 414 161 492 288
rect 414 127 436 161
rect 470 127 492 161
rect 414 0 492 127
rect 522 161 600 288
rect 522 127 544 161
rect 578 127 600 161
rect 522 0 600 127
rect 630 161 708 288
rect 630 127 652 161
rect 686 127 708 161
rect 630 0 708 127
rect 738 161 816 288
rect 738 127 760 161
rect 794 127 816 161
rect 738 0 816 127
rect 846 161 924 288
rect 846 127 868 161
rect 902 127 924 161
rect 846 0 924 127
rect 954 161 1032 288
rect 954 127 976 161
rect 1010 127 1032 161
rect 954 0 1032 127
rect 1062 161 1140 288
rect 1062 127 1084 161
rect 1118 127 1140 161
rect 1062 0 1140 127
rect 1170 161 1248 288
rect 1170 127 1192 161
rect 1226 127 1248 161
rect 1170 0 1248 127
rect 1278 161 1356 288
rect 1278 127 1300 161
rect 1334 127 1356 161
rect 1278 0 1356 127
rect 1386 161 1464 288
rect 1386 127 1408 161
rect 1442 127 1464 161
rect 1386 0 1464 127
rect 1494 161 1572 288
rect 1494 127 1516 161
rect 1550 127 1572 161
rect 1494 0 1572 127
rect 1602 161 1680 288
rect 1602 127 1624 161
rect 1658 127 1680 161
rect 1602 0 1680 127
rect 1710 161 1788 288
rect 1710 127 1732 161
rect 1766 127 1788 161
rect 1710 0 1788 127
rect 1818 161 1896 288
rect 1818 127 1840 161
rect 1874 127 1896 161
rect 1818 0 1896 127
rect 1926 161 2004 288
rect 1926 127 1948 161
rect 1982 127 2004 161
rect 1926 0 2004 127
rect 2034 161 2112 288
rect 2034 127 2056 161
rect 2090 127 2112 161
rect 2034 0 2112 127
rect 2142 161 2220 288
rect 2142 127 2164 161
rect 2198 127 2220 161
rect 2142 0 2220 127
rect 2250 161 2310 288
rect 2250 127 2268 161
rect 2302 127 2310 161
rect 2250 0 2310 127
<< pdiffc >>
rect 8 127 42 161
rect 112 127 146 161
rect 220 127 254 161
rect 328 127 362 161
rect 436 127 470 161
rect 544 127 578 161
rect 652 127 686 161
rect 760 127 794 161
rect 868 127 902 161
rect 976 127 1010 161
rect 1084 127 1118 161
rect 1192 127 1226 161
rect 1300 127 1334 161
rect 1408 127 1442 161
rect 1516 127 1550 161
rect 1624 127 1658 161
rect 1732 127 1766 161
rect 1840 127 1874 161
rect 1948 127 1982 161
rect 2056 127 2090 161
rect 2164 127 2198 161
rect 2268 127 2302 161
<< poly >>
rect 60 288 90 314
rect 168 288 198 314
rect 276 288 306 314
rect 384 288 414 314
rect 492 288 522 314
rect 600 288 630 314
rect 708 288 738 314
rect 816 288 846 314
rect 924 288 954 314
rect 1032 288 1062 314
rect 1140 288 1170 314
rect 1248 288 1278 314
rect 1356 288 1386 314
rect 1464 288 1494 314
rect 1572 288 1602 314
rect 1680 288 1710 314
rect 1788 288 1818 314
rect 1896 288 1926 314
rect 2004 288 2034 314
rect 2112 288 2142 314
rect 2220 288 2250 314
rect 60 -26 90 0
rect 168 -26 198 0
rect 276 -26 306 0
rect 384 -26 414 0
rect 492 -26 522 0
rect 600 -26 630 0
rect 708 -26 738 0
rect 816 -26 846 0
rect 924 -26 954 0
rect 1032 -26 1062 0
rect 1140 -26 1170 0
rect 1248 -26 1278 0
rect 1356 -26 1386 0
rect 1464 -26 1494 0
rect 1572 -26 1602 0
rect 1680 -26 1710 0
rect 1788 -26 1818 0
rect 1896 -26 1926 0
rect 2004 -26 2034 0
rect 2112 -26 2142 0
rect 2220 -26 2250 0
rect 60 -56 2250 -26
<< locali >>
rect 8 161 42 177
rect 8 111 42 127
rect 112 161 146 177
rect 112 77 146 127
rect 220 161 254 177
rect 220 111 254 127
rect 328 161 362 177
rect 328 77 362 127
rect 436 161 470 177
rect 436 111 470 127
rect 544 161 578 177
rect 544 77 578 127
rect 652 161 686 177
rect 652 111 686 127
rect 760 161 794 177
rect 760 77 794 127
rect 868 161 902 177
rect 868 111 902 127
rect 976 161 1010 177
rect 976 77 1010 127
rect 1084 161 1118 177
rect 1084 111 1118 127
rect 1192 161 1226 177
rect 1192 77 1226 127
rect 1300 161 1334 177
rect 1300 111 1334 127
rect 1408 161 1442 177
rect 1408 77 1442 127
rect 1516 161 1550 177
rect 1516 111 1550 127
rect 1624 161 1658 177
rect 1624 77 1658 127
rect 1732 161 1766 177
rect 1732 111 1766 127
rect 1840 161 1874 177
rect 1840 77 1874 127
rect 1948 161 1982 177
rect 1948 111 1982 127
rect 2056 161 2090 177
rect 2056 77 2090 127
rect 2164 161 2198 177
rect 2164 111 2198 127
rect 2268 161 2302 177
rect 2268 77 2302 127
rect 112 43 2302 77
use contact_9  contact_9_0
timestamp 1643671299
transform 1 0 2260 0 1 103
box 0 0 2 2
use contact_9  contact_9_1
timestamp 1643671299
transform 1 0 2156 0 1 103
box 0 0 2 2
use contact_9  contact_9_2
timestamp 1643671299
transform 1 0 2048 0 1 103
box 0 0 2 2
use contact_9  contact_9_3
timestamp 1643671299
transform 1 0 1940 0 1 103
box 0 0 2 2
use contact_9  contact_9_4
timestamp 1643671299
transform 1 0 1832 0 1 103
box 0 0 2 2
use contact_9  contact_9_5
timestamp 1643671299
transform 1 0 1724 0 1 103
box 0 0 2 2
use contact_9  contact_9_6
timestamp 1643671299
transform 1 0 1616 0 1 103
box 0 0 2 2
use contact_9  contact_9_7
timestamp 1643671299
transform 1 0 1508 0 1 103
box 0 0 2 2
use contact_9  contact_9_8
timestamp 1643671299
transform 1 0 1400 0 1 103
box 0 0 2 2
use contact_9  contact_9_9
timestamp 1643671299
transform 1 0 1292 0 1 103
box 0 0 2 2
use contact_9  contact_9_10
timestamp 1643671299
transform 1 0 1184 0 1 103
box 0 0 2 2
use contact_9  contact_9_11
timestamp 1643671299
transform 1 0 1076 0 1 103
box 0 0 2 2
use contact_9  contact_9_12
timestamp 1643671299
transform 1 0 968 0 1 103
box 0 0 2 2
use contact_9  contact_9_13
timestamp 1643671299
transform 1 0 860 0 1 103
box 0 0 2 2
use contact_9  contact_9_14
timestamp 1643671299
transform 1 0 752 0 1 103
box 0 0 2 2
use contact_9  contact_9_15
timestamp 1643671299
transform 1 0 644 0 1 103
box 0 0 2 2
use contact_9  contact_9_16
timestamp 1643671299
transform 1 0 536 0 1 103
box 0 0 2 2
use contact_9  contact_9_17
timestamp 1643671299
transform 1 0 428 0 1 103
box 0 0 2 2
use contact_9  contact_9_18
timestamp 1643671299
transform 1 0 320 0 1 103
box 0 0 2 2
use contact_9  contact_9_19
timestamp 1643671299
transform 1 0 212 0 1 103
box 0 0 2 2
use contact_9  contact_9_20
timestamp 1643671299
transform 1 0 104 0 1 103
box 0 0 2 2
use contact_9  contact_9_21
timestamp 1643671299
transform 1 0 0 0 1 103
box 0 0 2 2
<< labels >>
rlabel mvvaractor s 1155 -41 1155 -41 4 G
rlabel locali s 885 144 885 144 4 S
rlabel locali s 1749 144 1749 144 4 S
rlabel locali s 453 144 453 144 4 S
rlabel locali s 669 144 669 144 4 S
rlabel locali s 2181 144 2181 144 4 S
rlabel locali s 1533 144 1533 144 4 S
rlabel locali s 1317 144 1317 144 4 S
rlabel locali s 1965 144 1965 144 4 S
rlabel locali s 25 144 25 144 4 S
rlabel locali s 1101 144 1101 144 4 S
rlabel locali s 237 144 237 144 4 S
rlabel locali s 1207 60 1207 60 4 D
<< properties >>
string FIXED_BBOX -54 -56 2364 60
string GDS_FILE sram_0rw2r1w_16_32_sky130A.gds
string GDS_END 1205446
string GDS_START 1200634
<< end >>
