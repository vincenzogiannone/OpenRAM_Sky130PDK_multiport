magic
tech sky130A
magscale 1 2
timestamp 1644951705
<< checkpaint >>
rect -1260 -1302 7372 50518
<< viali >>
rect 2938 30047 2972 30081
rect 2938 28423 2972 28457
rect 2938 26967 2972 27001
rect 2938 25343 2972 25377
rect 2938 23887 2972 23921
rect 2938 22263 2972 22297
rect 2938 20807 2972 20841
rect 2938 19183 2972 19217
rect 2938 14651 2972 14685
rect 2938 13027 2972 13061
rect 2938 11571 2972 11605
rect 2938 9947 2972 9981
rect 2938 5415 2972 5449
rect 2938 3791 2972 3825
rect 2938 2335 2972 2369
rect 2938 711 2972 745
<< metal1 >>
rect 6014 49190 6020 49242
rect 6072 49190 6078 49242
rect 4268 48808 4274 48860
rect 4326 48848 4332 48860
rect 4326 48820 5526 48848
rect 4326 48808 4332 48820
rect 3764 48722 3770 48774
rect 3822 48762 3828 48774
rect 3822 48734 5430 48762
rect 3822 48722 3828 48734
rect 3344 48636 3350 48688
rect 3402 48676 3408 48688
rect 3402 48648 5334 48676
rect 3402 48636 3408 48648
rect 5666 48608 6032 48636
rect 4268 48550 4274 48602
rect 4326 48590 4332 48602
rect 4326 48562 5130 48590
rect 4326 48550 4332 48562
rect 3764 48464 3770 48516
rect 3822 48504 3828 48516
rect 3822 48476 5034 48504
rect 5748 48486 6032 48514
rect 3822 48464 3828 48476
rect 3260 48378 3266 48430
rect 3318 48418 3324 48430
rect 3318 48390 4938 48418
rect 3318 48378 3324 48390
rect 4268 48292 4274 48344
rect 4326 48332 4332 48344
rect 5956 48340 6032 48368
rect 4326 48304 4842 48332
rect 4326 48292 4332 48304
rect 3764 48206 3770 48258
rect 3822 48246 3828 48258
rect 3822 48218 4746 48246
rect 3822 48206 3828 48218
rect 3176 48120 3182 48172
rect 3234 48160 3240 48172
rect 3234 48132 4650 48160
rect 3234 48120 3240 48132
rect 6014 47652 6020 47704
rect 6072 47652 6078 47704
rect 3260 47184 3266 47236
rect 3318 47224 3324 47236
rect 3318 47196 4650 47224
rect 3318 47184 3324 47196
rect 3680 47098 3686 47150
rect 3738 47138 3744 47150
rect 3738 47110 4746 47138
rect 3738 47098 3744 47110
rect 4268 47012 4274 47064
rect 4326 47052 4332 47064
rect 4326 47024 4842 47052
rect 4326 47012 4332 47024
rect 5956 46988 6032 47016
rect 3344 46926 3350 46978
rect 3402 46966 3408 46978
rect 3402 46938 4938 46966
rect 3402 46926 3408 46938
rect 3680 46840 3686 46892
rect 3738 46880 3744 46892
rect 3738 46852 5034 46880
rect 3738 46840 3744 46852
rect 5748 46842 6032 46870
rect 4268 46754 4274 46806
rect 4326 46794 4332 46806
rect 4326 46766 5130 46794
rect 4326 46754 4332 46766
rect 5666 46720 6032 46748
rect 3428 46668 3434 46720
rect 3486 46708 3492 46720
rect 3486 46680 5334 46708
rect 3486 46668 3492 46680
rect 3680 46582 3686 46634
rect 3738 46622 3744 46634
rect 3738 46594 5430 46622
rect 3738 46582 3744 46594
rect 4268 46496 4274 46548
rect 4326 46536 4332 46548
rect 4326 46508 5526 46536
rect 4326 46496 4332 46508
rect 6014 46114 6020 46166
rect 6072 46114 6078 46166
rect 4268 45732 4274 45784
rect 4326 45772 4332 45784
rect 4326 45744 5526 45772
rect 4326 45732 4332 45744
rect 3680 45646 3686 45698
rect 3738 45686 3744 45698
rect 3738 45658 5430 45686
rect 3738 45646 3744 45658
rect 3176 45560 3182 45612
rect 3234 45600 3240 45612
rect 3234 45572 5334 45600
rect 3234 45560 3240 45572
rect 5666 45532 6032 45560
rect 4268 45474 4274 45526
rect 4326 45514 4332 45526
rect 4326 45486 5130 45514
rect 4326 45474 4332 45486
rect 3596 45388 3602 45440
rect 3654 45428 3660 45440
rect 3654 45400 5034 45428
rect 5748 45410 6032 45438
rect 3654 45388 3660 45400
rect 3428 45302 3434 45354
rect 3486 45342 3492 45354
rect 3486 45314 4938 45342
rect 3486 45302 3492 45314
rect 4268 45216 4274 45268
rect 4326 45256 4332 45268
rect 5956 45264 6032 45292
rect 4326 45228 4842 45256
rect 4326 45216 4332 45228
rect 3596 45130 3602 45182
rect 3654 45170 3660 45182
rect 3654 45142 4746 45170
rect 3654 45130 3660 45142
rect 3344 45044 3350 45096
rect 3402 45084 3408 45096
rect 3402 45056 4650 45084
rect 3402 45044 3408 45056
rect 6014 44576 6020 44628
rect 6072 44576 6078 44628
rect 3428 44108 3434 44160
rect 3486 44148 3492 44160
rect 3486 44120 4650 44148
rect 3486 44108 3492 44120
rect 3512 44022 3518 44074
rect 3570 44062 3576 44074
rect 3570 44034 4746 44062
rect 3570 44022 3576 44034
rect 4268 43936 4274 43988
rect 4326 43976 4332 43988
rect 4326 43948 4842 43976
rect 4326 43936 4332 43948
rect 5956 43912 6032 43940
rect 3176 43850 3182 43902
rect 3234 43890 3240 43902
rect 3234 43862 4938 43890
rect 3234 43850 3240 43862
rect 3596 43764 3602 43816
rect 3654 43804 3660 43816
rect 3654 43776 5034 43804
rect 3654 43764 3660 43776
rect 5748 43766 6032 43794
rect 4268 43678 4274 43730
rect 4326 43718 4332 43730
rect 4326 43690 5130 43718
rect 4326 43678 4332 43690
rect 5666 43644 6032 43672
rect 3260 43592 3266 43644
rect 3318 43632 3324 43644
rect 3318 43604 5334 43632
rect 3318 43592 3324 43604
rect 3596 43506 3602 43558
rect 3654 43546 3660 43558
rect 3654 43518 5430 43546
rect 3654 43506 3660 43518
rect 4268 43420 4274 43472
rect 4326 43460 4332 43472
rect 4326 43432 5526 43460
rect 4326 43420 4332 43432
rect 6014 43038 6020 43090
rect 6072 43038 6078 43090
rect 4268 42656 4274 42708
rect 4326 42696 4332 42708
rect 4326 42668 5526 42696
rect 4326 42656 4332 42668
rect 3512 42570 3518 42622
rect 3570 42610 3576 42622
rect 3570 42582 5430 42610
rect 3570 42570 3576 42582
rect 3344 42484 3350 42536
rect 3402 42524 3408 42536
rect 3402 42496 5334 42524
rect 3402 42484 3408 42496
rect 5666 42456 6032 42484
rect 4268 42398 4274 42450
rect 4326 42438 4332 42450
rect 4326 42410 5130 42438
rect 4326 42398 4332 42410
rect 3512 42312 3518 42364
rect 3570 42352 3576 42364
rect 3570 42324 5034 42352
rect 5748 42334 6032 42362
rect 3570 42312 3576 42324
rect 3260 42226 3266 42278
rect 3318 42266 3324 42278
rect 3318 42238 4938 42266
rect 3318 42226 3324 42238
rect 4268 42140 4274 42192
rect 4326 42180 4332 42192
rect 5956 42188 6032 42216
rect 4326 42152 4842 42180
rect 4326 42140 4332 42152
rect 3512 42054 3518 42106
rect 3570 42094 3576 42106
rect 3570 42066 4746 42094
rect 3570 42054 3576 42066
rect 3176 41968 3182 42020
rect 3234 42008 3240 42020
rect 3234 41980 4650 42008
rect 3234 41968 3240 41980
rect 6014 41500 6020 41552
rect 6072 41500 6078 41552
rect 3260 41032 3266 41084
rect 3318 41072 3324 41084
rect 3318 41044 4650 41072
rect 3318 41032 3324 41044
rect 3764 40946 3770 40998
rect 3822 40986 3828 40998
rect 3822 40958 4746 40986
rect 3822 40946 3828 40958
rect 4184 40860 4190 40912
rect 4242 40900 4248 40912
rect 4242 40872 4842 40900
rect 4242 40860 4248 40872
rect 5956 40836 6032 40864
rect 3344 40774 3350 40826
rect 3402 40814 3408 40826
rect 3402 40786 4938 40814
rect 3402 40774 3408 40786
rect 3764 40688 3770 40740
rect 3822 40728 3828 40740
rect 3822 40700 5034 40728
rect 3822 40688 3828 40700
rect 5748 40690 6032 40718
rect 4184 40602 4190 40654
rect 4242 40642 4248 40654
rect 4242 40614 5130 40642
rect 4242 40602 4248 40614
rect 5666 40568 6032 40596
rect 3428 40516 3434 40568
rect 3486 40556 3492 40568
rect 3486 40528 5334 40556
rect 3486 40516 3492 40528
rect 3764 40430 3770 40482
rect 3822 40470 3828 40482
rect 3822 40442 5430 40470
rect 3822 40430 3828 40442
rect 4184 40344 4190 40396
rect 4242 40384 4248 40396
rect 4242 40356 5526 40384
rect 4242 40344 4248 40356
rect 6014 39962 6020 40014
rect 6072 39962 6078 40014
rect 4184 39580 4190 39632
rect 4242 39620 4248 39632
rect 4242 39592 5526 39620
rect 4242 39580 4248 39592
rect 3764 39494 3770 39546
rect 3822 39534 3828 39546
rect 3822 39506 5430 39534
rect 3822 39494 3828 39506
rect 3176 39408 3182 39460
rect 3234 39448 3240 39460
rect 3234 39420 5334 39448
rect 3234 39408 3240 39420
rect 5666 39380 6032 39408
rect 4184 39322 4190 39374
rect 4242 39362 4248 39374
rect 4242 39334 5130 39362
rect 4242 39322 4248 39334
rect 3680 39236 3686 39288
rect 3738 39276 3744 39288
rect 3738 39248 5034 39276
rect 5748 39258 6032 39286
rect 3738 39236 3744 39248
rect 3428 39150 3434 39202
rect 3486 39190 3492 39202
rect 3486 39162 4938 39190
rect 3486 39150 3492 39162
rect 4184 39064 4190 39116
rect 4242 39104 4248 39116
rect 5956 39112 6032 39140
rect 4242 39076 4842 39104
rect 4242 39064 4248 39076
rect 3680 38978 3686 39030
rect 3738 39018 3744 39030
rect 3738 38990 4746 39018
rect 3738 38978 3744 38990
rect 3344 38892 3350 38944
rect 3402 38932 3408 38944
rect 3402 38904 4650 38932
rect 3402 38892 3408 38904
rect 6014 38424 6020 38476
rect 6072 38424 6078 38476
rect 3428 37956 3434 38008
rect 3486 37996 3492 38008
rect 3486 37968 4650 37996
rect 3486 37956 3492 37968
rect 3596 37870 3602 37922
rect 3654 37910 3660 37922
rect 3654 37882 4746 37910
rect 3654 37870 3660 37882
rect 4184 37784 4190 37836
rect 4242 37824 4248 37836
rect 4242 37796 4842 37824
rect 4242 37784 4248 37796
rect 5956 37760 6032 37788
rect 3176 37698 3182 37750
rect 3234 37738 3240 37750
rect 3234 37710 4938 37738
rect 3234 37698 3240 37710
rect 3680 37612 3686 37664
rect 3738 37652 3744 37664
rect 3738 37624 5034 37652
rect 3738 37612 3744 37624
rect 5748 37614 6032 37642
rect 4184 37526 4190 37578
rect 4242 37566 4248 37578
rect 4242 37538 5130 37566
rect 4242 37526 4248 37538
rect 5666 37492 6032 37520
rect 3260 37440 3266 37492
rect 3318 37480 3324 37492
rect 3318 37452 5334 37480
rect 3318 37440 3324 37452
rect 3680 37354 3686 37406
rect 3738 37394 3744 37406
rect 3738 37366 5430 37394
rect 3738 37354 3744 37366
rect 4184 37268 4190 37320
rect 4242 37308 4248 37320
rect 4242 37280 5526 37308
rect 4242 37268 4248 37280
rect 6014 36886 6020 36938
rect 6072 36886 6078 36938
rect 4184 36504 4190 36556
rect 4242 36544 4248 36556
rect 4242 36516 5526 36544
rect 4242 36504 4248 36516
rect 3596 36418 3602 36470
rect 3654 36458 3660 36470
rect 3654 36430 5430 36458
rect 3654 36418 3660 36430
rect 3344 36332 3350 36384
rect 3402 36372 3408 36384
rect 3402 36344 5334 36372
rect 3402 36332 3408 36344
rect 5666 36304 6032 36332
rect 4184 36246 4190 36298
rect 4242 36286 4248 36298
rect 4242 36258 5130 36286
rect 4242 36246 4248 36258
rect 3596 36160 3602 36212
rect 3654 36200 3660 36212
rect 3654 36172 5034 36200
rect 5748 36182 6032 36210
rect 3654 36160 3660 36172
rect 3260 36074 3266 36126
rect 3318 36114 3324 36126
rect 3318 36086 4938 36114
rect 3318 36074 3324 36086
rect 4184 35988 4190 36040
rect 4242 36028 4248 36040
rect 5956 36036 6032 36064
rect 4242 36000 4842 36028
rect 4242 35988 4248 36000
rect 3596 35902 3602 35954
rect 3654 35942 3660 35954
rect 3654 35914 4746 35942
rect 3654 35902 3660 35914
rect 3176 35816 3182 35868
rect 3234 35856 3240 35868
rect 3234 35828 4650 35856
rect 3234 35816 3240 35828
rect 6014 35348 6020 35400
rect 6072 35348 6078 35400
rect 3260 34880 3266 34932
rect 3318 34920 3324 34932
rect 3318 34892 4650 34920
rect 3318 34880 3324 34892
rect 3512 34794 3518 34846
rect 3570 34834 3576 34846
rect 3570 34806 4746 34834
rect 3570 34794 3576 34806
rect 4184 34708 4190 34760
rect 4242 34748 4248 34760
rect 4242 34720 4842 34748
rect 4242 34708 4248 34720
rect 5956 34684 6032 34712
rect 3344 34622 3350 34674
rect 3402 34662 3408 34674
rect 3402 34634 4938 34662
rect 3402 34622 3408 34634
rect 3512 34536 3518 34588
rect 3570 34576 3576 34588
rect 3570 34548 5034 34576
rect 3570 34536 3576 34548
rect 5748 34538 6032 34566
rect 4184 34450 4190 34502
rect 4242 34490 4248 34502
rect 4242 34462 5130 34490
rect 4242 34450 4248 34462
rect 5666 34416 6032 34444
rect 3428 34364 3434 34416
rect 3486 34404 3492 34416
rect 3486 34376 5334 34404
rect 3486 34364 3492 34376
rect 3512 34278 3518 34330
rect 3570 34318 3576 34330
rect 3570 34290 5430 34318
rect 3570 34278 3576 34290
rect 4184 34192 4190 34244
rect 4242 34232 4248 34244
rect 4242 34204 5526 34232
rect 4242 34192 4248 34204
rect 6014 33810 6020 33862
rect 6072 33810 6078 33862
rect 4184 33428 4190 33480
rect 4242 33468 4248 33480
rect 4242 33440 5526 33468
rect 4242 33428 4248 33440
rect 3512 33342 3518 33394
rect 3570 33382 3576 33394
rect 3570 33354 5430 33382
rect 3570 33342 3576 33354
rect 3176 33256 3182 33308
rect 3234 33296 3240 33308
rect 3234 33268 5334 33296
rect 3234 33256 3240 33268
rect 5666 33228 6032 33256
rect 4100 33170 4106 33222
rect 4158 33210 4164 33222
rect 4158 33182 5130 33210
rect 4158 33170 4164 33182
rect 3764 33084 3770 33136
rect 3822 33124 3828 33136
rect 3822 33096 5034 33124
rect 5748 33106 6032 33134
rect 3822 33084 3828 33096
rect 3428 32998 3434 33050
rect 3486 33038 3492 33050
rect 3486 33010 4938 33038
rect 3486 32998 3492 33010
rect 4100 32912 4106 32964
rect 4158 32952 4164 32964
rect 5956 32960 6032 32988
rect 4158 32924 4842 32952
rect 4158 32912 4164 32924
rect 3764 32826 3770 32878
rect 3822 32866 3828 32878
rect 3822 32838 4746 32866
rect 3822 32826 3828 32838
rect 3344 32740 3350 32792
rect 3402 32780 3408 32792
rect 3402 32752 4650 32780
rect 3402 32740 3408 32752
rect 6014 32272 6020 32324
rect 6072 32272 6078 32324
rect 3428 31804 3434 31856
rect 3486 31844 3492 31856
rect 3486 31816 4650 31844
rect 3486 31804 3492 31816
rect 3680 31718 3686 31770
rect 3738 31758 3744 31770
rect 3738 31730 4746 31758
rect 3738 31718 3744 31730
rect 4100 31632 4106 31684
rect 4158 31672 4164 31684
rect 4158 31644 4842 31672
rect 4158 31632 4164 31644
rect 5956 31608 6032 31636
rect 3176 31546 3182 31598
rect 3234 31586 3240 31598
rect 3234 31558 4938 31586
rect 3234 31546 3240 31558
rect 3764 31460 3770 31512
rect 3822 31500 3828 31512
rect 3822 31472 5034 31500
rect 3822 31460 3828 31472
rect 5748 31462 6032 31490
rect 4100 31374 4106 31426
rect 4158 31414 4164 31426
rect 4158 31386 5130 31414
rect 4158 31374 4164 31386
rect 5666 31340 6032 31368
rect 3260 31288 3266 31340
rect 3318 31328 3324 31340
rect 3318 31300 5334 31328
rect 3318 31288 3324 31300
rect 3764 31202 3770 31254
rect 3822 31242 3828 31254
rect 3822 31214 5430 31242
rect 3822 31202 3828 31214
rect 4100 31116 4106 31168
rect 4158 31156 4164 31168
rect 4158 31128 5526 31156
rect 4158 31116 4164 31128
rect 6014 30734 6020 30786
rect 6072 30734 6078 30786
rect 4100 30352 4106 30404
rect 4158 30392 4164 30404
rect 4158 30364 5526 30392
rect 4158 30352 4164 30364
rect 3680 30266 3686 30318
rect 3738 30306 3744 30318
rect 3738 30278 5430 30306
rect 3738 30266 3744 30278
rect 3344 30180 3350 30232
rect 3402 30220 3408 30232
rect 3402 30192 5334 30220
rect 3402 30180 3408 30192
rect 5666 30152 6032 30180
rect 4100 30094 4106 30146
rect 4158 30134 4164 30146
rect 4158 30106 5130 30134
rect 4158 30094 4164 30106
rect 2923 30038 2929 30090
rect 2981 30038 2987 30090
rect 3680 30008 3686 30060
rect 3738 30048 3744 30060
rect 3738 30020 5034 30048
rect 5748 30030 6032 30058
rect 3738 30008 3744 30020
rect 3260 29922 3266 29974
rect 3318 29962 3324 29974
rect 3318 29934 4938 29962
rect 3318 29922 3324 29934
rect 4100 29836 4106 29888
rect 4158 29876 4164 29888
rect 5956 29884 6032 29912
rect 4158 29848 4842 29876
rect 4158 29836 4164 29848
rect 3680 29750 3686 29802
rect 3738 29790 3744 29802
rect 3738 29762 4746 29790
rect 3738 29750 3744 29762
rect 3176 29664 3182 29716
rect 3234 29704 3240 29716
rect 3234 29676 4650 29704
rect 3234 29664 3240 29676
rect 6014 29196 6020 29248
rect 6072 29196 6078 29248
rect 3260 28728 3266 28780
rect 3318 28768 3324 28780
rect 3318 28740 4650 28768
rect 3318 28728 3324 28740
rect 3596 28642 3602 28694
rect 3654 28682 3660 28694
rect 3654 28654 4746 28682
rect 3654 28642 3660 28654
rect 4100 28556 4106 28608
rect 4158 28596 4164 28608
rect 4158 28568 4842 28596
rect 4158 28556 4164 28568
rect 5956 28532 6032 28560
rect 3344 28470 3350 28522
rect 3402 28510 3408 28522
rect 3402 28482 4938 28510
rect 3402 28470 3408 28482
rect 2923 28414 2929 28466
rect 2981 28414 2987 28466
rect 3596 28384 3602 28436
rect 3654 28424 3660 28436
rect 3654 28396 5034 28424
rect 3654 28384 3660 28396
rect 5748 28386 6032 28414
rect 4100 28298 4106 28350
rect 4158 28338 4164 28350
rect 4158 28310 5130 28338
rect 4158 28298 4164 28310
rect 5666 28264 6032 28292
rect 3428 28212 3434 28264
rect 3486 28252 3492 28264
rect 3486 28224 5334 28252
rect 3486 28212 3492 28224
rect 3596 28126 3602 28178
rect 3654 28166 3660 28178
rect 3654 28138 5430 28166
rect 3654 28126 3660 28138
rect 4100 28040 4106 28092
rect 4158 28080 4164 28092
rect 4158 28052 5526 28080
rect 4158 28040 4164 28052
rect 6014 27658 6020 27710
rect 6072 27658 6078 27710
rect 4100 27276 4106 27328
rect 4158 27316 4164 27328
rect 4158 27288 5526 27316
rect 4158 27276 4164 27288
rect 3596 27190 3602 27242
rect 3654 27230 3660 27242
rect 3654 27202 5430 27230
rect 3654 27190 3660 27202
rect 3176 27104 3182 27156
rect 3234 27144 3240 27156
rect 3234 27116 5334 27144
rect 3234 27104 3240 27116
rect 5666 27076 6032 27104
rect 4100 27018 4106 27070
rect 4158 27058 4164 27070
rect 4158 27030 5130 27058
rect 4158 27018 4164 27030
rect 2923 26958 2929 27010
rect 2981 26958 2987 27010
rect 3512 26932 3518 26984
rect 3570 26972 3576 26984
rect 3570 26944 5034 26972
rect 5748 26954 6032 26982
rect 3570 26932 3576 26944
rect 3428 26846 3434 26898
rect 3486 26886 3492 26898
rect 3486 26858 4938 26886
rect 3486 26846 3492 26858
rect 4100 26760 4106 26812
rect 4158 26800 4164 26812
rect 5956 26808 6032 26836
rect 4158 26772 4842 26800
rect 4158 26760 4164 26772
rect 3512 26674 3518 26726
rect 3570 26714 3576 26726
rect 3570 26686 4746 26714
rect 3570 26674 3576 26686
rect 3344 26588 3350 26640
rect 3402 26628 3408 26640
rect 3402 26600 4650 26628
rect 3402 26588 3408 26600
rect 6014 26120 6020 26172
rect 6072 26120 6078 26172
rect 3428 25652 3434 25704
rect 3486 25692 3492 25704
rect 3486 25664 4650 25692
rect 3486 25652 3492 25664
rect 3764 25566 3770 25618
rect 3822 25606 3828 25618
rect 3822 25578 4746 25606
rect 3822 25566 3828 25578
rect 4016 25480 4022 25532
rect 4074 25520 4080 25532
rect 4074 25492 4842 25520
rect 4074 25480 4080 25492
rect 5956 25456 6032 25484
rect 3176 25394 3182 25446
rect 3234 25434 3240 25446
rect 3234 25406 4938 25434
rect 3234 25394 3240 25406
rect 2923 25334 2929 25386
rect 2981 25334 2987 25386
rect 3512 25308 3518 25360
rect 3570 25348 3576 25360
rect 3570 25320 5034 25348
rect 3570 25308 3576 25320
rect 5748 25310 6032 25338
rect 4100 25222 4106 25274
rect 4158 25262 4164 25274
rect 4158 25234 5130 25262
rect 4158 25222 4164 25234
rect 5666 25188 6032 25216
rect 3260 25136 3266 25188
rect 3318 25176 3324 25188
rect 3318 25148 5334 25176
rect 3318 25136 3324 25148
rect 3512 25050 3518 25102
rect 3570 25090 3576 25102
rect 3570 25062 5430 25090
rect 3570 25050 3576 25062
rect 4100 24964 4106 25016
rect 4158 25004 4164 25016
rect 4158 24976 5526 25004
rect 4158 24964 4164 24976
rect 6014 24582 6020 24634
rect 6072 24582 6078 24634
rect 4016 24200 4022 24252
rect 4074 24240 4080 24252
rect 4074 24212 5526 24240
rect 4074 24200 4080 24212
rect 3764 24114 3770 24166
rect 3822 24154 3828 24166
rect 3822 24126 5430 24154
rect 3822 24114 3828 24126
rect 3344 24028 3350 24080
rect 3402 24068 3408 24080
rect 3402 24040 5334 24068
rect 3402 24028 3408 24040
rect 5666 24000 6032 24028
rect 4016 23942 4022 23994
rect 4074 23982 4080 23994
rect 4074 23954 5130 23982
rect 4074 23942 4080 23954
rect 2923 23878 2929 23930
rect 2981 23878 2987 23930
rect 3764 23856 3770 23908
rect 3822 23896 3828 23908
rect 3822 23868 5034 23896
rect 5748 23878 6032 23906
rect 3822 23856 3828 23868
rect 3260 23770 3266 23822
rect 3318 23810 3324 23822
rect 3318 23782 4938 23810
rect 3318 23770 3324 23782
rect 4016 23684 4022 23736
rect 4074 23724 4080 23736
rect 5956 23732 6032 23760
rect 4074 23696 4842 23724
rect 4074 23684 4080 23696
rect 3764 23598 3770 23650
rect 3822 23638 3828 23650
rect 3822 23610 4746 23638
rect 3822 23598 3828 23610
rect 3176 23512 3182 23564
rect 3234 23552 3240 23564
rect 3234 23524 4650 23552
rect 3234 23512 3240 23524
rect 6014 23044 6020 23096
rect 6072 23044 6078 23096
rect 3260 22576 3266 22628
rect 3318 22616 3324 22628
rect 3318 22588 4650 22616
rect 3318 22576 3324 22588
rect 3680 22490 3686 22542
rect 3738 22530 3744 22542
rect 3738 22502 4746 22530
rect 3738 22490 3744 22502
rect 4016 22404 4022 22456
rect 4074 22444 4080 22456
rect 4074 22416 4842 22444
rect 4074 22404 4080 22416
rect 5956 22380 6032 22408
rect 3344 22318 3350 22370
rect 3402 22358 3408 22370
rect 3402 22330 4938 22358
rect 3402 22318 3408 22330
rect 504 22254 510 22306
rect 562 22294 568 22306
rect 868 22294 874 22306
rect 562 22266 874 22294
rect 562 22254 568 22266
rect 868 22254 874 22266
rect 926 22254 932 22306
rect 2923 22254 2929 22306
rect 2981 22254 2987 22306
rect 3680 22232 3686 22284
rect 3738 22272 3744 22284
rect 3738 22244 5034 22272
rect 3738 22232 3744 22244
rect 5748 22234 6032 22262
rect 4016 22146 4022 22198
rect 4074 22186 4080 22198
rect 4074 22158 5130 22186
rect 4074 22146 4080 22158
rect 5666 22112 6032 22140
rect 3428 22060 3434 22112
rect 3486 22100 3492 22112
rect 3486 22072 5334 22100
rect 3486 22060 3492 22072
rect 3680 21974 3686 22026
rect 3738 22014 3744 22026
rect 3738 21986 5430 22014
rect 3738 21974 3744 21986
rect 4016 21888 4022 21940
rect 4074 21928 4080 21940
rect 4074 21900 5526 21928
rect 4074 21888 4080 21900
rect 6014 21506 6020 21558
rect 6072 21506 6078 21558
rect 4016 21124 4022 21176
rect 4074 21164 4080 21176
rect 4074 21136 5526 21164
rect 4074 21124 4080 21136
rect 3680 21038 3686 21090
rect 3738 21078 3744 21090
rect 3738 21050 5430 21078
rect 3738 21038 3744 21050
rect 3176 20952 3182 21004
rect 3234 20992 3240 21004
rect 3234 20964 5334 20992
rect 3234 20952 3240 20964
rect 5666 20924 6032 20952
rect 4016 20866 4022 20918
rect 4074 20906 4080 20918
rect 4074 20878 5130 20906
rect 4074 20866 4080 20878
rect 420 20798 426 20850
rect 478 20838 484 20850
rect 784 20838 790 20850
rect 478 20810 790 20838
rect 478 20798 484 20810
rect 784 20798 790 20810
rect 842 20798 848 20850
rect 2923 20798 2929 20850
rect 2981 20798 2987 20850
rect 3596 20780 3602 20832
rect 3654 20820 3660 20832
rect 3654 20792 5034 20820
rect 5748 20802 6032 20830
rect 3654 20780 3660 20792
rect 3428 20694 3434 20746
rect 3486 20734 3492 20746
rect 3486 20706 4938 20734
rect 3486 20694 3492 20706
rect 4016 20608 4022 20660
rect 4074 20648 4080 20660
rect 5956 20656 6032 20684
rect 4074 20620 4842 20648
rect 4074 20608 4080 20620
rect 3596 20522 3602 20574
rect 3654 20562 3660 20574
rect 3654 20534 4746 20562
rect 3654 20522 3660 20534
rect 3344 20436 3350 20488
rect 3402 20476 3408 20488
rect 3402 20448 4650 20476
rect 3402 20436 3408 20448
rect 6014 19968 6020 20020
rect 6072 19968 6078 20020
rect 3428 19500 3434 19552
rect 3486 19540 3492 19552
rect 3486 19512 4650 19540
rect 3486 19500 3492 19512
rect 3512 19414 3518 19466
rect 3570 19454 3576 19466
rect 3570 19426 4746 19454
rect 3570 19414 3576 19426
rect 4016 19328 4022 19380
rect 4074 19368 4080 19380
rect 4074 19340 4842 19368
rect 4074 19328 4080 19340
rect 5956 19304 6032 19332
rect 3176 19242 3182 19294
rect 3234 19282 3240 19294
rect 3234 19254 4938 19282
rect 3234 19242 3240 19254
rect 336 19174 342 19226
rect 394 19214 400 19226
rect 700 19214 706 19226
rect 394 19186 706 19214
rect 394 19174 400 19186
rect 700 19174 706 19186
rect 758 19174 764 19226
rect 2923 19174 2929 19226
rect 2981 19174 2987 19226
rect 3596 19156 3602 19208
rect 3654 19196 3660 19208
rect 3654 19168 5034 19196
rect 3654 19156 3660 19168
rect 5748 19158 6032 19186
rect 4016 19070 4022 19122
rect 4074 19110 4080 19122
rect 4074 19082 5130 19110
rect 4074 19070 4080 19082
rect 5666 19036 6032 19064
rect 3260 18984 3266 19036
rect 3318 19024 3324 19036
rect 3318 18996 5334 19024
rect 3318 18984 3324 18996
rect 3596 18898 3602 18950
rect 3654 18938 3660 18950
rect 3654 18910 5430 18938
rect 3654 18898 3660 18910
rect 4016 18812 4022 18864
rect 4074 18852 4080 18864
rect 4074 18824 5526 18852
rect 4074 18812 4080 18824
rect 6014 18430 6020 18482
rect 6072 18430 6078 18482
rect 4016 18048 4022 18100
rect 4074 18088 4080 18100
rect 4074 18060 5526 18088
rect 4074 18048 4080 18060
rect 3512 17962 3518 18014
rect 3570 18002 3576 18014
rect 3570 17974 5430 18002
rect 3570 17962 3576 17974
rect 3344 17876 3350 17928
rect 3402 17916 3408 17928
rect 3402 17888 5334 17916
rect 3402 17876 3408 17888
rect 5666 17848 6032 17876
rect 4016 17790 4022 17842
rect 4074 17830 4080 17842
rect 4074 17802 5130 17830
rect 4074 17790 4080 17802
rect 3512 17704 3518 17756
rect 3570 17744 3576 17756
rect 3570 17716 5034 17744
rect 5748 17726 6032 17754
rect 3570 17704 3576 17716
rect 3260 17618 3266 17670
rect 3318 17658 3324 17670
rect 3318 17630 4938 17658
rect 3318 17618 3324 17630
rect 4016 17532 4022 17584
rect 4074 17572 4080 17584
rect 5956 17580 6032 17608
rect 4074 17544 4842 17572
rect 4074 17532 4080 17544
rect 3512 17446 3518 17498
rect 3570 17486 3576 17498
rect 3570 17458 4746 17486
rect 3570 17446 3576 17458
rect 3176 17360 3182 17412
rect 3234 17400 3240 17412
rect 3234 17372 4650 17400
rect 3234 17360 3240 17372
rect 6014 16892 6020 16944
rect 6072 16892 6078 16944
rect 3260 16424 3266 16476
rect 3318 16464 3324 16476
rect 3318 16436 4650 16464
rect 3318 16424 3324 16436
rect 3764 16338 3770 16390
rect 3822 16378 3828 16390
rect 3822 16350 4746 16378
rect 3822 16338 3828 16350
rect 3932 16252 3938 16304
rect 3990 16292 3996 16304
rect 3990 16264 4842 16292
rect 3990 16252 3996 16264
rect 5956 16228 6032 16256
rect 3344 16166 3350 16218
rect 3402 16206 3408 16218
rect 3402 16178 4938 16206
rect 3402 16166 3408 16178
rect 3764 16080 3770 16132
rect 3822 16120 3828 16132
rect 3822 16092 5034 16120
rect 3822 16080 3828 16092
rect 5748 16082 6032 16110
rect 3932 15994 3938 16046
rect 3990 16034 3996 16046
rect 3990 16006 5130 16034
rect 3990 15994 3996 16006
rect 5666 15960 6032 15988
rect 3428 15908 3434 15960
rect 3486 15948 3492 15960
rect 3486 15920 5334 15948
rect 3486 15908 3492 15920
rect 3764 15822 3770 15874
rect 3822 15862 3828 15874
rect 3822 15834 5430 15862
rect 3822 15822 3828 15834
rect 3932 15736 3938 15788
rect 3990 15776 3996 15788
rect 3990 15748 5526 15776
rect 3990 15736 3996 15748
rect 6014 15354 6020 15406
rect 6072 15354 6078 15406
rect 3932 14972 3938 15024
rect 3990 15012 3996 15024
rect 3990 14984 5526 15012
rect 3990 14972 3996 14984
rect 3764 14886 3770 14938
rect 3822 14926 3828 14938
rect 3822 14898 5430 14926
rect 3822 14886 3828 14898
rect 3176 14800 3182 14852
rect 3234 14840 3240 14852
rect 3234 14812 5334 14840
rect 3234 14800 3240 14812
rect 5666 14772 6032 14800
rect 3932 14714 3938 14766
rect 3990 14754 3996 14766
rect 3990 14726 5130 14754
rect 3990 14714 3996 14726
rect 2923 14642 2929 14694
rect 2981 14642 2987 14694
rect 3680 14628 3686 14680
rect 3738 14668 3744 14680
rect 3738 14640 5034 14668
rect 5748 14650 6032 14678
rect 3738 14628 3744 14640
rect 3428 14542 3434 14594
rect 3486 14582 3492 14594
rect 3486 14554 4938 14582
rect 3486 14542 3492 14554
rect 3932 14456 3938 14508
rect 3990 14496 3996 14508
rect 5956 14504 6032 14532
rect 3990 14468 4842 14496
rect 3990 14456 3996 14468
rect 3680 14370 3686 14422
rect 3738 14410 3744 14422
rect 3738 14382 4746 14410
rect 3738 14370 3744 14382
rect 3344 14284 3350 14336
rect 3402 14324 3408 14336
rect 3402 14296 4650 14324
rect 3402 14284 3408 14296
rect 6014 13816 6020 13868
rect 6072 13816 6078 13868
rect 3428 13348 3434 13400
rect 3486 13388 3492 13400
rect 3486 13360 4650 13388
rect 3486 13348 3492 13360
rect 3596 13262 3602 13314
rect 3654 13302 3660 13314
rect 3654 13274 4746 13302
rect 3654 13262 3660 13274
rect 3932 13176 3938 13228
rect 3990 13216 3996 13228
rect 3990 13188 4842 13216
rect 3990 13176 3996 13188
rect 5956 13152 6032 13180
rect 3176 13090 3182 13142
rect 3234 13130 3240 13142
rect 3234 13102 4938 13130
rect 3234 13090 3240 13102
rect 2923 13018 2929 13070
rect 2981 13018 2987 13070
rect 3680 13004 3686 13056
rect 3738 13044 3744 13056
rect 3738 13016 5034 13044
rect 3738 13004 3744 13016
rect 5748 13006 6032 13034
rect 3932 12918 3938 12970
rect 3990 12958 3996 12970
rect 3990 12930 5130 12958
rect 3990 12918 3996 12930
rect 5666 12884 6032 12912
rect 3260 12832 3266 12884
rect 3318 12872 3324 12884
rect 3318 12844 5334 12872
rect 3318 12832 3324 12844
rect 3680 12746 3686 12798
rect 3738 12786 3744 12798
rect 3738 12758 5430 12786
rect 3738 12746 3744 12758
rect 3932 12660 3938 12712
rect 3990 12700 3996 12712
rect 3990 12672 5526 12700
rect 3990 12660 3996 12672
rect 6014 12278 6020 12330
rect 6072 12278 6078 12330
rect 3932 11896 3938 11948
rect 3990 11936 3996 11948
rect 3990 11908 5526 11936
rect 3990 11896 3996 11908
rect 3596 11810 3602 11862
rect 3654 11850 3660 11862
rect 3654 11822 5430 11850
rect 3654 11810 3660 11822
rect 3344 11724 3350 11776
rect 3402 11764 3408 11776
rect 3402 11736 5334 11764
rect 3402 11724 3408 11736
rect 5666 11696 6032 11724
rect 3932 11638 3938 11690
rect 3990 11678 3996 11690
rect 3990 11650 5130 11678
rect 3990 11638 3996 11650
rect 252 11562 258 11614
rect 310 11602 316 11614
rect 1216 11602 1222 11614
rect 310 11574 1222 11602
rect 310 11562 316 11574
rect 1216 11562 1222 11574
rect 1274 11562 1280 11614
rect 2923 11562 2929 11614
rect 2981 11562 2987 11614
rect 3596 11552 3602 11604
rect 3654 11592 3660 11604
rect 3654 11564 5034 11592
rect 5748 11574 6032 11602
rect 3654 11552 3660 11564
rect 3260 11466 3266 11518
rect 3318 11506 3324 11518
rect 3318 11478 4938 11506
rect 3318 11466 3324 11478
rect 3932 11380 3938 11432
rect 3990 11420 3996 11432
rect 5956 11428 6032 11456
rect 3990 11392 4842 11420
rect 3990 11380 3996 11392
rect 3596 11294 3602 11346
rect 3654 11334 3660 11346
rect 3654 11306 4746 11334
rect 3654 11294 3660 11306
rect 3176 11208 3182 11260
rect 3234 11248 3240 11260
rect 3234 11220 4650 11248
rect 3234 11208 3240 11220
rect 6014 10740 6020 10792
rect 6072 10740 6078 10792
rect 3260 10272 3266 10324
rect 3318 10312 3324 10324
rect 3318 10284 4650 10312
rect 3318 10272 3324 10284
rect 3512 10186 3518 10238
rect 3570 10226 3576 10238
rect 3570 10198 4746 10226
rect 3570 10186 3576 10198
rect 3932 10100 3938 10152
rect 3990 10140 3996 10152
rect 3990 10112 4842 10140
rect 3990 10100 3996 10112
rect 5956 10076 6032 10104
rect 3344 10014 3350 10066
rect 3402 10054 3408 10066
rect 3402 10026 4938 10054
rect 3402 10014 3408 10026
rect 168 9938 174 9990
rect 226 9978 232 9990
rect 1132 9978 1138 9990
rect 226 9950 1138 9978
rect 226 9938 232 9950
rect 1132 9938 1138 9950
rect 1190 9938 1196 9990
rect 2923 9938 2929 9990
rect 2981 9938 2987 9990
rect 3512 9928 3518 9980
rect 3570 9968 3576 9980
rect 3570 9940 5034 9968
rect 3570 9928 3576 9940
rect 5748 9930 6032 9958
rect 3932 9842 3938 9894
rect 3990 9882 3996 9894
rect 3990 9854 5130 9882
rect 3990 9842 3996 9854
rect 5666 9808 6032 9836
rect 3428 9756 3434 9808
rect 3486 9796 3492 9808
rect 3486 9768 5334 9796
rect 3486 9756 3492 9768
rect 3512 9670 3518 9722
rect 3570 9710 3576 9722
rect 3570 9682 5430 9710
rect 3570 9670 3576 9682
rect 3932 9584 3938 9636
rect 3990 9624 3996 9636
rect 3990 9596 5526 9624
rect 3990 9584 3996 9596
rect 6014 9202 6020 9254
rect 6072 9202 6078 9254
rect 3932 8820 3938 8872
rect 3990 8860 3996 8872
rect 3990 8832 5526 8860
rect 3990 8820 3996 8832
rect 3512 8734 3518 8786
rect 3570 8774 3576 8786
rect 3570 8746 5430 8774
rect 3570 8734 3576 8746
rect 3176 8648 3182 8700
rect 3234 8688 3240 8700
rect 3234 8660 5334 8688
rect 3234 8648 3240 8660
rect 5666 8620 6032 8648
rect 3848 8562 3854 8614
rect 3906 8602 3912 8614
rect 3906 8574 5130 8602
rect 3906 8562 3912 8574
rect 3764 8476 3770 8528
rect 3822 8516 3828 8528
rect 3822 8488 5034 8516
rect 5748 8498 6032 8526
rect 3822 8476 3828 8488
rect 3428 8390 3434 8442
rect 3486 8430 3492 8442
rect 3486 8402 4938 8430
rect 3486 8390 3492 8402
rect 3848 8304 3854 8356
rect 3906 8344 3912 8356
rect 5956 8352 6032 8380
rect 3906 8316 4842 8344
rect 3906 8304 3912 8316
rect 3764 8218 3770 8270
rect 3822 8258 3828 8270
rect 3822 8230 4746 8258
rect 3822 8218 3828 8230
rect 3344 8132 3350 8184
rect 3402 8172 3408 8184
rect 3402 8144 4650 8172
rect 3402 8132 3408 8144
rect 6014 7664 6020 7716
rect 6072 7664 6078 7716
rect 3428 7196 3434 7248
rect 3486 7236 3492 7248
rect 3486 7208 4650 7236
rect 3486 7196 3492 7208
rect 3680 7110 3686 7162
rect 3738 7150 3744 7162
rect 3738 7122 4746 7150
rect 3738 7110 3744 7122
rect 3848 7024 3854 7076
rect 3906 7064 3912 7076
rect 3906 7036 4842 7064
rect 3906 7024 3912 7036
rect 5956 7000 6032 7028
rect 3176 6938 3182 6990
rect 3234 6978 3240 6990
rect 3234 6950 4938 6978
rect 3234 6938 3240 6950
rect 3764 6852 3770 6904
rect 3822 6892 3828 6904
rect 3822 6864 5034 6892
rect 3822 6852 3828 6864
rect 5748 6854 6032 6882
rect 3848 6766 3854 6818
rect 3906 6806 3912 6818
rect 3906 6778 5130 6806
rect 3906 6766 3912 6778
rect 5666 6732 6032 6760
rect 3260 6680 3266 6732
rect 3318 6720 3324 6732
rect 3318 6692 5334 6720
rect 3318 6680 3324 6692
rect 3764 6594 3770 6646
rect 3822 6634 3828 6646
rect 3822 6606 5430 6634
rect 3822 6594 3828 6606
rect 3848 6508 3854 6560
rect 3906 6548 3912 6560
rect 3906 6520 5526 6548
rect 3906 6508 3912 6520
rect 6014 6126 6020 6178
rect 6072 6126 6078 6178
rect 3848 5744 3854 5796
rect 3906 5784 3912 5796
rect 3906 5756 5526 5784
rect 3906 5744 3912 5756
rect 3680 5658 3686 5710
rect 3738 5698 3744 5710
rect 3738 5670 5430 5698
rect 3738 5658 3744 5670
rect 3344 5572 3350 5624
rect 3402 5612 3408 5624
rect 3402 5584 5334 5612
rect 3402 5572 3408 5584
rect 5666 5544 6032 5572
rect 3848 5486 3854 5538
rect 3906 5526 3912 5538
rect 3906 5498 5130 5526
rect 3906 5486 3912 5498
rect 2923 5406 2929 5458
rect 2981 5406 2987 5458
rect 3680 5400 3686 5452
rect 3738 5440 3744 5452
rect 3738 5412 5034 5440
rect 5748 5422 6032 5450
rect 3738 5400 3744 5412
rect 3260 5314 3266 5366
rect 3318 5354 3324 5366
rect 3318 5326 4938 5354
rect 3318 5314 3324 5326
rect 3848 5228 3854 5280
rect 3906 5268 3912 5280
rect 5956 5276 6032 5304
rect 3906 5240 4842 5268
rect 3906 5228 3912 5240
rect 3680 5142 3686 5194
rect 3738 5182 3744 5194
rect 3738 5154 4746 5182
rect 3738 5142 3744 5154
rect 3176 5056 3182 5108
rect 3234 5096 3240 5108
rect 3234 5068 4650 5096
rect 3234 5056 3240 5068
rect 6014 4588 6020 4640
rect 6072 4588 6078 4640
rect 3260 4120 3266 4172
rect 3318 4160 3324 4172
rect 3318 4132 4650 4160
rect 3318 4120 3324 4132
rect 3596 4034 3602 4086
rect 3654 4074 3660 4086
rect 3654 4046 4746 4074
rect 3654 4034 3660 4046
rect 3848 3948 3854 4000
rect 3906 3988 3912 4000
rect 3906 3960 4842 3988
rect 3906 3948 3912 3960
rect 5956 3924 6032 3952
rect 3344 3862 3350 3914
rect 3402 3902 3408 3914
rect 3402 3874 4938 3902
rect 3402 3862 3408 3874
rect 2923 3782 2929 3834
rect 2981 3782 2987 3834
rect 3596 3776 3602 3828
rect 3654 3816 3660 3828
rect 3654 3788 5034 3816
rect 3654 3776 3660 3788
rect 5748 3778 6032 3806
rect 3848 3690 3854 3742
rect 3906 3730 3912 3742
rect 3906 3702 5130 3730
rect 3906 3690 3912 3702
rect 5666 3656 6032 3684
rect 3428 3604 3434 3656
rect 3486 3644 3492 3656
rect 3486 3616 5334 3644
rect 3486 3604 3492 3616
rect 3596 3518 3602 3570
rect 3654 3558 3660 3570
rect 3654 3530 5430 3558
rect 3654 3518 3660 3530
rect 3848 3432 3854 3484
rect 3906 3472 3912 3484
rect 3906 3444 5526 3472
rect 3906 3432 3912 3444
rect 6014 3050 6020 3102
rect 6072 3050 6078 3102
rect 3848 2668 3854 2720
rect 3906 2708 3912 2720
rect 3906 2680 5526 2708
rect 3906 2668 3912 2680
rect 3596 2582 3602 2634
rect 3654 2622 3660 2634
rect 3654 2594 5430 2622
rect 3654 2582 3660 2594
rect 3176 2496 3182 2548
rect 3234 2536 3240 2548
rect 3234 2508 5334 2536
rect 3234 2496 3240 2508
rect 5666 2468 6032 2496
rect 3848 2410 3854 2462
rect 3906 2450 3912 2462
rect 3906 2422 5130 2450
rect 3906 2410 3912 2422
rect 84 2326 90 2378
rect 142 2366 148 2378
rect 1216 2366 1222 2378
rect 142 2338 1222 2366
rect 142 2326 148 2338
rect 1216 2326 1222 2338
rect 1274 2326 1280 2378
rect 2923 2326 2929 2378
rect 2981 2326 2987 2378
rect 3512 2324 3518 2376
rect 3570 2364 3576 2376
rect 3570 2336 5034 2364
rect 5748 2346 6032 2374
rect 3570 2324 3576 2336
rect 3428 2238 3434 2290
rect 3486 2278 3492 2290
rect 3486 2250 4938 2278
rect 3486 2238 3492 2250
rect 3848 2152 3854 2204
rect 3906 2192 3912 2204
rect 5956 2200 6032 2228
rect 3906 2164 4842 2192
rect 3906 2152 3912 2164
rect 3512 2066 3518 2118
rect 3570 2106 3576 2118
rect 3570 2078 4746 2106
rect 3570 2066 3576 2078
rect 3344 1980 3350 2032
rect 3402 2020 3408 2032
rect 3402 1992 4650 2020
rect 3402 1980 3408 1992
rect 6014 1512 6020 1564
rect 6072 1512 6078 1564
rect 5956 848 6032 876
rect 3176 786 3182 838
rect 3234 826 3240 838
rect 3234 798 4938 826
rect 3234 786 3240 798
rect 0 702 6 754
rect 58 742 64 754
rect 1132 742 1138 754
rect 58 714 1138 742
rect 58 702 64 714
rect 1132 702 1138 714
rect 1190 702 1196 754
rect 2923 702 2929 754
rect 2981 702 2987 754
rect 3512 700 3518 752
rect 3570 740 3576 752
rect 3570 712 5034 740
rect 3570 700 3576 712
rect 5748 702 6032 730
rect 3848 614 3854 666
rect 3906 654 3912 666
rect 3906 626 5130 654
rect 3906 614 3912 626
rect 5666 580 6032 608
rect 3260 528 3266 580
rect 3318 568 3324 580
rect 3318 540 5334 568
rect 3318 528 3324 540
rect 3512 442 3518 494
rect 3570 482 3576 494
rect 3570 454 5430 482
rect 3570 442 3576 454
rect 3848 356 3854 408
rect 3906 396 3912 408
rect 3906 368 5526 396
rect 3906 356 3912 368
rect 6014 -26 6020 26
rect 6072 -26 6078 26
<< via1 >>
rect 6020 49190 6072 49242
rect 4274 48808 4326 48860
rect 3770 48722 3822 48774
rect 3350 48636 3402 48688
rect 4274 48550 4326 48602
rect 3770 48464 3822 48516
rect 3266 48378 3318 48430
rect 4274 48292 4326 48344
rect 3770 48206 3822 48258
rect 3182 48120 3234 48172
rect 6020 47652 6072 47704
rect 3266 47184 3318 47236
rect 3686 47098 3738 47150
rect 4274 47012 4326 47064
rect 3350 46926 3402 46978
rect 3686 46840 3738 46892
rect 4274 46754 4326 46806
rect 3434 46668 3486 46720
rect 3686 46582 3738 46634
rect 4274 46496 4326 46548
rect 6020 46114 6072 46166
rect 4274 45732 4326 45784
rect 3686 45646 3738 45698
rect 3182 45560 3234 45612
rect 4274 45474 4326 45526
rect 3602 45388 3654 45440
rect 3434 45302 3486 45354
rect 4274 45216 4326 45268
rect 3602 45130 3654 45182
rect 3350 45044 3402 45096
rect 6020 44576 6072 44628
rect 3434 44108 3486 44160
rect 3518 44022 3570 44074
rect 4274 43936 4326 43988
rect 3182 43850 3234 43902
rect 3602 43764 3654 43816
rect 4274 43678 4326 43730
rect 3266 43592 3318 43644
rect 3602 43506 3654 43558
rect 4274 43420 4326 43472
rect 6020 43038 6072 43090
rect 4274 42656 4326 42708
rect 3518 42570 3570 42622
rect 3350 42484 3402 42536
rect 4274 42398 4326 42450
rect 3518 42312 3570 42364
rect 3266 42226 3318 42278
rect 4274 42140 4326 42192
rect 3518 42054 3570 42106
rect 3182 41968 3234 42020
rect 6020 41500 6072 41552
rect 3266 41032 3318 41084
rect 3770 40946 3822 40998
rect 4190 40860 4242 40912
rect 3350 40774 3402 40826
rect 3770 40688 3822 40740
rect 4190 40602 4242 40654
rect 3434 40516 3486 40568
rect 3770 40430 3822 40482
rect 4190 40344 4242 40396
rect 6020 39962 6072 40014
rect 4190 39580 4242 39632
rect 3770 39494 3822 39546
rect 3182 39408 3234 39460
rect 4190 39322 4242 39374
rect 3686 39236 3738 39288
rect 3434 39150 3486 39202
rect 4190 39064 4242 39116
rect 3686 38978 3738 39030
rect 3350 38892 3402 38944
rect 6020 38424 6072 38476
rect 3434 37956 3486 38008
rect 3602 37870 3654 37922
rect 4190 37784 4242 37836
rect 3182 37698 3234 37750
rect 3686 37612 3738 37664
rect 4190 37526 4242 37578
rect 3266 37440 3318 37492
rect 3686 37354 3738 37406
rect 4190 37268 4242 37320
rect 6020 36886 6072 36938
rect 4190 36504 4242 36556
rect 3602 36418 3654 36470
rect 3350 36332 3402 36384
rect 4190 36246 4242 36298
rect 3602 36160 3654 36212
rect 3266 36074 3318 36126
rect 4190 35988 4242 36040
rect 3602 35902 3654 35954
rect 3182 35816 3234 35868
rect 6020 35348 6072 35400
rect 3266 34880 3318 34932
rect 3518 34794 3570 34846
rect 4190 34708 4242 34760
rect 3350 34622 3402 34674
rect 3518 34536 3570 34588
rect 4190 34450 4242 34502
rect 3434 34364 3486 34416
rect 3518 34278 3570 34330
rect 4190 34192 4242 34244
rect 6020 33810 6072 33862
rect 4190 33428 4242 33480
rect 3518 33342 3570 33394
rect 3182 33256 3234 33308
rect 4106 33170 4158 33222
rect 3770 33084 3822 33136
rect 3434 32998 3486 33050
rect 4106 32912 4158 32964
rect 3770 32826 3822 32878
rect 3350 32740 3402 32792
rect 6020 32272 6072 32324
rect 3434 31804 3486 31856
rect 3686 31718 3738 31770
rect 4106 31632 4158 31684
rect 3182 31546 3234 31598
rect 3770 31460 3822 31512
rect 4106 31374 4158 31426
rect 3266 31288 3318 31340
rect 3770 31202 3822 31254
rect 4106 31116 4158 31168
rect 6020 30734 6072 30786
rect 4106 30352 4158 30404
rect 3686 30266 3738 30318
rect 3350 30180 3402 30232
rect 4106 30094 4158 30146
rect 2929 30081 2981 30090
rect 2929 30047 2938 30081
rect 2938 30047 2972 30081
rect 2972 30047 2981 30081
rect 2929 30038 2981 30047
rect 3686 30008 3738 30060
rect 3266 29922 3318 29974
rect 4106 29836 4158 29888
rect 3686 29750 3738 29802
rect 3182 29664 3234 29716
rect 6020 29196 6072 29248
rect 3266 28728 3318 28780
rect 3602 28642 3654 28694
rect 4106 28556 4158 28608
rect 3350 28470 3402 28522
rect 2929 28457 2981 28466
rect 2929 28423 2938 28457
rect 2938 28423 2972 28457
rect 2972 28423 2981 28457
rect 2929 28414 2981 28423
rect 3602 28384 3654 28436
rect 4106 28298 4158 28350
rect 3434 28212 3486 28264
rect 3602 28126 3654 28178
rect 4106 28040 4158 28092
rect 6020 27658 6072 27710
rect 4106 27276 4158 27328
rect 3602 27190 3654 27242
rect 3182 27104 3234 27156
rect 4106 27018 4158 27070
rect 2929 27001 2981 27010
rect 2929 26967 2938 27001
rect 2938 26967 2972 27001
rect 2972 26967 2981 27001
rect 2929 26958 2981 26967
rect 3518 26932 3570 26984
rect 3434 26846 3486 26898
rect 4106 26760 4158 26812
rect 3518 26674 3570 26726
rect 3350 26588 3402 26640
rect 6020 26120 6072 26172
rect 3434 25652 3486 25704
rect 3770 25566 3822 25618
rect 4022 25480 4074 25532
rect 3182 25394 3234 25446
rect 2929 25377 2981 25386
rect 2929 25343 2938 25377
rect 2938 25343 2972 25377
rect 2972 25343 2981 25377
rect 2929 25334 2981 25343
rect 3518 25308 3570 25360
rect 4106 25222 4158 25274
rect 3266 25136 3318 25188
rect 3518 25050 3570 25102
rect 4106 24964 4158 25016
rect 6020 24582 6072 24634
rect 4022 24200 4074 24252
rect 3770 24114 3822 24166
rect 3350 24028 3402 24080
rect 4022 23942 4074 23994
rect 2929 23921 2981 23930
rect 2929 23887 2938 23921
rect 2938 23887 2972 23921
rect 2972 23887 2981 23921
rect 2929 23878 2981 23887
rect 3770 23856 3822 23908
rect 3266 23770 3318 23822
rect 4022 23684 4074 23736
rect 3770 23598 3822 23650
rect 3182 23512 3234 23564
rect 6020 23044 6072 23096
rect 3266 22576 3318 22628
rect 3686 22490 3738 22542
rect 4022 22404 4074 22456
rect 3350 22318 3402 22370
rect 510 22254 562 22306
rect 874 22254 926 22306
rect 2929 22297 2981 22306
rect 2929 22263 2938 22297
rect 2938 22263 2972 22297
rect 2972 22263 2981 22297
rect 2929 22254 2981 22263
rect 3686 22232 3738 22284
rect 4022 22146 4074 22198
rect 3434 22060 3486 22112
rect 3686 21974 3738 22026
rect 4022 21888 4074 21940
rect 6020 21506 6072 21558
rect 4022 21124 4074 21176
rect 3686 21038 3738 21090
rect 3182 20952 3234 21004
rect 4022 20866 4074 20918
rect 426 20798 478 20850
rect 790 20798 842 20850
rect 2929 20841 2981 20850
rect 2929 20807 2938 20841
rect 2938 20807 2972 20841
rect 2972 20807 2981 20841
rect 2929 20798 2981 20807
rect 3602 20780 3654 20832
rect 3434 20694 3486 20746
rect 4022 20608 4074 20660
rect 3602 20522 3654 20574
rect 3350 20436 3402 20488
rect 6020 19968 6072 20020
rect 3434 19500 3486 19552
rect 3518 19414 3570 19466
rect 4022 19328 4074 19380
rect 3182 19242 3234 19294
rect 342 19174 394 19226
rect 706 19174 758 19226
rect 2929 19217 2981 19226
rect 2929 19183 2938 19217
rect 2938 19183 2972 19217
rect 2972 19183 2981 19217
rect 2929 19174 2981 19183
rect 3602 19156 3654 19208
rect 4022 19070 4074 19122
rect 3266 18984 3318 19036
rect 3602 18898 3654 18950
rect 4022 18812 4074 18864
rect 6020 18430 6072 18482
rect 4022 18048 4074 18100
rect 3518 17962 3570 18014
rect 3350 17876 3402 17928
rect 4022 17790 4074 17842
rect 3518 17704 3570 17756
rect 3266 17618 3318 17670
rect 4022 17532 4074 17584
rect 3518 17446 3570 17498
rect 3182 17360 3234 17412
rect 6020 16892 6072 16944
rect 3266 16424 3318 16476
rect 3770 16338 3822 16390
rect 3938 16252 3990 16304
rect 3350 16166 3402 16218
rect 3770 16080 3822 16132
rect 3938 15994 3990 16046
rect 3434 15908 3486 15960
rect 3770 15822 3822 15874
rect 3938 15736 3990 15788
rect 6020 15354 6072 15406
rect 3938 14972 3990 15024
rect 3770 14886 3822 14938
rect 3182 14800 3234 14852
rect 3938 14714 3990 14766
rect 2929 14685 2981 14694
rect 2929 14651 2938 14685
rect 2938 14651 2972 14685
rect 2972 14651 2981 14685
rect 2929 14642 2981 14651
rect 3686 14628 3738 14680
rect 3434 14542 3486 14594
rect 3938 14456 3990 14508
rect 3686 14370 3738 14422
rect 3350 14284 3402 14336
rect 6020 13816 6072 13868
rect 3434 13348 3486 13400
rect 3602 13262 3654 13314
rect 3938 13176 3990 13228
rect 3182 13090 3234 13142
rect 2929 13061 2981 13070
rect 2929 13027 2938 13061
rect 2938 13027 2972 13061
rect 2972 13027 2981 13061
rect 2929 13018 2981 13027
rect 3686 13004 3738 13056
rect 3938 12918 3990 12970
rect 3266 12832 3318 12884
rect 3686 12746 3738 12798
rect 3938 12660 3990 12712
rect 6020 12278 6072 12330
rect 3938 11896 3990 11948
rect 3602 11810 3654 11862
rect 3350 11724 3402 11776
rect 3938 11638 3990 11690
rect 258 11562 310 11614
rect 1222 11562 1274 11614
rect 2929 11605 2981 11614
rect 2929 11571 2938 11605
rect 2938 11571 2972 11605
rect 2972 11571 2981 11605
rect 2929 11562 2981 11571
rect 3602 11552 3654 11604
rect 3266 11466 3318 11518
rect 3938 11380 3990 11432
rect 3602 11294 3654 11346
rect 3182 11208 3234 11260
rect 6020 10740 6072 10792
rect 3266 10272 3318 10324
rect 3518 10186 3570 10238
rect 3938 10100 3990 10152
rect 3350 10014 3402 10066
rect 174 9938 226 9990
rect 1138 9938 1190 9990
rect 2929 9981 2981 9990
rect 2929 9947 2938 9981
rect 2938 9947 2972 9981
rect 2972 9947 2981 9981
rect 2929 9938 2981 9947
rect 3518 9928 3570 9980
rect 3938 9842 3990 9894
rect 3434 9756 3486 9808
rect 3518 9670 3570 9722
rect 3938 9584 3990 9636
rect 6020 9202 6072 9254
rect 3938 8820 3990 8872
rect 3518 8734 3570 8786
rect 3182 8648 3234 8700
rect 3854 8562 3906 8614
rect 3770 8476 3822 8528
rect 3434 8390 3486 8442
rect 3854 8304 3906 8356
rect 3770 8218 3822 8270
rect 3350 8132 3402 8184
rect 6020 7664 6072 7716
rect 3434 7196 3486 7248
rect 3686 7110 3738 7162
rect 3854 7024 3906 7076
rect 3182 6938 3234 6990
rect 3770 6852 3822 6904
rect 3854 6766 3906 6818
rect 3266 6680 3318 6732
rect 3770 6594 3822 6646
rect 3854 6508 3906 6560
rect 6020 6126 6072 6178
rect 3854 5744 3906 5796
rect 3686 5658 3738 5710
rect 3350 5572 3402 5624
rect 3854 5486 3906 5538
rect 2929 5449 2981 5458
rect 2929 5415 2938 5449
rect 2938 5415 2972 5449
rect 2972 5415 2981 5449
rect 2929 5406 2981 5415
rect 3686 5400 3738 5452
rect 3266 5314 3318 5366
rect 3854 5228 3906 5280
rect 3686 5142 3738 5194
rect 3182 5056 3234 5108
rect 6020 4588 6072 4640
rect 3266 4120 3318 4172
rect 3602 4034 3654 4086
rect 3854 3948 3906 4000
rect 3350 3862 3402 3914
rect 2929 3825 2981 3834
rect 2929 3791 2938 3825
rect 2938 3791 2972 3825
rect 2972 3791 2981 3825
rect 2929 3782 2981 3791
rect 3602 3776 3654 3828
rect 3854 3690 3906 3742
rect 3434 3604 3486 3656
rect 3602 3518 3654 3570
rect 3854 3432 3906 3484
rect 6020 3050 6072 3102
rect 3854 2668 3906 2720
rect 3602 2582 3654 2634
rect 3182 2496 3234 2548
rect 3854 2410 3906 2462
rect 90 2326 142 2378
rect 1222 2326 1274 2378
rect 2929 2369 2981 2378
rect 2929 2335 2938 2369
rect 2938 2335 2972 2369
rect 2972 2335 2981 2369
rect 2929 2326 2981 2335
rect 3518 2324 3570 2376
rect 3434 2238 3486 2290
rect 3854 2152 3906 2204
rect 3518 2066 3570 2118
rect 3350 1980 3402 2032
rect 6020 1512 6072 1564
rect 3182 786 3234 838
rect 6 702 58 754
rect 1138 702 1190 754
rect 2929 745 2981 754
rect 2929 711 2938 745
rect 2938 711 2972 745
rect 2972 711 2981 745
rect 2929 702 2981 711
rect 3518 700 3570 752
rect 3854 614 3906 666
rect 3266 528 3318 580
rect 3518 442 3570 494
rect 3854 356 3906 408
rect 6020 -26 6072 26
<< metal2 >>
rect 6018 49244 6074 49253
rect 3194 48178 3222 49244
rect 3278 48436 3306 49244
rect 3362 48694 3390 49244
rect 3350 48688 3402 48694
rect 3350 48630 3402 48636
rect 3266 48430 3318 48436
rect 3266 48372 3318 48378
rect 3182 48172 3234 48178
rect 3182 48114 3234 48120
rect 3194 45618 3222 48114
rect 3278 47242 3306 48372
rect 3266 47236 3318 47242
rect 3266 47178 3318 47184
rect 3182 45612 3234 45618
rect 3182 45554 3234 45560
rect 3194 43908 3222 45554
rect 3182 43902 3234 43908
rect 3182 43844 3234 43850
rect 3194 42026 3222 43844
rect 3278 43650 3306 47178
rect 3362 46984 3390 48630
rect 3350 46978 3402 46984
rect 3350 46920 3402 46926
rect 3362 45102 3390 46920
rect 3446 46726 3474 49244
rect 3434 46720 3486 46726
rect 3434 46662 3486 46668
rect 3446 45360 3474 46662
rect 3434 45354 3486 45360
rect 3434 45296 3486 45302
rect 3350 45096 3402 45102
rect 3350 45038 3402 45044
rect 3266 43644 3318 43650
rect 3266 43586 3318 43592
rect 3278 42284 3306 43586
rect 3362 42542 3390 45038
rect 3446 44166 3474 45296
rect 3434 44160 3486 44166
rect 3434 44102 3486 44108
rect 3350 42536 3402 42542
rect 3350 42478 3402 42484
rect 3266 42278 3318 42284
rect 3266 42220 3318 42226
rect 3182 42020 3234 42026
rect 3182 41962 3234 41968
rect 3194 39466 3222 41962
rect 3278 41090 3306 42220
rect 3266 41084 3318 41090
rect 3266 41026 3318 41032
rect 3182 39460 3234 39466
rect 3182 39402 3234 39408
rect 3194 37756 3222 39402
rect 3182 37750 3234 37756
rect 3182 37692 3234 37698
rect 3194 35874 3222 37692
rect 3278 37498 3306 41026
rect 3362 40832 3390 42478
rect 3350 40826 3402 40832
rect 3350 40768 3402 40774
rect 3362 38950 3390 40768
rect 3446 40574 3474 44102
rect 3530 44080 3558 49244
rect 3614 45446 3642 49244
rect 3698 47156 3726 49244
rect 3782 48780 3810 49244
rect 3770 48774 3822 48780
rect 3770 48716 3822 48722
rect 3782 48522 3810 48716
rect 3770 48516 3822 48522
rect 3770 48458 3822 48464
rect 3782 48264 3810 48458
rect 3770 48258 3822 48264
rect 3770 48200 3822 48206
rect 3686 47150 3738 47156
rect 3686 47092 3738 47098
rect 3698 46898 3726 47092
rect 3686 46892 3738 46898
rect 3686 46834 3738 46840
rect 3698 46640 3726 46834
rect 3686 46634 3738 46640
rect 3686 46576 3738 46582
rect 3698 45704 3726 46576
rect 3686 45698 3738 45704
rect 3686 45640 3738 45646
rect 3602 45440 3654 45446
rect 3602 45382 3654 45388
rect 3614 45188 3642 45382
rect 3602 45182 3654 45188
rect 3602 45124 3654 45130
rect 3518 44074 3570 44080
rect 3518 44016 3570 44022
rect 3530 42628 3558 44016
rect 3614 43822 3642 45124
rect 3602 43816 3654 43822
rect 3602 43758 3654 43764
rect 3614 43564 3642 43758
rect 3602 43558 3654 43564
rect 3602 43500 3654 43506
rect 3518 42622 3570 42628
rect 3518 42564 3570 42570
rect 3530 42370 3558 42564
rect 3518 42364 3570 42370
rect 3518 42306 3570 42312
rect 3530 42112 3558 42306
rect 3518 42106 3570 42112
rect 3518 42048 3570 42054
rect 3434 40568 3486 40574
rect 3434 40510 3486 40516
rect 3446 39208 3474 40510
rect 3434 39202 3486 39208
rect 3434 39144 3486 39150
rect 3350 38944 3402 38950
rect 3350 38886 3402 38892
rect 3266 37492 3318 37498
rect 3266 37434 3318 37440
rect 3278 36132 3306 37434
rect 3362 36390 3390 38886
rect 3446 38014 3474 39144
rect 3434 38008 3486 38014
rect 3434 37950 3486 37956
rect 3350 36384 3402 36390
rect 3350 36326 3402 36332
rect 3266 36126 3318 36132
rect 3266 36068 3318 36074
rect 3182 35868 3234 35874
rect 3182 35810 3234 35816
rect 3194 33314 3222 35810
rect 3278 34938 3306 36068
rect 3266 34932 3318 34938
rect 3266 34874 3318 34880
rect 3182 33308 3234 33314
rect 3182 33250 3234 33256
rect 3194 31604 3222 33250
rect 3182 31598 3234 31604
rect 3182 31540 3234 31546
rect 18 760 46 30792
rect 102 2384 130 30792
rect 186 9996 214 30792
rect 270 11620 298 30792
rect 354 19232 382 30792
rect 438 20856 466 30792
rect 522 22312 550 30792
rect 2927 30092 2983 30101
rect 2927 30027 2983 30036
rect 3194 29722 3222 31540
rect 3278 31346 3306 34874
rect 3362 34680 3390 36326
rect 3350 34674 3402 34680
rect 3350 34616 3402 34622
rect 3362 32798 3390 34616
rect 3446 34422 3474 37950
rect 3530 34852 3558 42048
rect 3614 37928 3642 43500
rect 3698 39294 3726 45640
rect 3782 41004 3810 48200
rect 3770 40998 3822 41004
rect 3770 40940 3822 40946
rect 3782 40746 3810 40940
rect 3770 40740 3822 40746
rect 3770 40682 3822 40688
rect 3782 40488 3810 40682
rect 3770 40482 3822 40488
rect 3770 40424 3822 40430
rect 3782 39552 3810 40424
rect 3770 39546 3822 39552
rect 3770 39488 3822 39494
rect 3686 39288 3738 39294
rect 3686 39230 3738 39236
rect 3698 39036 3726 39230
rect 3686 39030 3738 39036
rect 3686 38972 3738 38978
rect 3602 37922 3654 37928
rect 3602 37864 3654 37870
rect 3614 36476 3642 37864
rect 3698 37670 3726 38972
rect 3686 37664 3738 37670
rect 3686 37606 3738 37612
rect 3698 37412 3726 37606
rect 3686 37406 3738 37412
rect 3686 37348 3738 37354
rect 3602 36470 3654 36476
rect 3602 36412 3654 36418
rect 3614 36218 3642 36412
rect 3602 36212 3654 36218
rect 3602 36154 3654 36160
rect 3614 35960 3642 36154
rect 3602 35954 3654 35960
rect 3602 35896 3654 35902
rect 3518 34846 3570 34852
rect 3518 34788 3570 34794
rect 3530 34594 3558 34788
rect 3518 34588 3570 34594
rect 3518 34530 3570 34536
rect 3434 34416 3486 34422
rect 3434 34358 3486 34364
rect 3446 33056 3474 34358
rect 3530 34336 3558 34530
rect 3518 34330 3570 34336
rect 3518 34272 3570 34278
rect 3530 33400 3558 34272
rect 3518 33394 3570 33400
rect 3518 33336 3570 33342
rect 3434 33050 3486 33056
rect 3434 32992 3486 32998
rect 3350 32792 3402 32798
rect 3350 32734 3402 32740
rect 3266 31340 3318 31346
rect 3266 31282 3318 31288
rect 3278 29980 3306 31282
rect 3362 30238 3390 32734
rect 3446 31862 3474 32992
rect 3434 31856 3486 31862
rect 3434 31798 3486 31804
rect 3350 30232 3402 30238
rect 3350 30174 3402 30180
rect 3266 29974 3318 29980
rect 3266 29916 3318 29922
rect 3182 29716 3234 29722
rect 3182 29658 3234 29664
rect 2927 28468 2983 28477
rect 2927 28403 2983 28412
rect 3194 27162 3222 29658
rect 3278 28786 3306 29916
rect 3266 28780 3318 28786
rect 3266 28722 3318 28728
rect 3182 27156 3234 27162
rect 3182 27098 3234 27104
rect 2927 27012 2983 27021
rect 2927 26947 2983 26956
rect 3194 25452 3222 27098
rect 3182 25446 3234 25452
rect 2927 25388 2983 25397
rect 3182 25388 3234 25394
rect 2927 25323 2983 25332
rect 2927 23932 2983 23941
rect 2927 23867 2983 23876
rect 3194 23570 3222 25388
rect 3278 25194 3306 28722
rect 3362 28528 3390 30174
rect 3350 28522 3402 28528
rect 3350 28464 3402 28470
rect 3362 26646 3390 28464
rect 3446 28270 3474 31798
rect 3434 28264 3486 28270
rect 3434 28206 3486 28212
rect 3446 26904 3474 28206
rect 3530 26990 3558 33336
rect 3614 28700 3642 35896
rect 3698 31776 3726 37348
rect 3782 33142 3810 39488
rect 3770 33136 3822 33142
rect 3770 33078 3822 33084
rect 3782 32884 3810 33078
rect 3770 32878 3822 32884
rect 3770 32820 3822 32826
rect 3686 31770 3738 31776
rect 3686 31712 3738 31718
rect 3698 30324 3726 31712
rect 3782 31518 3810 32820
rect 3770 31512 3822 31518
rect 3770 31454 3822 31460
rect 3782 31260 3810 31454
rect 3770 31254 3822 31260
rect 3770 31196 3822 31202
rect 3686 30318 3738 30324
rect 3686 30260 3738 30266
rect 3698 30066 3726 30260
rect 3686 30060 3738 30066
rect 3686 30002 3738 30008
rect 3698 29808 3726 30002
rect 3686 29802 3738 29808
rect 3686 29744 3738 29750
rect 3602 28694 3654 28700
rect 3602 28636 3654 28642
rect 3614 28442 3642 28636
rect 3602 28436 3654 28442
rect 3602 28378 3654 28384
rect 3614 28184 3642 28378
rect 3602 28178 3654 28184
rect 3602 28120 3654 28126
rect 3614 27248 3642 28120
rect 3602 27242 3654 27248
rect 3602 27184 3654 27190
rect 3518 26984 3570 26990
rect 3518 26926 3570 26932
rect 3434 26898 3486 26904
rect 3434 26840 3486 26846
rect 3350 26640 3402 26646
rect 3350 26582 3402 26588
rect 3266 25188 3318 25194
rect 3266 25130 3318 25136
rect 3278 23828 3306 25130
rect 3362 24086 3390 26582
rect 3446 25710 3474 26840
rect 3530 26732 3558 26926
rect 3518 26726 3570 26732
rect 3518 26668 3570 26674
rect 3434 25704 3486 25710
rect 3434 25646 3486 25652
rect 3350 24080 3402 24086
rect 3350 24022 3402 24028
rect 3266 23822 3318 23828
rect 3266 23764 3318 23770
rect 3182 23564 3234 23570
rect 3182 23506 3234 23512
rect 510 22306 562 22312
rect 510 22248 562 22254
rect 874 22306 926 22312
rect 874 22248 926 22254
rect 2927 22308 2983 22317
rect 426 20850 478 20856
rect 426 20792 478 20798
rect 342 19226 394 19232
rect 342 19168 394 19174
rect 258 11614 310 11620
rect 258 11556 310 11562
rect 174 9990 226 9996
rect 174 9932 226 9938
rect 90 2378 142 2384
rect 90 2320 142 2326
rect 6 754 58 760
rect 6 696 58 702
rect 18 0 46 696
rect 102 0 130 2320
rect 186 0 214 9932
rect 270 0 298 11556
rect 354 0 382 19168
rect 438 0 466 20792
rect 522 0 550 22248
rect 2927 22243 2983 22252
rect 3194 21010 3222 23506
rect 3278 22634 3306 23764
rect 3266 22628 3318 22634
rect 3266 22570 3318 22576
rect 3182 21004 3234 21010
rect 3182 20946 3234 20952
rect 790 20850 842 20856
rect 790 20792 842 20798
rect 2927 20852 2983 20861
rect 2927 20787 2983 20796
rect 3194 19300 3222 20946
rect 3182 19294 3234 19300
rect 706 19226 758 19232
rect 706 19168 758 19174
rect 2927 19228 2983 19237
rect 3182 19236 3234 19242
rect 2927 19163 2983 19172
rect 3194 17418 3222 19236
rect 3278 19042 3306 22570
rect 3362 22376 3390 24022
rect 3350 22370 3402 22376
rect 3350 22312 3402 22318
rect 3362 20494 3390 22312
rect 3446 22118 3474 25646
rect 3530 25366 3558 26668
rect 3518 25360 3570 25366
rect 3518 25302 3570 25308
rect 3530 25108 3558 25302
rect 3518 25102 3570 25108
rect 3518 25044 3570 25050
rect 3434 22112 3486 22118
rect 3434 22054 3486 22060
rect 3446 20752 3474 22054
rect 3434 20746 3486 20752
rect 3434 20688 3486 20694
rect 3350 20488 3402 20494
rect 3350 20430 3402 20436
rect 3266 19036 3318 19042
rect 3266 18978 3318 18984
rect 3278 17676 3306 18978
rect 3362 17934 3390 20430
rect 3446 19558 3474 20688
rect 3434 19552 3486 19558
rect 3434 19494 3486 19500
rect 3350 17928 3402 17934
rect 3350 17870 3402 17876
rect 3266 17670 3318 17676
rect 3266 17612 3318 17618
rect 3182 17412 3234 17418
rect 3182 17354 3234 17360
rect 3194 14858 3222 17354
rect 3278 16482 3306 17612
rect 3266 16476 3318 16482
rect 3266 16418 3318 16424
rect 3182 14852 3234 14858
rect 3182 14794 3234 14800
rect 2927 14696 2983 14705
rect 2927 14631 2983 14640
rect 3194 13148 3222 14794
rect 3182 13142 3234 13148
rect 3182 13084 3234 13090
rect 2927 13072 2983 13081
rect 2927 13007 2983 13016
rect 1222 11614 1274 11620
rect 1222 11556 1274 11562
rect 2927 11616 2983 11625
rect 2927 11551 2983 11560
rect 3194 11266 3222 13084
rect 3278 12890 3306 16418
rect 3362 16224 3390 17870
rect 3350 16218 3402 16224
rect 3350 16160 3402 16166
rect 3362 14342 3390 16160
rect 3446 15966 3474 19494
rect 3530 19472 3558 25044
rect 3614 20838 3642 27184
rect 3698 22548 3726 29744
rect 3782 25624 3810 31196
rect 3770 25618 3822 25624
rect 3770 25560 3822 25566
rect 3782 24172 3810 25560
rect 3770 24166 3822 24172
rect 3770 24108 3822 24114
rect 3782 23914 3810 24108
rect 3770 23908 3822 23914
rect 3770 23850 3822 23856
rect 3782 23656 3810 23850
rect 3770 23650 3822 23656
rect 3770 23592 3822 23598
rect 3686 22542 3738 22548
rect 3686 22484 3738 22490
rect 3698 22290 3726 22484
rect 3686 22284 3738 22290
rect 3686 22226 3738 22232
rect 3698 22032 3726 22226
rect 3686 22026 3738 22032
rect 3686 21968 3738 21974
rect 3698 21096 3726 21968
rect 3686 21090 3738 21096
rect 3686 21032 3738 21038
rect 3602 20832 3654 20838
rect 3602 20774 3654 20780
rect 3614 20580 3642 20774
rect 3602 20574 3654 20580
rect 3602 20516 3654 20522
rect 3518 19466 3570 19472
rect 3518 19408 3570 19414
rect 3530 18020 3558 19408
rect 3614 19214 3642 20516
rect 3602 19208 3654 19214
rect 3602 19150 3654 19156
rect 3614 18956 3642 19150
rect 3602 18950 3654 18956
rect 3602 18892 3654 18898
rect 3518 18014 3570 18020
rect 3518 17956 3570 17962
rect 3530 17762 3558 17956
rect 3518 17756 3570 17762
rect 3518 17698 3570 17704
rect 3530 17504 3558 17698
rect 3518 17498 3570 17504
rect 3518 17440 3570 17446
rect 3434 15960 3486 15966
rect 3434 15902 3486 15908
rect 3446 14600 3474 15902
rect 3434 14594 3486 14600
rect 3434 14536 3486 14542
rect 3350 14336 3402 14342
rect 3350 14278 3402 14284
rect 3266 12884 3318 12890
rect 3266 12826 3318 12832
rect 3278 11524 3306 12826
rect 3362 11782 3390 14278
rect 3446 13406 3474 14536
rect 3434 13400 3486 13406
rect 3434 13342 3486 13348
rect 3350 11776 3402 11782
rect 3350 11718 3402 11724
rect 3266 11518 3318 11524
rect 3266 11460 3318 11466
rect 3182 11260 3234 11266
rect 3182 11202 3234 11208
rect 1138 9990 1190 9996
rect 1138 9932 1190 9938
rect 2927 9992 2983 10001
rect 2927 9927 2983 9936
rect 3194 8706 3222 11202
rect 3278 10330 3306 11460
rect 3266 10324 3318 10330
rect 3266 10266 3318 10272
rect 3182 8700 3234 8706
rect 3182 8642 3234 8648
rect 3194 6996 3222 8642
rect 3182 6990 3234 6996
rect 3182 6932 3234 6938
rect 2927 5460 2983 5469
rect 2927 5395 2983 5404
rect 3194 5114 3222 6932
rect 3278 6738 3306 10266
rect 3362 10072 3390 11718
rect 3350 10066 3402 10072
rect 3350 10008 3402 10014
rect 3362 8190 3390 10008
rect 3446 9814 3474 13342
rect 3530 10244 3558 17440
rect 3614 13320 3642 18892
rect 3698 14686 3726 21032
rect 3782 16396 3810 23592
rect 3866 18509 3894 49244
rect 3950 20049 3978 49244
rect 4034 25538 4062 49244
rect 4118 33228 4146 49244
rect 4202 40918 4230 49244
rect 4286 48866 4314 49244
rect 4274 48860 4326 48866
rect 4274 48802 4326 48808
rect 4286 48608 4314 48802
rect 4274 48602 4326 48608
rect 4274 48544 4326 48550
rect 4286 48350 4314 48544
rect 4274 48344 4326 48350
rect 4274 48286 4326 48292
rect 4286 47070 4314 48286
rect 4274 47064 4326 47070
rect 4274 47006 4326 47012
rect 4286 46812 4314 47006
rect 4274 46806 4326 46812
rect 4274 46748 4326 46754
rect 4286 46554 4314 46748
rect 4274 46548 4326 46554
rect 4274 46490 4326 46496
rect 4286 45790 4314 46490
rect 4274 45784 4326 45790
rect 4274 45726 4326 45732
rect 4286 45532 4314 45726
rect 4274 45526 4326 45532
rect 4274 45468 4326 45474
rect 4286 45274 4314 45468
rect 4274 45268 4326 45274
rect 4274 45210 4326 45216
rect 4286 43994 4314 45210
rect 4274 43988 4326 43994
rect 4274 43930 4326 43936
rect 4286 43736 4314 43930
rect 4274 43730 4326 43736
rect 4274 43672 4326 43678
rect 4286 43478 4314 43672
rect 4274 43472 4326 43478
rect 4274 43414 4326 43420
rect 4286 42714 4314 43414
rect 4274 42708 4326 42714
rect 4274 42650 4326 42656
rect 4286 42456 4314 42650
rect 4274 42450 4326 42456
rect 4274 42392 4326 42398
rect 4286 42198 4314 42392
rect 4274 42192 4326 42198
rect 4274 42134 4326 42140
rect 4190 40912 4242 40918
rect 4190 40854 4242 40860
rect 4202 40660 4230 40854
rect 4190 40654 4242 40660
rect 4190 40596 4242 40602
rect 4202 40402 4230 40596
rect 4190 40396 4242 40402
rect 4190 40338 4242 40344
rect 4202 39638 4230 40338
rect 4190 39632 4242 39638
rect 4190 39574 4242 39580
rect 4202 39380 4230 39574
rect 4190 39374 4242 39380
rect 4190 39316 4242 39322
rect 4202 39122 4230 39316
rect 4190 39116 4242 39122
rect 4190 39058 4242 39064
rect 4202 37842 4230 39058
rect 4190 37836 4242 37842
rect 4190 37778 4242 37784
rect 4202 37584 4230 37778
rect 4190 37578 4242 37584
rect 4190 37520 4242 37526
rect 4202 37326 4230 37520
rect 4190 37320 4242 37326
rect 4190 37262 4242 37268
rect 4202 36562 4230 37262
rect 4190 36556 4242 36562
rect 4190 36498 4242 36504
rect 4202 36304 4230 36498
rect 4190 36298 4242 36304
rect 4190 36240 4242 36246
rect 4202 36046 4230 36240
rect 4190 36040 4242 36046
rect 4190 35982 4242 35988
rect 4202 34766 4230 35982
rect 4190 34760 4242 34766
rect 4190 34702 4242 34708
rect 4202 34508 4230 34702
rect 4190 34502 4242 34508
rect 4190 34444 4242 34450
rect 4202 34250 4230 34444
rect 4190 34244 4242 34250
rect 4190 34186 4242 34192
rect 4202 33486 4230 34186
rect 4190 33480 4242 33486
rect 4190 33422 4242 33428
rect 4106 33222 4158 33228
rect 4106 33164 4158 33170
rect 4118 32970 4146 33164
rect 4106 32964 4158 32970
rect 4106 32906 4158 32912
rect 4118 31690 4146 32906
rect 4106 31684 4158 31690
rect 4106 31626 4158 31632
rect 4118 31432 4146 31626
rect 4106 31426 4158 31432
rect 4106 31368 4158 31374
rect 4118 31174 4146 31368
rect 4106 31168 4158 31174
rect 4106 31110 4158 31116
rect 4118 30410 4146 31110
rect 4106 30404 4158 30410
rect 4106 30346 4158 30352
rect 4118 30152 4146 30346
rect 4106 30146 4158 30152
rect 4106 30088 4158 30094
rect 4118 29894 4146 30088
rect 4106 29888 4158 29894
rect 4106 29830 4158 29836
rect 4118 28614 4146 29830
rect 4106 28608 4158 28614
rect 4106 28550 4158 28556
rect 4118 28356 4146 28550
rect 4106 28350 4158 28356
rect 4106 28292 4158 28298
rect 4118 28098 4146 28292
rect 4106 28092 4158 28098
rect 4106 28034 4158 28040
rect 4118 27334 4146 28034
rect 4106 27328 4158 27334
rect 4106 27270 4158 27276
rect 4118 27076 4146 27270
rect 4106 27070 4158 27076
rect 4106 27012 4158 27018
rect 4118 26818 4146 27012
rect 4106 26812 4158 26818
rect 4106 26754 4158 26760
rect 4022 25532 4074 25538
rect 4022 25474 4074 25480
rect 4034 24258 4062 25474
rect 4118 25280 4146 26754
rect 4106 25274 4158 25280
rect 4106 25216 4158 25222
rect 4118 25022 4146 25216
rect 4106 25016 4158 25022
rect 4106 24958 4158 24964
rect 4022 24252 4074 24258
rect 4022 24194 4074 24200
rect 4034 24000 4062 24194
rect 4022 23994 4074 24000
rect 4022 23936 4074 23942
rect 4034 23742 4062 23936
rect 4022 23736 4074 23742
rect 4022 23678 4074 23684
rect 4034 22462 4062 23678
rect 4118 23129 4146 24958
rect 4202 24669 4230 33422
rect 4286 26209 4314 42134
rect 4370 27749 4398 49244
rect 4454 29289 4482 49244
rect 6018 49179 6074 49188
rect 6018 47706 6074 47715
rect 6018 47641 6074 47650
rect 6018 46168 6074 46177
rect 6018 46103 6074 46112
rect 6018 44630 6074 44639
rect 6018 44565 6074 44574
rect 6018 43092 6074 43101
rect 6018 43027 6074 43036
rect 6018 41554 6074 41563
rect 6018 41489 6074 41498
rect 6018 40016 6074 40025
rect 6018 39951 6074 39960
rect 6018 38478 6074 38487
rect 6018 38413 6074 38422
rect 6018 36940 6074 36949
rect 6018 36875 6074 36884
rect 6018 35402 6074 35411
rect 6018 35337 6074 35346
rect 6018 33864 6074 33873
rect 6018 33799 6074 33808
rect 6018 32326 6074 32335
rect 6018 32261 6074 32270
rect 6018 30788 6074 30797
rect 6018 30723 6074 30732
rect 4440 29280 4496 29289
rect 4440 29215 4496 29224
rect 6018 29250 6074 29259
rect 4356 27740 4412 27749
rect 4356 27675 4412 27684
rect 4272 26200 4328 26209
rect 4272 26135 4328 26144
rect 4188 24660 4244 24669
rect 4188 24595 4244 24604
rect 4104 23120 4160 23129
rect 4104 23055 4160 23064
rect 4022 22456 4074 22462
rect 4022 22398 4074 22404
rect 4034 22204 4062 22398
rect 4022 22198 4074 22204
rect 4022 22140 4074 22146
rect 4034 21946 4062 22140
rect 4022 21940 4074 21946
rect 4022 21882 4074 21888
rect 4034 21589 4062 21882
rect 4020 21580 4076 21589
rect 4020 21515 4076 21524
rect 4034 21182 4062 21515
rect 4022 21176 4074 21182
rect 4022 21118 4074 21124
rect 4034 20924 4062 21118
rect 4022 20918 4074 20924
rect 4022 20860 4074 20866
rect 4034 20666 4062 20860
rect 4022 20660 4074 20666
rect 4022 20602 4074 20608
rect 3936 20040 3992 20049
rect 3936 19975 3992 19984
rect 3852 18500 3908 18509
rect 3852 18435 3908 18444
rect 3770 16390 3822 16396
rect 3770 16332 3822 16338
rect 3782 16138 3810 16332
rect 3770 16132 3822 16138
rect 3770 16074 3822 16080
rect 3782 15880 3810 16074
rect 3770 15874 3822 15880
rect 3770 15816 3822 15822
rect 3782 14944 3810 15816
rect 3770 14938 3822 14944
rect 3770 14880 3822 14886
rect 3686 14680 3738 14686
rect 3686 14622 3738 14628
rect 3698 14428 3726 14622
rect 3686 14422 3738 14428
rect 3686 14364 3738 14370
rect 3602 13314 3654 13320
rect 3602 13256 3654 13262
rect 3614 11868 3642 13256
rect 3698 13062 3726 14364
rect 3782 13893 3810 14880
rect 3768 13884 3824 13893
rect 3768 13819 3824 13828
rect 3686 13056 3738 13062
rect 3686 12998 3738 13004
rect 3698 12804 3726 12998
rect 3686 12798 3738 12804
rect 3686 12740 3738 12746
rect 3698 12353 3726 12740
rect 3684 12344 3740 12353
rect 3684 12279 3740 12288
rect 3602 11862 3654 11868
rect 3602 11804 3654 11810
rect 3614 11610 3642 11804
rect 3602 11604 3654 11610
rect 3602 11546 3654 11552
rect 3614 11352 3642 11546
rect 3602 11346 3654 11352
rect 3602 11288 3654 11294
rect 3614 10813 3642 11288
rect 3600 10804 3656 10813
rect 3600 10739 3656 10748
rect 3518 10238 3570 10244
rect 3518 10180 3570 10186
rect 3530 9986 3558 10180
rect 3518 9980 3570 9986
rect 3518 9922 3570 9928
rect 3434 9808 3486 9814
rect 3434 9750 3486 9756
rect 3446 8448 3474 9750
rect 3530 9728 3558 9922
rect 3518 9722 3570 9728
rect 3518 9664 3570 9670
rect 3530 9273 3558 9664
rect 3516 9264 3572 9273
rect 3516 9199 3572 9208
rect 3530 8792 3558 9199
rect 3518 8786 3570 8792
rect 3518 8728 3570 8734
rect 3434 8442 3486 8448
rect 3434 8384 3486 8390
rect 3350 8184 3402 8190
rect 3350 8126 3402 8132
rect 3266 6732 3318 6738
rect 3266 6674 3318 6680
rect 3278 5372 3306 6674
rect 3362 5630 3390 8126
rect 3446 7254 3474 8384
rect 3434 7248 3486 7254
rect 3434 7190 3486 7196
rect 3350 5624 3402 5630
rect 3350 5566 3402 5572
rect 3266 5366 3318 5372
rect 3266 5308 3318 5314
rect 3182 5108 3234 5114
rect 3182 5050 3234 5056
rect 2927 3836 2983 3845
rect 2927 3771 2983 3780
rect 3194 2554 3222 5050
rect 3278 4178 3306 5308
rect 3266 4172 3318 4178
rect 3266 4114 3318 4120
rect 3182 2548 3234 2554
rect 3182 2490 3234 2496
rect 1222 2378 1274 2384
rect 1222 2320 1274 2326
rect 2927 2380 2983 2389
rect 2927 2315 2983 2324
rect 3194 844 3222 2490
rect 3278 1577 3306 4114
rect 3362 3920 3390 5566
rect 3446 4657 3474 7190
rect 3432 4648 3488 4657
rect 3432 4583 3488 4592
rect 3350 3914 3402 3920
rect 3350 3856 3402 3862
rect 3362 3117 3390 3856
rect 3446 3662 3474 4583
rect 3434 3656 3486 3662
rect 3434 3598 3486 3604
rect 3348 3108 3404 3117
rect 3348 3043 3404 3052
rect 3362 2038 3390 3043
rect 3446 2296 3474 3598
rect 3530 2382 3558 8728
rect 3614 4092 3642 10739
rect 3698 7168 3726 12279
rect 3782 8534 3810 13819
rect 3866 8620 3894 18435
rect 3950 16310 3978 19975
rect 4034 19386 4062 20602
rect 4022 19380 4074 19386
rect 4022 19322 4074 19328
rect 4034 19128 4062 19322
rect 4022 19122 4074 19128
rect 4022 19064 4074 19070
rect 4034 18870 4062 19064
rect 4022 18864 4074 18870
rect 4022 18806 4074 18812
rect 4034 18106 4062 18806
rect 4022 18100 4074 18106
rect 4022 18042 4074 18048
rect 4034 17848 4062 18042
rect 4022 17842 4074 17848
rect 4022 17784 4074 17790
rect 4034 17590 4062 17784
rect 4022 17584 4074 17590
rect 4022 17526 4074 17532
rect 3938 16304 3990 16310
rect 3938 16246 3990 16252
rect 3950 16052 3978 16246
rect 3938 16046 3990 16052
rect 3938 15988 3990 15994
rect 3950 15794 3978 15988
rect 3938 15788 3990 15794
rect 3938 15730 3990 15736
rect 3950 15030 3978 15730
rect 3938 15024 3990 15030
rect 3938 14966 3990 14972
rect 3950 14772 3978 14966
rect 3938 14766 3990 14772
rect 3938 14708 3990 14714
rect 3950 14514 3978 14708
rect 3938 14508 3990 14514
rect 3938 14450 3990 14456
rect 3950 13234 3978 14450
rect 3938 13228 3990 13234
rect 3938 13170 3990 13176
rect 3950 12976 3978 13170
rect 3938 12970 3990 12976
rect 3938 12912 3990 12918
rect 3950 12718 3978 12912
rect 3938 12712 3990 12718
rect 3938 12654 3990 12660
rect 3950 11954 3978 12654
rect 3938 11948 3990 11954
rect 3938 11890 3990 11896
rect 3950 11696 3978 11890
rect 3938 11690 3990 11696
rect 3938 11632 3990 11638
rect 3950 11438 3978 11632
rect 3938 11432 3990 11438
rect 3938 11374 3990 11380
rect 3950 10158 3978 11374
rect 3938 10152 3990 10158
rect 3938 10094 3990 10100
rect 3950 9900 3978 10094
rect 3938 9894 3990 9900
rect 3938 9836 3990 9842
rect 3950 9642 3978 9836
rect 3938 9636 3990 9642
rect 3938 9578 3990 9584
rect 3950 8878 3978 9578
rect 3938 8872 3990 8878
rect 3938 8814 3990 8820
rect 3854 8614 3906 8620
rect 3854 8556 3906 8562
rect 3770 8528 3822 8534
rect 3770 8470 3822 8476
rect 3782 8276 3810 8470
rect 3866 8362 3894 8556
rect 3854 8356 3906 8362
rect 3854 8298 3906 8304
rect 3770 8270 3822 8276
rect 3770 8212 3822 8218
rect 3686 7162 3738 7168
rect 3686 7104 3738 7110
rect 3698 5716 3726 7104
rect 3782 6910 3810 8212
rect 3866 7082 3894 8298
rect 3854 7076 3906 7082
rect 3854 7018 3906 7024
rect 3770 6904 3822 6910
rect 3770 6846 3822 6852
rect 3782 6652 3810 6846
rect 3866 6824 3894 7018
rect 3854 6818 3906 6824
rect 3854 6760 3906 6766
rect 3770 6646 3822 6652
rect 3770 6588 3822 6594
rect 3686 5710 3738 5716
rect 3686 5652 3738 5658
rect 3698 5458 3726 5652
rect 3686 5452 3738 5458
rect 3686 5394 3738 5400
rect 3698 5200 3726 5394
rect 3686 5194 3738 5200
rect 3686 5136 3738 5142
rect 3602 4086 3654 4092
rect 3602 4028 3654 4034
rect 3614 3834 3642 4028
rect 3602 3828 3654 3834
rect 3602 3770 3654 3776
rect 3614 3576 3642 3770
rect 3602 3570 3654 3576
rect 3602 3512 3654 3518
rect 3614 2640 3642 3512
rect 3602 2634 3654 2640
rect 3602 2576 3654 2582
rect 3518 2376 3570 2382
rect 3518 2318 3570 2324
rect 3434 2290 3486 2296
rect 3434 2232 3486 2238
rect 3350 2032 3402 2038
rect 3350 1974 3402 1980
rect 3264 1568 3320 1577
rect 3264 1503 3320 1512
rect 3182 838 3234 844
rect 3182 780 3234 786
rect 1138 754 1190 760
rect 1138 696 1190 702
rect 2927 756 2983 765
rect 2927 691 2983 700
rect 3194 37 3222 780
rect 3278 586 3306 1503
rect 3266 580 3318 586
rect 3266 522 3318 528
rect 3180 28 3236 37
rect 3278 0 3306 522
rect 3362 0 3390 1974
rect 3446 0 3474 2232
rect 3530 2124 3558 2318
rect 3518 2118 3570 2124
rect 3518 2060 3570 2066
rect 3530 758 3558 2060
rect 3518 752 3570 758
rect 3518 694 3570 700
rect 3530 500 3558 694
rect 3518 494 3570 500
rect 3518 436 3570 442
rect 3530 0 3558 436
rect 3614 0 3642 2576
rect 3698 0 3726 5136
rect 3782 0 3810 6588
rect 3866 6566 3894 6760
rect 3854 6560 3906 6566
rect 3854 6502 3906 6508
rect 3866 5802 3894 6502
rect 3854 5796 3906 5802
rect 3854 5738 3906 5744
rect 3866 5544 3894 5738
rect 3854 5538 3906 5544
rect 3854 5480 3906 5486
rect 3866 5286 3894 5480
rect 3854 5280 3906 5286
rect 3854 5222 3906 5228
rect 3866 4006 3894 5222
rect 3854 4000 3906 4006
rect 3854 3942 3906 3948
rect 3866 3748 3894 3942
rect 3854 3742 3906 3748
rect 3854 3684 3906 3690
rect 3866 3490 3894 3684
rect 3854 3484 3906 3490
rect 3854 3426 3906 3432
rect 3866 2726 3894 3426
rect 3854 2720 3906 2726
rect 3854 2662 3906 2668
rect 3866 2468 3894 2662
rect 3854 2462 3906 2468
rect 3854 2404 3906 2410
rect 3866 2210 3894 2404
rect 3854 2204 3906 2210
rect 3854 2146 3906 2152
rect 3866 672 3894 2146
rect 3854 666 3906 672
rect 3854 608 3906 614
rect 3866 414 3894 608
rect 3854 408 3906 414
rect 3854 350 3906 356
rect 3866 0 3894 350
rect 3950 0 3978 8814
rect 4034 0 4062 17526
rect 4118 0 4146 23055
rect 4202 0 4230 24595
rect 4286 0 4314 26135
rect 4370 0 4398 27675
rect 4454 0 4482 29215
rect 6018 29185 6074 29194
rect 6018 27712 6074 27721
rect 6018 27647 6074 27656
rect 6018 26174 6074 26183
rect 6018 26109 6074 26118
rect 6018 24636 6074 24645
rect 6018 24571 6074 24580
rect 6018 23098 6074 23107
rect 6018 23033 6074 23042
rect 6018 21560 6074 21569
rect 6018 21495 6074 21504
rect 6018 20022 6074 20031
rect 6018 19957 6074 19966
rect 6018 18484 6074 18493
rect 6018 18419 6074 18428
rect 6018 16946 6074 16955
rect 6018 16881 6074 16890
rect 6018 15408 6074 15417
rect 6018 15343 6074 15352
rect 6018 13870 6074 13879
rect 6018 13805 6074 13814
rect 6018 12332 6074 12341
rect 6018 12267 6074 12276
rect 6018 10794 6074 10803
rect 6018 10729 6074 10738
rect 6018 9256 6074 9265
rect 6018 9191 6074 9200
rect 6018 7718 6074 7727
rect 6018 7653 6074 7662
rect 6018 6180 6074 6189
rect 6018 6115 6074 6124
rect 6018 4642 6074 4651
rect 6018 4577 6074 4586
rect 6018 3104 6074 3113
rect 6018 3039 6074 3048
rect 6018 1566 6074 1575
rect 6018 1501 6074 1510
rect 6018 28 6074 37
rect 3180 -37 3236 -28
rect 6018 -37 6074 -28
<< via2 >>
rect 2927 30090 2983 30092
rect 2927 30038 2929 30090
rect 2929 30038 2981 30090
rect 2981 30038 2983 30090
rect 2927 30036 2983 30038
rect 2927 28466 2983 28468
rect 2927 28414 2929 28466
rect 2929 28414 2981 28466
rect 2981 28414 2983 28466
rect 2927 28412 2983 28414
rect 2927 27010 2983 27012
rect 2927 26958 2929 27010
rect 2929 26958 2981 27010
rect 2981 26958 2983 27010
rect 2927 26956 2983 26958
rect 2927 25386 2983 25388
rect 2927 25334 2929 25386
rect 2929 25334 2981 25386
rect 2981 25334 2983 25386
rect 2927 25332 2983 25334
rect 2927 23930 2983 23932
rect 2927 23878 2929 23930
rect 2929 23878 2981 23930
rect 2981 23878 2983 23930
rect 2927 23876 2983 23878
rect 2927 22306 2983 22308
rect 2927 22254 2929 22306
rect 2929 22254 2981 22306
rect 2981 22254 2983 22306
rect 2927 22252 2983 22254
rect 2927 20850 2983 20852
rect 2927 20798 2929 20850
rect 2929 20798 2981 20850
rect 2981 20798 2983 20850
rect 2927 20796 2983 20798
rect 2927 19226 2983 19228
rect 2927 19174 2929 19226
rect 2929 19174 2981 19226
rect 2981 19174 2983 19226
rect 2927 19172 2983 19174
rect 2927 14694 2983 14696
rect 2927 14642 2929 14694
rect 2929 14642 2981 14694
rect 2981 14642 2983 14694
rect 2927 14640 2983 14642
rect 2927 13070 2983 13072
rect 2927 13018 2929 13070
rect 2929 13018 2981 13070
rect 2981 13018 2983 13070
rect 2927 13016 2983 13018
rect 2927 11614 2983 11616
rect 2927 11562 2929 11614
rect 2929 11562 2981 11614
rect 2981 11562 2983 11614
rect 2927 11560 2983 11562
rect 2927 9990 2983 9992
rect 2927 9938 2929 9990
rect 2929 9938 2981 9990
rect 2981 9938 2983 9990
rect 2927 9936 2983 9938
rect 2927 5458 2983 5460
rect 2927 5406 2929 5458
rect 2929 5406 2981 5458
rect 2981 5406 2983 5458
rect 2927 5404 2983 5406
rect 6018 49242 6074 49244
rect 6018 49190 6020 49242
rect 6020 49190 6072 49242
rect 6072 49190 6074 49242
rect 6018 49188 6074 49190
rect 6018 47704 6074 47706
rect 6018 47652 6020 47704
rect 6020 47652 6072 47704
rect 6072 47652 6074 47704
rect 6018 47650 6074 47652
rect 6018 46166 6074 46168
rect 6018 46114 6020 46166
rect 6020 46114 6072 46166
rect 6072 46114 6074 46166
rect 6018 46112 6074 46114
rect 6018 44628 6074 44630
rect 6018 44576 6020 44628
rect 6020 44576 6072 44628
rect 6072 44576 6074 44628
rect 6018 44574 6074 44576
rect 6018 43090 6074 43092
rect 6018 43038 6020 43090
rect 6020 43038 6072 43090
rect 6072 43038 6074 43090
rect 6018 43036 6074 43038
rect 6018 41552 6074 41554
rect 6018 41500 6020 41552
rect 6020 41500 6072 41552
rect 6072 41500 6074 41552
rect 6018 41498 6074 41500
rect 6018 40014 6074 40016
rect 6018 39962 6020 40014
rect 6020 39962 6072 40014
rect 6072 39962 6074 40014
rect 6018 39960 6074 39962
rect 6018 38476 6074 38478
rect 6018 38424 6020 38476
rect 6020 38424 6072 38476
rect 6072 38424 6074 38476
rect 6018 38422 6074 38424
rect 6018 36938 6074 36940
rect 6018 36886 6020 36938
rect 6020 36886 6072 36938
rect 6072 36886 6074 36938
rect 6018 36884 6074 36886
rect 6018 35400 6074 35402
rect 6018 35348 6020 35400
rect 6020 35348 6072 35400
rect 6072 35348 6074 35400
rect 6018 35346 6074 35348
rect 6018 33862 6074 33864
rect 6018 33810 6020 33862
rect 6020 33810 6072 33862
rect 6072 33810 6074 33862
rect 6018 33808 6074 33810
rect 6018 32324 6074 32326
rect 6018 32272 6020 32324
rect 6020 32272 6072 32324
rect 6072 32272 6074 32324
rect 6018 32270 6074 32272
rect 6018 30786 6074 30788
rect 6018 30734 6020 30786
rect 6020 30734 6072 30786
rect 6072 30734 6074 30786
rect 6018 30732 6074 30734
rect 4440 29224 4496 29280
rect 6018 29248 6074 29250
rect 4356 27684 4412 27740
rect 4272 26144 4328 26200
rect 4188 24604 4244 24660
rect 4104 23064 4160 23120
rect 4020 21524 4076 21580
rect 3936 19984 3992 20040
rect 3852 18444 3908 18500
rect 3768 13828 3824 13884
rect 3684 12288 3740 12344
rect 3600 10748 3656 10804
rect 3516 9208 3572 9264
rect 2927 3834 2983 3836
rect 2927 3782 2929 3834
rect 2929 3782 2981 3834
rect 2981 3782 2983 3834
rect 2927 3780 2983 3782
rect 2927 2378 2983 2380
rect 2927 2326 2929 2378
rect 2929 2326 2981 2378
rect 2981 2326 2983 2378
rect 2927 2324 2983 2326
rect 3432 4592 3488 4648
rect 3348 3052 3404 3108
rect 3264 1512 3320 1568
rect 2927 754 2983 756
rect 2927 702 2929 754
rect 2929 702 2981 754
rect 2981 702 2983 754
rect 2927 700 2983 702
rect 3180 -28 3236 28
rect 6018 29196 6020 29248
rect 6020 29196 6072 29248
rect 6072 29196 6074 29248
rect 6018 29194 6074 29196
rect 6018 27710 6074 27712
rect 6018 27658 6020 27710
rect 6020 27658 6072 27710
rect 6072 27658 6074 27710
rect 6018 27656 6074 27658
rect 6018 26172 6074 26174
rect 6018 26120 6020 26172
rect 6020 26120 6072 26172
rect 6072 26120 6074 26172
rect 6018 26118 6074 26120
rect 6018 24634 6074 24636
rect 6018 24582 6020 24634
rect 6020 24582 6072 24634
rect 6072 24582 6074 24634
rect 6018 24580 6074 24582
rect 6018 23096 6074 23098
rect 6018 23044 6020 23096
rect 6020 23044 6072 23096
rect 6072 23044 6074 23096
rect 6018 23042 6074 23044
rect 6018 21558 6074 21560
rect 6018 21506 6020 21558
rect 6020 21506 6072 21558
rect 6072 21506 6074 21558
rect 6018 21504 6074 21506
rect 6018 20020 6074 20022
rect 6018 19968 6020 20020
rect 6020 19968 6072 20020
rect 6072 19968 6074 20020
rect 6018 19966 6074 19968
rect 6018 18482 6074 18484
rect 6018 18430 6020 18482
rect 6020 18430 6072 18482
rect 6072 18430 6074 18482
rect 6018 18428 6074 18430
rect 6018 16944 6074 16946
rect 6018 16892 6020 16944
rect 6020 16892 6072 16944
rect 6072 16892 6074 16944
rect 6018 16890 6074 16892
rect 6018 15406 6074 15408
rect 6018 15354 6020 15406
rect 6020 15354 6072 15406
rect 6072 15354 6074 15406
rect 6018 15352 6074 15354
rect 6018 13868 6074 13870
rect 6018 13816 6020 13868
rect 6020 13816 6072 13868
rect 6072 13816 6074 13868
rect 6018 13814 6074 13816
rect 6018 12330 6074 12332
rect 6018 12278 6020 12330
rect 6020 12278 6072 12330
rect 6072 12278 6074 12330
rect 6018 12276 6074 12278
rect 6018 10792 6074 10794
rect 6018 10740 6020 10792
rect 6020 10740 6072 10792
rect 6072 10740 6074 10792
rect 6018 10738 6074 10740
rect 6018 9254 6074 9256
rect 6018 9202 6020 9254
rect 6020 9202 6072 9254
rect 6072 9202 6074 9254
rect 6018 9200 6074 9202
rect 6018 7716 6074 7718
rect 6018 7664 6020 7716
rect 6020 7664 6072 7716
rect 6072 7664 6074 7716
rect 6018 7662 6074 7664
rect 6018 6178 6074 6180
rect 6018 6126 6020 6178
rect 6020 6126 6072 6178
rect 6072 6126 6074 6178
rect 6018 6124 6074 6126
rect 6018 4640 6074 4642
rect 6018 4588 6020 4640
rect 6020 4588 6072 4640
rect 6072 4588 6074 4640
rect 6018 4586 6074 4588
rect 6018 3102 6074 3104
rect 6018 3050 6020 3102
rect 6020 3050 6072 3102
rect 6072 3050 6074 3102
rect 6018 3048 6074 3050
rect 6018 1564 6074 1566
rect 6018 1512 6020 1564
rect 6020 1512 6072 1564
rect 6072 1512 6074 1564
rect 6018 1510 6074 1512
rect 6018 26 6074 28
rect 6018 -26 6020 26
rect 6020 -26 6072 26
rect 6072 -26 6074 26
rect 6018 -28 6074 -26
<< metal3 >>
rect 5980 49244 6112 49253
rect 5980 49188 6018 49244
rect 6074 49188 6112 49244
rect 5980 49179 6112 49188
rect 5980 47706 6112 47715
rect 5980 47650 6018 47706
rect 6074 47650 6112 47706
rect 5980 47641 6112 47650
rect 5980 46168 6112 46177
rect 5980 46112 6018 46168
rect 6074 46112 6112 46168
rect 5980 46103 6112 46112
rect 5980 44630 6112 44639
rect 5980 44574 6018 44630
rect 6074 44574 6112 44630
rect 5980 44565 6112 44574
rect 5980 43092 6112 43101
rect 5980 43036 6018 43092
rect 6074 43036 6112 43092
rect 5980 43027 6112 43036
rect 5980 41554 6112 41563
rect 5980 41498 6018 41554
rect 6074 41498 6112 41554
rect 5980 41489 6112 41498
rect 5980 40016 6112 40025
rect 5980 39960 6018 40016
rect 6074 39960 6112 40016
rect 5980 39951 6112 39960
rect 5980 38478 6112 38487
rect 5980 38422 6018 38478
rect 6074 38422 6112 38478
rect 5980 38413 6112 38422
rect 5980 36940 6112 36949
rect 5980 36884 6018 36940
rect 6074 36884 6112 36940
rect 5980 36875 6112 36884
rect 5980 35402 6112 35411
rect 5980 35346 6018 35402
rect 6074 35346 6112 35402
rect 5980 35337 6112 35346
rect 5980 33864 6112 33873
rect 5980 33808 6018 33864
rect 6074 33808 6112 33864
rect 5980 33799 6112 33808
rect 5980 32326 6112 32335
rect 5980 32270 6018 32326
rect 6074 32270 6112 32326
rect 5980 32261 6112 32270
rect 960 30755 1092 30829
rect 2000 30755 2132 30829
rect 5980 30788 6112 30797
rect 5980 30732 6018 30788
rect 6074 30732 6112 30788
rect 5980 30723 6112 30732
rect 2889 30092 3021 30097
rect 2889 30036 2927 30092
rect 2983 30036 3021 30092
rect 2889 30031 3021 30036
rect 960 29215 1092 29289
rect 2000 29215 2132 29289
rect 2925 29282 2985 30031
rect 4402 29282 4534 29285
rect 2925 29280 4534 29282
rect 2925 29224 4440 29280
rect 4496 29224 4534 29280
rect 2925 29222 4534 29224
rect 4402 29219 4534 29222
rect 5980 29250 6112 29259
rect 5980 29194 6018 29250
rect 6074 29194 6112 29250
rect 5980 29185 6112 29194
rect 2889 28468 3021 28473
rect 2889 28412 2927 28468
rect 2983 28412 3021 28468
rect 2889 28407 3021 28412
rect 960 27675 1092 27749
rect 2000 27675 2132 27749
rect 2925 27742 2985 28407
rect 4318 27742 4450 27745
rect 2925 27740 4450 27742
rect 2925 27684 4356 27740
rect 4412 27684 4450 27740
rect 2925 27682 4450 27684
rect 4318 27679 4450 27682
rect 5980 27712 6112 27721
rect 5980 27656 6018 27712
rect 6074 27656 6112 27712
rect 5980 27647 6112 27656
rect 2889 27012 3021 27017
rect 2889 26956 2927 27012
rect 2983 26956 3021 27012
rect 2889 26951 3021 26956
rect 960 26135 1092 26209
rect 2000 26135 2132 26209
rect 2925 26202 2985 26951
rect 4234 26202 4366 26205
rect 2925 26200 4366 26202
rect 2925 26144 4272 26200
rect 4328 26144 4366 26200
rect 2925 26142 4366 26144
rect 4234 26139 4366 26142
rect 5980 26174 6112 26183
rect 5980 26118 6018 26174
rect 6074 26118 6112 26174
rect 5980 26109 6112 26118
rect 2889 25388 3021 25393
rect 2889 25332 2927 25388
rect 2983 25332 3021 25388
rect 2889 25327 3021 25332
rect 960 24595 1092 24669
rect 2000 24595 2132 24669
rect 2925 24662 2985 25327
rect 4150 24662 4282 24665
rect 2925 24660 4282 24662
rect 2925 24604 4188 24660
rect 4244 24604 4282 24660
rect 2925 24602 4282 24604
rect 4150 24599 4282 24602
rect 5980 24636 6112 24645
rect 5980 24580 6018 24636
rect 6074 24580 6112 24636
rect 5980 24571 6112 24580
rect 2889 23932 3021 23937
rect 2889 23876 2927 23932
rect 2983 23876 3021 23932
rect 2889 23871 3021 23876
rect 960 23055 1092 23129
rect 2000 23055 2132 23129
rect 2925 23122 2985 23871
rect 4066 23122 4198 23125
rect 2925 23120 4198 23122
rect 2925 23064 4104 23120
rect 4160 23064 4198 23120
rect 2925 23062 4198 23064
rect 4066 23059 4198 23062
rect 5980 23098 6112 23107
rect 5980 23042 6018 23098
rect 6074 23042 6112 23098
rect 5980 23033 6112 23042
rect 2889 22308 3021 22313
rect 2889 22252 2927 22308
rect 2983 22252 3021 22308
rect 2889 22247 3021 22252
rect 960 21515 1092 21589
rect 2000 21515 2132 21589
rect 2925 21582 2985 22247
rect 3982 21582 4114 21585
rect 2925 21580 4114 21582
rect 2925 21524 4020 21580
rect 4076 21524 4114 21580
rect 2925 21522 4114 21524
rect 3982 21519 4114 21522
rect 5980 21560 6112 21569
rect 5980 21504 6018 21560
rect 6074 21504 6112 21560
rect 5980 21495 6112 21504
rect 2889 20852 3021 20857
rect 2889 20796 2927 20852
rect 2983 20796 3021 20852
rect 2889 20791 3021 20796
rect 960 19975 1092 20049
rect 2000 19975 2132 20049
rect 2925 20042 2985 20791
rect 3898 20042 4030 20045
rect 2925 20040 4030 20042
rect 2925 19984 3936 20040
rect 3992 19984 4030 20040
rect 2925 19982 4030 19984
rect 3898 19979 4030 19982
rect 5980 20022 6112 20031
rect 5980 19966 6018 20022
rect 6074 19966 6112 20022
rect 5980 19957 6112 19966
rect 2889 19228 3021 19233
rect 2889 19172 2927 19228
rect 2983 19172 3021 19228
rect 2889 19167 3021 19172
rect 960 18435 1092 18509
rect 2000 18435 2132 18509
rect 2925 18502 2985 19167
rect 3814 18502 3946 18505
rect 2925 18500 3946 18502
rect 2925 18444 3852 18500
rect 3908 18444 3946 18500
rect 2925 18442 3946 18444
rect 3814 18439 3946 18442
rect 5980 18484 6112 18493
rect 5980 18428 6018 18484
rect 6074 18428 6112 18484
rect 5980 18419 6112 18428
rect 5980 16946 6112 16955
rect 5980 16890 6018 16946
rect 6074 16890 6112 16946
rect 5980 16881 6112 16890
rect 1308 15359 1440 15433
rect 2180 15359 2312 15433
rect 5980 15408 6112 15417
rect 5980 15352 6018 15408
rect 6074 15352 6112 15408
rect 5980 15343 6112 15352
rect 2889 14696 3021 14701
rect 2889 14640 2927 14696
rect 2983 14640 3021 14696
rect 2889 14635 3021 14640
rect 1308 13819 1440 13893
rect 2180 13819 2312 13893
rect 2925 13886 2985 14635
rect 3730 13886 3862 13889
rect 2925 13884 3862 13886
rect 2925 13828 3768 13884
rect 3824 13828 3862 13884
rect 2925 13826 3862 13828
rect 3730 13823 3862 13826
rect 5980 13870 6112 13879
rect 5980 13814 6018 13870
rect 6074 13814 6112 13870
rect 5980 13805 6112 13814
rect 2889 13072 3021 13077
rect 2889 13016 2927 13072
rect 2983 13016 3021 13072
rect 2889 13011 3021 13016
rect 1308 12279 1440 12353
rect 2180 12279 2312 12353
rect 2925 12346 2985 13011
rect 3646 12346 3778 12349
rect 2925 12344 3778 12346
rect 2925 12288 3684 12344
rect 3740 12288 3778 12344
rect 2925 12286 3778 12288
rect 3646 12283 3778 12286
rect 5980 12332 6112 12341
rect 5980 12276 6018 12332
rect 6074 12276 6112 12332
rect 5980 12267 6112 12276
rect 2889 11616 3021 11621
rect 2889 11560 2927 11616
rect 2983 11560 3021 11616
rect 2889 11555 3021 11560
rect 1308 10739 1440 10813
rect 2180 10739 2312 10813
rect 2925 10806 2985 11555
rect 3562 10806 3694 10809
rect 2925 10804 3694 10806
rect 2925 10748 3600 10804
rect 3656 10748 3694 10804
rect 2925 10746 3694 10748
rect 3562 10743 3694 10746
rect 5980 10794 6112 10803
rect 5980 10738 6018 10794
rect 6074 10738 6112 10794
rect 5980 10729 6112 10738
rect 2889 9992 3021 9997
rect 2889 9936 2927 9992
rect 2983 9936 3021 9992
rect 2889 9931 3021 9936
rect 1308 9199 1440 9273
rect 2180 9199 2312 9273
rect 2925 9266 2985 9931
rect 3478 9266 3610 9269
rect 2925 9264 3610 9266
rect 2925 9208 3516 9264
rect 3572 9208 3610 9264
rect 2925 9206 3610 9208
rect 3478 9203 3610 9206
rect 5980 9256 6112 9265
rect 5980 9200 6018 9256
rect 6074 9200 6112 9256
rect 5980 9191 6112 9200
rect 5980 7718 6112 7727
rect 5980 7662 6018 7718
rect 6074 7662 6112 7718
rect 5980 7653 6112 7662
rect 1308 6123 1440 6197
rect 2180 6123 2312 6197
rect 5980 6180 6112 6189
rect 5980 6124 6018 6180
rect 6074 6124 6112 6180
rect 5980 6115 6112 6124
rect 2889 5460 3021 5465
rect 2889 5404 2927 5460
rect 2983 5404 3021 5460
rect 2889 5399 3021 5404
rect 1308 4583 1440 4657
rect 2180 4583 2312 4657
rect 2925 4650 2985 5399
rect 3394 4650 3526 4653
rect 2925 4648 3526 4650
rect 2925 4592 3432 4648
rect 3488 4592 3526 4648
rect 2925 4590 3526 4592
rect 3394 4587 3526 4590
rect 5980 4642 6112 4651
rect 5980 4586 6018 4642
rect 6074 4586 6112 4642
rect 5980 4577 6112 4586
rect 2889 3836 3021 3841
rect 2889 3780 2927 3836
rect 2983 3780 3021 3836
rect 2889 3775 3021 3780
rect 1308 3043 1440 3117
rect 2180 3043 2312 3117
rect 2925 3110 2985 3775
rect 3310 3110 3442 3113
rect 2925 3108 3442 3110
rect 2925 3052 3348 3108
rect 3404 3052 3442 3108
rect 2925 3050 3442 3052
rect 3310 3047 3442 3050
rect 5980 3104 6112 3113
rect 5980 3048 6018 3104
rect 6074 3048 6112 3104
rect 5980 3039 6112 3048
rect 2889 2380 3021 2385
rect 2889 2324 2927 2380
rect 2983 2324 3021 2380
rect 2889 2319 3021 2324
rect 1308 1503 1440 1577
rect 2180 1503 2312 1577
rect 2925 1570 2985 2319
rect 3226 1570 3358 1573
rect 2925 1568 3358 1570
rect 2925 1512 3264 1568
rect 3320 1512 3358 1568
rect 2925 1510 3358 1512
rect 3226 1507 3358 1510
rect 5980 1566 6112 1575
rect 5980 1510 6018 1566
rect 6074 1510 6112 1566
rect 5980 1501 6112 1510
rect 2889 756 3021 761
rect 2889 700 2927 756
rect 2983 700 3021 756
rect 2889 695 3021 700
rect 1308 -37 1440 37
rect 2180 -37 2312 37
rect 2925 30 2985 695
rect 3142 30 3274 33
rect 2925 28 3274 30
rect 2925 -28 3180 28
rect 3236 -28 3274 28
rect 2925 -30 3274 -28
rect 3142 -33 3274 -30
rect 5980 28 6112 37
rect 5980 -28 6018 28
rect 6074 -28 6112 28
rect 5980 -37 6112 -28
use contact_18  contact_18_0
timestamp 1644951705
transform 1 0 5980 0 1 49179
box 0 0 1 1
use contact_17  contact_17_0
timestamp 1644951705
transform 1 0 6014 0 1 49184
box 0 0 1 1
use contact_18  contact_18_1
timestamp 1644951705
transform 1 0 5980 0 1 47641
box 0 0 1 1
use contact_17  contact_17_1
timestamp 1644951705
transform 1 0 6014 0 1 47646
box 0 0 1 1
use contact_18  contact_18_2
timestamp 1644951705
transform 1 0 5980 0 1 46103
box 0 0 1 1
use contact_17  contact_17_2
timestamp 1644951705
transform 1 0 6014 0 1 46108
box 0 0 1 1
use contact_18  contact_18_3
timestamp 1644951705
transform 1 0 5980 0 1 47641
box 0 0 1 1
use contact_17  contact_17_3
timestamp 1644951705
transform 1 0 6014 0 1 47646
box 0 0 1 1
use contact_18  contact_18_4
timestamp 1644951705
transform 1 0 5980 0 1 46103
box 0 0 1 1
use contact_17  contact_17_4
timestamp 1644951705
transform 1 0 6014 0 1 46108
box 0 0 1 1
use contact_18  contact_18_5
timestamp 1644951705
transform 1 0 5980 0 1 44565
box 0 0 1 1
use contact_17  contact_17_5
timestamp 1644951705
transform 1 0 6014 0 1 44570
box 0 0 1 1
use contact_18  contact_18_6
timestamp 1644951705
transform 1 0 5980 0 1 43027
box 0 0 1 1
use contact_17  contact_17_6
timestamp 1644951705
transform 1 0 6014 0 1 43032
box 0 0 1 1
use contact_18  contact_18_7
timestamp 1644951705
transform 1 0 5980 0 1 44565
box 0 0 1 1
use contact_17  contact_17_7
timestamp 1644951705
transform 1 0 6014 0 1 44570
box 0 0 1 1
use contact_18  contact_18_8
timestamp 1644951705
transform 1 0 5980 0 1 43027
box 0 0 1 1
use contact_17  contact_17_8
timestamp 1644951705
transform 1 0 6014 0 1 43032
box 0 0 1 1
use contact_18  contact_18_9
timestamp 1644951705
transform 1 0 5980 0 1 41489
box 0 0 1 1
use contact_17  contact_17_9
timestamp 1644951705
transform 1 0 6014 0 1 41494
box 0 0 1 1
use contact_18  contact_18_10
timestamp 1644951705
transform 1 0 5980 0 1 39951
box 0 0 1 1
use contact_17  contact_17_10
timestamp 1644951705
transform 1 0 6014 0 1 39956
box 0 0 1 1
use contact_18  contact_18_11
timestamp 1644951705
transform 1 0 5980 0 1 41489
box 0 0 1 1
use contact_17  contact_17_11
timestamp 1644951705
transform 1 0 6014 0 1 41494
box 0 0 1 1
use contact_18  contact_18_12
timestamp 1644951705
transform 1 0 5980 0 1 39951
box 0 0 1 1
use contact_17  contact_17_12
timestamp 1644951705
transform 1 0 6014 0 1 39956
box 0 0 1 1
use contact_18  contact_18_13
timestamp 1644951705
transform 1 0 5980 0 1 38413
box 0 0 1 1
use contact_17  contact_17_13
timestamp 1644951705
transform 1 0 6014 0 1 38418
box 0 0 1 1
use contact_18  contact_18_14
timestamp 1644951705
transform 1 0 5980 0 1 36875
box 0 0 1 1
use contact_17  contact_17_14
timestamp 1644951705
transform 1 0 6014 0 1 36880
box 0 0 1 1
use contact_18  contact_18_15
timestamp 1644951705
transform 1 0 5980 0 1 38413
box 0 0 1 1
use contact_17  contact_17_15
timestamp 1644951705
transform 1 0 6014 0 1 38418
box 0 0 1 1
use contact_18  contact_18_16
timestamp 1644951705
transform 1 0 5980 0 1 36875
box 0 0 1 1
use contact_17  contact_17_16
timestamp 1644951705
transform 1 0 6014 0 1 36880
box 0 0 1 1
use contact_18  contact_18_17
timestamp 1644951705
transform 1 0 5980 0 1 35337
box 0 0 1 1
use contact_17  contact_17_17
timestamp 1644951705
transform 1 0 6014 0 1 35342
box 0 0 1 1
use contact_18  contact_18_18
timestamp 1644951705
transform 1 0 5980 0 1 33799
box 0 0 1 1
use contact_17  contact_17_18
timestamp 1644951705
transform 1 0 6014 0 1 33804
box 0 0 1 1
use contact_18  contact_18_19
timestamp 1644951705
transform 1 0 5980 0 1 35337
box 0 0 1 1
use contact_17  contact_17_19
timestamp 1644951705
transform 1 0 6014 0 1 35342
box 0 0 1 1
use contact_18  contact_18_20
timestamp 1644951705
transform 1 0 5980 0 1 33799
box 0 0 1 1
use contact_17  contact_17_20
timestamp 1644951705
transform 1 0 6014 0 1 33804
box 0 0 1 1
use contact_18  contact_18_21
timestamp 1644951705
transform 1 0 5980 0 1 32261
box 0 0 1 1
use contact_17  contact_17_21
timestamp 1644951705
transform 1 0 6014 0 1 32266
box 0 0 1 1
use contact_18  contact_18_22
timestamp 1644951705
transform 1 0 5980 0 1 30723
box 0 0 1 1
use contact_17  contact_17_22
timestamp 1644951705
transform 1 0 6014 0 1 30728
box 0 0 1 1
use contact_18  contact_18_23
timestamp 1644951705
transform 1 0 5980 0 1 32261
box 0 0 1 1
use contact_17  contact_17_23
timestamp 1644951705
transform 1 0 6014 0 1 32266
box 0 0 1 1
use contact_18  contact_18_24
timestamp 1644951705
transform 1 0 5980 0 1 30723
box 0 0 1 1
use contact_17  contact_17_24
timestamp 1644951705
transform 1 0 6014 0 1 30728
box 0 0 1 1
use contact_18  contact_18_25
timestamp 1644951705
transform 1 0 5980 0 1 29185
box 0 0 1 1
use contact_17  contact_17_25
timestamp 1644951705
transform 1 0 6014 0 1 29190
box 0 0 1 1
use contact_18  contact_18_26
timestamp 1644951705
transform 1 0 5980 0 1 27647
box 0 0 1 1
use contact_17  contact_17_26
timestamp 1644951705
transform 1 0 6014 0 1 27652
box 0 0 1 1
use contact_18  contact_18_27
timestamp 1644951705
transform 1 0 5980 0 1 29185
box 0 0 1 1
use contact_17  contact_17_27
timestamp 1644951705
transform 1 0 6014 0 1 29190
box 0 0 1 1
use contact_18  contact_18_28
timestamp 1644951705
transform 1 0 5980 0 1 27647
box 0 0 1 1
use contact_17  contact_17_28
timestamp 1644951705
transform 1 0 6014 0 1 27652
box 0 0 1 1
use contact_18  contact_18_29
timestamp 1644951705
transform 1 0 5980 0 1 26109
box 0 0 1 1
use contact_17  contact_17_29
timestamp 1644951705
transform 1 0 6014 0 1 26114
box 0 0 1 1
use contact_18  contact_18_30
timestamp 1644951705
transform 1 0 5980 0 1 24571
box 0 0 1 1
use contact_17  contact_17_30
timestamp 1644951705
transform 1 0 6014 0 1 24576
box 0 0 1 1
use contact_18  contact_18_31
timestamp 1644951705
transform 1 0 5980 0 1 26109
box 0 0 1 1
use contact_17  contact_17_31
timestamp 1644951705
transform 1 0 6014 0 1 26114
box 0 0 1 1
use contact_18  contact_18_32
timestamp 1644951705
transform 1 0 5980 0 1 24571
box 0 0 1 1
use contact_17  contact_17_32
timestamp 1644951705
transform 1 0 6014 0 1 24576
box 0 0 1 1
use contact_18  contact_18_33
timestamp 1644951705
transform 1 0 5980 0 1 23033
box 0 0 1 1
use contact_17  contact_17_33
timestamp 1644951705
transform 1 0 6014 0 1 23038
box 0 0 1 1
use contact_18  contact_18_34
timestamp 1644951705
transform 1 0 5980 0 1 21495
box 0 0 1 1
use contact_17  contact_17_34
timestamp 1644951705
transform 1 0 6014 0 1 21500
box 0 0 1 1
use contact_18  contact_18_35
timestamp 1644951705
transform 1 0 5980 0 1 23033
box 0 0 1 1
use contact_17  contact_17_35
timestamp 1644951705
transform 1 0 6014 0 1 23038
box 0 0 1 1
use contact_18  contact_18_36
timestamp 1644951705
transform 1 0 5980 0 1 21495
box 0 0 1 1
use contact_17  contact_17_36
timestamp 1644951705
transform 1 0 6014 0 1 21500
box 0 0 1 1
use contact_18  contact_18_37
timestamp 1644951705
transform 1 0 5980 0 1 19957
box 0 0 1 1
use contact_17  contact_17_37
timestamp 1644951705
transform 1 0 6014 0 1 19962
box 0 0 1 1
use contact_18  contact_18_38
timestamp 1644951705
transform 1 0 5980 0 1 18419
box 0 0 1 1
use contact_17  contact_17_38
timestamp 1644951705
transform 1 0 6014 0 1 18424
box 0 0 1 1
use contact_18  contact_18_39
timestamp 1644951705
transform 1 0 5980 0 1 19957
box 0 0 1 1
use contact_17  contact_17_39
timestamp 1644951705
transform 1 0 6014 0 1 19962
box 0 0 1 1
use contact_18  contact_18_40
timestamp 1644951705
transform 1 0 5980 0 1 18419
box 0 0 1 1
use contact_17  contact_17_40
timestamp 1644951705
transform 1 0 6014 0 1 18424
box 0 0 1 1
use contact_18  contact_18_41
timestamp 1644951705
transform 1 0 5980 0 1 16881
box 0 0 1 1
use contact_17  contact_17_41
timestamp 1644951705
transform 1 0 6014 0 1 16886
box 0 0 1 1
use contact_18  contact_18_42
timestamp 1644951705
transform 1 0 5980 0 1 15343
box 0 0 1 1
use contact_17  contact_17_42
timestamp 1644951705
transform 1 0 6014 0 1 15348
box 0 0 1 1
use contact_18  contact_18_43
timestamp 1644951705
transform 1 0 5980 0 1 16881
box 0 0 1 1
use contact_17  contact_17_43
timestamp 1644951705
transform 1 0 6014 0 1 16886
box 0 0 1 1
use contact_18  contact_18_44
timestamp 1644951705
transform 1 0 5980 0 1 15343
box 0 0 1 1
use contact_17  contact_17_44
timestamp 1644951705
transform 1 0 6014 0 1 15348
box 0 0 1 1
use contact_18  contact_18_45
timestamp 1644951705
transform 1 0 5980 0 1 13805
box 0 0 1 1
use contact_17  contact_17_45
timestamp 1644951705
transform 1 0 6014 0 1 13810
box 0 0 1 1
use contact_18  contact_18_46
timestamp 1644951705
transform 1 0 5980 0 1 12267
box 0 0 1 1
use contact_17  contact_17_46
timestamp 1644951705
transform 1 0 6014 0 1 12272
box 0 0 1 1
use contact_18  contact_18_47
timestamp 1644951705
transform 1 0 5980 0 1 13805
box 0 0 1 1
use contact_17  contact_17_47
timestamp 1644951705
transform 1 0 6014 0 1 13810
box 0 0 1 1
use contact_18  contact_18_48
timestamp 1644951705
transform 1 0 5980 0 1 12267
box 0 0 1 1
use contact_17  contact_17_48
timestamp 1644951705
transform 1 0 6014 0 1 12272
box 0 0 1 1
use contact_18  contact_18_49
timestamp 1644951705
transform 1 0 5980 0 1 10729
box 0 0 1 1
use contact_17  contact_17_49
timestamp 1644951705
transform 1 0 6014 0 1 10734
box 0 0 1 1
use contact_18  contact_18_50
timestamp 1644951705
transform 1 0 5980 0 1 9191
box 0 0 1 1
use contact_17  contact_17_50
timestamp 1644951705
transform 1 0 6014 0 1 9196
box 0 0 1 1
use contact_18  contact_18_51
timestamp 1644951705
transform 1 0 5980 0 1 10729
box 0 0 1 1
use contact_17  contact_17_51
timestamp 1644951705
transform 1 0 6014 0 1 10734
box 0 0 1 1
use contact_18  contact_18_52
timestamp 1644951705
transform 1 0 5980 0 1 9191
box 0 0 1 1
use contact_17  contact_17_52
timestamp 1644951705
transform 1 0 6014 0 1 9196
box 0 0 1 1
use contact_18  contact_18_53
timestamp 1644951705
transform 1 0 5980 0 1 7653
box 0 0 1 1
use contact_17  contact_17_53
timestamp 1644951705
transform 1 0 6014 0 1 7658
box 0 0 1 1
use contact_18  contact_18_54
timestamp 1644951705
transform 1 0 5980 0 1 6115
box 0 0 1 1
use contact_17  contact_17_54
timestamp 1644951705
transform 1 0 6014 0 1 6120
box 0 0 1 1
use contact_18  contact_18_55
timestamp 1644951705
transform 1 0 5980 0 1 7653
box 0 0 1 1
use contact_17  contact_17_55
timestamp 1644951705
transform 1 0 6014 0 1 7658
box 0 0 1 1
use contact_18  contact_18_56
timestamp 1644951705
transform 1 0 5980 0 1 6115
box 0 0 1 1
use contact_17  contact_17_56
timestamp 1644951705
transform 1 0 6014 0 1 6120
box 0 0 1 1
use contact_18  contact_18_57
timestamp 1644951705
transform 1 0 5980 0 1 4577
box 0 0 1 1
use contact_17  contact_17_57
timestamp 1644951705
transform 1 0 6014 0 1 4582
box 0 0 1 1
use contact_18  contact_18_58
timestamp 1644951705
transform 1 0 5980 0 1 3039
box 0 0 1 1
use contact_17  contact_17_58
timestamp 1644951705
transform 1 0 6014 0 1 3044
box 0 0 1 1
use contact_18  contact_18_59
timestamp 1644951705
transform 1 0 5980 0 1 4577
box 0 0 1 1
use contact_17  contact_17_59
timestamp 1644951705
transform 1 0 6014 0 1 4582
box 0 0 1 1
use contact_18  contact_18_60
timestamp 1644951705
transform 1 0 5980 0 1 3039
box 0 0 1 1
use contact_17  contact_17_60
timestamp 1644951705
transform 1 0 6014 0 1 3044
box 0 0 1 1
use contact_18  contact_18_61
timestamp 1644951705
transform 1 0 5980 0 1 1501
box 0 0 1 1
use contact_17  contact_17_61
timestamp 1644951705
transform 1 0 6014 0 1 1506
box 0 0 1 1
use contact_18  contact_18_62
timestamp 1644951705
transform 1 0 5980 0 1 -37
box 0 0 1 1
use contact_17  contact_17_62
timestamp 1644951705
transform 1 0 6014 0 1 -32
box 0 0 1 1
use contact_18  contact_18_63
timestamp 1644951705
transform 1 0 5980 0 1 1501
box 0 0 1 1
use contact_17  contact_17_63
timestamp 1644951705
transform 1 0 6014 0 1 1506
box 0 0 1 1
use contact_20  contact_20_0
timestamp 1644951705
transform 1 0 4402 0 1 29215
box 0 0 1 1
use contact_18  contact_18_64
timestamp 1644951705
transform 1 0 2889 0 1 30027
box 0 0 1 1
use contact_17  contact_17_64
timestamp 1644951705
transform 1 0 2923 0 1 30032
box 0 0 1 1
use contact_13  contact_13_0
timestamp 1644951705
transform 1 0 2926 0 1 30041
box 0 0 1 1
use contact_20  contact_20_1
timestamp 1644951705
transform 1 0 4318 0 1 27675
box 0 0 1 1
use contact_18  contact_18_65
timestamp 1644951705
transform 1 0 2889 0 1 28403
box 0 0 1 1
use contact_17  contact_17_65
timestamp 1644951705
transform 1 0 2923 0 1 28408
box 0 0 1 1
use contact_13  contact_13_1
timestamp 1644951705
transform 1 0 2926 0 1 28417
box 0 0 1 1
use contact_20  contact_20_2
timestamp 1644951705
transform 1 0 4234 0 1 26135
box 0 0 1 1
use contact_18  contact_18_66
timestamp 1644951705
transform 1 0 2889 0 1 26947
box 0 0 1 1
use contact_17  contact_17_66
timestamp 1644951705
transform 1 0 2923 0 1 26952
box 0 0 1 1
use contact_13  contact_13_2
timestamp 1644951705
transform 1 0 2926 0 1 26961
box 0 0 1 1
use contact_20  contact_20_3
timestamp 1644951705
transform 1 0 4150 0 1 24595
box 0 0 1 1
use contact_18  contact_18_67
timestamp 1644951705
transform 1 0 2889 0 1 25323
box 0 0 1 1
use contact_17  contact_17_67
timestamp 1644951705
transform 1 0 2923 0 1 25328
box 0 0 1 1
use contact_13  contact_13_3
timestamp 1644951705
transform 1 0 2926 0 1 25337
box 0 0 1 1
use contact_20  contact_20_4
timestamp 1644951705
transform 1 0 4066 0 1 23055
box 0 0 1 1
use contact_18  contact_18_68
timestamp 1644951705
transform 1 0 2889 0 1 23867
box 0 0 1 1
use contact_17  contact_17_68
timestamp 1644951705
transform 1 0 2923 0 1 23872
box 0 0 1 1
use contact_13  contact_13_4
timestamp 1644951705
transform 1 0 2926 0 1 23881
box 0 0 1 1
use contact_20  contact_20_5
timestamp 1644951705
transform 1 0 3982 0 1 21515
box 0 0 1 1
use contact_18  contact_18_69
timestamp 1644951705
transform 1 0 2889 0 1 22243
box 0 0 1 1
use contact_17  contact_17_69
timestamp 1644951705
transform 1 0 2923 0 1 22248
box 0 0 1 1
use contact_13  contact_13_5
timestamp 1644951705
transform 1 0 2926 0 1 22257
box 0 0 1 1
use contact_20  contact_20_6
timestamp 1644951705
transform 1 0 3898 0 1 19975
box 0 0 1 1
use contact_18  contact_18_70
timestamp 1644951705
transform 1 0 2889 0 1 20787
box 0 0 1 1
use contact_17  contact_17_70
timestamp 1644951705
transform 1 0 2923 0 1 20792
box 0 0 1 1
use contact_13  contact_13_6
timestamp 1644951705
transform 1 0 2926 0 1 20801
box 0 0 1 1
use contact_20  contact_20_7
timestamp 1644951705
transform 1 0 3814 0 1 18435
box 0 0 1 1
use contact_18  contact_18_71
timestamp 1644951705
transform 1 0 2889 0 1 19163
box 0 0 1 1
use contact_17  contact_17_71
timestamp 1644951705
transform 1 0 2923 0 1 19168
box 0 0 1 1
use contact_13  contact_13_7
timestamp 1644951705
transform 1 0 2926 0 1 19177
box 0 0 1 1
use contact_20  contact_20_8
timestamp 1644951705
transform 1 0 3730 0 1 13819
box 0 0 1 1
use contact_18  contact_18_72
timestamp 1644951705
transform 1 0 2889 0 1 14631
box 0 0 1 1
use contact_17  contact_17_72
timestamp 1644951705
transform 1 0 2923 0 1 14636
box 0 0 1 1
use contact_13  contact_13_8
timestamp 1644951705
transform 1 0 2926 0 1 14645
box 0 0 1 1
use contact_20  contact_20_9
timestamp 1644951705
transform 1 0 3646 0 1 12279
box 0 0 1 1
use contact_18  contact_18_73
timestamp 1644951705
transform 1 0 2889 0 1 13007
box 0 0 1 1
use contact_17  contact_17_73
timestamp 1644951705
transform 1 0 2923 0 1 13012
box 0 0 1 1
use contact_13  contact_13_9
timestamp 1644951705
transform 1 0 2926 0 1 13021
box 0 0 1 1
use contact_20  contact_20_10
timestamp 1644951705
transform 1 0 3562 0 1 10739
box 0 0 1 1
use contact_18  contact_18_74
timestamp 1644951705
transform 1 0 2889 0 1 11551
box 0 0 1 1
use contact_17  contact_17_74
timestamp 1644951705
transform 1 0 2923 0 1 11556
box 0 0 1 1
use contact_13  contact_13_10
timestamp 1644951705
transform 1 0 2926 0 1 11565
box 0 0 1 1
use contact_20  contact_20_11
timestamp 1644951705
transform 1 0 3478 0 1 9199
box 0 0 1 1
use contact_18  contact_18_75
timestamp 1644951705
transform 1 0 2889 0 1 9927
box 0 0 1 1
use contact_17  contact_17_75
timestamp 1644951705
transform 1 0 2923 0 1 9932
box 0 0 1 1
use contact_13  contact_13_11
timestamp 1644951705
transform 1 0 2926 0 1 9941
box 0 0 1 1
use contact_20  contact_20_12
timestamp 1644951705
transform 1 0 3394 0 1 4583
box 0 0 1 1
use contact_18  contact_18_76
timestamp 1644951705
transform 1 0 2889 0 1 5395
box 0 0 1 1
use contact_17  contact_17_76
timestamp 1644951705
transform 1 0 2923 0 1 5400
box 0 0 1 1
use contact_13  contact_13_12
timestamp 1644951705
transform 1 0 2926 0 1 5409
box 0 0 1 1
use contact_20  contact_20_13
timestamp 1644951705
transform 1 0 3310 0 1 3043
box 0 0 1 1
use contact_18  contact_18_77
timestamp 1644951705
transform 1 0 2889 0 1 3771
box 0 0 1 1
use contact_17  contact_17_77
timestamp 1644951705
transform 1 0 2923 0 1 3776
box 0 0 1 1
use contact_13  contact_13_13
timestamp 1644951705
transform 1 0 2926 0 1 3785
box 0 0 1 1
use contact_20  contact_20_14
timestamp 1644951705
transform 1 0 3226 0 1 1503
box 0 0 1 1
use contact_18  contact_18_78
timestamp 1644951705
transform 1 0 2889 0 1 2315
box 0 0 1 1
use contact_17  contact_17_78
timestamp 1644951705
transform 1 0 2923 0 1 2320
box 0 0 1 1
use contact_13  contact_13_14
timestamp 1644951705
transform 1 0 2926 0 1 2329
box 0 0 1 1
use contact_20  contact_20_15
timestamp 1644951705
transform 1 0 3142 0 1 -37
box 0 0 1 1
use contact_18  contact_18_79
timestamp 1644951705
transform 1 0 2889 0 1 691
box 0 0 1 1
use contact_17  contact_17_79
timestamp 1644951705
transform 1 0 2923 0 1 696
box 0 0 1 1
use contact_13  contact_13_15
timestamp 1644951705
transform 1 0 2926 0 1 705
box 0 0 1 1
use contact_14  contact_14_0
timestamp 1644951705
transform 1 0 4268 0 1 48802
box 0 0 1 1
use contact_14  contact_14_1
timestamp 1644951705
transform 1 0 3764 0 1 48716
box 0 0 1 1
use contact_14  contact_14_2
timestamp 1644951705
transform 1 0 3344 0 1 48630
box 0 0 1 1
use contact_14  contact_14_3
timestamp 1644951705
transform 1 0 4268 0 1 48544
box 0 0 1 1
use contact_14  contact_14_4
timestamp 1644951705
transform 1 0 3764 0 1 48458
box 0 0 1 1
use contact_14  contact_14_5
timestamp 1644951705
transform 1 0 3260 0 1 48372
box 0 0 1 1
use contact_14  contact_14_6
timestamp 1644951705
transform 1 0 4268 0 1 48286
box 0 0 1 1
use contact_14  contact_14_7
timestamp 1644951705
transform 1 0 3764 0 1 48200
box 0 0 1 1
use contact_14  contact_14_8
timestamp 1644951705
transform 1 0 3176 0 1 48114
box 0 0 1 1
use contact_14  contact_14_9
timestamp 1644951705
transform 1 0 4268 0 1 46490
box 0 0 1 1
use contact_14  contact_14_10
timestamp 1644951705
transform 1 0 3680 0 1 46576
box 0 0 1 1
use contact_14  contact_14_11
timestamp 1644951705
transform 1 0 3428 0 1 46662
box 0 0 1 1
use contact_14  contact_14_12
timestamp 1644951705
transform 1 0 4268 0 1 46748
box 0 0 1 1
use contact_14  contact_14_13
timestamp 1644951705
transform 1 0 3680 0 1 46834
box 0 0 1 1
use contact_14  contact_14_14
timestamp 1644951705
transform 1 0 3344 0 1 46920
box 0 0 1 1
use contact_14  contact_14_15
timestamp 1644951705
transform 1 0 4268 0 1 47006
box 0 0 1 1
use contact_14  contact_14_16
timestamp 1644951705
transform 1 0 3680 0 1 47092
box 0 0 1 1
use contact_14  contact_14_17
timestamp 1644951705
transform 1 0 3260 0 1 47178
box 0 0 1 1
use contact_14  contact_14_18
timestamp 1644951705
transform 1 0 4268 0 1 45726
box 0 0 1 1
use contact_14  contact_14_19
timestamp 1644951705
transform 1 0 3680 0 1 45640
box 0 0 1 1
use contact_14  contact_14_20
timestamp 1644951705
transform 1 0 3176 0 1 45554
box 0 0 1 1
use contact_14  contact_14_21
timestamp 1644951705
transform 1 0 4268 0 1 45468
box 0 0 1 1
use contact_14  contact_14_22
timestamp 1644951705
transform 1 0 3596 0 1 45382
box 0 0 1 1
use contact_14  contact_14_23
timestamp 1644951705
transform 1 0 3428 0 1 45296
box 0 0 1 1
use contact_14  contact_14_24
timestamp 1644951705
transform 1 0 4268 0 1 45210
box 0 0 1 1
use contact_14  contact_14_25
timestamp 1644951705
transform 1 0 3596 0 1 45124
box 0 0 1 1
use contact_14  contact_14_26
timestamp 1644951705
transform 1 0 3344 0 1 45038
box 0 0 1 1
use contact_14  contact_14_27
timestamp 1644951705
transform 1 0 4268 0 1 43414
box 0 0 1 1
use contact_14  contact_14_28
timestamp 1644951705
transform 1 0 3596 0 1 43500
box 0 0 1 1
use contact_14  contact_14_29
timestamp 1644951705
transform 1 0 3260 0 1 43586
box 0 0 1 1
use contact_14  contact_14_30
timestamp 1644951705
transform 1 0 4268 0 1 43672
box 0 0 1 1
use contact_14  contact_14_31
timestamp 1644951705
transform 1 0 3596 0 1 43758
box 0 0 1 1
use contact_14  contact_14_32
timestamp 1644951705
transform 1 0 3176 0 1 43844
box 0 0 1 1
use contact_14  contact_14_33
timestamp 1644951705
transform 1 0 4268 0 1 43930
box 0 0 1 1
use contact_14  contact_14_34
timestamp 1644951705
transform 1 0 3512 0 1 44016
box 0 0 1 1
use contact_14  contact_14_35
timestamp 1644951705
transform 1 0 3428 0 1 44102
box 0 0 1 1
use contact_14  contact_14_36
timestamp 1644951705
transform 1 0 4268 0 1 42650
box 0 0 1 1
use contact_14  contact_14_37
timestamp 1644951705
transform 1 0 3512 0 1 42564
box 0 0 1 1
use contact_14  contact_14_38
timestamp 1644951705
transform 1 0 3344 0 1 42478
box 0 0 1 1
use contact_14  contact_14_39
timestamp 1644951705
transform 1 0 4268 0 1 42392
box 0 0 1 1
use contact_14  contact_14_40
timestamp 1644951705
transform 1 0 3512 0 1 42306
box 0 0 1 1
use contact_14  contact_14_41
timestamp 1644951705
transform 1 0 3260 0 1 42220
box 0 0 1 1
use contact_14  contact_14_42
timestamp 1644951705
transform 1 0 4268 0 1 42134
box 0 0 1 1
use contact_14  contact_14_43
timestamp 1644951705
transform 1 0 3512 0 1 42048
box 0 0 1 1
use contact_14  contact_14_44
timestamp 1644951705
transform 1 0 3176 0 1 41962
box 0 0 1 1
use contact_14  contact_14_45
timestamp 1644951705
transform 1 0 4184 0 1 40338
box 0 0 1 1
use contact_14  contact_14_46
timestamp 1644951705
transform 1 0 3764 0 1 40424
box 0 0 1 1
use contact_14  contact_14_47
timestamp 1644951705
transform 1 0 3428 0 1 40510
box 0 0 1 1
use contact_14  contact_14_48
timestamp 1644951705
transform 1 0 4184 0 1 40596
box 0 0 1 1
use contact_14  contact_14_49
timestamp 1644951705
transform 1 0 3764 0 1 40682
box 0 0 1 1
use contact_14  contact_14_50
timestamp 1644951705
transform 1 0 3344 0 1 40768
box 0 0 1 1
use contact_14  contact_14_51
timestamp 1644951705
transform 1 0 4184 0 1 40854
box 0 0 1 1
use contact_14  contact_14_52
timestamp 1644951705
transform 1 0 3764 0 1 40940
box 0 0 1 1
use contact_14  contact_14_53
timestamp 1644951705
transform 1 0 3260 0 1 41026
box 0 0 1 1
use contact_14  contact_14_54
timestamp 1644951705
transform 1 0 4184 0 1 39574
box 0 0 1 1
use contact_14  contact_14_55
timestamp 1644951705
transform 1 0 3764 0 1 39488
box 0 0 1 1
use contact_14  contact_14_56
timestamp 1644951705
transform 1 0 3176 0 1 39402
box 0 0 1 1
use contact_14  contact_14_57
timestamp 1644951705
transform 1 0 4184 0 1 39316
box 0 0 1 1
use contact_14  contact_14_58
timestamp 1644951705
transform 1 0 3680 0 1 39230
box 0 0 1 1
use contact_14  contact_14_59
timestamp 1644951705
transform 1 0 3428 0 1 39144
box 0 0 1 1
use contact_14  contact_14_60
timestamp 1644951705
transform 1 0 4184 0 1 39058
box 0 0 1 1
use contact_14  contact_14_61
timestamp 1644951705
transform 1 0 3680 0 1 38972
box 0 0 1 1
use contact_14  contact_14_62
timestamp 1644951705
transform 1 0 3344 0 1 38886
box 0 0 1 1
use contact_14  contact_14_63
timestamp 1644951705
transform 1 0 4184 0 1 37262
box 0 0 1 1
use contact_14  contact_14_64
timestamp 1644951705
transform 1 0 3680 0 1 37348
box 0 0 1 1
use contact_14  contact_14_65
timestamp 1644951705
transform 1 0 3260 0 1 37434
box 0 0 1 1
use contact_14  contact_14_66
timestamp 1644951705
transform 1 0 4184 0 1 37520
box 0 0 1 1
use contact_14  contact_14_67
timestamp 1644951705
transform 1 0 3680 0 1 37606
box 0 0 1 1
use contact_14  contact_14_68
timestamp 1644951705
transform 1 0 3176 0 1 37692
box 0 0 1 1
use contact_14  contact_14_69
timestamp 1644951705
transform 1 0 4184 0 1 37778
box 0 0 1 1
use contact_14  contact_14_70
timestamp 1644951705
transform 1 0 3596 0 1 37864
box 0 0 1 1
use contact_14  contact_14_71
timestamp 1644951705
transform 1 0 3428 0 1 37950
box 0 0 1 1
use contact_14  contact_14_72
timestamp 1644951705
transform 1 0 4184 0 1 36498
box 0 0 1 1
use contact_14  contact_14_73
timestamp 1644951705
transform 1 0 3596 0 1 36412
box 0 0 1 1
use contact_14  contact_14_74
timestamp 1644951705
transform 1 0 3344 0 1 36326
box 0 0 1 1
use contact_14  contact_14_75
timestamp 1644951705
transform 1 0 4184 0 1 36240
box 0 0 1 1
use contact_14  contact_14_76
timestamp 1644951705
transform 1 0 3596 0 1 36154
box 0 0 1 1
use contact_14  contact_14_77
timestamp 1644951705
transform 1 0 3260 0 1 36068
box 0 0 1 1
use contact_14  contact_14_78
timestamp 1644951705
transform 1 0 4184 0 1 35982
box 0 0 1 1
use contact_14  contact_14_79
timestamp 1644951705
transform 1 0 3596 0 1 35896
box 0 0 1 1
use contact_14  contact_14_80
timestamp 1644951705
transform 1 0 3176 0 1 35810
box 0 0 1 1
use contact_14  contact_14_81
timestamp 1644951705
transform 1 0 4184 0 1 34186
box 0 0 1 1
use contact_14  contact_14_82
timestamp 1644951705
transform 1 0 3512 0 1 34272
box 0 0 1 1
use contact_14  contact_14_83
timestamp 1644951705
transform 1 0 3428 0 1 34358
box 0 0 1 1
use contact_14  contact_14_84
timestamp 1644951705
transform 1 0 4184 0 1 34444
box 0 0 1 1
use contact_14  contact_14_85
timestamp 1644951705
transform 1 0 3512 0 1 34530
box 0 0 1 1
use contact_14  contact_14_86
timestamp 1644951705
transform 1 0 3344 0 1 34616
box 0 0 1 1
use contact_14  contact_14_87
timestamp 1644951705
transform 1 0 4184 0 1 34702
box 0 0 1 1
use contact_14  contact_14_88
timestamp 1644951705
transform 1 0 3512 0 1 34788
box 0 0 1 1
use contact_14  contact_14_89
timestamp 1644951705
transform 1 0 3260 0 1 34874
box 0 0 1 1
use contact_14  contact_14_90
timestamp 1644951705
transform 1 0 4184 0 1 33422
box 0 0 1 1
use contact_14  contact_14_91
timestamp 1644951705
transform 1 0 3512 0 1 33336
box 0 0 1 1
use contact_14  contact_14_92
timestamp 1644951705
transform 1 0 3176 0 1 33250
box 0 0 1 1
use contact_14  contact_14_93
timestamp 1644951705
transform 1 0 4100 0 1 33164
box 0 0 1 1
use contact_14  contact_14_94
timestamp 1644951705
transform 1 0 3764 0 1 33078
box 0 0 1 1
use contact_14  contact_14_95
timestamp 1644951705
transform 1 0 3428 0 1 32992
box 0 0 1 1
use contact_14  contact_14_96
timestamp 1644951705
transform 1 0 4100 0 1 32906
box 0 0 1 1
use contact_14  contact_14_97
timestamp 1644951705
transform 1 0 3764 0 1 32820
box 0 0 1 1
use contact_14  contact_14_98
timestamp 1644951705
transform 1 0 3344 0 1 32734
box 0 0 1 1
use contact_14  contact_14_99
timestamp 1644951705
transform 1 0 4100 0 1 31110
box 0 0 1 1
use contact_14  contact_14_100
timestamp 1644951705
transform 1 0 3764 0 1 31196
box 0 0 1 1
use contact_14  contact_14_101
timestamp 1644951705
transform 1 0 3260 0 1 31282
box 0 0 1 1
use contact_14  contact_14_102
timestamp 1644951705
transform 1 0 4100 0 1 31368
box 0 0 1 1
use contact_14  contact_14_103
timestamp 1644951705
transform 1 0 3764 0 1 31454
box 0 0 1 1
use contact_14  contact_14_104
timestamp 1644951705
transform 1 0 3176 0 1 31540
box 0 0 1 1
use contact_14  contact_14_105
timestamp 1644951705
transform 1 0 4100 0 1 31626
box 0 0 1 1
use contact_14  contact_14_106
timestamp 1644951705
transform 1 0 3680 0 1 31712
box 0 0 1 1
use contact_14  contact_14_107
timestamp 1644951705
transform 1 0 3428 0 1 31798
box 0 0 1 1
use contact_14  contact_14_108
timestamp 1644951705
transform 1 0 4100 0 1 30346
box 0 0 1 1
use contact_14  contact_14_109
timestamp 1644951705
transform 1 0 3680 0 1 30260
box 0 0 1 1
use contact_14  contact_14_110
timestamp 1644951705
transform 1 0 3344 0 1 30174
box 0 0 1 1
use contact_14  contact_14_111
timestamp 1644951705
transform 1 0 4100 0 1 30088
box 0 0 1 1
use contact_14  contact_14_112
timestamp 1644951705
transform 1 0 3680 0 1 30002
box 0 0 1 1
use contact_14  contact_14_113
timestamp 1644951705
transform 1 0 3260 0 1 29916
box 0 0 1 1
use contact_14  contact_14_114
timestamp 1644951705
transform 1 0 4100 0 1 29830
box 0 0 1 1
use contact_14  contact_14_115
timestamp 1644951705
transform 1 0 3680 0 1 29744
box 0 0 1 1
use contact_14  contact_14_116
timestamp 1644951705
transform 1 0 3176 0 1 29658
box 0 0 1 1
use contact_14  contact_14_117
timestamp 1644951705
transform 1 0 4100 0 1 28034
box 0 0 1 1
use contact_14  contact_14_118
timestamp 1644951705
transform 1 0 3596 0 1 28120
box 0 0 1 1
use contact_14  contact_14_119
timestamp 1644951705
transform 1 0 3428 0 1 28206
box 0 0 1 1
use contact_14  contact_14_120
timestamp 1644951705
transform 1 0 4100 0 1 28292
box 0 0 1 1
use contact_14  contact_14_121
timestamp 1644951705
transform 1 0 3596 0 1 28378
box 0 0 1 1
use contact_14  contact_14_122
timestamp 1644951705
transform 1 0 3344 0 1 28464
box 0 0 1 1
use contact_14  contact_14_123
timestamp 1644951705
transform 1 0 4100 0 1 28550
box 0 0 1 1
use contact_14  contact_14_124
timestamp 1644951705
transform 1 0 3596 0 1 28636
box 0 0 1 1
use contact_14  contact_14_125
timestamp 1644951705
transform 1 0 3260 0 1 28722
box 0 0 1 1
use contact_14  contact_14_126
timestamp 1644951705
transform 1 0 4100 0 1 27270
box 0 0 1 1
use contact_14  contact_14_127
timestamp 1644951705
transform 1 0 3596 0 1 27184
box 0 0 1 1
use contact_14  contact_14_128
timestamp 1644951705
transform 1 0 3176 0 1 27098
box 0 0 1 1
use contact_14  contact_14_129
timestamp 1644951705
transform 1 0 4100 0 1 27012
box 0 0 1 1
use contact_14  contact_14_130
timestamp 1644951705
transform 1 0 3512 0 1 26926
box 0 0 1 1
use contact_14  contact_14_131
timestamp 1644951705
transform 1 0 3428 0 1 26840
box 0 0 1 1
use contact_14  contact_14_132
timestamp 1644951705
transform 1 0 4100 0 1 26754
box 0 0 1 1
use contact_14  contact_14_133
timestamp 1644951705
transform 1 0 3512 0 1 26668
box 0 0 1 1
use contact_14  contact_14_134
timestamp 1644951705
transform 1 0 3344 0 1 26582
box 0 0 1 1
use contact_14  contact_14_135
timestamp 1644951705
transform 1 0 4100 0 1 24958
box 0 0 1 1
use contact_14  contact_14_136
timestamp 1644951705
transform 1 0 3512 0 1 25044
box 0 0 1 1
use contact_14  contact_14_137
timestamp 1644951705
transform 1 0 3260 0 1 25130
box 0 0 1 1
use contact_14  contact_14_138
timestamp 1644951705
transform 1 0 4100 0 1 25216
box 0 0 1 1
use contact_14  contact_14_139
timestamp 1644951705
transform 1 0 3512 0 1 25302
box 0 0 1 1
use contact_14  contact_14_140
timestamp 1644951705
transform 1 0 3176 0 1 25388
box 0 0 1 1
use contact_14  contact_14_141
timestamp 1644951705
transform 1 0 4016 0 1 25474
box 0 0 1 1
use contact_14  contact_14_142
timestamp 1644951705
transform 1 0 3764 0 1 25560
box 0 0 1 1
use contact_14  contact_14_143
timestamp 1644951705
transform 1 0 3428 0 1 25646
box 0 0 1 1
use contact_14  contact_14_144
timestamp 1644951705
transform 1 0 4016 0 1 24194
box 0 0 1 1
use contact_14  contact_14_145
timestamp 1644951705
transform 1 0 3764 0 1 24108
box 0 0 1 1
use contact_14  contact_14_146
timestamp 1644951705
transform 1 0 3344 0 1 24022
box 0 0 1 1
use contact_14  contact_14_147
timestamp 1644951705
transform 1 0 4016 0 1 23936
box 0 0 1 1
use contact_14  contact_14_148
timestamp 1644951705
transform 1 0 3764 0 1 23850
box 0 0 1 1
use contact_14  contact_14_149
timestamp 1644951705
transform 1 0 3260 0 1 23764
box 0 0 1 1
use contact_14  contact_14_150
timestamp 1644951705
transform 1 0 4016 0 1 23678
box 0 0 1 1
use contact_14  contact_14_151
timestamp 1644951705
transform 1 0 3764 0 1 23592
box 0 0 1 1
use contact_14  contact_14_152
timestamp 1644951705
transform 1 0 3176 0 1 23506
box 0 0 1 1
use contact_14  contact_14_153
timestamp 1644951705
transform 1 0 4016 0 1 21882
box 0 0 1 1
use contact_14  contact_14_154
timestamp 1644951705
transform 1 0 3680 0 1 21968
box 0 0 1 1
use contact_14  contact_14_155
timestamp 1644951705
transform 1 0 3428 0 1 22054
box 0 0 1 1
use contact_14  contact_14_156
timestamp 1644951705
transform 1 0 4016 0 1 22140
box 0 0 1 1
use contact_14  contact_14_157
timestamp 1644951705
transform 1 0 3680 0 1 22226
box 0 0 1 1
use contact_14  contact_14_158
timestamp 1644951705
transform 1 0 3344 0 1 22312
box 0 0 1 1
use contact_14  contact_14_159
timestamp 1644951705
transform 1 0 4016 0 1 22398
box 0 0 1 1
use contact_14  contact_14_160
timestamp 1644951705
transform 1 0 3680 0 1 22484
box 0 0 1 1
use contact_14  contact_14_161
timestamp 1644951705
transform 1 0 3260 0 1 22570
box 0 0 1 1
use contact_14  contact_14_162
timestamp 1644951705
transform 1 0 4016 0 1 21118
box 0 0 1 1
use contact_14  contact_14_163
timestamp 1644951705
transform 1 0 3680 0 1 21032
box 0 0 1 1
use contact_14  contact_14_164
timestamp 1644951705
transform 1 0 3176 0 1 20946
box 0 0 1 1
use contact_14  contact_14_165
timestamp 1644951705
transform 1 0 4016 0 1 20860
box 0 0 1 1
use contact_14  contact_14_166
timestamp 1644951705
transform 1 0 3596 0 1 20774
box 0 0 1 1
use contact_14  contact_14_167
timestamp 1644951705
transform 1 0 3428 0 1 20688
box 0 0 1 1
use contact_14  contact_14_168
timestamp 1644951705
transform 1 0 4016 0 1 20602
box 0 0 1 1
use contact_14  contact_14_169
timestamp 1644951705
transform 1 0 3596 0 1 20516
box 0 0 1 1
use contact_14  contact_14_170
timestamp 1644951705
transform 1 0 3344 0 1 20430
box 0 0 1 1
use contact_14  contact_14_171
timestamp 1644951705
transform 1 0 4016 0 1 18806
box 0 0 1 1
use contact_14  contact_14_172
timestamp 1644951705
transform 1 0 3596 0 1 18892
box 0 0 1 1
use contact_14  contact_14_173
timestamp 1644951705
transform 1 0 3260 0 1 18978
box 0 0 1 1
use contact_14  contact_14_174
timestamp 1644951705
transform 1 0 4016 0 1 19064
box 0 0 1 1
use contact_14  contact_14_175
timestamp 1644951705
transform 1 0 3596 0 1 19150
box 0 0 1 1
use contact_14  contact_14_176
timestamp 1644951705
transform 1 0 3176 0 1 19236
box 0 0 1 1
use contact_14  contact_14_177
timestamp 1644951705
transform 1 0 4016 0 1 19322
box 0 0 1 1
use contact_14  contact_14_178
timestamp 1644951705
transform 1 0 3512 0 1 19408
box 0 0 1 1
use contact_14  contact_14_179
timestamp 1644951705
transform 1 0 3428 0 1 19494
box 0 0 1 1
use contact_14  contact_14_180
timestamp 1644951705
transform 1 0 4016 0 1 18042
box 0 0 1 1
use contact_14  contact_14_181
timestamp 1644951705
transform 1 0 3512 0 1 17956
box 0 0 1 1
use contact_14  contact_14_182
timestamp 1644951705
transform 1 0 3344 0 1 17870
box 0 0 1 1
use contact_14  contact_14_183
timestamp 1644951705
transform 1 0 4016 0 1 17784
box 0 0 1 1
use contact_14  contact_14_184
timestamp 1644951705
transform 1 0 3512 0 1 17698
box 0 0 1 1
use contact_14  contact_14_185
timestamp 1644951705
transform 1 0 3260 0 1 17612
box 0 0 1 1
use contact_14  contact_14_186
timestamp 1644951705
transform 1 0 4016 0 1 17526
box 0 0 1 1
use contact_14  contact_14_187
timestamp 1644951705
transform 1 0 3512 0 1 17440
box 0 0 1 1
use contact_14  contact_14_188
timestamp 1644951705
transform 1 0 3176 0 1 17354
box 0 0 1 1
use contact_14  contact_14_189
timestamp 1644951705
transform 1 0 3932 0 1 15730
box 0 0 1 1
use contact_14  contact_14_190
timestamp 1644951705
transform 1 0 3764 0 1 15816
box 0 0 1 1
use contact_14  contact_14_191
timestamp 1644951705
transform 1 0 3428 0 1 15902
box 0 0 1 1
use contact_14  contact_14_192
timestamp 1644951705
transform 1 0 3932 0 1 15988
box 0 0 1 1
use contact_14  contact_14_193
timestamp 1644951705
transform 1 0 3764 0 1 16074
box 0 0 1 1
use contact_14  contact_14_194
timestamp 1644951705
transform 1 0 3344 0 1 16160
box 0 0 1 1
use contact_14  contact_14_195
timestamp 1644951705
transform 1 0 3932 0 1 16246
box 0 0 1 1
use contact_14  contact_14_196
timestamp 1644951705
transform 1 0 3764 0 1 16332
box 0 0 1 1
use contact_14  contact_14_197
timestamp 1644951705
transform 1 0 3260 0 1 16418
box 0 0 1 1
use contact_14  contact_14_198
timestamp 1644951705
transform 1 0 3932 0 1 14966
box 0 0 1 1
use contact_14  contact_14_199
timestamp 1644951705
transform 1 0 3764 0 1 14880
box 0 0 1 1
use contact_14  contact_14_200
timestamp 1644951705
transform 1 0 3176 0 1 14794
box 0 0 1 1
use contact_14  contact_14_201
timestamp 1644951705
transform 1 0 3932 0 1 14708
box 0 0 1 1
use contact_14  contact_14_202
timestamp 1644951705
transform 1 0 3680 0 1 14622
box 0 0 1 1
use contact_14  contact_14_203
timestamp 1644951705
transform 1 0 3428 0 1 14536
box 0 0 1 1
use contact_14  contact_14_204
timestamp 1644951705
transform 1 0 3932 0 1 14450
box 0 0 1 1
use contact_14  contact_14_205
timestamp 1644951705
transform 1 0 3680 0 1 14364
box 0 0 1 1
use contact_14  contact_14_206
timestamp 1644951705
transform 1 0 3344 0 1 14278
box 0 0 1 1
use contact_14  contact_14_207
timestamp 1644951705
transform 1 0 3932 0 1 12654
box 0 0 1 1
use contact_14  contact_14_208
timestamp 1644951705
transform 1 0 3680 0 1 12740
box 0 0 1 1
use contact_14  contact_14_209
timestamp 1644951705
transform 1 0 3260 0 1 12826
box 0 0 1 1
use contact_14  contact_14_210
timestamp 1644951705
transform 1 0 3932 0 1 12912
box 0 0 1 1
use contact_14  contact_14_211
timestamp 1644951705
transform 1 0 3680 0 1 12998
box 0 0 1 1
use contact_14  contact_14_212
timestamp 1644951705
transform 1 0 3176 0 1 13084
box 0 0 1 1
use contact_14  contact_14_213
timestamp 1644951705
transform 1 0 3932 0 1 13170
box 0 0 1 1
use contact_14  contact_14_214
timestamp 1644951705
transform 1 0 3596 0 1 13256
box 0 0 1 1
use contact_14  contact_14_215
timestamp 1644951705
transform 1 0 3428 0 1 13342
box 0 0 1 1
use contact_14  contact_14_216
timestamp 1644951705
transform 1 0 3932 0 1 11890
box 0 0 1 1
use contact_14  contact_14_217
timestamp 1644951705
transform 1 0 3596 0 1 11804
box 0 0 1 1
use contact_14  contact_14_218
timestamp 1644951705
transform 1 0 3344 0 1 11718
box 0 0 1 1
use contact_14  contact_14_219
timestamp 1644951705
transform 1 0 3932 0 1 11632
box 0 0 1 1
use contact_14  contact_14_220
timestamp 1644951705
transform 1 0 3596 0 1 11546
box 0 0 1 1
use contact_14  contact_14_221
timestamp 1644951705
transform 1 0 3260 0 1 11460
box 0 0 1 1
use contact_14  contact_14_222
timestamp 1644951705
transform 1 0 3932 0 1 11374
box 0 0 1 1
use contact_14  contact_14_223
timestamp 1644951705
transform 1 0 3596 0 1 11288
box 0 0 1 1
use contact_14  contact_14_224
timestamp 1644951705
transform 1 0 3176 0 1 11202
box 0 0 1 1
use contact_14  contact_14_225
timestamp 1644951705
transform 1 0 3932 0 1 9578
box 0 0 1 1
use contact_14  contact_14_226
timestamp 1644951705
transform 1 0 3512 0 1 9664
box 0 0 1 1
use contact_14  contact_14_227
timestamp 1644951705
transform 1 0 3428 0 1 9750
box 0 0 1 1
use contact_14  contact_14_228
timestamp 1644951705
transform 1 0 3932 0 1 9836
box 0 0 1 1
use contact_14  contact_14_229
timestamp 1644951705
transform 1 0 3512 0 1 9922
box 0 0 1 1
use contact_14  contact_14_230
timestamp 1644951705
transform 1 0 3344 0 1 10008
box 0 0 1 1
use contact_14  contact_14_231
timestamp 1644951705
transform 1 0 3932 0 1 10094
box 0 0 1 1
use contact_14  contact_14_232
timestamp 1644951705
transform 1 0 3512 0 1 10180
box 0 0 1 1
use contact_14  contact_14_233
timestamp 1644951705
transform 1 0 3260 0 1 10266
box 0 0 1 1
use contact_14  contact_14_234
timestamp 1644951705
transform 1 0 3932 0 1 8814
box 0 0 1 1
use contact_14  contact_14_235
timestamp 1644951705
transform 1 0 3512 0 1 8728
box 0 0 1 1
use contact_14  contact_14_236
timestamp 1644951705
transform 1 0 3176 0 1 8642
box 0 0 1 1
use contact_14  contact_14_237
timestamp 1644951705
transform 1 0 3848 0 1 8556
box 0 0 1 1
use contact_14  contact_14_238
timestamp 1644951705
transform 1 0 3764 0 1 8470
box 0 0 1 1
use contact_14  contact_14_239
timestamp 1644951705
transform 1 0 3428 0 1 8384
box 0 0 1 1
use contact_14  contact_14_240
timestamp 1644951705
transform 1 0 3848 0 1 8298
box 0 0 1 1
use contact_14  contact_14_241
timestamp 1644951705
transform 1 0 3764 0 1 8212
box 0 0 1 1
use contact_14  contact_14_242
timestamp 1644951705
transform 1 0 3344 0 1 8126
box 0 0 1 1
use contact_14  contact_14_243
timestamp 1644951705
transform 1 0 3848 0 1 6502
box 0 0 1 1
use contact_14  contact_14_244
timestamp 1644951705
transform 1 0 3764 0 1 6588
box 0 0 1 1
use contact_14  contact_14_245
timestamp 1644951705
transform 1 0 3260 0 1 6674
box 0 0 1 1
use contact_14  contact_14_246
timestamp 1644951705
transform 1 0 3848 0 1 6760
box 0 0 1 1
use contact_14  contact_14_247
timestamp 1644951705
transform 1 0 3764 0 1 6846
box 0 0 1 1
use contact_14  contact_14_248
timestamp 1644951705
transform 1 0 3176 0 1 6932
box 0 0 1 1
use contact_14  contact_14_249
timestamp 1644951705
transform 1 0 3848 0 1 7018
box 0 0 1 1
use contact_14  contact_14_250
timestamp 1644951705
transform 1 0 3680 0 1 7104
box 0 0 1 1
use contact_14  contact_14_251
timestamp 1644951705
transform 1 0 3428 0 1 7190
box 0 0 1 1
use contact_14  contact_14_252
timestamp 1644951705
transform 1 0 3848 0 1 5738
box 0 0 1 1
use contact_14  contact_14_253
timestamp 1644951705
transform 1 0 3680 0 1 5652
box 0 0 1 1
use contact_14  contact_14_254
timestamp 1644951705
transform 1 0 3344 0 1 5566
box 0 0 1 1
use contact_14  contact_14_255
timestamp 1644951705
transform 1 0 3848 0 1 5480
box 0 0 1 1
use contact_14  contact_14_256
timestamp 1644951705
transform 1 0 3680 0 1 5394
box 0 0 1 1
use contact_14  contact_14_257
timestamp 1644951705
transform 1 0 3260 0 1 5308
box 0 0 1 1
use contact_14  contact_14_258
timestamp 1644951705
transform 1 0 3848 0 1 5222
box 0 0 1 1
use contact_14  contact_14_259
timestamp 1644951705
transform 1 0 3680 0 1 5136
box 0 0 1 1
use contact_14  contact_14_260
timestamp 1644951705
transform 1 0 3176 0 1 5050
box 0 0 1 1
use contact_14  contact_14_261
timestamp 1644951705
transform 1 0 3848 0 1 3426
box 0 0 1 1
use contact_14  contact_14_262
timestamp 1644951705
transform 1 0 3596 0 1 3512
box 0 0 1 1
use contact_14  contact_14_263
timestamp 1644951705
transform 1 0 3428 0 1 3598
box 0 0 1 1
use contact_14  contact_14_264
timestamp 1644951705
transform 1 0 3848 0 1 3684
box 0 0 1 1
use contact_14  contact_14_265
timestamp 1644951705
transform 1 0 3596 0 1 3770
box 0 0 1 1
use contact_14  contact_14_266
timestamp 1644951705
transform 1 0 3344 0 1 3856
box 0 0 1 1
use contact_14  contact_14_267
timestamp 1644951705
transform 1 0 3848 0 1 3942
box 0 0 1 1
use contact_14  contact_14_268
timestamp 1644951705
transform 1 0 3596 0 1 4028
box 0 0 1 1
use contact_14  contact_14_269
timestamp 1644951705
transform 1 0 3260 0 1 4114
box 0 0 1 1
use contact_14  contact_14_270
timestamp 1644951705
transform 1 0 3848 0 1 2662
box 0 0 1 1
use contact_14  contact_14_271
timestamp 1644951705
transform 1 0 3596 0 1 2576
box 0 0 1 1
use contact_14  contact_14_272
timestamp 1644951705
transform 1 0 3176 0 1 2490
box 0 0 1 1
use contact_14  contact_14_273
timestamp 1644951705
transform 1 0 3848 0 1 2404
box 0 0 1 1
use contact_14  contact_14_274
timestamp 1644951705
transform 1 0 3512 0 1 2318
box 0 0 1 1
use contact_14  contact_14_275
timestamp 1644951705
transform 1 0 3428 0 1 2232
box 0 0 1 1
use contact_14  contact_14_276
timestamp 1644951705
transform 1 0 3848 0 1 2146
box 0 0 1 1
use contact_14  contact_14_277
timestamp 1644951705
transform 1 0 3512 0 1 2060
box 0 0 1 1
use contact_14  contact_14_278
timestamp 1644951705
transform 1 0 3344 0 1 1974
box 0 0 1 1
use contact_14  contact_14_279
timestamp 1644951705
transform 1 0 3848 0 1 350
box 0 0 1 1
use contact_14  contact_14_280
timestamp 1644951705
transform 1 0 3512 0 1 436
box 0 0 1 1
use contact_14  contact_14_281
timestamp 1644951705
transform 1 0 3260 0 1 522
box 0 0 1 1
use contact_14  contact_14_282
timestamp 1644951705
transform 1 0 3848 0 1 608
box 0 0 1 1
use contact_14  contact_14_283
timestamp 1644951705
transform 1 0 3512 0 1 694
box 0 0 1 1
use contact_14  contact_14_284
timestamp 1644951705
transform 1 0 3176 0 1 780
box 0 0 1 1
use contact_14  contact_14_285
timestamp 1644951705
transform 1 0 504 0 1 22248
box 0 0 1 1
use contact_17  contact_17_80
timestamp 1644951705
transform 1 0 868 0 1 22248
box 0 0 1 1
use contact_14  contact_14_286
timestamp 1644951705
transform 1 0 420 0 1 20792
box 0 0 1 1
use contact_17  contact_17_81
timestamp 1644951705
transform 1 0 784 0 1 20792
box 0 0 1 1
use contact_14  contact_14_287
timestamp 1644951705
transform 1 0 336 0 1 19168
box 0 0 1 1
use contact_17  contact_17_82
timestamp 1644951705
transform 1 0 700 0 1 19168
box 0 0 1 1
use contact_14  contact_14_288
timestamp 1644951705
transform 1 0 252 0 1 11556
box 0 0 1 1
use contact_17  contact_17_83
timestamp 1644951705
transform 1 0 1216 0 1 11556
box 0 0 1 1
use contact_14  contact_14_289
timestamp 1644951705
transform 1 0 168 0 1 9932
box 0 0 1 1
use contact_17  contact_17_84
timestamp 1644951705
transform 1 0 1132 0 1 9932
box 0 0 1 1
use contact_14  contact_14_290
timestamp 1644951705
transform 1 0 84 0 1 2320
box 0 0 1 1
use contact_17  contact_17_85
timestamp 1644951705
transform 1 0 1216 0 1 2320
box 0 0 1 1
use contact_14  contact_14_291
timestamp 1644951705
transform 1 0 0 0 1 696
box 0 0 1 1
use contact_17  contact_17_86
timestamp 1644951705
transform 1 0 1132 0 1 696
box 0 0 1 1
use dec_cell3_2r1w  dec_cell3_2r1w_0
timestamp 1644951705
transform 1 0 4538 0 -1 49216
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_1
timestamp 1644951705
transform 1 0 4538 0 1 46140
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_2
timestamp 1644951705
transform 1 0 4538 0 -1 46140
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_3
timestamp 1644951705
transform 1 0 4538 0 1 43064
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_4
timestamp 1644951705
transform 1 0 4538 0 -1 43064
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_5
timestamp 1644951705
transform 1 0 4538 0 1 39988
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_6
timestamp 1644951705
transform 1 0 4538 0 -1 39988
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_7
timestamp 1644951705
transform 1 0 4538 0 1 36912
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_8
timestamp 1644951705
transform 1 0 4538 0 -1 36912
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_9
timestamp 1644951705
transform 1 0 4538 0 1 33836
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_10
timestamp 1644951705
transform 1 0 4538 0 -1 33836
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_11
timestamp 1644951705
transform 1 0 4538 0 1 30760
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_12
timestamp 1644951705
transform 1 0 4538 0 -1 30760
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_13
timestamp 1644951705
transform 1 0 4538 0 1 27684
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_14
timestamp 1644951705
transform 1 0 4538 0 -1 27684
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_15
timestamp 1644951705
transform 1 0 4538 0 1 24608
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_16
timestamp 1644951705
transform 1 0 4538 0 -1 24608
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_17
timestamp 1644951705
transform 1 0 4538 0 1 21532
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_18
timestamp 1644951705
transform 1 0 4538 0 -1 21532
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_19
timestamp 1644951705
transform 1 0 4538 0 1 18456
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_20
timestamp 1644951705
transform 1 0 4538 0 -1 18456
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_21
timestamp 1644951705
transform 1 0 4538 0 1 15380
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_22
timestamp 1644951705
transform 1 0 4538 0 -1 15380
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_23
timestamp 1644951705
transform 1 0 4538 0 1 12304
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_24
timestamp 1644951705
transform 1 0 4538 0 -1 12304
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_25
timestamp 1644951705
transform 1 0 4538 0 1 9228
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_26
timestamp 1644951705
transform 1 0 4538 0 -1 9228
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_27
timestamp 1644951705
transform 1 0 4538 0 1 6152
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_28
timestamp 1644951705
transform 1 0 4538 0 -1 6152
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_29
timestamp 1644951705
transform 1 0 4538 0 1 3076
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_30
timestamp 1644951705
transform 1 0 4538 0 -1 3076
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_31
timestamp 1644951705
transform 1 0 4538 0 1 0
box 0 -42 1494 1616
use hierarchical_predecode3x8  hierarchical_predecode3x8_0
timestamp 1644951705
transform 1 0 634 0 1 18472
box 0 -37 2512 12357
use hierarchical_predecode2x4  hierarchical_predecode2x4_0
timestamp 1644951705
transform 1 0 1066 0 1 9236
box 0 -37 2080 6197
use hierarchical_predecode2x4  hierarchical_predecode2x4_1
timestamp 1644951705
transform 1 0 1066 0 1 0
box 0 -37 2080 6197
<< labels >>
rlabel metal2 s 18 0 46 30792 4 addr_0
rlabel metal2 s 102 0 130 30792 4 addr_1
rlabel metal2 s 186 0 214 30792 4 addr_2
rlabel metal2 s 270 0 298 30792 4 addr_3
rlabel metal2 s 354 0 382 30792 4 addr_4
rlabel metal2 s 438 0 466 30792 4 addr_5
rlabel metal2 s 522 0 550 30792 4 addr_6
rlabel metal1 s 5956 848 6032 876 4 decode0_0
rlabel metal1 s 5748 702 6032 730 4 decode1_0
rlabel metal1 s 5666 580 6032 608 4 decode2_0
rlabel metal1 s 5956 2200 6032 2228 4 decode0_1
rlabel metal1 s 5748 2346 6032 2374 4 decode1_1
rlabel metal1 s 5666 2468 6032 2496 4 decode2_1
rlabel metal1 s 5956 3924 6032 3952 4 decode0_2
rlabel metal1 s 5748 3778 6032 3806 4 decode1_2
rlabel metal1 s 5666 3656 6032 3684 4 decode2_2
rlabel metal1 s 5956 5276 6032 5304 4 decode0_3
rlabel metal1 s 5748 5422 6032 5450 4 decode1_3
rlabel metal1 s 5666 5544 6032 5572 4 decode2_3
rlabel metal1 s 5956 7000 6032 7028 4 decode0_4
rlabel metal1 s 5748 6854 6032 6882 4 decode1_4
rlabel metal1 s 5666 6732 6032 6760 4 decode2_4
rlabel metal1 s 5956 8352 6032 8380 4 decode0_5
rlabel metal1 s 5748 8498 6032 8526 4 decode1_5
rlabel metal1 s 5666 8620 6032 8648 4 decode2_5
rlabel metal1 s 5956 10076 6032 10104 4 decode0_6
rlabel metal1 s 5748 9930 6032 9958 4 decode1_6
rlabel metal1 s 5666 9808 6032 9836 4 decode2_6
rlabel metal1 s 5956 11428 6032 11456 4 decode0_7
rlabel metal1 s 5748 11574 6032 11602 4 decode1_7
rlabel metal1 s 5666 11696 6032 11724 4 decode2_7
rlabel metal1 s 5956 13152 6032 13180 4 decode0_8
rlabel metal1 s 5748 13006 6032 13034 4 decode1_8
rlabel metal1 s 5666 12884 6032 12912 4 decode2_8
rlabel metal1 s 5956 14504 6032 14532 4 decode0_9
rlabel metal1 s 5748 14650 6032 14678 4 decode1_9
rlabel metal1 s 5666 14772 6032 14800 4 decode2_9
rlabel metal1 s 5956 16228 6032 16256 4 decode0_10
rlabel metal1 s 5748 16082 6032 16110 4 decode1_10
rlabel metal1 s 5666 15960 6032 15988 4 decode2_10
rlabel metal1 s 5956 17580 6032 17608 4 decode0_11
rlabel metal1 s 5748 17726 6032 17754 4 decode1_11
rlabel metal1 s 5666 17848 6032 17876 4 decode2_11
rlabel metal1 s 5956 19304 6032 19332 4 decode0_12
rlabel metal1 s 5748 19158 6032 19186 4 decode1_12
rlabel metal1 s 5666 19036 6032 19064 4 decode2_12
rlabel metal1 s 5956 20656 6032 20684 4 decode0_13
rlabel metal1 s 5748 20802 6032 20830 4 decode1_13
rlabel metal1 s 5666 20924 6032 20952 4 decode2_13
rlabel metal1 s 5956 22380 6032 22408 4 decode0_14
rlabel metal1 s 5748 22234 6032 22262 4 decode1_14
rlabel metal1 s 5666 22112 6032 22140 4 decode2_14
rlabel metal1 s 5956 23732 6032 23760 4 decode0_15
rlabel metal1 s 5748 23878 6032 23906 4 decode1_15
rlabel metal1 s 5666 24000 6032 24028 4 decode2_15
rlabel metal1 s 5956 25456 6032 25484 4 decode0_16
rlabel metal1 s 5748 25310 6032 25338 4 decode1_16
rlabel metal1 s 5666 25188 6032 25216 4 decode2_16
rlabel metal1 s 5956 26808 6032 26836 4 decode0_17
rlabel metal1 s 5748 26954 6032 26982 4 decode1_17
rlabel metal1 s 5666 27076 6032 27104 4 decode2_17
rlabel metal1 s 5956 28532 6032 28560 4 decode0_18
rlabel metal1 s 5748 28386 6032 28414 4 decode1_18
rlabel metal1 s 5666 28264 6032 28292 4 decode2_18
rlabel metal1 s 5956 29884 6032 29912 4 decode0_19
rlabel metal1 s 5748 30030 6032 30058 4 decode1_19
rlabel metal1 s 5666 30152 6032 30180 4 decode2_19
rlabel metal1 s 5956 31608 6032 31636 4 decode0_20
rlabel metal1 s 5748 31462 6032 31490 4 decode1_20
rlabel metal1 s 5666 31340 6032 31368 4 decode2_20
rlabel metal1 s 5956 32960 6032 32988 4 decode0_21
rlabel metal1 s 5748 33106 6032 33134 4 decode1_21
rlabel metal1 s 5666 33228 6032 33256 4 decode2_21
rlabel metal1 s 5956 34684 6032 34712 4 decode0_22
rlabel metal1 s 5748 34538 6032 34566 4 decode1_22
rlabel metal1 s 5666 34416 6032 34444 4 decode2_22
rlabel metal1 s 5956 36036 6032 36064 4 decode0_23
rlabel metal1 s 5748 36182 6032 36210 4 decode1_23
rlabel metal1 s 5666 36304 6032 36332 4 decode2_23
rlabel metal1 s 5956 37760 6032 37788 4 decode0_24
rlabel metal1 s 5748 37614 6032 37642 4 decode1_24
rlabel metal1 s 5666 37492 6032 37520 4 decode2_24
rlabel metal1 s 5956 39112 6032 39140 4 decode0_25
rlabel metal1 s 5748 39258 6032 39286 4 decode1_25
rlabel metal1 s 5666 39380 6032 39408 4 decode2_25
rlabel metal1 s 5956 40836 6032 40864 4 decode0_26
rlabel metal1 s 5748 40690 6032 40718 4 decode1_26
rlabel metal1 s 5666 40568 6032 40596 4 decode2_26
rlabel metal1 s 5956 42188 6032 42216 4 decode0_27
rlabel metal1 s 5748 42334 6032 42362 4 decode1_27
rlabel metal1 s 5666 42456 6032 42484 4 decode2_27
rlabel metal1 s 5956 43912 6032 43940 4 decode0_28
rlabel metal1 s 5748 43766 6032 43794 4 decode1_28
rlabel metal1 s 5666 43644 6032 43672 4 decode2_28
rlabel metal1 s 5956 45264 6032 45292 4 decode0_29
rlabel metal1 s 5748 45410 6032 45438 4 decode1_29
rlabel metal1 s 5666 45532 6032 45560 4 decode2_29
rlabel metal1 s 5956 46988 6032 47016 4 decode0_30
rlabel metal1 s 5748 46842 6032 46870 4 decode1_30
rlabel metal1 s 5666 46720 6032 46748 4 decode2_30
rlabel metal1 s 5956 48340 6032 48368 4 decode0_31
rlabel metal1 s 5748 48486 6032 48514 4 decode1_31
rlabel metal1 s 5666 48608 6032 48636 4 decode2_31
rlabel metal2 s 3194 0 3222 49244 4 predecode_0
rlabel metal2 s 3278 0 3306 49244 4 predecode_1
rlabel metal2 s 3362 0 3390 49244 4 predecode_2
rlabel metal2 s 3446 0 3474 49244 4 predecode_3
rlabel metal2 s 3530 0 3558 49244 4 predecode_4
rlabel metal2 s 3614 0 3642 49244 4 predecode_5
rlabel metal2 s 3698 0 3726 49244 4 predecode_6
rlabel metal2 s 3782 0 3810 49244 4 predecode_7
rlabel metal2 s 3866 0 3894 49244 4 predecode_8
rlabel metal2 s 3950 0 3978 49244 4 predecode_9
rlabel metal2 s 4034 0 4062 49244 4 predecode_10
rlabel metal2 s 4118 0 4146 49244 4 predecode_11
rlabel metal2 s 4202 0 4230 49244 4 predecode_12
rlabel metal2 s 4286 0 4314 49244 4 predecode_13
rlabel metal2 s 4370 0 4398 49244 4 predecode_14
rlabel metal2 s 4454 0 4482 49244 4 predecode_15
rlabel metal3 s 960 29215 1092 29289 4 vdd
rlabel metal3 s 5980 38413 6112 38487 4 vdd
rlabel metal3 s 1308 4583 1440 4657 4 vdd
rlabel metal3 s 960 26135 1092 26209 4 vdd
rlabel metal3 s 5980 19957 6112 20031 4 vdd
rlabel metal3 s 5980 16881 6112 16955 4 vdd
rlabel metal3 s 5980 29185 6112 29259 4 vdd
rlabel metal3 s 5980 13805 6112 13879 4 vdd
rlabel metal3 s 5980 41489 6112 41563 4 vdd
rlabel metal3 s 5980 35337 6112 35411 4 vdd
rlabel metal3 s 5980 44565 6112 44639 4 vdd
rlabel metal3 s 6046 44602 6046 44602 4 vdd
rlabel metal3 s 1308 1503 1440 1577 4 vdd
rlabel metal3 s 960 19975 1092 20049 4 vdd
rlabel metal3 s 5980 47641 6112 47715 4 vdd
rlabel metal3 s 2180 4583 2312 4657 4 vdd
rlabel metal3 s 2180 1503 2312 1577 4 vdd
rlabel metal3 s 1308 10739 1440 10813 4 vdd
rlabel metal3 s 960 23055 1092 23129 4 vdd
rlabel metal3 s 2180 13819 2312 13893 4 vdd
rlabel metal3 s 5980 10729 6112 10803 4 vdd
rlabel metal3 s 6046 10766 6046 10766 4 vdd
rlabel metal3 s 5980 4577 6112 4651 4 vdd
rlabel metal3 s 1308 13819 1440 13893 4 vdd
rlabel metal3 s 2180 10739 2312 10813 4 vdd
rlabel metal3 s 5980 26109 6112 26183 4 vdd
rlabel metal3 s 2000 19975 2132 20049 4 vdd
rlabel metal3 s 5980 1501 6112 1575 4 vdd
rlabel metal3 s 6046 1538 6046 1538 4 vdd
rlabel metal3 s 5980 32261 6112 32335 4 vdd
rlabel metal3 s 2000 23055 2132 23129 4 vdd
rlabel metal3 s 5980 23033 6112 23107 4 vdd
rlabel metal3 s 2000 26135 2132 26209 4 vdd
rlabel metal3 s 2000 29215 2132 29289 4 vdd
rlabel metal3 s 5980 7653 6112 7727 4 vdd
rlabel metal3 s 2000 30755 2132 30829 4 gnd
rlabel metal3 s 5980 21495 6112 21569 4 gnd
rlabel metal3 s 960 18435 1092 18509 4 gnd
rlabel metal3 s 2180 9199 2312 9273 4 gnd
rlabel metal3 s 5980 30723 6112 30797 4 gnd
rlabel metal3 s 5980 46103 6112 46177 4 gnd
rlabel metal3 s 1308 6123 1440 6197 4 gnd
rlabel metal3 s 5980 36875 6112 36949 4 gnd
rlabel metal3 s 5980 9191 6112 9265 4 gnd
rlabel metal3 s 2000 27675 2132 27749 4 gnd
rlabel metal3 s 5980 18419 6112 18493 4 gnd
rlabel metal3 s 5980 15343 6112 15417 4 gnd
rlabel metal3 s 5980 33799 6112 33873 4 gnd
rlabel metal3 s 5980 3039 6112 3113 4 gnd
rlabel metal3 s 960 21515 1092 21589 4 gnd
rlabel metal3 s 1308 3043 1440 3117 4 gnd
rlabel metal3 s 2000 21515 2132 21589 4 gnd
rlabel metal3 s 1308 12279 1440 12353 4 gnd
rlabel metal3 s 1308 9199 1440 9273 4 gnd
rlabel metal3 s 2180 12279 2312 12353 4 gnd
rlabel metal3 s 2180 3043 2312 3117 4 gnd
rlabel metal3 s 5980 24571 6112 24645 4 gnd
rlabel metal3 s 960 30755 1092 30829 4 gnd
rlabel metal3 s 5980 27647 6112 27721 4 gnd
rlabel metal3 s 2180 -37 2312 37 4 gnd
rlabel metal3 s 2000 18435 2132 18509 4 gnd
rlabel metal3 s 2000 24595 2132 24669 4 gnd
rlabel metal3 s 5980 43027 6112 43101 4 gnd
rlabel metal3 s 2180 6123 2312 6197 4 gnd
rlabel metal3 s 960 24595 1092 24669 4 gnd
rlabel metal3 s 5980 49179 6112 49253 4 gnd
rlabel metal3 s 5980 6115 6112 6189 4 gnd
rlabel metal3 s 1308 15359 1440 15433 4 gnd
rlabel metal3 s 5980 39951 6112 40025 4 gnd
rlabel metal3 s 5980 -37 6112 37 4 gnd
rlabel metal3 s 1308 -37 1440 37 4 gnd
rlabel metal3 s 2180 15359 2312 15433 4 gnd
rlabel metal3 s 5980 12267 6112 12341 4 gnd
rlabel metal3 s 960 27675 1092 27749 4 gnd
<< properties >>
string FIXED_BBOX 5980 -37 6112 0
string GDS_FILE sram_0rw2r1w_16_128_sky130A.gds
string GDS_END 1772100
string GDS_START 1667992
<< end >>
