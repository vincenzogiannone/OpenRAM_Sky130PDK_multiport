VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO sram_0rw2r1w_32_128_sky130A
   CLASS BLOCK ;
   SIZE 397.2 BY 564.68 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  106.0 0.0 106.76 1.82 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  113.42 0.0 114.18 1.82 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  120.84 0.0 121.6 1.82 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  128.26 0.0 129.02 1.82 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  136.74 0.0 137.5 1.82 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  144.16 0.0 144.92 1.82 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  150.52 0.0 151.28 1.82 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  159.0 0.0 159.76 1.82 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  165.36 0.0 166.12 1.82 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  173.84 0.0 174.6 1.82 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  181.26 0.0 182.02 1.82 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  188.68 0.0 189.44 1.82 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  196.1 0.0 196.86 1.82 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  202.46 0.0 203.22 1.82 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  209.88 0.0 210.64 1.82 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  217.3 0.0 218.06 1.82 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  224.72 0.0 225.48 1.82 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  232.14 0.0 232.9 1.82 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  239.56 0.0 240.32 1.82 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  246.98 0.0 247.74 1.82 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  254.4 0.0 255.16 1.82 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  261.82 0.0 262.58 1.82 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  269.24 0.0 270.0 1.82 ;
      END
   END din0[22]
   PIN din0[23]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  276.66 0.0 277.42 1.82 ;
      END
   END din0[23]
   PIN din0[24]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  284.08 0.0 284.84 1.82 ;
      END
   END din0[24]
   PIN din0[25]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  290.44 0.0 291.2 1.82 ;
      END
   END din0[25]
   PIN din0[26]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  298.92 0.0 299.68 1.82 ;
      END
   END din0[26]
   PIN din0[27]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  306.34 0.0 307.1 1.82 ;
      END
   END din0[27]
   PIN din0[28]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  312.7 0.0 313.46 1.82 ;
      END
   END din0[28]
   PIN din0[29]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  321.18 0.0 321.94 1.82 ;
      END
   END din0[29]
   PIN din0[30]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  328.6 0.0 329.36 1.82 ;
      END
   END din0[30]
   PIN din0[31]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  336.02 0.0 336.78 1.82 ;
      END
   END din0[31]
   PIN addr[0]
      DIRECTION INPUT ;
      PORT
      END
   END addr[0]
   PIN addr[1]
      DIRECTION INPUT ;
      PORT
      END
   END addr[1]
   PIN addr[2]
      DIRECTION INPUT ;
      PORT
      END
   END addr[2]
   PIN addr[3]
      DIRECTION INPUT ;
      PORT
      END
   END addr[3]
   PIN addr[4]
      DIRECTION INPUT ;
      PORT
      END
   END addr[4]
   PIN addr[5]
      DIRECTION INPUT ;
      PORT
      END
   END addr[5]
   PIN addr[6]
      DIRECTION INPUT ;
      PORT
      END
   END addr[6]
   PIN addr[7]
      DIRECTION INPUT ;
      PORT
      END
   END addr[7]
   PIN addr[8]
      DIRECTION INPUT ;
      PORT
      END
   END addr[8]
   PIN csb
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  13.765 37.895 14.425 38.265 ;
      END
   END csb
   PIN web
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  13.765 31.975 14.425 32.345 ;
      END
   END web
   PIN clk
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 36.04 1.82 36.8 ;
      END
   END clk
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  134.62 0.0 135.38 1.82 ;
      END
   END dout0[0]
   PIN dout1[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  134.355 53.235 135.015 53.605 ;
      END
   END dout1[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  135.68 0.0 136.44 1.82 ;
      END
   END dout0[1]
   PIN dout1[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  135.715 53.235 136.375 53.605 ;
      END
   END dout1[1]
   PIN dout0[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  142.04 0.0 142.8 1.82 ;
      END
   END dout0[2]
   PIN dout1[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  142.135 53.235 142.795 53.605 ;
      END
   END dout1[2]
   PIN dout0[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  143.1 0.0 143.86 1.82 ;
      END
   END dout0[3]
   PIN dout1[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  143.495 53.235 144.155 53.605 ;
      END
   END dout1[3]
   PIN dout0[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  149.46 0.0 150.22 1.82 ;
      END
   END dout0[4]
   PIN dout1[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  149.915 53.235 150.575 53.605 ;
      END
   END dout1[4]
   PIN dout0[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  151.58 0.0 152.34 1.82 ;
      END
   END dout0[5]
   PIN dout1[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  151.275 53.235 151.935 53.605 ;
      END
   END dout1[5]
   PIN dout0[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  157.94 0.0 158.7 1.82 ;
      END
   END dout0[6]
   PIN dout1[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  157.695 53.235 158.355 53.605 ;
      END
   END dout1[6]
   PIN dout0[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  160.06 0.0 160.82 1.82 ;
      END
   END dout0[7]
   PIN dout1[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  159.055 53.235 159.715 53.605 ;
      END
   END dout1[7]
   PIN dout0[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  166.42 0.0 167.18 1.82 ;
      END
   END dout0[8]
   PIN dout1[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  165.475 53.235 166.135 53.605 ;
      END
   END dout1[8]
   PIN dout0[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  167.48 0.0 168.24 1.82 ;
      END
   END dout0[9]
   PIN dout1[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  166.835 53.235 167.495 53.605 ;
      END
   END dout1[9]
   PIN dout0[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  172.78 0.0 173.54 1.82 ;
      END
   END dout0[10]
   PIN dout1[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  173.255 53.235 173.915 53.605 ;
      END
   END dout1[10]
   PIN dout0[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  174.9 0.0 175.66 1.82 ;
      END
   END dout0[11]
   PIN dout1[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  174.615 53.235 175.275 53.605 ;
      END
   END dout1[11]
   PIN dout0[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  180.2 0.0 180.96 1.82 ;
      END
   END dout0[12]
   PIN dout1[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  181.035 53.235 181.695 53.605 ;
      END
   END dout1[12]
   PIN dout0[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  182.32 0.0 183.08 1.82 ;
      END
   END dout0[13]
   PIN dout1[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  182.395 53.235 183.055 53.605 ;
      END
   END dout1[13]
   PIN dout0[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  189.74 0.0 190.5 1.82 ;
      END
   END dout0[14]
   PIN dout1[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  188.815 53.235 189.475 53.605 ;
      END
   END dout1[14]
   PIN dout0[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  190.8 0.0 191.56 1.82 ;
      END
   END dout0[15]
   PIN dout1[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  190.175 53.235 190.835 53.605 ;
      END
   END dout1[15]
   PIN dout0[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  197.16 0.0 197.92 1.82 ;
      END
   END dout0[16]
   PIN dout1[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  196.595 53.235 197.255 53.605 ;
      END
   END dout1[16]
   PIN dout0[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  198.22 0.0 198.98 1.82 ;
      END
   END dout0[17]
   PIN dout1[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  197.955 53.235 198.615 53.605 ;
      END
   END dout1[17]
   PIN dout0[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  203.52 0.0 204.28 1.82 ;
      END
   END dout0[18]
   PIN dout1[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  204.375 53.235 205.035 53.605 ;
      END
   END dout1[18]
   PIN dout0[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  205.64 0.0 206.4 1.82 ;
      END
   END dout0[19]
   PIN dout1[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  205.735 53.235 206.395 53.605 ;
      END
   END dout1[19]
   PIN dout0[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  212.0 0.0 212.76 1.82 ;
      END
   END dout0[20]
   PIN dout1[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  212.155 53.235 212.815 53.605 ;
      END
   END dout1[20]
   PIN dout0[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  213.06 0.0 213.82 1.82 ;
      END
   END dout0[21]
   PIN dout1[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  213.515 53.235 214.175 53.605 ;
      END
   END dout1[21]
   PIN dout0[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  220.48 0.0 221.24 1.82 ;
      END
   END dout0[22]
   PIN dout1[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  219.935 53.235 220.595 53.605 ;
      END
   END dout1[22]
   PIN dout0[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  221.54 0.0 222.3 1.82 ;
      END
   END dout0[23]
   PIN dout1[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  221.295 53.235 221.955 53.605 ;
      END
   END dout1[23]
   PIN dout0[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  226.84 0.0 227.6 1.82 ;
      END
   END dout0[24]
   PIN dout1[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  227.715 53.235 228.375 53.605 ;
      END
   END dout1[24]
   PIN dout0[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  230.02 0.0 230.78 1.82 ;
      END
   END dout0[25]
   PIN dout1[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  229.075 53.235 229.735 53.605 ;
      END
   END dout1[25]
   PIN dout0[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  235.32 0.0 236.08 1.82 ;
      END
   END dout0[26]
   PIN dout1[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  235.495 53.235 236.155 53.605 ;
      END
   END dout1[26]
   PIN dout0[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  236.38 0.0 237.14 1.82 ;
      END
   END dout0[27]
   PIN dout1[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  236.855 53.235 237.515 53.605 ;
      END
   END dout1[27]
   PIN dout0[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  243.8 0.0 244.56 1.82 ;
      END
   END dout0[28]
   PIN dout1[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  243.275 53.235 243.935 53.605 ;
      END
   END dout1[28]
   PIN dout0[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  244.86 0.0 245.62 1.82 ;
      END
   END dout0[29]
   PIN dout1[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  244.635 53.235 245.295 53.605 ;
      END
   END dout1[29]
   PIN dout0[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  250.16 0.0 250.92 1.82 ;
      END
   END dout0[30]
   PIN dout1[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  251.055 53.235 251.715 53.605 ;
      END
   END dout1[30]
   PIN dout0[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  252.28 0.0 253.04 1.82 ;
      END
   END dout0[31]
   PIN dout1[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  252.415 53.235 253.075 53.605 ;
      END
   END dout1[31]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met3 ;
         RECT  7.42 7.42 391.9 10.3 ;
         LAYER met4 ;
         RECT  389.02 7.42 391.9 559.38 ;
         LAYER met3 ;
         RECT  7.42 556.5 391.9 559.38 ;
         LAYER met4 ;
         RECT  7.42 7.42 10.3 559.38 ;
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met3 ;
         RECT  2.12 2.12 397.2 5.0 ;
         LAYER met4 ;
         RECT  2.12 2.12 5.0 564.68 ;
         LAYER met3 ;
         RECT  2.12 561.8 397.2 564.68 ;
         LAYER met4 ;
         RECT  394.32 2.12 397.2 564.68 ;
      END
   END gnd
   OBS
   LAYER  met1 ;
      RECT  0.62 0.62 396.58 564.06 ;
   LAYER  met2 ;
      RECT  0.62 0.62 396.58 564.06 ;
   LAYER  met3 ;
      RECT  15.025 37.295 396.58 38.865 ;
      RECT  13.165 32.945 15.025 37.295 ;
      RECT  2.42 35.44 13.165 37.295 ;
      RECT  0.62 37.4 2.42 38.865 ;
      RECT  2.42 37.295 13.165 37.4 ;
      RECT  2.42 37.4 13.165 38.865 ;
      RECT  15.025 38.865 133.755 52.635 ;
      RECT  15.025 52.635 133.755 54.205 ;
      RECT  133.755 38.865 135.615 52.635 ;
      RECT  135.615 38.865 396.58 52.635 ;
      RECT  136.975 52.635 141.535 54.205 ;
      RECT  144.755 52.635 149.315 54.205 ;
      RECT  152.535 52.635 157.095 54.205 ;
      RECT  160.315 52.635 164.875 54.205 ;
      RECT  168.095 52.635 172.655 54.205 ;
      RECT  175.875 52.635 180.435 54.205 ;
      RECT  183.655 52.635 188.215 54.205 ;
      RECT  191.435 52.635 195.995 54.205 ;
      RECT  199.215 52.635 203.775 54.205 ;
      RECT  206.995 52.635 211.555 54.205 ;
      RECT  214.775 52.635 219.335 54.205 ;
      RECT  222.555 52.635 227.115 54.205 ;
      RECT  230.335 52.635 234.895 54.205 ;
      RECT  238.115 52.635 242.675 54.205 ;
      RECT  245.895 52.635 250.455 54.205 ;
      RECT  253.675 52.635 396.58 54.205 ;
      RECT  15.025 10.9 392.5 37.295 ;
      RECT  392.5 6.82 396.58 10.9 ;
      RECT  392.5 10.9 396.58 37.295 ;
      RECT  13.165 10.9 15.025 31.375 ;
      RECT  2.42 6.82 6.82 10.9 ;
      RECT  2.42 10.9 6.82 35.44 ;
      RECT  6.82 10.9 13.165 35.44 ;
      RECT  0.62 38.865 6.82 555.9 ;
      RECT  0.62 555.9 6.82 559.98 ;
      RECT  6.82 38.865 13.165 555.9 ;
      RECT  13.165 38.865 15.025 555.9 ;
      RECT  15.025 54.205 133.755 555.9 ;
      RECT  133.755 54.205 135.615 555.9 ;
      RECT  135.615 54.205 392.5 555.9 ;
      RECT  392.5 54.205 396.58 555.9 ;
      RECT  392.5 555.9 396.58 559.98 ;
      RECT  0.62 0.62 1.52 1.52 ;
      RECT  0.62 1.52 1.52 5.6 ;
      RECT  0.62 5.6 1.52 35.44 ;
      RECT  1.52 0.62 2.42 1.52 ;
      RECT  1.52 5.6 2.42 35.44 ;
      RECT  15.025 0.62 392.5 1.52 ;
      RECT  15.025 5.6 392.5 6.82 ;
      RECT  392.5 0.62 396.58 1.52 ;
      RECT  392.5 5.6 396.58 6.82 ;
      RECT  13.165 0.62 15.025 1.52 ;
      RECT  13.165 5.6 15.025 6.82 ;
      RECT  2.42 0.62 6.82 1.52 ;
      RECT  2.42 5.6 6.82 6.82 ;
      RECT  6.82 0.62 13.165 1.52 ;
      RECT  6.82 5.6 13.165 6.82 ;
      RECT  0.62 559.98 1.52 561.2 ;
      RECT  0.62 561.2 1.52 564.06 ;
      RECT  1.52 559.98 6.82 561.2 ;
      RECT  6.82 559.98 13.165 561.2 ;
      RECT  13.165 559.98 15.025 561.2 ;
      RECT  15.025 559.98 133.755 561.2 ;
      RECT  133.755 559.98 135.615 561.2 ;
      RECT  135.615 559.98 392.5 561.2 ;
      RECT  392.5 559.98 396.58 561.2 ;
   LAYER  met4 ;
      RECT  105.4 2.42 107.36 564.06 ;
      RECT  107.36 0.62 112.82 2.42 ;
      RECT  114.78 0.62 120.24 2.42 ;
      RECT  122.2 0.62 127.66 2.42 ;
      RECT  255.76 0.62 261.22 2.42 ;
      RECT  263.18 0.62 268.64 2.42 ;
      RECT  270.6 0.62 276.06 2.42 ;
      RECT  278.02 0.62 283.48 2.42 ;
      RECT  285.44 0.62 289.84 2.42 ;
      RECT  291.8 0.62 298.32 2.42 ;
      RECT  300.28 0.62 305.74 2.42 ;
      RECT  307.7 0.62 312.1 2.42 ;
      RECT  314.06 0.62 320.58 2.42 ;
      RECT  322.54 0.62 328.0 2.42 ;
      RECT  329.96 0.62 335.42 2.42 ;
      RECT  129.62 0.62 134.02 2.42 ;
      RECT  138.1 0.62 141.44 2.42 ;
      RECT  145.52 0.62 148.86 2.42 ;
      RECT  152.94 0.62 157.34 2.42 ;
      RECT  161.42 0.62 164.76 2.42 ;
      RECT  168.84 0.62 172.18 2.42 ;
      RECT  176.26 0.62 179.6 2.42 ;
      RECT  183.68 0.62 188.08 2.42 ;
      RECT  192.16 0.62 195.5 2.42 ;
      RECT  199.58 0.62 201.86 2.42 ;
      RECT  204.88 0.62 205.04 2.42 ;
      RECT  207.0 0.62 209.28 2.42 ;
      RECT  211.24 0.62 211.4 2.42 ;
      RECT  214.42 0.62 216.7 2.42 ;
      RECT  218.66 0.62 219.88 2.42 ;
      RECT  222.9 0.62 224.12 2.42 ;
      RECT  226.08 0.62 226.24 2.42 ;
      RECT  228.2 0.62 229.42 2.42 ;
      RECT  231.38 0.62 231.54 2.42 ;
      RECT  233.5 0.62 234.72 2.42 ;
      RECT  237.74 0.62 238.96 2.42 ;
      RECT  240.92 0.62 243.2 2.42 ;
      RECT  246.22 0.62 246.38 2.42 ;
      RECT  248.34 0.62 249.56 2.42 ;
      RECT  251.52 0.62 251.68 2.42 ;
      RECT  253.64 0.62 253.8 2.42 ;
      RECT  107.36 2.42 388.42 6.82 ;
      RECT  107.36 6.82 388.42 559.98 ;
      RECT  107.36 559.98 388.42 564.06 ;
      RECT  388.42 2.42 392.5 6.82 ;
      RECT  388.42 559.98 392.5 564.06 ;
      RECT  6.82 2.42 10.9 6.82 ;
      RECT  6.82 559.98 10.9 564.06 ;
      RECT  10.9 2.42 105.4 6.82 ;
      RECT  10.9 6.82 105.4 559.98 ;
      RECT  10.9 559.98 105.4 564.06 ;
      RECT  0.62 0.62 1.52 1.52 ;
      RECT  0.62 1.52 1.52 2.42 ;
      RECT  1.52 0.62 5.6 1.52 ;
      RECT  5.6 0.62 105.4 1.52 ;
      RECT  5.6 1.52 105.4 2.42 ;
      RECT  0.62 2.42 1.52 6.82 ;
      RECT  5.6 2.42 6.82 6.82 ;
      RECT  0.62 6.82 1.52 559.98 ;
      RECT  5.6 6.82 6.82 559.98 ;
      RECT  0.62 559.98 1.52 564.06 ;
      RECT  5.6 559.98 6.82 564.06 ;
      RECT  337.38 0.62 393.72 1.52 ;
      RECT  337.38 1.52 393.72 2.42 ;
      RECT  393.72 0.62 396.58 1.52 ;
      RECT  392.5 2.42 393.72 6.82 ;
      RECT  392.5 6.82 393.72 559.98 ;
      RECT  392.5 559.98 393.72 564.06 ;
   END
END    sram_0rw2r1w_32_128_sky130A
END    LIBRARY
