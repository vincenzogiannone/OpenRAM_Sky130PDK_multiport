magic
tech sky130A
magscale 1 2
timestamp 1643593061
<< checkpaint >>
rect -1260 -1302 6486 25922
<< viali >>
rect 2422 23887 2456 23921
rect 2422 22263 2456 22297
rect 2422 20807 2456 20841
rect 2422 19183 2456 19217
rect 2422 14651 2456 14685
rect 2422 13027 2456 13061
rect 2422 11571 2456 11605
rect 2422 9947 2456 9981
rect 2422 5415 2456 5449
rect 2422 3791 2456 3825
rect 2422 2335 2456 2369
rect 2422 711 2456 745
<< metal1 >>
rect 5162 24198 5168 24250
rect 5220 24198 5226 24250
rect 2407 23878 2413 23930
rect 2465 23878 2471 23930
rect 3500 23718 3506 23770
rect 3558 23758 3564 23770
rect 3558 23730 4674 23758
rect 3558 23718 3564 23730
rect 3248 23662 3254 23714
rect 3306 23702 3312 23714
rect 3306 23674 4578 23702
rect 3306 23662 3312 23674
rect 2828 23606 2834 23658
rect 2886 23646 2892 23658
rect 2886 23618 4482 23646
rect 2886 23606 2892 23618
rect 4814 23616 5180 23644
rect 3500 23550 3506 23602
rect 3558 23590 3564 23602
rect 3558 23562 4278 23590
rect 3558 23550 3564 23562
rect 3248 23494 3254 23546
rect 3306 23534 3312 23546
rect 3306 23506 4182 23534
rect 3306 23494 3312 23506
rect 4896 23494 5180 23522
rect 2744 23438 2750 23490
rect 2802 23478 2808 23490
rect 2802 23450 4086 23478
rect 2802 23438 2808 23450
rect 3500 23382 3506 23434
rect 3558 23422 3564 23434
rect 3558 23394 3990 23422
rect 3558 23382 3564 23394
rect 3248 23326 3254 23378
rect 3306 23366 3312 23378
rect 3306 23338 3894 23366
rect 5104 23348 5180 23376
rect 3306 23326 3312 23338
rect 2660 23270 2666 23322
rect 2718 23310 2724 23322
rect 2718 23282 3798 23310
rect 2718 23270 2724 23282
rect 5162 22684 5168 22736
rect 5220 22684 5226 22736
rect 2407 22254 2413 22306
rect 2465 22254 2471 22306
rect 2744 22098 2750 22150
rect 2802 22138 2808 22150
rect 2802 22110 3798 22138
rect 2802 22098 2808 22110
rect 3164 22042 3170 22094
rect 3222 22082 3228 22094
rect 3222 22054 3894 22082
rect 3222 22042 3228 22054
rect 5104 22044 5180 22072
rect 3500 21986 3506 22038
rect 3558 22026 3564 22038
rect 3558 21998 3990 22026
rect 3558 21986 3564 21998
rect 2828 21930 2834 21982
rect 2886 21970 2892 21982
rect 2886 21942 4086 21970
rect 2886 21930 2892 21942
rect 3164 21874 3170 21926
rect 3222 21914 3228 21926
rect 3222 21886 4182 21914
rect 4896 21898 5180 21926
rect 3222 21874 3228 21886
rect 3500 21818 3506 21870
rect 3558 21858 3564 21870
rect 3558 21830 4278 21858
rect 3558 21818 3564 21830
rect 2912 21762 2918 21814
rect 2970 21802 2976 21814
rect 2970 21774 4482 21802
rect 4814 21776 5180 21804
rect 2970 21762 2976 21774
rect 3164 21706 3170 21758
rect 3222 21746 3228 21758
rect 3222 21718 4578 21746
rect 3222 21706 3228 21718
rect 3500 21650 3506 21702
rect 3558 21690 3564 21702
rect 3558 21662 4674 21690
rect 3558 21650 3564 21662
rect 5162 21170 5168 21222
rect 5220 21170 5226 21222
rect 420 20798 426 20850
rect 478 20838 484 20850
rect 700 20838 706 20850
rect 478 20810 706 20838
rect 478 20798 484 20810
rect 700 20798 706 20810
rect 758 20798 764 20850
rect 2407 20798 2413 20850
rect 2465 20798 2471 20850
rect 3500 20690 3506 20742
rect 3558 20730 3564 20742
rect 3558 20702 4674 20730
rect 3558 20690 3564 20702
rect 3164 20634 3170 20686
rect 3222 20674 3228 20686
rect 3222 20646 4578 20674
rect 3222 20634 3228 20646
rect 2660 20578 2666 20630
rect 2718 20618 2724 20630
rect 2718 20590 4482 20618
rect 2718 20578 2724 20590
rect 4814 20588 5180 20616
rect 3500 20522 3506 20574
rect 3558 20562 3564 20574
rect 3558 20534 4278 20562
rect 3558 20522 3564 20534
rect 3080 20466 3086 20518
rect 3138 20506 3144 20518
rect 3138 20478 4182 20506
rect 3138 20466 3144 20478
rect 4896 20466 5180 20494
rect 2912 20410 2918 20462
rect 2970 20450 2976 20462
rect 2970 20422 4086 20450
rect 2970 20410 2976 20422
rect 3500 20354 3506 20406
rect 3558 20394 3564 20406
rect 3558 20366 3990 20394
rect 3558 20354 3564 20366
rect 3080 20298 3086 20350
rect 3138 20338 3144 20350
rect 3138 20310 3894 20338
rect 5104 20320 5180 20348
rect 3138 20298 3144 20310
rect 2828 20242 2834 20294
rect 2886 20282 2892 20294
rect 2886 20254 3798 20282
rect 2886 20242 2892 20254
rect 5162 19656 5168 19708
rect 5220 19656 5226 19708
rect 336 19174 342 19226
rect 394 19214 400 19226
rect 616 19214 622 19226
rect 394 19186 622 19214
rect 394 19174 400 19186
rect 616 19174 622 19186
rect 674 19174 680 19226
rect 2407 19174 2413 19226
rect 2465 19174 2471 19226
rect 2912 19070 2918 19122
rect 2970 19110 2976 19122
rect 2970 19082 3798 19110
rect 2970 19070 2976 19082
rect 2996 19014 3002 19066
rect 3054 19054 3060 19066
rect 3054 19026 3894 19054
rect 3054 19014 3060 19026
rect 5104 19016 5180 19044
rect 3500 18958 3506 19010
rect 3558 18998 3564 19010
rect 3558 18970 3990 18998
rect 3558 18958 3564 18970
rect 2660 18902 2666 18954
rect 2718 18942 2724 18954
rect 2718 18914 4086 18942
rect 2718 18902 2724 18914
rect 3080 18846 3086 18898
rect 3138 18886 3144 18898
rect 3138 18858 4182 18886
rect 4896 18870 5180 18898
rect 3138 18846 3144 18858
rect 3500 18790 3506 18842
rect 3558 18830 3564 18842
rect 3558 18802 4278 18830
rect 3558 18790 3564 18802
rect 2744 18734 2750 18786
rect 2802 18774 2808 18786
rect 2802 18746 4482 18774
rect 4814 18748 5180 18776
rect 2802 18734 2808 18746
rect 3080 18678 3086 18730
rect 3138 18718 3144 18730
rect 3138 18690 4578 18718
rect 3138 18678 3144 18690
rect 3500 18622 3506 18674
rect 3558 18662 3564 18674
rect 3558 18634 4674 18662
rect 3558 18622 3564 18634
rect 5162 18142 5168 18194
rect 5220 18142 5226 18194
rect 3500 17662 3506 17714
rect 3558 17702 3564 17714
rect 3558 17674 4674 17702
rect 3558 17662 3564 17674
rect 2996 17606 3002 17658
rect 3054 17646 3060 17658
rect 3054 17618 4578 17646
rect 3054 17606 3060 17618
rect 2828 17550 2834 17602
rect 2886 17590 2892 17602
rect 2886 17562 4482 17590
rect 2886 17550 2892 17562
rect 4814 17560 5180 17588
rect 3500 17494 3506 17546
rect 3558 17534 3564 17546
rect 3558 17506 4278 17534
rect 3558 17494 3564 17506
rect 2996 17438 3002 17490
rect 3054 17478 3060 17490
rect 3054 17450 4182 17478
rect 3054 17438 3060 17450
rect 4896 17438 5180 17466
rect 2744 17382 2750 17434
rect 2802 17422 2808 17434
rect 2802 17394 4086 17422
rect 2802 17382 2808 17394
rect 3500 17326 3506 17378
rect 3558 17366 3564 17378
rect 3558 17338 3990 17366
rect 3558 17326 3564 17338
rect 2996 17270 3002 17322
rect 3054 17310 3060 17322
rect 3054 17282 3894 17310
rect 5104 17292 5180 17320
rect 3054 17270 3060 17282
rect 2660 17214 2666 17266
rect 2718 17254 2724 17266
rect 2718 17226 3798 17254
rect 2718 17214 2724 17226
rect 5162 16628 5168 16680
rect 5220 16628 5226 16680
rect 2744 16042 2750 16094
rect 2802 16082 2808 16094
rect 2802 16054 3798 16082
rect 2802 16042 2808 16054
rect 3248 15986 3254 16038
rect 3306 16026 3312 16038
rect 3306 15998 3894 16026
rect 3306 15986 3312 15998
rect 5104 15988 5180 16016
rect 3416 15930 3422 15982
rect 3474 15970 3480 15982
rect 3474 15942 3990 15970
rect 3474 15930 3480 15942
rect 2828 15874 2834 15926
rect 2886 15914 2892 15926
rect 2886 15886 4086 15914
rect 2886 15874 2892 15886
rect 3248 15818 3254 15870
rect 3306 15858 3312 15870
rect 3306 15830 4182 15858
rect 4896 15842 5180 15870
rect 3306 15818 3312 15830
rect 3416 15762 3422 15814
rect 3474 15802 3480 15814
rect 3474 15774 4278 15802
rect 3474 15762 3480 15774
rect 2912 15706 2918 15758
rect 2970 15746 2976 15758
rect 2970 15718 4482 15746
rect 4814 15720 5180 15748
rect 2970 15706 2976 15718
rect 3248 15650 3254 15702
rect 3306 15690 3312 15702
rect 3306 15662 4578 15690
rect 3306 15650 3312 15662
rect 3416 15594 3422 15646
rect 3474 15634 3480 15646
rect 3474 15606 4674 15634
rect 3474 15594 3480 15606
rect 5162 15114 5168 15166
rect 5220 15114 5226 15166
rect 2407 14642 2413 14694
rect 2465 14642 2471 14694
rect 3416 14634 3422 14686
rect 3474 14674 3480 14686
rect 3474 14646 4674 14674
rect 3474 14634 3480 14646
rect 3248 14578 3254 14630
rect 3306 14618 3312 14630
rect 3306 14590 4578 14618
rect 3306 14578 3312 14590
rect 2660 14522 2666 14574
rect 2718 14562 2724 14574
rect 2718 14534 4482 14562
rect 2718 14522 2724 14534
rect 4814 14532 5180 14560
rect 3416 14466 3422 14518
rect 3474 14506 3480 14518
rect 3474 14478 4278 14506
rect 3474 14466 3480 14478
rect 3164 14410 3170 14462
rect 3222 14450 3228 14462
rect 3222 14422 4182 14450
rect 3222 14410 3228 14422
rect 4896 14410 5180 14438
rect 2912 14354 2918 14406
rect 2970 14394 2976 14406
rect 2970 14366 4086 14394
rect 2970 14354 2976 14366
rect 3416 14298 3422 14350
rect 3474 14338 3480 14350
rect 3474 14310 3990 14338
rect 3474 14298 3480 14310
rect 3164 14242 3170 14294
rect 3222 14282 3228 14294
rect 3222 14254 3894 14282
rect 5104 14264 5180 14292
rect 3222 14242 3228 14254
rect 2828 14186 2834 14238
rect 2886 14226 2892 14238
rect 2886 14198 3798 14226
rect 2886 14186 2892 14198
rect 5162 13600 5168 13652
rect 5220 13600 5226 13652
rect 2407 13018 2413 13070
rect 2465 13018 2471 13070
rect 2912 13014 2918 13066
rect 2970 13054 2976 13066
rect 2970 13026 3798 13054
rect 2970 13014 2976 13026
rect 3080 12958 3086 13010
rect 3138 12998 3144 13010
rect 3138 12970 3894 12998
rect 3138 12958 3144 12970
rect 5104 12960 5180 12988
rect 3416 12902 3422 12954
rect 3474 12942 3480 12954
rect 3474 12914 3990 12942
rect 3474 12902 3480 12914
rect 2660 12846 2666 12898
rect 2718 12886 2724 12898
rect 2718 12858 4086 12886
rect 2718 12846 2724 12858
rect 3164 12790 3170 12842
rect 3222 12830 3228 12842
rect 3222 12802 4182 12830
rect 4896 12814 5180 12842
rect 3222 12790 3228 12802
rect 3416 12734 3422 12786
rect 3474 12774 3480 12786
rect 3474 12746 4278 12774
rect 3474 12734 3480 12746
rect 2744 12678 2750 12730
rect 2802 12718 2808 12730
rect 2802 12690 4482 12718
rect 4814 12692 5180 12720
rect 2802 12678 2808 12690
rect 3164 12622 3170 12674
rect 3222 12662 3228 12674
rect 3222 12634 4578 12662
rect 3222 12622 3228 12634
rect 3416 12566 3422 12618
rect 3474 12606 3480 12618
rect 3474 12578 4674 12606
rect 3474 12566 3480 12578
rect 5162 12086 5168 12138
rect 5220 12086 5226 12138
rect 252 11562 258 11614
rect 310 11602 316 11614
rect 700 11602 706 11614
rect 310 11574 706 11602
rect 310 11562 316 11574
rect 700 11562 706 11574
rect 758 11562 764 11614
rect 2407 11562 2413 11614
rect 2465 11562 2471 11614
rect 3416 11606 3422 11658
rect 3474 11646 3480 11658
rect 3474 11618 4674 11646
rect 3474 11606 3480 11618
rect 3080 11550 3086 11602
rect 3138 11590 3144 11602
rect 3138 11562 4578 11590
rect 3138 11550 3144 11562
rect 2828 11494 2834 11546
rect 2886 11534 2892 11546
rect 2886 11506 4482 11534
rect 2886 11494 2892 11506
rect 4814 11504 5180 11532
rect 3416 11438 3422 11490
rect 3474 11478 3480 11490
rect 3474 11450 4278 11478
rect 3474 11438 3480 11450
rect 3080 11382 3086 11434
rect 3138 11422 3144 11434
rect 3138 11394 4182 11422
rect 3138 11382 3144 11394
rect 4896 11382 5180 11410
rect 2744 11326 2750 11378
rect 2802 11366 2808 11378
rect 2802 11338 4086 11366
rect 2802 11326 2808 11338
rect 3416 11270 3422 11322
rect 3474 11310 3480 11322
rect 3474 11282 3990 11310
rect 3474 11270 3480 11282
rect 3080 11214 3086 11266
rect 3138 11254 3144 11266
rect 3138 11226 3894 11254
rect 5104 11236 5180 11264
rect 3138 11214 3144 11226
rect 2660 11158 2666 11210
rect 2718 11198 2724 11210
rect 2718 11170 3798 11198
rect 2718 11158 2724 11170
rect 5162 10572 5168 10624
rect 5220 10572 5226 10624
rect 168 9938 174 9990
rect 226 9978 232 9990
rect 616 9978 622 9990
rect 226 9950 622 9978
rect 226 9938 232 9950
rect 616 9938 622 9950
rect 674 9938 680 9990
rect 2407 9938 2413 9990
rect 2465 9938 2471 9990
rect 2744 9986 2750 10038
rect 2802 10026 2808 10038
rect 2802 9998 3798 10026
rect 2802 9986 2808 9998
rect 2996 9930 3002 9982
rect 3054 9970 3060 9982
rect 3054 9942 3894 9970
rect 3054 9930 3060 9942
rect 5104 9932 5180 9960
rect 3416 9874 3422 9926
rect 3474 9914 3480 9926
rect 3474 9886 3990 9914
rect 3474 9874 3480 9886
rect 2828 9818 2834 9870
rect 2886 9858 2892 9870
rect 2886 9830 4086 9858
rect 2886 9818 2892 9830
rect 2996 9762 3002 9814
rect 3054 9802 3060 9814
rect 3054 9774 4182 9802
rect 4896 9786 5180 9814
rect 3054 9762 3060 9774
rect 3416 9706 3422 9758
rect 3474 9746 3480 9758
rect 3474 9718 4278 9746
rect 3474 9706 3480 9718
rect 2912 9650 2918 9702
rect 2970 9690 2976 9702
rect 2970 9662 4482 9690
rect 4814 9664 5180 9692
rect 2970 9650 2976 9662
rect 2996 9594 3002 9646
rect 3054 9634 3060 9646
rect 3054 9606 4578 9634
rect 3054 9594 3060 9606
rect 3416 9538 3422 9590
rect 3474 9578 3480 9590
rect 3474 9550 4674 9578
rect 3474 9538 3480 9550
rect 5162 9058 5168 9110
rect 5220 9058 5226 9110
rect 3416 8578 3422 8630
rect 3474 8618 3480 8630
rect 3474 8590 4674 8618
rect 3474 8578 3480 8590
rect 2996 8522 3002 8574
rect 3054 8562 3060 8574
rect 3054 8534 4578 8562
rect 3054 8522 3060 8534
rect 2660 8466 2666 8518
rect 2718 8506 2724 8518
rect 2718 8478 4482 8506
rect 2718 8466 2724 8478
rect 4814 8476 5180 8504
rect 3332 8410 3338 8462
rect 3390 8450 3396 8462
rect 3390 8422 4278 8450
rect 3390 8410 3396 8422
rect 3248 8354 3254 8406
rect 3306 8394 3312 8406
rect 3306 8366 4182 8394
rect 3306 8354 3312 8366
rect 4896 8354 5180 8382
rect 2912 8298 2918 8350
rect 2970 8338 2976 8350
rect 2970 8310 4086 8338
rect 2970 8298 2976 8310
rect 3332 8242 3338 8294
rect 3390 8282 3396 8294
rect 3390 8254 3990 8282
rect 3390 8242 3396 8254
rect 3248 8186 3254 8238
rect 3306 8226 3312 8238
rect 3306 8198 3894 8226
rect 5104 8208 5180 8236
rect 3306 8186 3312 8198
rect 2828 8130 2834 8182
rect 2886 8170 2892 8182
rect 2886 8142 3798 8170
rect 2886 8130 2892 8142
rect 5162 7544 5168 7596
rect 5220 7544 5226 7596
rect 2912 6958 2918 7010
rect 2970 6998 2976 7010
rect 2970 6970 3798 6998
rect 2970 6958 2976 6970
rect 3164 6902 3170 6954
rect 3222 6942 3228 6954
rect 3222 6914 3894 6942
rect 3222 6902 3228 6914
rect 5104 6904 5180 6932
rect 3332 6846 3338 6898
rect 3390 6886 3396 6898
rect 3390 6858 3990 6886
rect 3390 6846 3396 6858
rect 2660 6790 2666 6842
rect 2718 6830 2724 6842
rect 2718 6802 4086 6830
rect 2718 6790 2724 6802
rect 3248 6734 3254 6786
rect 3306 6774 3312 6786
rect 3306 6746 4182 6774
rect 4896 6758 5180 6786
rect 3306 6734 3312 6746
rect 3332 6678 3338 6730
rect 3390 6718 3396 6730
rect 3390 6690 4278 6718
rect 3390 6678 3396 6690
rect 2744 6622 2750 6674
rect 2802 6662 2808 6674
rect 2802 6634 4482 6662
rect 4814 6636 5180 6664
rect 2802 6622 2808 6634
rect 3248 6566 3254 6618
rect 3306 6606 3312 6618
rect 3306 6578 4578 6606
rect 3306 6566 3312 6578
rect 3332 6510 3338 6562
rect 3390 6550 3396 6562
rect 3390 6522 4674 6550
rect 3390 6510 3396 6522
rect 5162 6030 5168 6082
rect 5220 6030 5226 6082
rect 3332 5550 3338 5602
rect 3390 5590 3396 5602
rect 3390 5562 4674 5590
rect 3390 5550 3396 5562
rect 3164 5494 3170 5546
rect 3222 5534 3228 5546
rect 3222 5506 4578 5534
rect 3222 5494 3228 5506
rect 2407 5406 2413 5458
rect 2465 5406 2471 5458
rect 2828 5438 2834 5490
rect 2886 5478 2892 5490
rect 2886 5450 4482 5478
rect 2886 5438 2892 5450
rect 4814 5448 5180 5476
rect 3332 5382 3338 5434
rect 3390 5422 3396 5434
rect 3390 5394 4278 5422
rect 3390 5382 3396 5394
rect 3164 5326 3170 5378
rect 3222 5366 3228 5378
rect 3222 5338 4182 5366
rect 3222 5326 3228 5338
rect 4896 5326 5180 5354
rect 2744 5270 2750 5322
rect 2802 5310 2808 5322
rect 2802 5282 4086 5310
rect 2802 5270 2808 5282
rect 3332 5214 3338 5266
rect 3390 5254 3396 5266
rect 3390 5226 3990 5254
rect 3390 5214 3396 5226
rect 3164 5158 3170 5210
rect 3222 5198 3228 5210
rect 3222 5170 3894 5198
rect 5104 5180 5180 5208
rect 3222 5158 3228 5170
rect 2660 5102 2666 5154
rect 2718 5142 2724 5154
rect 2718 5114 3798 5142
rect 2718 5102 2724 5114
rect 5162 4516 5168 4568
rect 5220 4516 5226 4568
rect 2744 3930 2750 3982
rect 2802 3970 2808 3982
rect 2802 3942 3798 3970
rect 2802 3930 2808 3942
rect 3080 3874 3086 3926
rect 3138 3914 3144 3926
rect 3138 3886 3894 3914
rect 3138 3874 3144 3886
rect 5104 3876 5180 3904
rect 2407 3782 2413 3834
rect 2465 3782 2471 3834
rect 3332 3818 3338 3870
rect 3390 3858 3396 3870
rect 3390 3830 3990 3858
rect 3390 3818 3396 3830
rect 2828 3762 2834 3814
rect 2886 3802 2892 3814
rect 2886 3774 4086 3802
rect 2886 3762 2892 3774
rect 3080 3706 3086 3758
rect 3138 3746 3144 3758
rect 3138 3718 4182 3746
rect 4896 3730 5180 3758
rect 3138 3706 3144 3718
rect 3332 3650 3338 3702
rect 3390 3690 3396 3702
rect 3390 3662 4278 3690
rect 3390 3650 3396 3662
rect 2912 3594 2918 3646
rect 2970 3634 2976 3646
rect 2970 3606 4482 3634
rect 4814 3608 5180 3636
rect 2970 3594 2976 3606
rect 3080 3538 3086 3590
rect 3138 3578 3144 3590
rect 3138 3550 4578 3578
rect 3138 3538 3144 3550
rect 3332 3482 3338 3534
rect 3390 3522 3396 3534
rect 3390 3494 4674 3522
rect 3390 3482 3396 3494
rect 5162 3002 5168 3054
rect 5220 3002 5226 3054
rect 3332 2522 3338 2574
rect 3390 2562 3396 2574
rect 3390 2534 4674 2562
rect 3390 2522 3396 2534
rect 3080 2466 3086 2518
rect 3138 2506 3144 2518
rect 3138 2478 4578 2506
rect 3138 2466 3144 2478
rect 2660 2410 2666 2462
rect 2718 2450 2724 2462
rect 2718 2422 4482 2450
rect 2718 2410 2724 2422
rect 4814 2420 5180 2448
rect 84 2326 90 2378
rect 142 2366 148 2378
rect 700 2366 706 2378
rect 142 2338 706 2366
rect 142 2326 148 2338
rect 700 2326 706 2338
rect 758 2326 764 2378
rect 2407 2326 2413 2378
rect 2465 2326 2471 2378
rect 3332 2354 3338 2406
rect 3390 2394 3396 2406
rect 3390 2366 4278 2394
rect 3390 2354 3396 2366
rect 2996 2298 3002 2350
rect 3054 2338 3060 2350
rect 3054 2310 4182 2338
rect 3054 2298 3060 2310
rect 4896 2298 5180 2326
rect 2912 2242 2918 2294
rect 2970 2282 2976 2294
rect 2970 2254 4086 2282
rect 2970 2242 2976 2254
rect 3332 2186 3338 2238
rect 3390 2226 3396 2238
rect 3390 2198 3990 2226
rect 3390 2186 3396 2198
rect 2996 2130 3002 2182
rect 3054 2170 3060 2182
rect 3054 2142 3894 2170
rect 5104 2152 5180 2180
rect 3054 2130 3060 2142
rect 2828 2074 2834 2126
rect 2886 2114 2892 2126
rect 2886 2086 3798 2114
rect 2886 2074 2892 2086
rect 5162 1488 5168 1540
rect 5220 1488 5226 1540
rect 2912 942 2918 954
rect 2678 914 2918 942
rect 2912 902 2918 914
rect 2970 902 2976 954
rect 3248 886 3254 898
rect 2774 858 3254 886
rect 3248 846 3254 858
rect 3306 846 3312 898
rect 5104 848 5180 876
rect 3500 830 3506 842
rect 2870 802 3506 830
rect 3500 790 3506 802
rect 3558 790 3564 842
rect 0 702 6 754
rect 58 742 64 754
rect 616 742 622 754
rect 58 714 622 742
rect 58 702 64 714
rect 616 702 622 714
rect 674 702 680 754
rect 2407 702 2413 754
rect 2465 702 2471 754
rect 2660 734 2666 786
rect 2718 774 2724 786
rect 2718 746 4086 774
rect 2718 734 2724 746
rect 2996 678 3002 730
rect 3054 718 3060 730
rect 3054 690 4182 718
rect 4896 702 5180 730
rect 3054 678 3060 690
rect 3332 622 3338 674
rect 3390 662 3396 674
rect 3390 634 4278 662
rect 3390 622 3396 634
rect 2744 566 2750 618
rect 2802 606 2808 618
rect 2802 578 4482 606
rect 4814 580 5180 608
rect 2802 566 2808 578
rect 2996 510 3002 562
rect 3054 550 3060 562
rect 3054 522 4578 550
rect 3054 510 3060 522
rect 3332 454 3338 506
rect 3390 494 3396 506
rect 3390 466 4674 494
rect 3390 454 3396 466
rect 5162 -26 5168 26
rect 5220 -26 5226 26
<< via1 >>
rect 5168 24198 5220 24250
rect 2413 23921 2465 23930
rect 2413 23887 2422 23921
rect 2422 23887 2456 23921
rect 2456 23887 2465 23921
rect 2413 23878 2465 23887
rect 3506 23718 3558 23770
rect 3254 23662 3306 23714
rect 2834 23606 2886 23658
rect 3506 23550 3558 23602
rect 3254 23494 3306 23546
rect 2750 23438 2802 23490
rect 3506 23382 3558 23434
rect 3254 23326 3306 23378
rect 2666 23270 2718 23322
rect 5168 22684 5220 22736
rect 2413 22297 2465 22306
rect 2413 22263 2422 22297
rect 2422 22263 2456 22297
rect 2456 22263 2465 22297
rect 2413 22254 2465 22263
rect 2750 22098 2802 22150
rect 3170 22042 3222 22094
rect 3506 21986 3558 22038
rect 2834 21930 2886 21982
rect 3170 21874 3222 21926
rect 3506 21818 3558 21870
rect 2918 21762 2970 21814
rect 3170 21706 3222 21758
rect 3506 21650 3558 21702
rect 5168 21170 5220 21222
rect 426 20798 478 20850
rect 706 20798 758 20850
rect 2413 20841 2465 20850
rect 2413 20807 2422 20841
rect 2422 20807 2456 20841
rect 2456 20807 2465 20841
rect 2413 20798 2465 20807
rect 3506 20690 3558 20742
rect 3170 20634 3222 20686
rect 2666 20578 2718 20630
rect 3506 20522 3558 20574
rect 3086 20466 3138 20518
rect 2918 20410 2970 20462
rect 3506 20354 3558 20406
rect 3086 20298 3138 20350
rect 2834 20242 2886 20294
rect 5168 19656 5220 19708
rect 342 19174 394 19226
rect 622 19174 674 19226
rect 2413 19217 2465 19226
rect 2413 19183 2422 19217
rect 2422 19183 2456 19217
rect 2456 19183 2465 19217
rect 2413 19174 2465 19183
rect 2918 19070 2970 19122
rect 3002 19014 3054 19066
rect 3506 18958 3558 19010
rect 2666 18902 2718 18954
rect 3086 18846 3138 18898
rect 3506 18790 3558 18842
rect 2750 18734 2802 18786
rect 3086 18678 3138 18730
rect 3506 18622 3558 18674
rect 5168 18142 5220 18194
rect 3506 17662 3558 17714
rect 3002 17606 3054 17658
rect 2834 17550 2886 17602
rect 3506 17494 3558 17546
rect 3002 17438 3054 17490
rect 2750 17382 2802 17434
rect 3506 17326 3558 17378
rect 3002 17270 3054 17322
rect 2666 17214 2718 17266
rect 5168 16628 5220 16680
rect 2750 16042 2802 16094
rect 3254 15986 3306 16038
rect 3422 15930 3474 15982
rect 2834 15874 2886 15926
rect 3254 15818 3306 15870
rect 3422 15762 3474 15814
rect 2918 15706 2970 15758
rect 3254 15650 3306 15702
rect 3422 15594 3474 15646
rect 5168 15114 5220 15166
rect 2413 14685 2465 14694
rect 2413 14651 2422 14685
rect 2422 14651 2456 14685
rect 2456 14651 2465 14685
rect 2413 14642 2465 14651
rect 3422 14634 3474 14686
rect 3254 14578 3306 14630
rect 2666 14522 2718 14574
rect 3422 14466 3474 14518
rect 3170 14410 3222 14462
rect 2918 14354 2970 14406
rect 3422 14298 3474 14350
rect 3170 14242 3222 14294
rect 2834 14186 2886 14238
rect 5168 13600 5220 13652
rect 2413 13061 2465 13070
rect 2413 13027 2422 13061
rect 2422 13027 2456 13061
rect 2456 13027 2465 13061
rect 2413 13018 2465 13027
rect 2918 13014 2970 13066
rect 3086 12958 3138 13010
rect 3422 12902 3474 12954
rect 2666 12846 2718 12898
rect 3170 12790 3222 12842
rect 3422 12734 3474 12786
rect 2750 12678 2802 12730
rect 3170 12622 3222 12674
rect 3422 12566 3474 12618
rect 5168 12086 5220 12138
rect 258 11562 310 11614
rect 706 11562 758 11614
rect 2413 11605 2465 11614
rect 2413 11571 2422 11605
rect 2422 11571 2456 11605
rect 2456 11571 2465 11605
rect 2413 11562 2465 11571
rect 3422 11606 3474 11658
rect 3086 11550 3138 11602
rect 2834 11494 2886 11546
rect 3422 11438 3474 11490
rect 3086 11382 3138 11434
rect 2750 11326 2802 11378
rect 3422 11270 3474 11322
rect 3086 11214 3138 11266
rect 2666 11158 2718 11210
rect 5168 10572 5220 10624
rect 174 9938 226 9990
rect 622 9938 674 9990
rect 2413 9981 2465 9990
rect 2413 9947 2422 9981
rect 2422 9947 2456 9981
rect 2456 9947 2465 9981
rect 2413 9938 2465 9947
rect 2750 9986 2802 10038
rect 3002 9930 3054 9982
rect 3422 9874 3474 9926
rect 2834 9818 2886 9870
rect 3002 9762 3054 9814
rect 3422 9706 3474 9758
rect 2918 9650 2970 9702
rect 3002 9594 3054 9646
rect 3422 9538 3474 9590
rect 5168 9058 5220 9110
rect 3422 8578 3474 8630
rect 3002 8522 3054 8574
rect 2666 8466 2718 8518
rect 3338 8410 3390 8462
rect 3254 8354 3306 8406
rect 2918 8298 2970 8350
rect 3338 8242 3390 8294
rect 3254 8186 3306 8238
rect 2834 8130 2886 8182
rect 5168 7544 5220 7596
rect 2918 6958 2970 7010
rect 3170 6902 3222 6954
rect 3338 6846 3390 6898
rect 2666 6790 2718 6842
rect 3254 6734 3306 6786
rect 3338 6678 3390 6730
rect 2750 6622 2802 6674
rect 3254 6566 3306 6618
rect 3338 6510 3390 6562
rect 5168 6030 5220 6082
rect 3338 5550 3390 5602
rect 3170 5494 3222 5546
rect 2413 5449 2465 5458
rect 2413 5415 2422 5449
rect 2422 5415 2456 5449
rect 2456 5415 2465 5449
rect 2413 5406 2465 5415
rect 2834 5438 2886 5490
rect 3338 5382 3390 5434
rect 3170 5326 3222 5378
rect 2750 5270 2802 5322
rect 3338 5214 3390 5266
rect 3170 5158 3222 5210
rect 2666 5102 2718 5154
rect 5168 4516 5220 4568
rect 2750 3930 2802 3982
rect 3086 3874 3138 3926
rect 2413 3825 2465 3834
rect 2413 3791 2422 3825
rect 2422 3791 2456 3825
rect 2456 3791 2465 3825
rect 2413 3782 2465 3791
rect 3338 3818 3390 3870
rect 2834 3762 2886 3814
rect 3086 3706 3138 3758
rect 3338 3650 3390 3702
rect 2918 3594 2970 3646
rect 3086 3538 3138 3590
rect 3338 3482 3390 3534
rect 5168 3002 5220 3054
rect 3338 2522 3390 2574
rect 3086 2466 3138 2518
rect 2666 2410 2718 2462
rect 90 2326 142 2378
rect 706 2326 758 2378
rect 2413 2369 2465 2378
rect 2413 2335 2422 2369
rect 2422 2335 2456 2369
rect 2456 2335 2465 2369
rect 2413 2326 2465 2335
rect 3338 2354 3390 2406
rect 3002 2298 3054 2350
rect 2918 2242 2970 2294
rect 3338 2186 3390 2238
rect 3002 2130 3054 2182
rect 2834 2074 2886 2126
rect 5168 1488 5220 1540
rect 2918 902 2970 954
rect 3254 846 3306 898
rect 3506 790 3558 842
rect 6 702 58 754
rect 622 702 674 754
rect 2413 745 2465 754
rect 2413 711 2422 745
rect 2422 711 2456 745
rect 2456 711 2465 745
rect 2413 702 2465 711
rect 2666 734 2718 786
rect 3002 678 3054 730
rect 3338 622 3390 674
rect 2750 566 2802 618
rect 3002 510 3054 562
rect 3338 454 3390 506
rect 5168 -26 5220 26
<< metal2 >>
rect 18 754 46 24632
rect 102 2378 130 24632
rect 186 9990 214 24632
rect 270 11614 298 24632
rect 354 19226 382 24632
rect 438 20850 466 24632
rect 2678 23322 2706 24660
rect 2762 23490 2790 24660
rect 2846 23658 2874 24660
rect 18 0 46 702
rect 102 0 130 2326
rect 186 0 214 9938
rect 270 0 298 11562
rect 354 0 382 19174
rect 438 0 466 20798
rect 2678 20630 2706 23270
rect 2762 22150 2790 23438
rect 2678 18954 2706 20578
rect 2678 17266 2706 18902
rect 2762 18786 2790 22098
rect 2846 21982 2874 23606
rect 2846 20294 2874 21930
rect 2930 21814 2958 24660
rect 2930 20462 2958 21762
rect 2762 17434 2790 18734
rect 2846 17602 2874 20242
rect 2930 19122 2958 20410
rect 2678 14574 2706 17214
rect 2762 16094 2790 17382
rect 2678 12898 2706 14522
rect 2678 11210 2706 12846
rect 2762 12730 2790 16042
rect 2846 15926 2874 17550
rect 2846 14238 2874 15874
rect 2930 15758 2958 19070
rect 3014 19066 3042 24660
rect 3098 20518 3126 24660
rect 3182 22094 3210 24660
rect 3266 23714 3294 24660
rect 3266 23546 3294 23662
rect 3266 23378 3294 23494
rect 3182 21926 3210 22042
rect 3182 21758 3210 21874
rect 3182 20686 3210 21706
rect 3098 20350 3126 20466
rect 3014 17658 3042 19014
rect 3098 18898 3126 20298
rect 3098 18730 3126 18846
rect 3014 17490 3042 17606
rect 3014 17322 3042 17438
rect 2930 14406 2958 15706
rect 2762 11378 2790 12678
rect 2846 11546 2874 14186
rect 2930 13066 2958 14354
rect 2678 8518 2706 11158
rect 2762 10038 2790 11326
rect 2678 6842 2706 8466
rect 2678 5154 2706 6790
rect 2762 6674 2790 9986
rect 2846 9870 2874 11494
rect 2846 8182 2874 9818
rect 2930 9702 2958 13014
rect 3014 9982 3042 17270
rect 3098 13010 3126 18678
rect 3182 14462 3210 20634
rect 3266 16038 3294 23326
rect 3350 18500 3378 24660
rect 3434 20040 3462 24660
rect 3518 23770 3546 24660
rect 3518 23602 3546 23718
rect 3518 23434 3546 23550
rect 3518 22038 3546 23382
rect 3602 23120 3630 24660
rect 3518 21870 3546 21986
rect 3518 21702 3546 21818
rect 3518 21580 3546 21650
rect 3518 20742 3546 21524
rect 3518 20574 3546 20690
rect 3518 20406 3546 20522
rect 3266 15870 3294 15986
rect 3266 15702 3294 15818
rect 3266 14630 3294 15650
rect 3182 14294 3210 14410
rect 3098 11602 3126 12958
rect 3182 12842 3210 14242
rect 3266 13884 3294 14578
rect 3182 12674 3210 12790
rect 3182 12344 3210 12622
rect 3098 11434 3126 11550
rect 3098 11266 3126 11382
rect 3098 10804 3126 11214
rect 3014 9814 3042 9930
rect 2930 8350 2958 9650
rect 3014 9646 3042 9762
rect 3014 9264 3042 9594
rect 3014 8574 3042 9208
rect 2762 5322 2790 6622
rect 2846 5490 2874 8130
rect 2930 7010 2958 8298
rect 2678 2462 2706 5102
rect 2762 3982 2790 5270
rect 2678 786 2706 2410
rect 2762 1568 2790 3930
rect 2846 3814 2874 5438
rect 2930 4648 2958 6958
rect 2846 3108 2874 3762
rect 2930 3646 2958 4592
rect 2846 2126 2874 3052
rect 2930 2294 2958 3594
rect 3014 2350 3042 8522
rect 3098 3926 3126 10748
rect 3182 6954 3210 12288
rect 3266 8406 3294 13828
rect 3350 8462 3378 18444
rect 3434 15982 3462 19984
rect 3518 19010 3546 20354
rect 3518 18842 3546 18958
rect 3518 18674 3546 18790
rect 3518 17714 3546 18622
rect 3518 17546 3546 17662
rect 3518 17378 3546 17494
rect 3434 15814 3462 15930
rect 3434 15646 3462 15762
rect 3434 14686 3462 15594
rect 3434 14518 3462 14634
rect 3434 14350 3462 14466
rect 3434 12954 3462 14298
rect 3434 12786 3462 12902
rect 3434 12618 3462 12734
rect 3434 11658 3462 12566
rect 3434 11490 3462 11606
rect 3434 11322 3462 11438
rect 3434 9926 3462 11270
rect 3434 9758 3462 9874
rect 3434 9590 3462 9706
rect 3434 8630 3462 9538
rect 3266 8238 3294 8354
rect 3350 8294 3378 8410
rect 3182 5546 3210 6902
rect 3266 6786 3294 8186
rect 3350 6898 3378 8242
rect 3266 6618 3294 6734
rect 3350 6730 3378 6846
rect 3182 5378 3210 5494
rect 3182 5210 3210 5326
rect 3098 3758 3126 3874
rect 3098 3590 3126 3706
rect 3098 2518 3126 3538
rect 2678 28 2706 734
rect 2762 618 2790 1512
rect 2762 0 2790 566
rect 2846 0 2874 2074
rect 2930 954 2958 2242
rect 3014 2182 3042 2298
rect 2930 0 2958 902
rect 3014 730 3042 2130
rect 3014 562 3042 678
rect 3014 0 3042 510
rect 3098 0 3126 2466
rect 3182 0 3210 5158
rect 3266 898 3294 6566
rect 3350 6562 3378 6678
rect 3350 5602 3378 6510
rect 3350 5434 3378 5550
rect 3350 5266 3378 5382
rect 3350 3870 3378 5214
rect 3350 3702 3378 3818
rect 3350 3534 3378 3650
rect 3350 2574 3378 3482
rect 3350 2406 3378 2522
rect 3350 2238 3378 2354
rect 3266 0 3294 846
rect 3350 674 3378 2186
rect 3350 506 3378 622
rect 3350 0 3378 454
rect 3434 0 3462 8578
rect 3518 842 3546 17326
rect 3518 0 3546 790
rect 3602 0 3630 23064
<< via2 >>
rect 2411 23930 2467 23932
rect 2411 23878 2413 23930
rect 2413 23878 2465 23930
rect 2465 23878 2467 23930
rect 2411 23876 2467 23878
rect 2411 22306 2467 22308
rect 2411 22254 2413 22306
rect 2413 22254 2465 22306
rect 2465 22254 2467 22306
rect 2411 22252 2467 22254
rect 2411 20850 2467 20852
rect 2411 20798 2413 20850
rect 2413 20798 2465 20850
rect 2465 20798 2467 20850
rect 2411 20796 2467 20798
rect 2411 19226 2467 19228
rect 2411 19174 2413 19226
rect 2413 19174 2465 19226
rect 2465 19174 2467 19226
rect 2411 19172 2467 19174
rect 2411 14694 2467 14696
rect 2411 14642 2413 14694
rect 2413 14642 2465 14694
rect 2465 14642 2467 14694
rect 2411 14640 2467 14642
rect 2411 13070 2467 13072
rect 2411 13018 2413 13070
rect 2413 13018 2465 13070
rect 2465 13018 2467 13070
rect 2411 13016 2467 13018
rect 2411 11614 2467 11616
rect 2411 11562 2413 11614
rect 2413 11562 2465 11614
rect 2465 11562 2467 11614
rect 2411 11560 2467 11562
rect 2411 9990 2467 9992
rect 2411 9938 2413 9990
rect 2413 9938 2465 9990
rect 2465 9938 2467 9990
rect 2411 9936 2467 9938
rect 2411 5458 2467 5460
rect 2411 5406 2413 5458
rect 2413 5406 2465 5458
rect 2465 5406 2467 5458
rect 2411 5404 2467 5406
rect 5166 24250 5222 24252
rect 5166 24198 5168 24250
rect 5168 24198 5220 24250
rect 5220 24198 5222 24250
rect 5166 24196 5222 24198
rect 3588 23064 3644 23120
rect 3504 21524 3560 21580
rect 3420 19984 3476 20040
rect 3336 18444 3392 18500
rect 3252 13828 3308 13884
rect 3168 12288 3224 12344
rect 3084 10748 3140 10804
rect 3000 9208 3056 9264
rect 2411 3834 2467 3836
rect 2411 3782 2413 3834
rect 2413 3782 2465 3834
rect 2465 3782 2467 3834
rect 2411 3780 2467 3782
rect 2411 2378 2467 2380
rect 2411 2326 2413 2378
rect 2413 2326 2465 2378
rect 2465 2326 2467 2378
rect 2411 2324 2467 2326
rect 2916 4592 2972 4648
rect 2832 3052 2888 3108
rect 2748 1512 2804 1568
rect 2411 754 2467 756
rect 2411 702 2413 754
rect 2413 702 2465 754
rect 2465 702 2467 754
rect 2411 700 2467 702
rect 2664 -28 2720 28
rect 5166 22736 5222 22738
rect 5166 22684 5168 22736
rect 5168 22684 5220 22736
rect 5220 22684 5222 22736
rect 5166 22682 5222 22684
rect 5166 21222 5222 21224
rect 5166 21170 5168 21222
rect 5168 21170 5220 21222
rect 5220 21170 5222 21222
rect 5166 21168 5222 21170
rect 5166 19708 5222 19710
rect 5166 19656 5168 19708
rect 5168 19656 5220 19708
rect 5220 19656 5222 19708
rect 5166 19654 5222 19656
rect 5166 18194 5222 18196
rect 5166 18142 5168 18194
rect 5168 18142 5220 18194
rect 5220 18142 5222 18194
rect 5166 18140 5222 18142
rect 5166 16680 5222 16682
rect 5166 16628 5168 16680
rect 5168 16628 5220 16680
rect 5220 16628 5222 16680
rect 5166 16626 5222 16628
rect 5166 15166 5222 15168
rect 5166 15114 5168 15166
rect 5168 15114 5220 15166
rect 5220 15114 5222 15166
rect 5166 15112 5222 15114
rect 5166 13652 5222 13654
rect 5166 13600 5168 13652
rect 5168 13600 5220 13652
rect 5220 13600 5222 13652
rect 5166 13598 5222 13600
rect 5166 12138 5222 12140
rect 5166 12086 5168 12138
rect 5168 12086 5220 12138
rect 5220 12086 5222 12138
rect 5166 12084 5222 12086
rect 5166 10624 5222 10626
rect 5166 10572 5168 10624
rect 5168 10572 5220 10624
rect 5220 10572 5222 10624
rect 5166 10570 5222 10572
rect 5166 9110 5222 9112
rect 5166 9058 5168 9110
rect 5168 9058 5220 9110
rect 5220 9058 5222 9110
rect 5166 9056 5222 9058
rect 5166 7596 5222 7598
rect 5166 7544 5168 7596
rect 5168 7544 5220 7596
rect 5220 7544 5222 7596
rect 5166 7542 5222 7544
rect 5166 6082 5222 6084
rect 5166 6030 5168 6082
rect 5168 6030 5220 6082
rect 5220 6030 5222 6082
rect 5166 6028 5222 6030
rect 5166 4568 5222 4570
rect 5166 4516 5168 4568
rect 5168 4516 5220 4568
rect 5220 4516 5222 4568
rect 5166 4514 5222 4516
rect 5166 3054 5222 3056
rect 5166 3002 5168 3054
rect 5168 3002 5220 3054
rect 5220 3002 5222 3054
rect 5166 3000 5222 3002
rect 5166 1540 5222 1542
rect 5166 1488 5168 1540
rect 5168 1488 5220 1540
rect 5220 1488 5222 1540
rect 5166 1486 5222 1488
rect 5166 26 5222 28
rect 5166 -26 5168 26
rect 5168 -26 5220 26
rect 5220 -26 5222 26
rect 5166 -28 5222 -26
<< metal3 >>
rect 828 24602 888 24662
rect 1700 24602 1760 24662
rect 5164 24252 5224 24254
rect 5164 24196 5166 24252
rect 5222 24196 5224 24252
rect 5164 24194 5224 24196
rect 2409 23932 2469 23934
rect 2409 23876 2411 23932
rect 2467 23876 2469 23932
rect 2409 23122 2469 23876
rect 828 23062 888 23122
rect 1700 23062 1760 23122
rect 2409 23120 3646 23122
rect 2409 23064 3588 23120
rect 3644 23064 3646 23120
rect 2409 23062 3646 23064
rect 5164 22738 5224 22740
rect 5164 22682 5166 22738
rect 5222 22682 5224 22738
rect 5164 22680 5224 22682
rect 2409 22308 2469 22310
rect 2409 22252 2411 22308
rect 2467 22252 2469 22308
rect 2409 21582 2469 22252
rect 828 21522 888 21582
rect 1700 21522 1760 21582
rect 2409 21580 3562 21582
rect 2409 21524 3504 21580
rect 3560 21524 3562 21580
rect 2409 21522 3562 21524
rect 5164 21224 5224 21226
rect 5164 21168 5166 21224
rect 5222 21168 5224 21224
rect 5164 21166 5224 21168
rect 2409 20852 2469 20854
rect 2409 20796 2411 20852
rect 2467 20796 2469 20852
rect 2409 20042 2469 20796
rect 828 19982 888 20042
rect 1700 19982 1760 20042
rect 2409 20040 3478 20042
rect 2409 19984 3420 20040
rect 3476 19984 3478 20040
rect 2409 19982 3478 19984
rect 5164 19710 5224 19712
rect 5164 19654 5166 19710
rect 5222 19654 5224 19710
rect 5164 19652 5224 19654
rect 2409 19228 2469 19230
rect 2409 19172 2411 19228
rect 2467 19172 2469 19228
rect 2409 18502 2469 19172
rect 828 18442 888 18502
rect 1700 18442 1760 18502
rect 2409 18500 3394 18502
rect 2409 18444 3336 18500
rect 3392 18444 3394 18500
rect 2409 18442 3394 18444
rect 5164 18196 5224 18198
rect 5164 18140 5166 18196
rect 5222 18140 5224 18196
rect 5164 18138 5224 18140
rect 5164 16682 5224 16684
rect 5164 16626 5166 16682
rect 5222 16626 5224 16682
rect 5164 16624 5224 16626
rect 828 15366 888 15426
rect 1700 15366 1760 15426
rect 5164 15168 5224 15170
rect 5164 15112 5166 15168
rect 5222 15112 5224 15168
rect 5164 15110 5224 15112
rect 2409 14696 2469 14698
rect 2409 14640 2411 14696
rect 2467 14640 2469 14696
rect 2409 13886 2469 14640
rect 828 13826 888 13886
rect 1700 13826 1760 13886
rect 2409 13884 3310 13886
rect 2409 13828 3252 13884
rect 3308 13828 3310 13884
rect 2409 13826 3310 13828
rect 5164 13654 5224 13656
rect 5164 13598 5166 13654
rect 5222 13598 5224 13654
rect 5164 13596 5224 13598
rect 2409 13072 2469 13074
rect 2409 13016 2411 13072
rect 2467 13016 2469 13072
rect 2409 12346 2469 13016
rect 828 12286 888 12346
rect 1700 12286 1760 12346
rect 2409 12344 3226 12346
rect 2409 12288 3168 12344
rect 3224 12288 3226 12344
rect 2409 12286 3226 12288
rect 5164 12140 5224 12142
rect 5164 12084 5166 12140
rect 5222 12084 5224 12140
rect 5164 12082 5224 12084
rect 2409 11616 2469 11618
rect 2409 11560 2411 11616
rect 2467 11560 2469 11616
rect 2409 10806 2469 11560
rect 828 10746 888 10806
rect 1700 10746 1760 10806
rect 2409 10804 3142 10806
rect 2409 10748 3084 10804
rect 3140 10748 3142 10804
rect 2409 10746 3142 10748
rect 5164 10626 5224 10628
rect 5164 10570 5166 10626
rect 5222 10570 5224 10626
rect 5164 10568 5224 10570
rect 2409 9992 2469 9994
rect 2409 9936 2411 9992
rect 2467 9936 2469 9992
rect 2409 9266 2469 9936
rect 828 9206 888 9266
rect 1700 9206 1760 9266
rect 2409 9264 3058 9266
rect 2409 9208 3000 9264
rect 3056 9208 3058 9264
rect 2409 9206 3058 9208
rect 5164 9112 5224 9114
rect 5164 9056 5166 9112
rect 5222 9056 5224 9112
rect 5164 9054 5224 9056
rect 5164 7598 5224 7600
rect 5164 7542 5166 7598
rect 5222 7542 5224 7598
rect 5164 7540 5224 7542
rect 828 6130 888 6190
rect 1700 6130 1760 6190
rect 5164 6084 5224 6086
rect 5164 6028 5166 6084
rect 5222 6028 5224 6084
rect 5164 6026 5224 6028
rect 2409 5460 2469 5462
rect 2409 5404 2411 5460
rect 2467 5404 2469 5460
rect 2409 4650 2469 5404
rect 828 4590 888 4650
rect 1700 4590 1760 4650
rect 2409 4648 2974 4650
rect 2409 4592 2916 4648
rect 2972 4592 2974 4648
rect 2409 4590 2974 4592
rect 5164 4570 5224 4572
rect 5164 4514 5166 4570
rect 5222 4514 5224 4570
rect 5164 4512 5224 4514
rect 2409 3836 2469 3838
rect 2409 3780 2411 3836
rect 2467 3780 2469 3836
rect 2409 3110 2469 3780
rect 828 3050 888 3110
rect 1700 3050 1760 3110
rect 2409 3108 2890 3110
rect 2409 3052 2832 3108
rect 2888 3052 2890 3108
rect 2409 3050 2890 3052
rect 5164 3056 5224 3058
rect 5164 3000 5166 3056
rect 5222 3000 5224 3056
rect 5164 2998 5224 3000
rect 2409 2380 2469 2382
rect 2409 2324 2411 2380
rect 2467 2324 2469 2380
rect 2409 1570 2469 2324
rect 828 1510 888 1570
rect 1700 1510 1760 1570
rect 2409 1568 2806 1570
rect 2409 1512 2748 1568
rect 2804 1512 2806 1568
rect 2409 1510 2806 1512
rect 5164 1542 5224 1544
rect 5164 1486 5166 1542
rect 5222 1486 5224 1542
rect 5164 1484 5224 1486
rect 2409 756 2469 758
rect 2409 700 2411 756
rect 2467 700 2469 756
rect 2409 30 2469 700
rect 828 -30 888 30
rect 1700 -30 1760 30
rect 2409 28 2722 30
rect 2409 -28 2664 28
rect 2720 -28 2722 28
rect 2409 -30 2722 -28
rect 5164 28 5224 30
rect 5164 -28 5166 28
rect 5222 -28 5224 28
rect 5164 -30 5224 -28
use contact_18  contact_18_0
timestamp 1643593061
transform 1 0 5164 0 1 -30
box 0 0 1 1
use contact_17  contact_17_0
timestamp 1643593061
transform 1 0 5162 0 1 -26
box 0 0 1 1
use contact_18  contact_18_1
timestamp 1643593061
transform 1 0 5164 0 1 1484
box 0 0 1 1
use contact_17  contact_17_1
timestamp 1643593061
transform 1 0 5162 0 1 1488
box 0 0 1 1
use contact_18  contact_18_2
timestamp 1643593061
transform 1 0 5164 0 1 -30
box 0 0 1 1
use contact_17  contact_17_2
timestamp 1643593061
transform 1 0 5162 0 1 -26
box 0 0 1 1
use contact_18  contact_18_3
timestamp 1643593061
transform 1 0 5164 0 1 1484
box 0 0 1 1
use contact_17  contact_17_3
timestamp 1643593061
transform 1 0 5162 0 1 1488
box 0 0 1 1
use contact_18  contact_18_4
timestamp 1643593061
transform 1 0 5164 0 1 -30
box 0 0 1 1
use contact_17  contact_17_4
timestamp 1643593061
transform 1 0 5162 0 1 -26
box 0 0 1 1
use contact_18  contact_18_5
timestamp 1643593061
transform 1 0 5164 0 1 1484
box 0 0 1 1
use contact_17  contact_17_5
timestamp 1643593061
transform 1 0 5162 0 1 1488
box 0 0 1 1
use contact_18  contact_18_6
timestamp 1643593061
transform 1 0 5164 0 1 -30
box 0 0 1 1
use contact_17  contact_17_6
timestamp 1643593061
transform 1 0 5162 0 1 -26
box 0 0 1 1
use contact_18  contact_18_7
timestamp 1643593061
transform 1 0 5164 0 1 1484
box 0 0 1 1
use contact_17  contact_17_7
timestamp 1643593061
transform 1 0 5162 0 1 1488
box 0 0 1 1
use contact_18  contact_18_8
timestamp 1643593061
transform 1 0 5164 0 1 -30
box 0 0 1 1
use contact_17  contact_17_8
timestamp 1643593061
transform 1 0 5162 0 1 -26
box 0 0 1 1
use contact_18  contact_18_9
timestamp 1643593061
transform 1 0 5164 0 1 1484
box 0 0 1 1
use contact_17  contact_17_9
timestamp 1643593061
transform 1 0 5162 0 1 1488
box 0 0 1 1
use contact_18  contact_18_10
timestamp 1643593061
transform 1 0 5164 0 1 -30
box 0 0 1 1
use contact_17  contact_17_10
timestamp 1643593061
transform 1 0 5162 0 1 -26
box 0 0 1 1
use contact_18  contact_18_11
timestamp 1643593061
transform 1 0 5164 0 1 1484
box 0 0 1 1
use contact_17  contact_17_11
timestamp 1643593061
transform 1 0 5162 0 1 1488
box 0 0 1 1
use contact_18  contact_18_12
timestamp 1643593061
transform 1 0 5164 0 1 -30
box 0 0 1 1
use contact_17  contact_17_12
timestamp 1643593061
transform 1 0 5162 0 1 -26
box 0 0 1 1
use contact_18  contact_18_13
timestamp 1643593061
transform 1 0 5164 0 1 1484
box 0 0 1 1
use contact_17  contact_17_13
timestamp 1643593061
transform 1 0 5162 0 1 1488
box 0 0 1 1
use contact_18  contact_18_14
timestamp 1643593061
transform 1 0 5164 0 1 -30
box 0 0 1 1
use contact_17  contact_17_14
timestamp 1643593061
transform 1 0 5162 0 1 -26
box 0 0 1 1
use contact_18  contact_18_15
timestamp 1643593061
transform 1 0 5164 0 1 1484
box 0 0 1 1
use contact_17  contact_17_15
timestamp 1643593061
transform 1 0 5162 0 1 1488
box 0 0 1 1
use contact_18  contact_18_16
timestamp 1643593061
transform 1 0 5164 0 1 -30
box 0 0 1 1
use contact_17  contact_17_16
timestamp 1643593061
transform 1 0 5162 0 1 -26
box 0 0 1 1
use contact_18  contact_18_17
timestamp 1643593061
transform 1 0 5164 0 1 1484
box 0 0 1 1
use contact_17  contact_17_17
timestamp 1643593061
transform 1 0 5162 0 1 1488
box 0 0 1 1
use contact_18  contact_18_18
timestamp 1643593061
transform 1 0 5164 0 1 -30
box 0 0 1 1
use contact_17  contact_17_18
timestamp 1643593061
transform 1 0 5162 0 1 -26
box 0 0 1 1
use contact_18  contact_18_19
timestamp 1643593061
transform 1 0 5164 0 1 1484
box 0 0 1 1
use contact_17  contact_17_19
timestamp 1643593061
transform 1 0 5162 0 1 1488
box 0 0 1 1
use contact_18  contact_18_20
timestamp 1643593061
transform 1 0 5164 0 1 -30
box 0 0 1 1
use contact_17  contact_17_20
timestamp 1643593061
transform 1 0 5162 0 1 -26
box 0 0 1 1
use contact_18  contact_18_21
timestamp 1643593061
transform 1 0 5164 0 1 1484
box 0 0 1 1
use contact_17  contact_17_21
timestamp 1643593061
transform 1 0 5162 0 1 1488
box 0 0 1 1
use contact_18  contact_18_22
timestamp 1643593061
transform 1 0 5164 0 1 -30
box 0 0 1 1
use contact_17  contact_17_22
timestamp 1643593061
transform 1 0 5162 0 1 -26
box 0 0 1 1
use contact_18  contact_18_23
timestamp 1643593061
transform 1 0 5164 0 1 1484
box 0 0 1 1
use contact_17  contact_17_23
timestamp 1643593061
transform 1 0 5162 0 1 1488
box 0 0 1 1
use contact_18  contact_18_24
timestamp 1643593061
transform 1 0 5164 0 1 -30
box 0 0 1 1
use contact_17  contact_17_24
timestamp 1643593061
transform 1 0 5162 0 1 -26
box 0 0 1 1
use contact_18  contact_18_25
timestamp 1643593061
transform 1 0 5164 0 1 1484
box 0 0 1 1
use contact_17  contact_17_25
timestamp 1643593061
transform 1 0 5162 0 1 1488
box 0 0 1 1
use contact_18  contact_18_26
timestamp 1643593061
transform 1 0 5164 0 1 -30
box 0 0 1 1
use contact_17  contact_17_26
timestamp 1643593061
transform 1 0 5162 0 1 -26
box 0 0 1 1
use contact_18  contact_18_27
timestamp 1643593061
transform 1 0 5164 0 1 1484
box 0 0 1 1
use contact_17  contact_17_27
timestamp 1643593061
transform 1 0 5162 0 1 1488
box 0 0 1 1
use contact_18  contact_18_28
timestamp 1643593061
transform 1 0 5164 0 1 -30
box 0 0 1 1
use contact_17  contact_17_28
timestamp 1643593061
transform 1 0 5162 0 1 -26
box 0 0 1 1
use contact_18  contact_18_29
timestamp 1643593061
transform 1 0 5164 0 1 1484
box 0 0 1 1
use contact_17  contact_17_29
timestamp 1643593061
transform 1 0 5162 0 1 1488
box 0 0 1 1
use contact_18  contact_18_30
timestamp 1643593061
transform 1 0 5164 0 1 -30
box 0 0 1 1
use contact_17  contact_17_30
timestamp 1643593061
transform 1 0 5162 0 1 -26
box 0 0 1 1
use contact_18  contact_18_31
timestamp 1643593061
transform 1 0 5164 0 1 1484
box 0 0 1 1
use contact_17  contact_17_31
timestamp 1643593061
transform 1 0 5162 0 1 1488
box 0 0 1 1
use contact_18  contact_18_32
timestamp 1643593061
transform 1 0 5164 0 1 -30
box 0 0 1 1
use contact_17  contact_17_32
timestamp 1643593061
transform 1 0 5162 0 1 -26
box 0 0 1 1
use contact_18  contact_18_33
timestamp 1643593061
transform 1 0 5164 0 1 1484
box 0 0 1 1
use contact_17  contact_17_33
timestamp 1643593061
transform 1 0 5162 0 1 1488
box 0 0 1 1
use contact_18  contact_18_34
timestamp 1643593061
transform 1 0 5164 0 1 -30
box 0 0 1 1
use contact_17  contact_17_34
timestamp 1643593061
transform 1 0 5162 0 1 -26
box 0 0 1 1
use contact_18  contact_18_35
timestamp 1643593061
transform 1 0 5164 0 1 1484
box 0 0 1 1
use contact_17  contact_17_35
timestamp 1643593061
transform 1 0 5162 0 1 1488
box 0 0 1 1
use contact_18  contact_18_36
timestamp 1643593061
transform 1 0 5164 0 1 -30
box 0 0 1 1
use contact_17  contact_17_36
timestamp 1643593061
transform 1 0 5162 0 1 -26
box 0 0 1 1
use contact_18  contact_18_37
timestamp 1643593061
transform 1 0 5164 0 1 1484
box 0 0 1 1
use contact_17  contact_17_37
timestamp 1643593061
transform 1 0 5162 0 1 1488
box 0 0 1 1
use contact_18  contact_18_38
timestamp 1643593061
transform 1 0 5164 0 1 -30
box 0 0 1 1
use contact_17  contact_17_38
timestamp 1643593061
transform 1 0 5162 0 1 -26
box 0 0 1 1
use contact_18  contact_18_39
timestamp 1643593061
transform 1 0 5164 0 1 1484
box 0 0 1 1
use contact_17  contact_17_39
timestamp 1643593061
transform 1 0 5162 0 1 1488
box 0 0 1 1
use contact_18  contact_18_40
timestamp 1643593061
transform 1 0 5164 0 1 -30
box 0 0 1 1
use contact_17  contact_17_40
timestamp 1643593061
transform 1 0 5162 0 1 -26
box 0 0 1 1
use contact_18  contact_18_41
timestamp 1643593061
transform 1 0 5164 0 1 1484
box 0 0 1 1
use contact_17  contact_17_41
timestamp 1643593061
transform 1 0 5162 0 1 1488
box 0 0 1 1
use contact_18  contact_18_42
timestamp 1643593061
transform 1 0 5164 0 1 -30
box 0 0 1 1
use contact_17  contact_17_42
timestamp 1643593061
transform 1 0 5162 0 1 -26
box 0 0 1 1
use contact_18  contact_18_43
timestamp 1643593061
transform 1 0 5164 0 1 1484
box 0 0 1 1
use contact_17  contact_17_43
timestamp 1643593061
transform 1 0 5162 0 1 1488
box 0 0 1 1
use contact_18  contact_18_44
timestamp 1643593061
transform 1 0 5164 0 1 -30
box 0 0 1 1
use contact_17  contact_17_44
timestamp 1643593061
transform 1 0 5162 0 1 -26
box 0 0 1 1
use contact_18  contact_18_45
timestamp 1643593061
transform 1 0 5164 0 1 1484
box 0 0 1 1
use contact_17  contact_17_45
timestamp 1643593061
transform 1 0 5162 0 1 1488
box 0 0 1 1
use contact_18  contact_18_46
timestamp 1643593061
transform 1 0 5164 0 1 -30
box 0 0 1 1
use contact_17  contact_17_46
timestamp 1643593061
transform 1 0 5162 0 1 -26
box 0 0 1 1
use contact_18  contact_18_47
timestamp 1643593061
transform 1 0 5164 0 1 1484
box 0 0 1 1
use contact_17  contact_17_47
timestamp 1643593061
transform 1 0 5162 0 1 1488
box 0 0 1 1
use contact_18  contact_18_48
timestamp 1643593061
transform 1 0 5164 0 1 -30
box 0 0 1 1
use contact_17  contact_17_48
timestamp 1643593061
transform 1 0 5162 0 1 -26
box 0 0 1 1
use contact_18  contact_18_49
timestamp 1643593061
transform 1 0 5164 0 1 1484
box 0 0 1 1
use contact_17  contact_17_49
timestamp 1643593061
transform 1 0 5162 0 1 1488
box 0 0 1 1
use contact_18  contact_18_50
timestamp 1643593061
transform 1 0 5164 0 1 -30
box 0 0 1 1
use contact_17  contact_17_50
timestamp 1643593061
transform 1 0 5162 0 1 -26
box 0 0 1 1
use contact_18  contact_18_51
timestamp 1643593061
transform 1 0 5164 0 1 1484
box 0 0 1 1
use contact_17  contact_17_51
timestamp 1643593061
transform 1 0 5162 0 1 1488
box 0 0 1 1
use contact_18  contact_18_52
timestamp 1643593061
transform 1 0 5164 0 1 -30
box 0 0 1 1
use contact_17  contact_17_52
timestamp 1643593061
transform 1 0 5162 0 1 -26
box 0 0 1 1
use contact_18  contact_18_53
timestamp 1643593061
transform 1 0 5164 0 1 1484
box 0 0 1 1
use contact_17  contact_17_53
timestamp 1643593061
transform 1 0 5162 0 1 1488
box 0 0 1 1
use contact_18  contact_18_54
timestamp 1643593061
transform 1 0 5164 0 1 -30
box 0 0 1 1
use contact_17  contact_17_54
timestamp 1643593061
transform 1 0 5162 0 1 -26
box 0 0 1 1
use contact_18  contact_18_55
timestamp 1643593061
transform 1 0 5164 0 1 1484
box 0 0 1 1
use contact_17  contact_17_55
timestamp 1643593061
transform 1 0 5162 0 1 1488
box 0 0 1 1
use contact_18  contact_18_56
timestamp 1643593061
transform 1 0 5164 0 1 -30
box 0 0 1 1
use contact_17  contact_17_56
timestamp 1643593061
transform 1 0 5162 0 1 -26
box 0 0 1 1
use contact_18  contact_18_57
timestamp 1643593061
transform 1 0 5164 0 1 1484
box 0 0 1 1
use contact_17  contact_17_57
timestamp 1643593061
transform 1 0 5162 0 1 1488
box 0 0 1 1
use contact_18  contact_18_58
timestamp 1643593061
transform 1 0 5164 0 1 -30
box 0 0 1 1
use contact_17  contact_17_58
timestamp 1643593061
transform 1 0 5162 0 1 -26
box 0 0 1 1
use contact_18  contact_18_59
timestamp 1643593061
transform 1 0 5164 0 1 1484
box 0 0 1 1
use contact_17  contact_17_59
timestamp 1643593061
transform 1 0 5162 0 1 1488
box 0 0 1 1
use contact_18  contact_18_60
timestamp 1643593061
transform 1 0 5164 0 1 -30
box 0 0 1 1
use contact_17  contact_17_60
timestamp 1643593061
transform 1 0 5162 0 1 -26
box 0 0 1 1
use contact_18  contact_18_61
timestamp 1643593061
transform 1 0 5164 0 1 1484
box 0 0 1 1
use contact_17  contact_17_61
timestamp 1643593061
transform 1 0 5162 0 1 1488
box 0 0 1 1
use contact_18  contact_18_62
timestamp 1643593061
transform 1 0 5164 0 1 -30
box 0 0 1 1
use contact_17  contact_17_62
timestamp 1643593061
transform 1 0 5162 0 1 -26
box 0 0 1 1
use contact_18  contact_18_63
timestamp 1643593061
transform 1 0 5164 0 1 1484
box 0 0 1 1
use contact_17  contact_17_63
timestamp 1643593061
transform 1 0 5162 0 1 1488
box 0 0 1 1
use contact_18  contact_18_64
timestamp 1643593061
transform 1 0 5164 0 1 24194
box 0 0 1 1
use contact_17  contact_17_64
timestamp 1643593061
transform 1 0 5162 0 1 24198
box 0 0 1 1
use contact_18  contact_18_65
timestamp 1643593061
transform 1 0 5164 0 1 22680
box 0 0 1 1
use contact_17  contact_17_65
timestamp 1643593061
transform 1 0 5162 0 1 22684
box 0 0 1 1
use contact_18  contact_18_66
timestamp 1643593061
transform 1 0 5164 0 1 21166
box 0 0 1 1
use contact_17  contact_17_66
timestamp 1643593061
transform 1 0 5162 0 1 21170
box 0 0 1 1
use contact_18  contact_18_67
timestamp 1643593061
transform 1 0 5164 0 1 22680
box 0 0 1 1
use contact_17  contact_17_67
timestamp 1643593061
transform 1 0 5162 0 1 22684
box 0 0 1 1
use contact_18  contact_18_68
timestamp 1643593061
transform 1 0 5164 0 1 21166
box 0 0 1 1
use contact_17  contact_17_68
timestamp 1643593061
transform 1 0 5162 0 1 21170
box 0 0 1 1
use contact_18  contact_18_69
timestamp 1643593061
transform 1 0 5164 0 1 19652
box 0 0 1 1
use contact_17  contact_17_69
timestamp 1643593061
transform 1 0 5162 0 1 19656
box 0 0 1 1
use contact_18  contact_18_70
timestamp 1643593061
transform 1 0 5164 0 1 18138
box 0 0 1 1
use contact_17  contact_17_70
timestamp 1643593061
transform 1 0 5162 0 1 18142
box 0 0 1 1
use contact_18  contact_18_71
timestamp 1643593061
transform 1 0 5164 0 1 19652
box 0 0 1 1
use contact_17  contact_17_71
timestamp 1643593061
transform 1 0 5162 0 1 19656
box 0 0 1 1
use contact_18  contact_18_72
timestamp 1643593061
transform 1 0 5164 0 1 18138
box 0 0 1 1
use contact_17  contact_17_72
timestamp 1643593061
transform 1 0 5162 0 1 18142
box 0 0 1 1
use contact_18  contact_18_73
timestamp 1643593061
transform 1 0 5164 0 1 16624
box 0 0 1 1
use contact_17  contact_17_73
timestamp 1643593061
transform 1 0 5162 0 1 16628
box 0 0 1 1
use contact_18  contact_18_74
timestamp 1643593061
transform 1 0 5164 0 1 15110
box 0 0 1 1
use contact_17  contact_17_74
timestamp 1643593061
transform 1 0 5162 0 1 15114
box 0 0 1 1
use contact_18  contact_18_75
timestamp 1643593061
transform 1 0 5164 0 1 16624
box 0 0 1 1
use contact_17  contact_17_75
timestamp 1643593061
transform 1 0 5162 0 1 16628
box 0 0 1 1
use contact_18  contact_18_76
timestamp 1643593061
transform 1 0 5164 0 1 15110
box 0 0 1 1
use contact_17  contact_17_76
timestamp 1643593061
transform 1 0 5162 0 1 15114
box 0 0 1 1
use contact_18  contact_18_77
timestamp 1643593061
transform 1 0 5164 0 1 13596
box 0 0 1 1
use contact_17  contact_17_77
timestamp 1643593061
transform 1 0 5162 0 1 13600
box 0 0 1 1
use contact_18  contact_18_78
timestamp 1643593061
transform 1 0 5164 0 1 12082
box 0 0 1 1
use contact_17  contact_17_78
timestamp 1643593061
transform 1 0 5162 0 1 12086
box 0 0 1 1
use contact_18  contact_18_79
timestamp 1643593061
transform 1 0 5164 0 1 13596
box 0 0 1 1
use contact_17  contact_17_79
timestamp 1643593061
transform 1 0 5162 0 1 13600
box 0 0 1 1
use contact_18  contact_18_80
timestamp 1643593061
transform 1 0 5164 0 1 12082
box 0 0 1 1
use contact_17  contact_17_80
timestamp 1643593061
transform 1 0 5162 0 1 12086
box 0 0 1 1
use contact_18  contact_18_81
timestamp 1643593061
transform 1 0 5164 0 1 10568
box 0 0 1 1
use contact_17  contact_17_81
timestamp 1643593061
transform 1 0 5162 0 1 10572
box 0 0 1 1
use contact_18  contact_18_82
timestamp 1643593061
transform 1 0 5164 0 1 9054
box 0 0 1 1
use contact_17  contact_17_82
timestamp 1643593061
transform 1 0 5162 0 1 9058
box 0 0 1 1
use contact_18  contact_18_83
timestamp 1643593061
transform 1 0 5164 0 1 10568
box 0 0 1 1
use contact_17  contact_17_83
timestamp 1643593061
transform 1 0 5162 0 1 10572
box 0 0 1 1
use contact_18  contact_18_84
timestamp 1643593061
transform 1 0 5164 0 1 9054
box 0 0 1 1
use contact_17  contact_17_84
timestamp 1643593061
transform 1 0 5162 0 1 9058
box 0 0 1 1
use contact_18  contact_18_85
timestamp 1643593061
transform 1 0 5164 0 1 7540
box 0 0 1 1
use contact_17  contact_17_85
timestamp 1643593061
transform 1 0 5162 0 1 7544
box 0 0 1 1
use contact_18  contact_18_86
timestamp 1643593061
transform 1 0 5164 0 1 6026
box 0 0 1 1
use contact_17  contact_17_86
timestamp 1643593061
transform 1 0 5162 0 1 6030
box 0 0 1 1
use contact_18  contact_18_87
timestamp 1643593061
transform 1 0 5164 0 1 7540
box 0 0 1 1
use contact_17  contact_17_87
timestamp 1643593061
transform 1 0 5162 0 1 7544
box 0 0 1 1
use contact_18  contact_18_88
timestamp 1643593061
transform 1 0 5164 0 1 6026
box 0 0 1 1
use contact_17  contact_17_88
timestamp 1643593061
transform 1 0 5162 0 1 6030
box 0 0 1 1
use contact_18  contact_18_89
timestamp 1643593061
transform 1 0 5164 0 1 4512
box 0 0 1 1
use contact_17  contact_17_89
timestamp 1643593061
transform 1 0 5162 0 1 4516
box 0 0 1 1
use contact_18  contact_18_90
timestamp 1643593061
transform 1 0 5164 0 1 2998
box 0 0 1 1
use contact_17  contact_17_90
timestamp 1643593061
transform 1 0 5162 0 1 3002
box 0 0 1 1
use contact_18  contact_18_91
timestamp 1643593061
transform 1 0 5164 0 1 4512
box 0 0 1 1
use contact_17  contact_17_91
timestamp 1643593061
transform 1 0 5162 0 1 4516
box 0 0 1 1
use contact_18  contact_18_92
timestamp 1643593061
transform 1 0 5164 0 1 2998
box 0 0 1 1
use contact_17  contact_17_92
timestamp 1643593061
transform 1 0 5162 0 1 3002
box 0 0 1 1
use contact_18  contact_18_93
timestamp 1643593061
transform 1 0 5164 0 1 1484
box 0 0 1 1
use contact_17  contact_17_93
timestamp 1643593061
transform 1 0 5162 0 1 1488
box 0 0 1 1
use contact_18  contact_18_94
timestamp 1643593061
transform 1 0 5164 0 1 -30
box 0 0 1 1
use contact_17  contact_17_94
timestamp 1643593061
transform 1 0 5162 0 1 -26
box 0 0 1 1
use contact_18  contact_18_95
timestamp 1643593061
transform 1 0 5164 0 1 1484
box 0 0 1 1
use contact_17  contact_17_95
timestamp 1643593061
transform 1 0 5162 0 1 1488
box 0 0 1 1
use contact_20  contact_20_0
timestamp 1643593061
transform 1 0 3586 0 1 23062
box 0 0 1 1
use contact_18  contact_18_96
timestamp 1643593061
transform 1 0 2409 0 1 23874
box 0 0 1 1
use contact_17  contact_17_96
timestamp 1643593061
transform 1 0 2407 0 1 23878
box 0 0 1 1
use contact_13  contact_13_0
timestamp 1643593061
transform 1 0 2410 0 1 23881
box 0 0 1 1
use contact_20  contact_20_1
timestamp 1643593061
transform 1 0 3502 0 1 21522
box 0 0 1 1
use contact_18  contact_18_97
timestamp 1643593061
transform 1 0 2409 0 1 22250
box 0 0 1 1
use contact_17  contact_17_97
timestamp 1643593061
transform 1 0 2407 0 1 22254
box 0 0 1 1
use contact_13  contact_13_1
timestamp 1643593061
transform 1 0 2410 0 1 22257
box 0 0 1 1
use contact_20  contact_20_2
timestamp 1643593061
transform 1 0 3418 0 1 19982
box 0 0 1 1
use contact_18  contact_18_98
timestamp 1643593061
transform 1 0 2409 0 1 20794
box 0 0 1 1
use contact_17  contact_17_98
timestamp 1643593061
transform 1 0 2407 0 1 20798
box 0 0 1 1
use contact_13  contact_13_2
timestamp 1643593061
transform 1 0 2410 0 1 20801
box 0 0 1 1
use contact_20  contact_20_3
timestamp 1643593061
transform 1 0 3334 0 1 18442
box 0 0 1 1
use contact_18  contact_18_99
timestamp 1643593061
transform 1 0 2409 0 1 19170
box 0 0 1 1
use contact_17  contact_17_99
timestamp 1643593061
transform 1 0 2407 0 1 19174
box 0 0 1 1
use contact_13  contact_13_3
timestamp 1643593061
transform 1 0 2410 0 1 19177
box 0 0 1 1
use contact_20  contact_20_4
timestamp 1643593061
transform 1 0 3250 0 1 13826
box 0 0 1 1
use contact_18  contact_18_100
timestamp 1643593061
transform 1 0 2409 0 1 14638
box 0 0 1 1
use contact_17  contact_17_100
timestamp 1643593061
transform 1 0 2407 0 1 14642
box 0 0 1 1
use contact_13  contact_13_4
timestamp 1643593061
transform 1 0 2410 0 1 14645
box 0 0 1 1
use contact_20  contact_20_5
timestamp 1643593061
transform 1 0 3166 0 1 12286
box 0 0 1 1
use contact_18  contact_18_101
timestamp 1643593061
transform 1 0 2409 0 1 13014
box 0 0 1 1
use contact_17  contact_17_101
timestamp 1643593061
transform 1 0 2407 0 1 13018
box 0 0 1 1
use contact_13  contact_13_5
timestamp 1643593061
transform 1 0 2410 0 1 13021
box 0 0 1 1
use contact_20  contact_20_6
timestamp 1643593061
transform 1 0 3082 0 1 10746
box 0 0 1 1
use contact_18  contact_18_102
timestamp 1643593061
transform 1 0 2409 0 1 11558
box 0 0 1 1
use contact_17  contact_17_102
timestamp 1643593061
transform 1 0 2407 0 1 11562
box 0 0 1 1
use contact_13  contact_13_6
timestamp 1643593061
transform 1 0 2410 0 1 11565
box 0 0 1 1
use contact_20  contact_20_7
timestamp 1643593061
transform 1 0 2998 0 1 9206
box 0 0 1 1
use contact_18  contact_18_103
timestamp 1643593061
transform 1 0 2409 0 1 9934
box 0 0 1 1
use contact_17  contact_17_103
timestamp 1643593061
transform 1 0 2407 0 1 9938
box 0 0 1 1
use contact_13  contact_13_7
timestamp 1643593061
transform 1 0 2410 0 1 9941
box 0 0 1 1
use contact_20  contact_20_8
timestamp 1643593061
transform 1 0 2914 0 1 4590
box 0 0 1 1
use contact_18  contact_18_104
timestamp 1643593061
transform 1 0 2409 0 1 5402
box 0 0 1 1
use contact_17  contact_17_104
timestamp 1643593061
transform 1 0 2407 0 1 5406
box 0 0 1 1
use contact_13  contact_13_8
timestamp 1643593061
transform 1 0 2410 0 1 5409
box 0 0 1 1
use contact_20  contact_20_9
timestamp 1643593061
transform 1 0 2830 0 1 3050
box 0 0 1 1
use contact_18  contact_18_105
timestamp 1643593061
transform 1 0 2409 0 1 3778
box 0 0 1 1
use contact_17  contact_17_105
timestamp 1643593061
transform 1 0 2407 0 1 3782
box 0 0 1 1
use contact_13  contact_13_9
timestamp 1643593061
transform 1 0 2410 0 1 3785
box 0 0 1 1
use contact_20  contact_20_10
timestamp 1643593061
transform 1 0 2746 0 1 1510
box 0 0 1 1
use contact_18  contact_18_106
timestamp 1643593061
transform 1 0 2409 0 1 2322
box 0 0 1 1
use contact_17  contact_17_106
timestamp 1643593061
transform 1 0 2407 0 1 2326
box 0 0 1 1
use contact_13  contact_13_10
timestamp 1643593061
transform 1 0 2410 0 1 2329
box 0 0 1 1
use contact_20  contact_20_11
timestamp 1643593061
transform 1 0 2662 0 1 -30
box 0 0 1 1
use contact_18  contact_18_107
timestamp 1643593061
transform 1 0 2409 0 1 698
box 0 0 1 1
use contact_17  contact_17_107
timestamp 1643593061
transform 1 0 2407 0 1 702
box 0 0 1 1
use contact_13  contact_13_11
timestamp 1643593061
transform 1 0 2410 0 1 705
box 0 0 1 1
use contact_14  contact_14_0
timestamp 1643593061
transform 1 0 3500 0 1 790
box 0 0 1 1
use contact_14  contact_14_1
timestamp 1643593061
transform 1 0 3248 0 1 846
box 0 0 1 1
use contact_14  contact_14_2
timestamp 1643593061
transform 1 0 2912 0 1 902
box 0 0 1 1
use contact_14  contact_14_3
timestamp 1643593061
transform 1 0 3500 0 1 23718
box 0 0 1 1
use contact_14  contact_14_4
timestamp 1643593061
transform 1 0 3248 0 1 23662
box 0 0 1 1
use contact_14  contact_14_5
timestamp 1643593061
transform 1 0 2828 0 1 23606
box 0 0 1 1
use contact_14  contact_14_6
timestamp 1643593061
transform 1 0 3500 0 1 23550
box 0 0 1 1
use contact_14  contact_14_7
timestamp 1643593061
transform 1 0 3248 0 1 23494
box 0 0 1 1
use contact_14  contact_14_8
timestamp 1643593061
transform 1 0 2744 0 1 23438
box 0 0 1 1
use contact_14  contact_14_9
timestamp 1643593061
transform 1 0 3500 0 1 23382
box 0 0 1 1
use contact_14  contact_14_10
timestamp 1643593061
transform 1 0 3248 0 1 23326
box 0 0 1 1
use contact_14  contact_14_11
timestamp 1643593061
transform 1 0 2660 0 1 23270
box 0 0 1 1
use contact_14  contact_14_12
timestamp 1643593061
transform 1 0 3500 0 1 21650
box 0 0 1 1
use contact_14  contact_14_13
timestamp 1643593061
transform 1 0 3164 0 1 21706
box 0 0 1 1
use contact_14  contact_14_14
timestamp 1643593061
transform 1 0 2912 0 1 21762
box 0 0 1 1
use contact_14  contact_14_15
timestamp 1643593061
transform 1 0 3500 0 1 21818
box 0 0 1 1
use contact_14  contact_14_16
timestamp 1643593061
transform 1 0 3164 0 1 21874
box 0 0 1 1
use contact_14  contact_14_17
timestamp 1643593061
transform 1 0 2828 0 1 21930
box 0 0 1 1
use contact_14  contact_14_18
timestamp 1643593061
transform 1 0 3500 0 1 21986
box 0 0 1 1
use contact_14  contact_14_19
timestamp 1643593061
transform 1 0 3164 0 1 22042
box 0 0 1 1
use contact_14  contact_14_20
timestamp 1643593061
transform 1 0 2744 0 1 22098
box 0 0 1 1
use contact_14  contact_14_21
timestamp 1643593061
transform 1 0 3500 0 1 20690
box 0 0 1 1
use contact_14  contact_14_22
timestamp 1643593061
transform 1 0 3164 0 1 20634
box 0 0 1 1
use contact_14  contact_14_23
timestamp 1643593061
transform 1 0 2660 0 1 20578
box 0 0 1 1
use contact_14  contact_14_24
timestamp 1643593061
transform 1 0 3500 0 1 20522
box 0 0 1 1
use contact_14  contact_14_25
timestamp 1643593061
transform 1 0 3080 0 1 20466
box 0 0 1 1
use contact_14  contact_14_26
timestamp 1643593061
transform 1 0 2912 0 1 20410
box 0 0 1 1
use contact_14  contact_14_27
timestamp 1643593061
transform 1 0 3500 0 1 20354
box 0 0 1 1
use contact_14  contact_14_28
timestamp 1643593061
transform 1 0 3080 0 1 20298
box 0 0 1 1
use contact_14  contact_14_29
timestamp 1643593061
transform 1 0 2828 0 1 20242
box 0 0 1 1
use contact_14  contact_14_30
timestamp 1643593061
transform 1 0 3500 0 1 18622
box 0 0 1 1
use contact_14  contact_14_31
timestamp 1643593061
transform 1 0 3080 0 1 18678
box 0 0 1 1
use contact_14  contact_14_32
timestamp 1643593061
transform 1 0 2744 0 1 18734
box 0 0 1 1
use contact_14  contact_14_33
timestamp 1643593061
transform 1 0 3500 0 1 18790
box 0 0 1 1
use contact_14  contact_14_34
timestamp 1643593061
transform 1 0 3080 0 1 18846
box 0 0 1 1
use contact_14  contact_14_35
timestamp 1643593061
transform 1 0 2660 0 1 18902
box 0 0 1 1
use contact_14  contact_14_36
timestamp 1643593061
transform 1 0 3500 0 1 18958
box 0 0 1 1
use contact_14  contact_14_37
timestamp 1643593061
transform 1 0 2996 0 1 19014
box 0 0 1 1
use contact_14  contact_14_38
timestamp 1643593061
transform 1 0 2912 0 1 19070
box 0 0 1 1
use contact_14  contact_14_39
timestamp 1643593061
transform 1 0 3500 0 1 17662
box 0 0 1 1
use contact_14  contact_14_40
timestamp 1643593061
transform 1 0 2996 0 1 17606
box 0 0 1 1
use contact_14  contact_14_41
timestamp 1643593061
transform 1 0 2828 0 1 17550
box 0 0 1 1
use contact_14  contact_14_42
timestamp 1643593061
transform 1 0 3500 0 1 17494
box 0 0 1 1
use contact_14  contact_14_43
timestamp 1643593061
transform 1 0 2996 0 1 17438
box 0 0 1 1
use contact_14  contact_14_44
timestamp 1643593061
transform 1 0 2744 0 1 17382
box 0 0 1 1
use contact_14  contact_14_45
timestamp 1643593061
transform 1 0 3500 0 1 17326
box 0 0 1 1
use contact_14  contact_14_46
timestamp 1643593061
transform 1 0 2996 0 1 17270
box 0 0 1 1
use contact_14  contact_14_47
timestamp 1643593061
transform 1 0 2660 0 1 17214
box 0 0 1 1
use contact_14  contact_14_48
timestamp 1643593061
transform 1 0 3416 0 1 15594
box 0 0 1 1
use contact_14  contact_14_49
timestamp 1643593061
transform 1 0 3248 0 1 15650
box 0 0 1 1
use contact_14  contact_14_50
timestamp 1643593061
transform 1 0 2912 0 1 15706
box 0 0 1 1
use contact_14  contact_14_51
timestamp 1643593061
transform 1 0 3416 0 1 15762
box 0 0 1 1
use contact_14  contact_14_52
timestamp 1643593061
transform 1 0 3248 0 1 15818
box 0 0 1 1
use contact_14  contact_14_53
timestamp 1643593061
transform 1 0 2828 0 1 15874
box 0 0 1 1
use contact_14  contact_14_54
timestamp 1643593061
transform 1 0 3416 0 1 15930
box 0 0 1 1
use contact_14  contact_14_55
timestamp 1643593061
transform 1 0 3248 0 1 15986
box 0 0 1 1
use contact_14  contact_14_56
timestamp 1643593061
transform 1 0 2744 0 1 16042
box 0 0 1 1
use contact_14  contact_14_57
timestamp 1643593061
transform 1 0 3416 0 1 14634
box 0 0 1 1
use contact_14  contact_14_58
timestamp 1643593061
transform 1 0 3248 0 1 14578
box 0 0 1 1
use contact_14  contact_14_59
timestamp 1643593061
transform 1 0 2660 0 1 14522
box 0 0 1 1
use contact_14  contact_14_60
timestamp 1643593061
transform 1 0 3416 0 1 14466
box 0 0 1 1
use contact_14  contact_14_61
timestamp 1643593061
transform 1 0 3164 0 1 14410
box 0 0 1 1
use contact_14  contact_14_62
timestamp 1643593061
transform 1 0 2912 0 1 14354
box 0 0 1 1
use contact_14  contact_14_63
timestamp 1643593061
transform 1 0 3416 0 1 14298
box 0 0 1 1
use contact_14  contact_14_64
timestamp 1643593061
transform 1 0 3164 0 1 14242
box 0 0 1 1
use contact_14  contact_14_65
timestamp 1643593061
transform 1 0 2828 0 1 14186
box 0 0 1 1
use contact_14  contact_14_66
timestamp 1643593061
transform 1 0 3416 0 1 12566
box 0 0 1 1
use contact_14  contact_14_67
timestamp 1643593061
transform 1 0 3164 0 1 12622
box 0 0 1 1
use contact_14  contact_14_68
timestamp 1643593061
transform 1 0 2744 0 1 12678
box 0 0 1 1
use contact_14  contact_14_69
timestamp 1643593061
transform 1 0 3416 0 1 12734
box 0 0 1 1
use contact_14  contact_14_70
timestamp 1643593061
transform 1 0 3164 0 1 12790
box 0 0 1 1
use contact_14  contact_14_71
timestamp 1643593061
transform 1 0 2660 0 1 12846
box 0 0 1 1
use contact_14  contact_14_72
timestamp 1643593061
transform 1 0 3416 0 1 12902
box 0 0 1 1
use contact_14  contact_14_73
timestamp 1643593061
transform 1 0 3080 0 1 12958
box 0 0 1 1
use contact_14  contact_14_74
timestamp 1643593061
transform 1 0 2912 0 1 13014
box 0 0 1 1
use contact_14  contact_14_75
timestamp 1643593061
transform 1 0 3416 0 1 11606
box 0 0 1 1
use contact_14  contact_14_76
timestamp 1643593061
transform 1 0 3080 0 1 11550
box 0 0 1 1
use contact_14  contact_14_77
timestamp 1643593061
transform 1 0 2828 0 1 11494
box 0 0 1 1
use contact_14  contact_14_78
timestamp 1643593061
transform 1 0 3416 0 1 11438
box 0 0 1 1
use contact_14  contact_14_79
timestamp 1643593061
transform 1 0 3080 0 1 11382
box 0 0 1 1
use contact_14  contact_14_80
timestamp 1643593061
transform 1 0 2744 0 1 11326
box 0 0 1 1
use contact_14  contact_14_81
timestamp 1643593061
transform 1 0 3416 0 1 11270
box 0 0 1 1
use contact_14  contact_14_82
timestamp 1643593061
transform 1 0 3080 0 1 11214
box 0 0 1 1
use contact_14  contact_14_83
timestamp 1643593061
transform 1 0 2660 0 1 11158
box 0 0 1 1
use contact_14  contact_14_84
timestamp 1643593061
transform 1 0 3416 0 1 9538
box 0 0 1 1
use contact_14  contact_14_85
timestamp 1643593061
transform 1 0 2996 0 1 9594
box 0 0 1 1
use contact_14  contact_14_86
timestamp 1643593061
transform 1 0 2912 0 1 9650
box 0 0 1 1
use contact_14  contact_14_87
timestamp 1643593061
transform 1 0 3416 0 1 9706
box 0 0 1 1
use contact_14  contact_14_88
timestamp 1643593061
transform 1 0 2996 0 1 9762
box 0 0 1 1
use contact_14  contact_14_89
timestamp 1643593061
transform 1 0 2828 0 1 9818
box 0 0 1 1
use contact_14  contact_14_90
timestamp 1643593061
transform 1 0 3416 0 1 9874
box 0 0 1 1
use contact_14  contact_14_91
timestamp 1643593061
transform 1 0 2996 0 1 9930
box 0 0 1 1
use contact_14  contact_14_92
timestamp 1643593061
transform 1 0 2744 0 1 9986
box 0 0 1 1
use contact_14  contact_14_93
timestamp 1643593061
transform 1 0 3416 0 1 8578
box 0 0 1 1
use contact_14  contact_14_94
timestamp 1643593061
transform 1 0 2996 0 1 8522
box 0 0 1 1
use contact_14  contact_14_95
timestamp 1643593061
transform 1 0 2660 0 1 8466
box 0 0 1 1
use contact_14  contact_14_96
timestamp 1643593061
transform 1 0 3332 0 1 8410
box 0 0 1 1
use contact_14  contact_14_97
timestamp 1643593061
transform 1 0 3248 0 1 8354
box 0 0 1 1
use contact_14  contact_14_98
timestamp 1643593061
transform 1 0 2912 0 1 8298
box 0 0 1 1
use contact_14  contact_14_99
timestamp 1643593061
transform 1 0 3332 0 1 8242
box 0 0 1 1
use contact_14  contact_14_100
timestamp 1643593061
transform 1 0 3248 0 1 8186
box 0 0 1 1
use contact_14  contact_14_101
timestamp 1643593061
transform 1 0 2828 0 1 8130
box 0 0 1 1
use contact_14  contact_14_102
timestamp 1643593061
transform 1 0 3332 0 1 6510
box 0 0 1 1
use contact_14  contact_14_103
timestamp 1643593061
transform 1 0 3248 0 1 6566
box 0 0 1 1
use contact_14  contact_14_104
timestamp 1643593061
transform 1 0 2744 0 1 6622
box 0 0 1 1
use contact_14  contact_14_105
timestamp 1643593061
transform 1 0 3332 0 1 6678
box 0 0 1 1
use contact_14  contact_14_106
timestamp 1643593061
transform 1 0 3248 0 1 6734
box 0 0 1 1
use contact_14  contact_14_107
timestamp 1643593061
transform 1 0 2660 0 1 6790
box 0 0 1 1
use contact_14  contact_14_108
timestamp 1643593061
transform 1 0 3332 0 1 6846
box 0 0 1 1
use contact_14  contact_14_109
timestamp 1643593061
transform 1 0 3164 0 1 6902
box 0 0 1 1
use contact_14  contact_14_110
timestamp 1643593061
transform 1 0 2912 0 1 6958
box 0 0 1 1
use contact_14  contact_14_111
timestamp 1643593061
transform 1 0 3332 0 1 5550
box 0 0 1 1
use contact_14  contact_14_112
timestamp 1643593061
transform 1 0 3164 0 1 5494
box 0 0 1 1
use contact_14  contact_14_113
timestamp 1643593061
transform 1 0 2828 0 1 5438
box 0 0 1 1
use contact_14  contact_14_114
timestamp 1643593061
transform 1 0 3332 0 1 5382
box 0 0 1 1
use contact_14  contact_14_115
timestamp 1643593061
transform 1 0 3164 0 1 5326
box 0 0 1 1
use contact_14  contact_14_116
timestamp 1643593061
transform 1 0 2744 0 1 5270
box 0 0 1 1
use contact_14  contact_14_117
timestamp 1643593061
transform 1 0 3332 0 1 5214
box 0 0 1 1
use contact_14  contact_14_118
timestamp 1643593061
transform 1 0 3164 0 1 5158
box 0 0 1 1
use contact_14  contact_14_119
timestamp 1643593061
transform 1 0 2660 0 1 5102
box 0 0 1 1
use contact_14  contact_14_120
timestamp 1643593061
transform 1 0 3332 0 1 3482
box 0 0 1 1
use contact_14  contact_14_121
timestamp 1643593061
transform 1 0 3080 0 1 3538
box 0 0 1 1
use contact_14  contact_14_122
timestamp 1643593061
transform 1 0 2912 0 1 3594
box 0 0 1 1
use contact_14  contact_14_123
timestamp 1643593061
transform 1 0 3332 0 1 3650
box 0 0 1 1
use contact_14  contact_14_124
timestamp 1643593061
transform 1 0 3080 0 1 3706
box 0 0 1 1
use contact_14  contact_14_125
timestamp 1643593061
transform 1 0 2828 0 1 3762
box 0 0 1 1
use contact_14  contact_14_126
timestamp 1643593061
transform 1 0 3332 0 1 3818
box 0 0 1 1
use contact_14  contact_14_127
timestamp 1643593061
transform 1 0 3080 0 1 3874
box 0 0 1 1
use contact_14  contact_14_128
timestamp 1643593061
transform 1 0 2744 0 1 3930
box 0 0 1 1
use contact_14  contact_14_129
timestamp 1643593061
transform 1 0 3332 0 1 2522
box 0 0 1 1
use contact_14  contact_14_130
timestamp 1643593061
transform 1 0 3080 0 1 2466
box 0 0 1 1
use contact_14  contact_14_131
timestamp 1643593061
transform 1 0 2660 0 1 2410
box 0 0 1 1
use contact_14  contact_14_132
timestamp 1643593061
transform 1 0 3332 0 1 2354
box 0 0 1 1
use contact_14  contact_14_133
timestamp 1643593061
transform 1 0 2996 0 1 2298
box 0 0 1 1
use contact_14  contact_14_134
timestamp 1643593061
transform 1 0 2912 0 1 2242
box 0 0 1 1
use contact_14  contact_14_135
timestamp 1643593061
transform 1 0 3332 0 1 2186
box 0 0 1 1
use contact_14  contact_14_136
timestamp 1643593061
transform 1 0 2996 0 1 2130
box 0 0 1 1
use contact_14  contact_14_137
timestamp 1643593061
transform 1 0 2828 0 1 2074
box 0 0 1 1
use contact_14  contact_14_138
timestamp 1643593061
transform 1 0 3332 0 1 454
box 0 0 1 1
use contact_14  contact_14_139
timestamp 1643593061
transform 1 0 2996 0 1 510
box 0 0 1 1
use contact_14  contact_14_140
timestamp 1643593061
transform 1 0 2744 0 1 566
box 0 0 1 1
use contact_14  contact_14_141
timestamp 1643593061
transform 1 0 3332 0 1 622
box 0 0 1 1
use contact_14  contact_14_142
timestamp 1643593061
transform 1 0 2996 0 1 678
box 0 0 1 1
use contact_14  contact_14_143
timestamp 1643593061
transform 1 0 2660 0 1 734
box 0 0 1 1
use contact_14  contact_14_144
timestamp 1643593061
transform 1 0 420 0 1 20798
box 0 0 1 1
use contact_17  contact_17_108
timestamp 1643593061
transform 1 0 700 0 1 20798
box 0 0 1 1
use contact_14  contact_14_145
timestamp 1643593061
transform 1 0 336 0 1 19174
box 0 0 1 1
use contact_17  contact_17_109
timestamp 1643593061
transform 1 0 616 0 1 19174
box 0 0 1 1
use contact_14  contact_14_146
timestamp 1643593061
transform 1 0 252 0 1 11562
box 0 0 1 1
use contact_17  contact_17_110
timestamp 1643593061
transform 1 0 700 0 1 11562
box 0 0 1 1
use contact_14  contact_14_147
timestamp 1643593061
transform 1 0 168 0 1 9938
box 0 0 1 1
use contact_17  contact_17_111
timestamp 1643593061
transform 1 0 616 0 1 9938
box 0 0 1 1
use contact_14  contact_14_148
timestamp 1643593061
transform 1 0 84 0 1 2326
box 0 0 1 1
use contact_17  contact_17_112
timestamp 1643593061
transform 1 0 700 0 1 2326
box 0 0 1 1
use contact_14  contact_14_149
timestamp 1643593061
transform 1 0 0 0 1 702
box 0 0 1 1
use contact_17  contact_17_113
timestamp 1643593061
transform 1 0 616 0 1 702
box 0 0 1 1
use dec_cell3_2r1w  dec_cell3_2r1w_0
timestamp 1643593061
transform 1 0 2594 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_1
timestamp 1643593061
transform 1 0 2594 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_2
timestamp 1643593061
transform 1 0 2594 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_3
timestamp 1643593061
transform 1 0 2594 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_4
timestamp 1643593061
transform 1 0 2594 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_5
timestamp 1643593061
transform 1 0 2594 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_6
timestamp 1643593061
transform 1 0 2594 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_7
timestamp 1643593061
transform 1 0 2594 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_8
timestamp 1643593061
transform 1 0 2594 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_9
timestamp 1643593061
transform 1 0 2594 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_10
timestamp 1643593061
transform 1 0 2594 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_11
timestamp 1643593061
transform 1 0 2594 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_12
timestamp 1643593061
transform 1 0 2594 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_13
timestamp 1643593061
transform 1 0 2594 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_14
timestamp 1643593061
transform 1 0 2594 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_15
timestamp 1643593061
transform 1 0 2594 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_16
timestamp 1643593061
transform 1 0 2594 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_17
timestamp 1643593061
transform 1 0 2594 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_18
timestamp 1643593061
transform 1 0 2594 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_19
timestamp 1643593061
transform 1 0 2594 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_20
timestamp 1643593061
transform 1 0 2594 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_21
timestamp 1643593061
transform 1 0 2594 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_22
timestamp 1643593061
transform 1 0 2594 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_23
timestamp 1643593061
transform 1 0 2594 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_24
timestamp 1643593061
transform 1 0 2594 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_25
timestamp 1643593061
transform 1 0 2594 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_26
timestamp 1643593061
transform 1 0 2594 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_27
timestamp 1643593061
transform 1 0 2594 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_28
timestamp 1643593061
transform 1 0 2594 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_29
timestamp 1643593061
transform 1 0 2594 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_30
timestamp 1643593061
transform 1 0 2594 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_31
timestamp 1643593061
transform 1 0 2594 0 1 0
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_32
timestamp 1643593061
transform 1 0 3686 0 -1 24224
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_33
timestamp 1643593061
transform 1 0 3686 0 1 21196
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_34
timestamp 1643593061
transform 1 0 3686 0 -1 21196
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_35
timestamp 1643593061
transform 1 0 3686 0 1 18168
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_36
timestamp 1643593061
transform 1 0 3686 0 -1 18168
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_37
timestamp 1643593061
transform 1 0 3686 0 1 15140
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_38
timestamp 1643593061
transform 1 0 3686 0 -1 15140
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_39
timestamp 1643593061
transform 1 0 3686 0 1 12112
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_40
timestamp 1643593061
transform 1 0 3686 0 -1 12112
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_41
timestamp 1643593061
transform 1 0 3686 0 1 9084
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_42
timestamp 1643593061
transform 1 0 3686 0 -1 9084
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_43
timestamp 1643593061
transform 1 0 3686 0 1 6056
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_44
timestamp 1643593061
transform 1 0 3686 0 -1 6056
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_45
timestamp 1643593061
transform 1 0 3686 0 1 3028
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_46
timestamp 1643593061
transform 1 0 3686 0 -1 3028
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_47
timestamp 1643593061
transform 1 0 3686 0 1 0
box 0 -42 1494 1616
use hierarchical_predecode2x4  hierarchical_predecode2x4_0
timestamp 1643593061
transform 1 0 550 0 1 18472
box 0 -30 2080 6190
use hierarchical_predecode2x4  hierarchical_predecode2x4_1
timestamp 1643593061
transform 1 0 550 0 1 9236
box 0 -30 2080 6190
use hierarchical_predecode2x4  hierarchical_predecode2x4_2
timestamp 1643593061
transform 1 0 550 0 1 0
box 0 -30 2080 6190
<< labels >>
rlabel metal2 s 18 0 46 24632 4 addr_0
rlabel metal2 s 102 0 130 24632 4 addr_1
rlabel metal2 s 186 0 214 24632 4 addr_2
rlabel metal2 s 270 0 298 24632 4 addr_3
rlabel metal2 s 354 0 382 24632 4 addr_4
rlabel metal2 s 438 0 466 24632 4 addr_5
rlabel metal1 s 4896 702 5180 730 4 decode0_0
rlabel metal1 s 5104 848 5180 876 4 decode1_0
rlabel metal1 s 4814 580 5180 608 4 decode2_0
rlabel metal1 s 4896 2298 5180 2326 4 decode0_1
rlabel metal1 s 5104 2152 5180 2180 4 decode1_1
rlabel metal1 s 4814 2420 5180 2448 4 decode2_1
rlabel metal1 s 4896 3730 5180 3758 4 decode0_2
rlabel metal1 s 5104 3876 5180 3904 4 decode1_2
rlabel metal1 s 4814 3608 5180 3636 4 decode2_2
rlabel metal1 s 4896 5326 5180 5354 4 decode0_3
rlabel metal1 s 5104 5180 5180 5208 4 decode1_3
rlabel metal1 s 4814 5448 5180 5476 4 decode2_3
rlabel metal1 s 4896 6758 5180 6786 4 decode0_4
rlabel metal1 s 5104 6904 5180 6932 4 decode1_4
rlabel metal1 s 4814 6636 5180 6664 4 decode2_4
rlabel metal1 s 4896 8354 5180 8382 4 decode0_5
rlabel metal1 s 5104 8208 5180 8236 4 decode1_5
rlabel metal1 s 4814 8476 5180 8504 4 decode2_5
rlabel metal1 s 4896 9786 5180 9814 4 decode0_6
rlabel metal1 s 5104 9932 5180 9960 4 decode1_6
rlabel metal1 s 4814 9664 5180 9692 4 decode2_6
rlabel metal1 s 4896 11382 5180 11410 4 decode0_7
rlabel metal1 s 5104 11236 5180 11264 4 decode1_7
rlabel metal1 s 4814 11504 5180 11532 4 decode2_7
rlabel metal1 s 4896 12814 5180 12842 4 decode0_8
rlabel metal1 s 5104 12960 5180 12988 4 decode1_8
rlabel metal1 s 4814 12692 5180 12720 4 decode2_8
rlabel metal1 s 4896 14410 5180 14438 4 decode0_9
rlabel metal1 s 5104 14264 5180 14292 4 decode1_9
rlabel metal1 s 4814 14532 5180 14560 4 decode2_9
rlabel metal1 s 4896 15842 5180 15870 4 decode0_10
rlabel metal1 s 5104 15988 5180 16016 4 decode1_10
rlabel metal1 s 4814 15720 5180 15748 4 decode2_10
rlabel metal1 s 4896 17438 5180 17466 4 decode0_11
rlabel metal1 s 5104 17292 5180 17320 4 decode1_11
rlabel metal1 s 4814 17560 5180 17588 4 decode2_11
rlabel metal1 s 4896 18870 5180 18898 4 decode0_12
rlabel metal1 s 5104 19016 5180 19044 4 decode1_12
rlabel metal1 s 4814 18748 5180 18776 4 decode2_12
rlabel metal1 s 4896 20466 5180 20494 4 decode0_13
rlabel metal1 s 5104 20320 5180 20348 4 decode1_13
rlabel metal1 s 4814 20588 5180 20616 4 decode2_13
rlabel metal1 s 4896 21898 5180 21926 4 decode0_14
rlabel metal1 s 5104 22044 5180 22072 4 decode1_14
rlabel metal1 s 4814 21776 5180 21804 4 decode2_14
rlabel metal1 s 4896 23494 5180 23522 4 decode0_15
rlabel metal1 s 5104 23348 5180 23376 4 decode1_15
rlabel metal1 s 4814 23616 5180 23644 4 decode2_15
rlabel metal2 s 2678 0 2706 24660 4 predecode_0
rlabel metal2 s 2762 0 2790 24660 4 predecode_1
rlabel metal2 s 2846 0 2874 24660 4 predecode_2
rlabel metal2 s 2930 0 2958 24660 4 predecode_3
rlabel metal2 s 3014 0 3042 24660 4 predecode_4
rlabel metal2 s 3098 0 3126 24660 4 predecode_5
rlabel metal2 s 3182 0 3210 24660 4 predecode_6
rlabel metal2 s 3266 0 3294 24660 4 predecode_7
rlabel metal2 s 3350 0 3378 24660 4 predecode_8
rlabel metal2 s 3434 0 3462 24660 4 predecode_9
rlabel metal2 s 3518 0 3546 24660 4 predecode_10
rlabel metal2 s 3602 0 3630 24660 4 predecode_11
rlabel metal3 s 1700 23062 1760 23122 4 vdd
rlabel metal3 s 828 10746 888 10806 4 vdd
rlabel metal3 s 5164 16624 5224 16684 4 vdd
rlabel metal3 s 5164 13596 5224 13656 4 vdd
rlabel metal3 s 1700 13826 1760 13886 4 vdd
rlabel metal3 s 1700 1510 1760 1570 4 vdd
rlabel metal3 s 828 13826 888 13886 4 vdd
rlabel metal3 s 828 23062 888 23122 4 vdd
rlabel metal3 s 828 1510 888 1570 4 vdd
rlabel metal3 s 1700 19982 1760 20042 4 vdd
rlabel metal3 s 1700 10746 1760 10806 4 vdd
rlabel metal3 s 5164 10568 5224 10628 4 vdd
rlabel metal3 s 5164 1484 5224 1544 4 vdd
rlabel metal3 s 5164 22680 5224 22740 4 vdd
rlabel metal3 s 828 4590 888 4650 4 vdd
rlabel metal3 s 5164 7540 5224 7600 4 vdd
rlabel metal3 s 5164 19652 5224 19712 4 vdd
rlabel metal3 s 5164 4512 5224 4572 4 vdd
rlabel metal3 s 1700 4590 1760 4650 4 vdd
rlabel metal3 s 828 19982 888 20042 4 vdd
rlabel metal3 s 1700 15366 1760 15426 4 gnd
rlabel metal3 s 828 24602 888 24662 4 gnd
rlabel metal3 s 828 21522 888 21582 4 gnd
rlabel metal3 s 1700 9206 1760 9266 4 gnd
rlabel metal3 s 5164 2998 5224 3058 4 gnd
rlabel metal3 s 1700 6130 1760 6190 4 gnd
rlabel metal3 s 828 18442 888 18502 4 gnd
rlabel metal3 s 5164 9054 5224 9114 4 gnd
rlabel metal3 s 828 3050 888 3110 4 gnd
rlabel metal3 s 828 12286 888 12346 4 gnd
rlabel metal3 s 5164 24194 5224 24254 4 gnd
rlabel metal3 s 5164 18138 5224 18198 4 gnd
rlabel metal3 s 1700 18442 1760 18502 4 gnd
rlabel metal3 s 1700 12286 1760 12346 4 gnd
rlabel metal3 s 5164 15110 5224 15170 4 gnd
rlabel metal3 s 828 15366 888 15426 4 gnd
rlabel metal3 s 5164 6026 5224 6086 4 gnd
rlabel metal3 s 5164 21166 5224 21226 4 gnd
rlabel metal3 s 1700 21522 1760 21582 4 gnd
rlabel metal3 s 828 -30 888 30 4 gnd
rlabel metal3 s 828 9206 888 9266 4 gnd
rlabel metal3 s 1700 -30 1760 30 4 gnd
rlabel metal3 s 1700 3050 1760 3110 4 gnd
rlabel metal3 s 828 6130 888 6190 4 gnd
rlabel metal3 s 5164 -30 5224 30 4 gnd
rlabel metal3 s 5164 12082 5224 12142 4 gnd
rlabel metal3 s 1700 24602 1760 24662 4 gnd
<< properties >>
string FIXED_BBOX 5164 -30 5224 -26
string GDS_FILE sram_0rw2r1w_2_16_sky130A.gds
string GDS_END 386616
string GDS_START 318150
<< end >>
