magic
tech sky130A
timestamp 1648462787
<< nwell >>
rect 0 362 389 1007
<< nmos >>
rect 54 195 69 237
rect 110 195 125 237
rect 264 69 279 237
rect 320 69 335 237
<< pmos >>
rect 54 380 69 515
rect 110 380 125 515
rect 264 380 279 920
rect 320 380 335 920
<< ndiff >>
rect 18 224 54 237
rect 18 207 25 224
rect 42 207 54 224
rect 18 195 54 207
rect 69 224 110 237
rect 69 207 81 224
rect 98 207 110 224
rect 69 195 110 207
rect 125 224 161 237
rect 125 207 137 224
rect 154 207 161 224
rect 125 195 161 207
rect 228 224 264 237
rect 228 207 235 224
rect 252 207 264 224
rect 228 183 264 207
rect 228 166 235 183
rect 252 166 264 183
rect 228 140 264 166
rect 228 123 235 140
rect 252 123 264 140
rect 228 99 264 123
rect 228 82 235 99
rect 252 82 264 99
rect 228 69 264 82
rect 279 69 320 237
rect 335 224 371 237
rect 335 207 347 224
rect 364 207 371 224
rect 335 183 371 207
rect 335 166 347 183
rect 364 166 371 183
rect 335 140 371 166
rect 335 123 347 140
rect 364 123 371 140
rect 335 99 371 123
rect 335 82 347 99
rect 364 82 371 99
rect 335 69 371 82
<< pdiff >>
rect 228 898 264 920
rect 228 881 235 898
rect 252 881 264 898
rect 228 858 264 881
rect 228 841 235 858
rect 252 841 264 858
rect 228 818 264 841
rect 228 801 235 818
rect 252 801 264 818
rect 228 778 264 801
rect 228 761 235 778
rect 252 761 264 778
rect 228 738 264 761
rect 228 721 235 738
rect 252 721 264 738
rect 228 698 264 721
rect 228 681 235 698
rect 252 681 264 698
rect 228 658 264 681
rect 228 641 235 658
rect 252 641 264 658
rect 228 618 264 641
rect 228 601 235 618
rect 252 601 264 618
rect 228 578 264 601
rect 228 561 235 578
rect 252 561 264 578
rect 228 538 264 561
rect 228 521 235 538
rect 252 521 264 538
rect 18 494 54 515
rect 18 477 25 494
rect 42 477 54 494
rect 18 456 54 477
rect 18 439 25 456
rect 42 439 54 456
rect 18 418 54 439
rect 18 401 25 418
rect 42 401 54 418
rect 18 380 54 401
rect 69 494 110 515
rect 69 477 81 494
rect 98 477 110 494
rect 69 456 110 477
rect 69 439 81 456
rect 98 439 110 456
rect 69 418 110 439
rect 69 401 81 418
rect 98 401 110 418
rect 69 380 110 401
rect 125 494 161 515
rect 125 477 137 494
rect 154 477 161 494
rect 125 456 161 477
rect 125 439 137 456
rect 154 439 161 456
rect 125 418 161 439
rect 125 401 137 418
rect 154 401 161 418
rect 125 380 161 401
rect 228 498 264 521
rect 228 481 235 498
rect 252 481 264 498
rect 228 458 264 481
rect 228 441 235 458
rect 252 441 264 458
rect 228 418 264 441
rect 228 401 235 418
rect 252 401 264 418
rect 228 380 264 401
rect 279 380 320 920
rect 335 898 371 920
rect 335 881 347 898
rect 364 881 371 898
rect 335 858 371 881
rect 335 841 347 858
rect 364 841 371 858
rect 335 818 371 841
rect 335 801 347 818
rect 364 801 371 818
rect 335 778 371 801
rect 335 761 347 778
rect 364 761 371 778
rect 335 738 371 761
rect 335 721 347 738
rect 364 721 371 738
rect 335 698 371 721
rect 335 681 347 698
rect 364 681 371 698
rect 335 658 371 681
rect 335 641 347 658
rect 364 641 371 658
rect 335 618 371 641
rect 335 601 347 618
rect 364 601 371 618
rect 335 578 371 601
rect 335 561 347 578
rect 364 561 371 578
rect 335 538 371 561
rect 335 521 347 538
rect 364 521 371 538
rect 335 498 371 521
rect 335 481 347 498
rect 364 481 371 498
rect 335 458 371 481
rect 335 441 347 458
rect 364 441 371 458
rect 335 418 371 441
rect 335 401 347 418
rect 364 401 371 418
rect 335 380 371 401
<< ndiffc >>
rect 25 207 42 224
rect 81 207 98 224
rect 137 207 154 224
rect 235 207 252 224
rect 235 166 252 183
rect 235 123 252 140
rect 235 82 252 99
rect 347 207 364 224
rect 347 166 364 183
rect 347 123 364 140
rect 347 82 364 99
<< pdiffc >>
rect 235 881 252 898
rect 235 841 252 858
rect 235 801 252 818
rect 235 761 252 778
rect 235 721 252 738
rect 235 681 252 698
rect 235 641 252 658
rect 235 601 252 618
rect 235 561 252 578
rect 235 521 252 538
rect 25 477 42 494
rect 25 439 42 456
rect 25 401 42 418
rect 81 477 98 494
rect 81 439 98 456
rect 81 401 98 418
rect 137 477 154 494
rect 137 439 154 456
rect 137 401 154 418
rect 235 481 252 498
rect 235 441 252 458
rect 235 401 252 418
rect 347 881 364 898
rect 347 841 364 858
rect 347 801 364 818
rect 347 761 364 778
rect 347 721 364 738
rect 347 681 364 698
rect 347 641 364 658
rect 347 601 364 618
rect 347 561 364 578
rect 347 521 364 538
rect 347 481 364 498
rect 347 441 364 458
rect 347 401 364 418
<< psubdiff >>
rect 81 30 117 42
rect 81 12 90 30
rect 108 12 117 30
rect 81 0 117 12
rect 177 30 213 42
rect 177 12 186 30
rect 204 12 213 30
rect 177 0 213 12
rect 273 30 309 42
rect 273 12 282 30
rect 300 12 309 30
rect 273 0 309 12
<< nsubdiff >>
rect 81 977 117 989
rect 81 959 90 977
rect 108 959 117 977
rect 81 947 117 959
rect 177 977 213 989
rect 177 959 186 977
rect 204 959 213 977
rect 177 947 213 959
rect 273 977 309 989
rect 273 959 282 977
rect 300 959 309 977
rect 273 947 309 959
<< psubdiffcont >>
rect 90 12 108 30
rect 186 12 204 30
rect 282 12 300 30
<< nsubdiffcont >>
rect 90 959 108 977
rect 186 959 204 977
rect 282 959 300 977
<< poly >>
rect 264 920 279 933
rect 320 920 335 933
rect 54 515 69 528
rect 110 515 125 528
rect 54 329 69 380
rect 4 321 69 329
rect 4 304 9 321
rect 26 314 69 321
rect 26 304 31 314
rect 4 296 31 304
rect 54 237 69 314
rect 110 287 125 380
rect 264 363 279 380
rect 320 363 335 380
rect 252 355 279 363
rect 252 338 257 355
rect 274 338 279 355
rect 252 330 279 338
rect 308 355 335 363
rect 308 338 313 355
rect 330 338 335 355
rect 308 330 335 338
rect 98 279 125 287
rect 98 262 103 279
rect 120 262 125 279
rect 98 254 125 262
rect 110 237 125 254
rect 264 237 279 330
rect 308 279 335 287
rect 308 262 313 279
rect 330 262 335 279
rect 308 254 335 262
rect 320 237 335 254
rect 54 182 69 195
rect 110 182 125 195
rect 264 56 279 69
rect 320 56 335 69
<< polycont >>
rect 9 304 26 321
rect 257 338 274 355
rect 313 338 330 355
rect 103 262 120 279
rect 313 262 330 279
<< locali >>
rect 88 977 108 985
rect 88 959 90 977
rect 88 951 108 959
rect 186 977 204 985
rect 282 977 300 985
rect 204 959 245 968
rect 186 951 245 959
rect 282 951 300 959
rect 88 515 105 951
rect 228 920 245 951
rect 228 898 259 920
rect 228 881 235 898
rect 252 881 259 898
rect 228 858 259 881
rect 228 841 235 858
rect 252 841 259 858
rect 228 818 259 841
rect 228 801 235 818
rect 252 801 259 818
rect 228 778 259 801
rect 228 761 235 778
rect 252 761 259 778
rect 228 738 259 761
rect 228 721 235 738
rect 252 721 259 738
rect 228 698 259 721
rect 228 681 235 698
rect 252 681 259 698
rect 228 658 259 681
rect 228 641 235 658
rect 252 641 259 658
rect 228 618 259 641
rect 228 601 235 618
rect 252 601 259 618
rect 228 578 259 601
rect 228 561 235 578
rect 252 561 259 578
rect 228 538 259 561
rect 228 521 235 538
rect 252 521 259 538
rect 18 494 49 515
rect 18 477 25 494
rect 42 477 49 494
rect 18 456 49 477
rect 18 439 25 456
rect 42 439 49 456
rect 18 418 49 439
rect 18 401 25 418
rect 42 401 49 418
rect 18 380 49 401
rect 74 494 105 515
rect 74 477 81 494
rect 98 477 105 494
rect 74 456 105 477
rect 74 439 81 456
rect 98 439 105 456
rect 74 418 105 439
rect 74 401 81 418
rect 98 401 105 418
rect 74 380 105 401
rect 130 494 161 515
rect 130 477 137 494
rect 154 477 161 494
rect 130 456 161 477
rect 130 439 137 456
rect 154 439 161 456
rect 130 418 161 439
rect 130 401 137 418
rect 154 401 161 418
rect 130 380 161 401
rect 228 498 259 521
rect 228 481 235 498
rect 252 481 259 498
rect 228 458 259 481
rect 228 441 235 458
rect 252 441 259 458
rect 228 418 259 441
rect 228 401 235 418
rect 252 401 259 418
rect 228 380 259 401
rect 340 898 371 920
rect 340 881 347 898
rect 364 881 371 898
rect 340 858 371 881
rect 340 841 347 858
rect 364 841 371 858
rect 340 818 371 841
rect 340 801 347 818
rect 364 801 371 818
rect 340 778 371 801
rect 340 761 347 778
rect 364 761 371 778
rect 340 738 371 761
rect 340 721 347 738
rect 364 721 371 738
rect 340 698 371 721
rect 340 681 347 698
rect 364 681 371 698
rect 340 658 371 681
rect 340 641 347 658
rect 364 641 371 658
rect 340 618 371 641
rect 340 601 347 618
rect 364 601 371 618
rect 340 578 371 601
rect 340 561 347 578
rect 364 561 371 578
rect 340 538 371 561
rect 340 521 347 538
rect 364 521 371 538
rect 340 498 371 521
rect 340 481 347 498
rect 364 481 371 498
rect 340 458 371 481
rect 340 441 347 458
rect 364 441 371 458
rect 340 418 371 441
rect 340 401 347 418
rect 364 401 371 418
rect 340 380 371 401
rect 32 363 49 380
rect 32 346 69 363
rect 9 321 26 329
rect 9 296 26 304
rect 52 273 69 346
rect 144 356 161 380
rect 257 356 274 363
rect 144 355 274 356
rect 144 338 257 355
rect 32 255 69 273
rect 103 279 120 287
rect 32 237 49 255
rect 103 254 120 262
rect 144 237 161 338
rect 257 330 274 338
rect 313 355 330 363
rect 313 330 330 338
rect 313 279 330 287
rect 313 254 330 262
rect 354 279 371 380
rect 354 237 371 262
rect 18 224 49 237
rect 18 207 25 224
rect 42 207 49 224
rect 18 195 49 207
rect 74 224 105 237
rect 74 207 81 224
rect 98 207 105 224
rect 74 195 105 207
rect 130 224 161 237
rect 130 207 137 224
rect 154 207 161 224
rect 130 195 161 207
rect 228 224 259 237
rect 228 207 235 224
rect 252 207 259 224
rect 88 38 105 195
rect 228 183 259 207
rect 228 166 235 183
rect 252 166 259 183
rect 228 140 259 166
rect 228 123 235 140
rect 252 123 259 140
rect 228 99 259 123
rect 228 82 235 99
rect 252 82 259 99
rect 228 69 259 82
rect 340 224 371 237
rect 340 207 347 224
rect 364 207 371 224
rect 340 183 371 207
rect 340 166 347 183
rect 364 166 371 183
rect 340 140 371 166
rect 340 123 347 140
rect 364 123 371 140
rect 340 99 371 123
rect 340 82 347 99
rect 364 82 371 99
rect 340 69 371 82
rect 228 38 245 69
rect 88 30 108 38
rect 88 12 90 30
rect 88 4 108 12
rect 186 30 245 38
rect 204 21 245 30
rect 282 30 300 38
rect 186 4 204 12
rect 282 4 300 12
<< viali >>
rect 90 959 108 977
rect 186 959 204 977
rect 282 959 300 977
rect 25 401 42 418
rect 9 304 26 321
rect 103 262 120 279
rect 313 338 330 355
rect 313 262 330 279
rect 354 262 371 279
rect 90 12 108 30
rect 186 12 204 30
rect 282 12 300 30
<< metal1 >>
rect 0 977 389 983
rect 0 959 90 977
rect 108 959 186 977
rect 204 959 282 977
rect 300 959 389 977
rect 0 953 389 959
rect 22 418 45 424
rect 22 401 25 418
rect 42 409 45 418
rect 42 401 324 409
rect 22 395 324 401
rect 310 361 324 395
rect 310 355 333 361
rect 310 338 313 355
rect 330 338 333 355
rect 310 332 333 338
rect 5 321 31 328
rect 5 318 9 321
rect 4 304 9 318
rect 26 318 31 321
rect 26 304 241 318
rect 5 296 31 304
rect 98 283 125 286
rect 98 257 99 283
rect 227 285 241 304
rect 227 279 333 285
rect 227 271 313 279
rect 98 254 125 257
rect 310 262 313 271
rect 330 262 333 279
rect 310 256 333 262
rect 349 284 375 287
rect 349 255 375 258
rect 0 30 389 36
rect 0 12 90 30
rect 108 12 186 30
rect 204 12 282 30
rect 300 12 389 30
rect 0 6 389 12
<< via1 >>
rect 99 279 125 283
rect 99 262 103 279
rect 103 262 120 279
rect 120 262 125 279
rect 99 257 125 262
rect 349 279 375 284
rect 349 262 354 279
rect 354 262 371 279
rect 371 262 375 279
rect 349 258 375 262
<< metal2 >>
rect 355 287 369 1007
rect 99 283 125 286
rect 98 262 99 276
rect 99 254 125 257
rect 349 284 375 287
rect 349 255 375 258
rect 355 0 369 255
<< labels >>
flabel metal2 98 269 98 269 0 FreeSans 80 0 0 0 din
port 1 nsew
flabel locali 38 261 38 261 0 FreeSans 80 0 0 0 enb
flabel locali 153 284 153 284 0 FreeSans 80 0 0 0 net1
flabel metal1 4 310 4 310 0 FreeSans 80 0 0 0 en
port 5 nsew
flabel metal2 361 310 361 310 0 FreeSans 80 0 0 0 wbl
port 6 nsew
flabel ndiff 298 213 298 213 0 FreeSans 80 0 0 0 net3
flabel pdiff 300 458 300 458 0 FreeSans 80 0 0 0 net2
flabel metal1 144 20 144 20 0 FreeSans 80 0 0 0 gnd
port 4 nsew
flabel metal1 144 968 144 968 0 FreeSans 80 0 0 0 vdd
port 3 nsew
<< properties >>
string FIXED_BBOX 0 0 389 1007
<< end >>
