magic
tech sky130A
magscale 1 2
timestamp 1643671299
<< checkpaint >>
rect -1296 -1277 3807 2155
<< nwell >>
rect -36 402 2547 895
<< locali >>
rect 0 821 2511 855
rect 48 338 114 404
rect 1261 354 1295 388
rect 0 -17 2511 17
use pinv_11  pinv_11_0
timestamp 1643671299
transform 1 0 0 0 1 0
box -36 -17 2547 895
<< labels >>
rlabel locali s 1278 371 1278 371 4 Z
rlabel locali s 81 371 81 371 4 A
rlabel locali s 1255 0 1255 0 4 gnd
rlabel locali s 1255 838 1255 838 4 vdd
<< properties >>
string FIXED_BBOX 0 0 2511 838
string GDS_FILE sram_0rw2r1w_16_32_sky130A.gds
string GDS_END 1197762
string GDS_START 1196916
<< end >>
