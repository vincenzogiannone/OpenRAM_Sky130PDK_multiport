magic
tech sky130A
magscale 1 2
timestamp 1644969367
<< checkpaint >>
rect -1296 -1277 8144 2155
<< nwell >>
rect -36 402 6884 895
<< pwell >>
rect 6738 51 6788 133
<< psubdiff >>
rect 6738 109 6788 133
rect 6738 75 6746 109
rect 6780 75 6788 109
rect 6738 51 6788 75
<< nsubdiff >>
rect 6738 763 6788 787
rect 6738 729 6746 763
rect 6780 729 6788 763
rect 6738 705 6788 729
<< psubdiffcont >>
rect 6746 75 6780 109
<< nsubdiffcont >>
rect 6746 729 6780 763
<< poly >>
rect 114 402 144 434
rect 48 386 144 402
rect 48 352 64 386
rect 98 352 144 386
rect 48 336 144 352
rect 114 206 144 336
<< polycont >>
rect 64 352 98 386
<< locali >>
rect 0 821 6848 855
rect 62 606 96 821
rect 274 606 308 821
rect 490 606 524 821
rect 706 606 740 821
rect 922 606 956 821
rect 1138 606 1172 821
rect 1354 606 1388 821
rect 1570 606 1604 821
rect 1786 606 1820 821
rect 2002 606 2036 821
rect 2218 606 2252 821
rect 2434 606 2468 821
rect 2650 606 2684 821
rect 2866 606 2900 821
rect 3082 606 3116 821
rect 3298 606 3332 821
rect 3514 606 3548 821
rect 3730 606 3764 821
rect 3946 606 3980 821
rect 4162 606 4196 821
rect 4378 606 4412 821
rect 4594 606 4628 821
rect 4810 606 4844 821
rect 5026 606 5060 821
rect 5242 606 5276 821
rect 5458 606 5492 821
rect 5674 606 5708 821
rect 5890 606 5924 821
rect 6106 606 6140 821
rect 6322 606 6356 821
rect 6538 606 6572 821
rect 6746 763 6780 821
rect 6746 713 6780 729
rect 48 386 114 402
rect 48 352 64 386
rect 98 352 114 386
rect 48 336 114 352
rect 3404 386 3438 572
rect 3404 352 3455 386
rect 3404 167 3438 352
rect 6746 109 6780 125
rect 62 17 96 67
rect 274 17 308 67
rect 490 17 524 67
rect 706 17 740 67
rect 922 17 956 67
rect 1138 17 1172 67
rect 1354 17 1388 67
rect 1570 17 1604 67
rect 1786 17 1820 67
rect 2002 17 2036 67
rect 2218 17 2252 67
rect 2434 17 2468 67
rect 2650 17 2684 67
rect 2866 17 2900 67
rect 3082 17 3116 67
rect 3298 17 3332 67
rect 3514 17 3548 67
rect 3730 17 3764 67
rect 3946 17 3980 67
rect 4162 17 4196 67
rect 4378 17 4412 67
rect 4594 17 4628 67
rect 4810 17 4844 67
rect 5026 17 5060 67
rect 5242 17 5276 67
rect 5458 17 5492 67
rect 5674 17 5708 67
rect 5890 17 5924 67
rect 6106 17 6140 67
rect 6322 17 6356 67
rect 6538 17 6572 67
rect 6746 17 6780 75
rect 0 -17 6848 17
use contact_12  contact_12_0
timestamp 1644969367
transform 1 0 48 0 1 336
box 0 0 1 1
use contact_11  contact_11_0
timestamp 1644969367
transform 1 0 6738 0 1 51
box 0 0 1 1
use contact_10  contact_10_0
timestamp 1644969367
transform 1 0 6738 0 1 705
box 0 0 1 1
use nmos_m61_w0_495_sli_dli_da_p  nmos_m61_w0_495_sli_dli_da_p_0
timestamp 1644969367
transform 1 0 54 0 1 51
box 0 -26 6630 155
use pmos_m61_w1_485_sli_dli_da_p  pmos_m61_w1_485_sli_dli_da_p_0
timestamp 1644969367
transform 1 0 54 0 1 490
box -59 -56 6689 351
<< labels >>
rlabel locali s 81 369 81 369 4 A
rlabel locali s 3438 369 3438 369 4 Z
rlabel locali s 3424 0 3424 0 4 gnd
rlabel locali s 3424 838 3424 838 4 vdd
<< properties >>
string FIXED_BBOX 0 0 6848 838
string GDS_FILE sram_0rw2r1w_32_128_sky130A.gds
string GDS_END 3335020
string GDS_START 3329688
<< end >>
