magic
tech sky130A
magscale 1 2
timestamp 1643593061
<< checkpaint >>
rect -1260 -1022 8096 5056
<< metal1 >>
rect 0 3412 1476 3440
rect 0 1251 2334 1279
<< metal2 >>
rect 196 3496 250 3524
rect 974 3496 1028 3524
rect 630 2844 658 3474
rect 4750 2352 4778 2592
rect 5210 2352 5238 2592
rect 70 252 98 1290
rect 532 252 560 1290
rect 848 252 876 1290
rect 1310 252 1338 1290
<< metal3 >>
rect 319 3724 379 3784
rect 1097 3724 1157 3784
rect 319 2892 379 2952
rect 1097 2892 1157 2952
rect 4654 2528 4714 2588
rect 5114 2528 5174 2588
rect 6210 2528 6270 2588
rect 6670 2528 6730 2588
rect 4654 1582 4714 1642
rect 5114 1582 5174 1642
rect 6210 1582 6270 1642
rect 6670 1582 6730 1642
rect 163 332 223 392
rect 941 332 1001 392
rect 1719 332 1779 392
use write_driver_array  write_driver_array_0
timestamp 1643593061
transform 1 0 0 0 -1 3796
box 0 0 1476 952
use sense_amp_array  sense_amp_array_0
timestamp 1643593061
transform 1 0 0 0 -1 2592
box 4548 0 6836 1050
use precharge_array_multiport  precharge_array_multiport_0
timestamp 1643593061
transform 1 0 0 0 -1 1290
box 0 -8 2334 1052
<< labels >>
rlabel metal2 s 196 3496 250 3524 4 din0_0
rlabel metal2 s 974 3496 1028 3524 4 din0_1
rlabel metal2 s 4750 2352 4778 2592 4 dout0_0
rlabel metal2 s 4764 2472 4764 2472 4 dout1_0
rlabel metal2 s 5210 2352 5238 2592 4 dout0_1
rlabel metal2 s 5224 2472 5224 2472 4 dout1_1
rlabel metal2 s 70 252 98 1290 4 rbl0_0
rlabel metal2 s 532 252 560 1290 4 rbl1_0
rlabel metal2 s 848 252 876 1290 4 rbl0_1
rlabel metal2 s 1310 252 1338 1290 4 rbl1_1
rlabel metal2 s 630 2844 658 3474 4 wbl0_0
rlabel metal1 s 0 1250 2334 1278 4 p_en_bar
rlabel metal1 s 0 3412 1476 3440 4 w_en
rlabel metal3 s 5114 1582 5174 1642 4 vdd
rlabel metal3 s 4654 1582 4714 1642 4 vdd
rlabel metal3 s 318 2892 378 2952 4 vdd
rlabel metal3 s 1718 332 1778 392 4 vdd
rlabel metal3 s 162 332 222 392 4 vdd
rlabel metal3 s 6670 1582 6730 1642 4 vdd
rlabel metal3 s 6210 1582 6270 1642 4 vdd
rlabel metal3 s 1096 2892 1156 2952 4 vdd
rlabel metal3 s 940 332 1000 392 4 vdd
rlabel metal3 s 5114 2528 5174 2588 4 gnd
rlabel metal3 s 6210 2528 6270 2588 4 gnd
rlabel metal3 s 6670 2528 6730 2588 4 gnd
rlabel metal3 s 4654 2528 4714 2588 4 gnd
rlabel metal3 s 318 3724 378 3784 4 gnd
rlabel metal3 s 1096 3724 1156 3784 4 gnd
<< properties >>
string FIXED_BBOX 0 0 6836 3796
string GDS_FILE sram_0rw2r1w_2_16_sky130A.gds
string GDS_END 242100
string GDS_START 236576
<< end >>
