magic
tech sky130A
magscale 1 2
timestamp 1644969367
<< checkpaint >>
rect -1260 -1297 3772 13617
<< locali >>
rect 0 12303 375 12337
rect 409 12303 1415 12337
rect 1449 12303 2476 12337
rect 2287 11575 2321 11609
rect 0 10763 375 10797
rect 409 10763 1415 10797
rect 1449 10763 2476 10797
rect 2287 9951 2321 9985
rect 0 9223 375 9257
rect 409 9223 1415 9257
rect 1449 9223 2476 9257
rect 2287 8495 2321 8529
rect 0 7683 375 7717
rect 409 7683 1415 7717
rect 1449 7683 2476 7717
rect 2287 6871 2321 6905
rect 0 6143 375 6177
rect 409 6143 1415 6177
rect 1449 6143 2476 6177
rect 2287 5415 2321 5449
rect 0 4603 375 4637
rect 409 4603 1415 4637
rect 1449 4603 2476 4637
rect 2287 3791 2321 3825
rect 0 3063 375 3097
rect 409 3063 1415 3097
rect 1449 3063 2476 3097
rect 2287 2335 2321 2369
rect 0 1523 375 1557
rect 409 1523 1415 1557
rect 1449 1523 2476 1557
rect 2287 711 2321 745
rect 0 -17 375 17
rect 409 -17 1415 17
rect 1449 -17 2476 17
<< viali >>
rect 375 12303 409 12337
rect 1415 12303 1449 12337
rect 1539 12013 1573 12047
rect 1672 11889 1706 11923
rect 1805 11765 1839 11799
rect 375 10763 409 10797
rect 1415 10763 1449 10797
rect 1805 9761 1839 9795
rect 1672 9637 1706 9671
rect 1539 9513 1573 9547
rect 375 9223 409 9257
rect 1415 9223 1449 9257
rect 1539 8933 1573 8967
rect 1672 8809 1706 8843
rect 1805 8685 1839 8719
rect 375 7683 409 7717
rect 1415 7683 1449 7717
rect 1805 6681 1839 6715
rect 1672 6557 1706 6591
rect 1539 6433 1573 6467
rect 375 6143 409 6177
rect 1415 6143 1449 6177
rect 1539 5853 1573 5887
rect 1672 5729 1706 5763
rect 1805 5605 1839 5639
rect 375 4603 409 4637
rect 1415 4603 1449 4637
rect 484 3791 518 3825
rect 616 3791 650 3825
rect 1805 3601 1839 3635
rect 1672 3477 1706 3511
rect 1539 3353 1573 3387
rect 375 3063 409 3097
rect 1415 3063 1449 3097
rect 1539 2773 1573 2807
rect 1672 2649 1706 2683
rect 1805 2525 1839 2559
rect 484 2335 518 2369
rect 616 2335 650 2369
rect 375 1523 409 1557
rect 1415 1523 1449 1557
rect 484 711 518 745
rect 616 711 650 745
rect 1805 521 1839 555
rect 1672 397 1706 431
rect 1539 273 1573 307
rect 375 -17 409 17
rect 1415 -17 1449 17
<< metal1 >>
rect 360 12294 366 12346
rect 418 12294 424 12346
rect 1400 12294 1406 12346
rect 1458 12294 1464 12346
rect 66 12004 72 12056
rect 124 12044 130 12056
rect 1106 12044 1112 12056
rect 124 12016 1112 12044
rect 124 12004 130 12016
rect 1106 12004 1112 12016
rect 1164 12044 1170 12056
rect 1527 12047 1585 12053
rect 1527 12044 1539 12047
rect 1164 12016 1539 12044
rect 1164 12004 1170 12016
rect 1527 12013 1539 12016
rect 1573 12013 1585 12047
rect 1527 12007 1585 12013
rect 150 11880 156 11932
rect 208 11920 214 11932
rect 1190 11920 1196 11932
rect 208 11892 1196 11920
rect 208 11880 214 11892
rect 1190 11880 1196 11892
rect 1248 11920 1254 11932
rect 1660 11923 1718 11929
rect 1660 11920 1672 11923
rect 1248 11892 1672 11920
rect 1248 11880 1254 11892
rect 1660 11889 1672 11892
rect 1706 11889 1718 11923
rect 1660 11883 1718 11889
rect 234 11756 240 11808
rect 292 11796 298 11808
rect 1274 11796 1280 11808
rect 292 11768 1280 11796
rect 292 11756 298 11768
rect 1274 11756 1280 11768
rect 1332 11796 1338 11808
rect 1793 11799 1851 11805
rect 1793 11796 1805 11799
rect 1332 11768 1805 11796
rect 1332 11756 1338 11768
rect 1793 11765 1805 11768
rect 1839 11765 1851 11799
rect 1793 11759 1851 11765
rect 360 10754 366 10806
rect 418 10754 424 10806
rect 1400 10754 1406 10806
rect 1458 10754 1464 10806
rect 1274 9752 1280 9804
rect 1332 9792 1338 9804
rect 1793 9795 1851 9801
rect 1793 9792 1805 9795
rect 1332 9764 1805 9792
rect 1332 9752 1338 9764
rect 1793 9761 1805 9764
rect 1839 9761 1851 9795
rect 1793 9755 1851 9761
rect 1190 9628 1196 9680
rect 1248 9668 1254 9680
rect 1660 9671 1718 9677
rect 1660 9668 1672 9671
rect 1248 9640 1672 9668
rect 1248 9628 1254 9640
rect 1660 9637 1672 9640
rect 1706 9637 1718 9671
rect 1660 9631 1718 9637
rect 854 9504 860 9556
rect 912 9544 918 9556
rect 1527 9547 1585 9553
rect 1527 9544 1539 9547
rect 912 9516 1539 9544
rect 912 9504 918 9516
rect 1527 9513 1539 9516
rect 1573 9513 1585 9547
rect 1527 9507 1585 9513
rect 360 9214 366 9266
rect 418 9214 424 9266
rect 1400 9214 1406 9266
rect 1458 9214 1464 9266
rect 1106 8924 1112 8976
rect 1164 8964 1170 8976
rect 1527 8967 1585 8973
rect 1527 8964 1539 8967
rect 1164 8936 1539 8964
rect 1164 8924 1170 8936
rect 1527 8933 1539 8936
rect 1573 8933 1585 8967
rect 1527 8927 1585 8933
rect 938 8800 944 8852
rect 996 8840 1002 8852
rect 1660 8843 1718 8849
rect 1660 8840 1672 8843
rect 996 8812 1672 8840
rect 996 8800 1002 8812
rect 1660 8809 1672 8812
rect 1706 8809 1718 8843
rect 1660 8803 1718 8809
rect 1274 8676 1280 8728
rect 1332 8716 1338 8728
rect 1793 8719 1851 8725
rect 1793 8716 1805 8719
rect 1332 8688 1805 8716
rect 1332 8676 1338 8688
rect 1793 8685 1805 8688
rect 1839 8685 1851 8719
rect 1793 8679 1851 8685
rect 360 7674 366 7726
rect 418 7674 424 7726
rect 1400 7674 1406 7726
rect 1458 7674 1464 7726
rect 1274 6672 1280 6724
rect 1332 6712 1338 6724
rect 1793 6715 1851 6721
rect 1793 6712 1805 6715
rect 1332 6684 1805 6712
rect 1332 6672 1338 6684
rect 1793 6681 1805 6684
rect 1839 6681 1851 6715
rect 1793 6675 1851 6681
rect 938 6548 944 6600
rect 996 6588 1002 6600
rect 1660 6591 1718 6597
rect 1660 6588 1672 6591
rect 996 6560 1672 6588
rect 996 6548 1002 6560
rect 1660 6557 1672 6560
rect 1706 6557 1718 6591
rect 1660 6551 1718 6557
rect 854 6424 860 6476
rect 912 6464 918 6476
rect 1527 6467 1585 6473
rect 1527 6464 1539 6467
rect 912 6436 1539 6464
rect 912 6424 918 6436
rect 1527 6433 1539 6436
rect 1573 6433 1585 6467
rect 1527 6427 1585 6433
rect 360 6134 366 6186
rect 418 6134 424 6186
rect 1400 6134 1406 6186
rect 1458 6134 1464 6186
rect 1106 5844 1112 5896
rect 1164 5884 1170 5896
rect 1527 5887 1585 5893
rect 1527 5884 1539 5887
rect 1164 5856 1539 5884
rect 1164 5844 1170 5856
rect 1527 5853 1539 5856
rect 1573 5853 1585 5887
rect 1527 5847 1585 5853
rect 1190 5720 1196 5772
rect 1248 5760 1254 5772
rect 1660 5763 1718 5769
rect 1660 5760 1672 5763
rect 1248 5732 1672 5760
rect 1248 5720 1254 5732
rect 1660 5729 1672 5732
rect 1706 5729 1718 5763
rect 1660 5723 1718 5729
rect 1022 5596 1028 5648
rect 1080 5636 1086 5648
rect 1793 5639 1851 5645
rect 1793 5636 1805 5639
rect 1080 5608 1805 5636
rect 1080 5596 1086 5608
rect 1793 5605 1805 5608
rect 1839 5605 1851 5639
rect 1793 5599 1851 5605
rect 360 4594 366 4646
rect 418 4594 424 4646
rect 1400 4594 1406 4646
rect 1458 4594 1464 4646
rect 1022 4554 1028 4566
rect 774 4526 1028 4554
rect 234 3782 240 3834
rect 292 3822 298 3834
rect 472 3825 530 3831
rect 472 3822 484 3825
rect 292 3794 484 3822
rect 292 3782 298 3794
rect 472 3791 484 3794
rect 518 3791 530 3825
rect 472 3785 530 3791
rect 604 3825 662 3831
rect 604 3791 616 3825
rect 650 3822 662 3825
rect 774 3822 802 4526
rect 1022 4514 1028 4526
rect 1080 4514 1086 4566
rect 650 3794 802 3822
rect 650 3791 662 3794
rect 604 3785 662 3791
rect 1022 3592 1028 3644
rect 1080 3632 1086 3644
rect 1793 3635 1851 3641
rect 1793 3632 1805 3635
rect 1080 3604 1805 3632
rect 1080 3592 1086 3604
rect 1793 3601 1805 3604
rect 1839 3601 1851 3635
rect 1793 3595 1851 3601
rect 1190 3468 1196 3520
rect 1248 3508 1254 3520
rect 1660 3511 1718 3517
rect 1660 3508 1672 3511
rect 1248 3480 1672 3508
rect 1248 3468 1254 3480
rect 1660 3477 1672 3480
rect 1706 3477 1718 3511
rect 1660 3471 1718 3477
rect 854 3344 860 3396
rect 912 3384 918 3396
rect 1527 3387 1585 3393
rect 1527 3384 1539 3387
rect 912 3356 1539 3384
rect 912 3344 918 3356
rect 1527 3353 1539 3356
rect 1573 3353 1585 3387
rect 1527 3347 1585 3353
rect 360 3054 366 3106
rect 418 3054 424 3106
rect 1400 3054 1406 3106
rect 1458 3054 1464 3106
rect 938 3014 944 3026
rect 774 2986 944 3014
rect 150 2326 156 2378
rect 208 2366 214 2378
rect 472 2369 530 2375
rect 472 2366 484 2369
rect 208 2338 484 2366
rect 208 2326 214 2338
rect 472 2335 484 2338
rect 518 2335 530 2369
rect 472 2329 530 2335
rect 604 2369 662 2375
rect 604 2335 616 2369
rect 650 2366 662 2369
rect 774 2366 802 2986
rect 938 2974 944 2986
rect 996 2974 1002 3026
rect 1106 2764 1112 2816
rect 1164 2804 1170 2816
rect 1527 2807 1585 2813
rect 1527 2804 1539 2807
rect 1164 2776 1539 2804
rect 1164 2764 1170 2776
rect 1527 2773 1539 2776
rect 1573 2773 1585 2807
rect 1527 2767 1585 2773
rect 938 2640 944 2692
rect 996 2680 1002 2692
rect 1660 2683 1718 2689
rect 1660 2680 1672 2683
rect 996 2652 1672 2680
rect 996 2640 1002 2652
rect 1660 2649 1672 2652
rect 1706 2649 1718 2683
rect 1660 2643 1718 2649
rect 1022 2516 1028 2568
rect 1080 2556 1086 2568
rect 1793 2559 1851 2565
rect 1793 2556 1805 2559
rect 1080 2528 1805 2556
rect 1080 2516 1086 2528
rect 1793 2525 1805 2528
rect 1839 2525 1851 2559
rect 1793 2519 1851 2525
rect 650 2338 802 2366
rect 650 2335 662 2338
rect 604 2329 662 2335
rect 360 1514 366 1566
rect 418 1514 424 1566
rect 1400 1514 1406 1566
rect 1458 1514 1464 1566
rect 854 1474 860 1486
rect 774 1446 860 1474
rect 66 702 72 754
rect 124 742 130 754
rect 472 745 530 751
rect 472 742 484 745
rect 124 714 484 742
rect 124 702 130 714
rect 472 711 484 714
rect 518 711 530 745
rect 472 705 530 711
rect 604 745 662 751
rect 604 711 616 745
rect 650 742 662 745
rect 774 742 802 1446
rect 854 1434 860 1446
rect 912 1434 918 1486
rect 650 714 802 742
rect 650 711 662 714
rect 604 705 662 711
rect 1022 512 1028 564
rect 1080 552 1086 564
rect 1793 555 1851 561
rect 1793 552 1805 555
rect 1080 524 1805 552
rect 1080 512 1086 524
rect 1793 521 1805 524
rect 1839 521 1851 555
rect 1793 515 1851 521
rect 938 388 944 440
rect 996 428 1002 440
rect 1660 431 1718 437
rect 1660 428 1672 431
rect 996 400 1672 428
rect 996 388 1002 400
rect 1660 397 1672 400
rect 1706 397 1718 431
rect 1660 391 1718 397
rect 854 264 860 316
rect 912 304 918 316
rect 1527 307 1585 313
rect 1527 304 1539 307
rect 912 276 1539 304
rect 912 264 918 276
rect 1527 273 1539 276
rect 1573 273 1585 307
rect 1527 267 1585 273
rect 360 -26 366 26
rect 418 -26 424 26
rect 1400 -26 1406 26
rect 1458 -26 1464 26
<< via1 >>
rect 366 12337 418 12346
rect 366 12303 375 12337
rect 375 12303 409 12337
rect 409 12303 418 12337
rect 366 12294 418 12303
rect 1406 12337 1458 12346
rect 1406 12303 1415 12337
rect 1415 12303 1449 12337
rect 1449 12303 1458 12337
rect 1406 12294 1458 12303
rect 72 12004 124 12056
rect 1112 12004 1164 12056
rect 156 11880 208 11932
rect 1196 11880 1248 11932
rect 240 11756 292 11808
rect 1280 11756 1332 11808
rect 366 10797 418 10806
rect 366 10763 375 10797
rect 375 10763 409 10797
rect 409 10763 418 10797
rect 366 10754 418 10763
rect 1406 10797 1458 10806
rect 1406 10763 1415 10797
rect 1415 10763 1449 10797
rect 1449 10763 1458 10797
rect 1406 10754 1458 10763
rect 1280 9752 1332 9804
rect 1196 9628 1248 9680
rect 860 9504 912 9556
rect 366 9257 418 9266
rect 366 9223 375 9257
rect 375 9223 409 9257
rect 409 9223 418 9257
rect 366 9214 418 9223
rect 1406 9257 1458 9266
rect 1406 9223 1415 9257
rect 1415 9223 1449 9257
rect 1449 9223 1458 9257
rect 1406 9214 1458 9223
rect 1112 8924 1164 8976
rect 944 8800 996 8852
rect 1280 8676 1332 8728
rect 366 7717 418 7726
rect 366 7683 375 7717
rect 375 7683 409 7717
rect 409 7683 418 7717
rect 366 7674 418 7683
rect 1406 7717 1458 7726
rect 1406 7683 1415 7717
rect 1415 7683 1449 7717
rect 1449 7683 1458 7717
rect 1406 7674 1458 7683
rect 1280 6672 1332 6724
rect 944 6548 996 6600
rect 860 6424 912 6476
rect 366 6177 418 6186
rect 366 6143 375 6177
rect 375 6143 409 6177
rect 409 6143 418 6177
rect 366 6134 418 6143
rect 1406 6177 1458 6186
rect 1406 6143 1415 6177
rect 1415 6143 1449 6177
rect 1449 6143 1458 6177
rect 1406 6134 1458 6143
rect 1112 5844 1164 5896
rect 1196 5720 1248 5772
rect 1028 5596 1080 5648
rect 366 4637 418 4646
rect 366 4603 375 4637
rect 375 4603 409 4637
rect 409 4603 418 4637
rect 366 4594 418 4603
rect 1406 4637 1458 4646
rect 1406 4603 1415 4637
rect 1415 4603 1449 4637
rect 1449 4603 1458 4637
rect 1406 4594 1458 4603
rect 240 3782 292 3834
rect 1028 4514 1080 4566
rect 1028 3592 1080 3644
rect 1196 3468 1248 3520
rect 860 3344 912 3396
rect 366 3097 418 3106
rect 366 3063 375 3097
rect 375 3063 409 3097
rect 409 3063 418 3097
rect 366 3054 418 3063
rect 1406 3097 1458 3106
rect 1406 3063 1415 3097
rect 1415 3063 1449 3097
rect 1449 3063 1458 3097
rect 1406 3054 1458 3063
rect 156 2326 208 2378
rect 944 2974 996 3026
rect 1112 2764 1164 2816
rect 944 2640 996 2692
rect 1028 2516 1080 2568
rect 366 1557 418 1566
rect 366 1523 375 1557
rect 375 1523 409 1557
rect 409 1523 418 1557
rect 366 1514 418 1523
rect 1406 1557 1458 1566
rect 1406 1523 1415 1557
rect 1415 1523 1449 1557
rect 1449 1523 1458 1557
rect 1406 1514 1458 1523
rect 72 702 124 754
rect 860 1434 912 1486
rect 1028 512 1080 564
rect 944 388 996 440
rect 860 264 912 316
rect 366 17 418 26
rect 366 -17 375 17
rect 375 -17 409 17
rect 409 -17 418 17
rect 366 -26 418 -17
rect 1406 17 1458 26
rect 1406 -17 1415 17
rect 1415 -17 1449 17
rect 1449 -17 1458 17
rect 1406 -26 1458 -17
<< metal2 >>
rect 364 12348 420 12357
rect 84 12062 112 12320
rect 72 12056 124 12062
rect 72 11998 124 12004
rect 84 760 112 11998
rect 168 11938 196 12320
rect 156 11932 208 11938
rect 156 11874 208 11880
rect 168 2384 196 11874
rect 252 11814 280 12320
rect 1404 12348 1460 12357
rect 364 12283 420 12292
rect 240 11808 292 11814
rect 240 11750 292 11756
rect 252 3840 280 11750
rect 364 10808 420 10817
rect 364 10743 420 10752
rect 872 9562 900 12320
rect 860 9556 912 9562
rect 860 9498 912 9504
rect 364 9268 420 9277
rect 364 9203 420 9212
rect 364 7728 420 7737
rect 364 7663 420 7672
rect 872 6482 900 9498
rect 956 8858 984 12320
rect 944 8852 996 8858
rect 944 8794 996 8800
rect 956 6606 984 8794
rect 944 6600 996 6606
rect 944 6542 996 6548
rect 860 6476 912 6482
rect 860 6418 912 6424
rect 364 6188 420 6197
rect 364 6123 420 6132
rect 364 4648 420 4657
rect 364 4583 420 4592
rect 240 3834 292 3840
rect 240 3776 292 3782
rect 156 2378 208 2384
rect 156 2320 208 2326
rect 72 754 124 760
rect 72 696 124 702
rect 84 84 112 696
rect 168 84 196 2320
rect 252 84 280 3776
rect 872 3402 900 6418
rect 860 3396 912 3402
rect 860 3338 912 3344
rect 364 3108 420 3117
rect 364 3043 420 3052
rect 364 1568 420 1577
rect 364 1503 420 1512
rect 872 1492 900 3338
rect 956 3032 984 6542
rect 1040 5654 1068 12320
rect 1124 12062 1152 12320
rect 1112 12056 1164 12062
rect 1112 11998 1164 12004
rect 1124 8982 1152 11998
rect 1208 11938 1236 12320
rect 1196 11932 1248 11938
rect 1196 11874 1248 11880
rect 1208 9686 1236 11874
rect 1292 11814 1320 12320
rect 1404 12283 1460 12292
rect 1280 11808 1332 11814
rect 1280 11750 1332 11756
rect 1292 9810 1320 11750
rect 1404 10808 1460 10817
rect 1404 10743 1460 10752
rect 1280 9804 1332 9810
rect 1280 9746 1332 9752
rect 1196 9680 1248 9686
rect 1196 9622 1248 9628
rect 1112 8976 1164 8982
rect 1112 8918 1164 8924
rect 1124 5902 1152 8918
rect 1112 5896 1164 5902
rect 1112 5838 1164 5844
rect 1028 5648 1080 5654
rect 1028 5590 1080 5596
rect 1040 4572 1068 5590
rect 1028 4566 1080 4572
rect 1028 4508 1080 4514
rect 1040 3650 1068 4508
rect 1028 3644 1080 3650
rect 1028 3586 1080 3592
rect 944 3026 996 3032
rect 944 2968 996 2974
rect 956 2698 984 2968
rect 944 2692 996 2698
rect 944 2634 996 2640
rect 860 1486 912 1492
rect 860 1428 912 1434
rect 872 322 900 1428
rect 956 446 984 2634
rect 1040 2574 1068 3586
rect 1124 2822 1152 5838
rect 1208 5778 1236 9622
rect 1292 8734 1320 9746
rect 1404 9268 1460 9277
rect 1404 9203 1460 9212
rect 1280 8728 1332 8734
rect 1280 8670 1332 8676
rect 1292 6730 1320 8670
rect 1404 7728 1460 7737
rect 1404 7663 1460 7672
rect 1280 6724 1332 6730
rect 1280 6666 1332 6672
rect 1196 5772 1248 5778
rect 1196 5714 1248 5720
rect 1208 3526 1236 5714
rect 1196 3520 1248 3526
rect 1196 3462 1248 3468
rect 1112 2816 1164 2822
rect 1112 2758 1164 2764
rect 1028 2568 1080 2574
rect 1028 2510 1080 2516
rect 1040 570 1068 2510
rect 1028 564 1080 570
rect 1028 506 1080 512
rect 944 440 996 446
rect 944 382 996 388
rect 860 316 912 322
rect 860 258 912 264
rect 872 84 900 258
rect 956 84 984 382
rect 1040 84 1068 506
rect 1124 84 1152 2758
rect 1208 84 1236 3462
rect 1292 84 1320 6666
rect 1404 6188 1460 6197
rect 1404 6123 1460 6132
rect 1404 4648 1460 4657
rect 1404 4583 1460 4592
rect 1404 3108 1460 3117
rect 1404 3043 1460 3052
rect 1404 1568 1460 1577
rect 1404 1503 1460 1512
rect 364 28 420 37
rect 364 -37 420 -28
rect 1404 28 1460 37
rect 1404 -37 1460 -28
<< via2 >>
rect 364 12346 420 12348
rect 364 12294 366 12346
rect 366 12294 418 12346
rect 418 12294 420 12346
rect 1404 12346 1460 12348
rect 364 12292 420 12294
rect 364 10806 420 10808
rect 364 10754 366 10806
rect 366 10754 418 10806
rect 418 10754 420 10806
rect 364 10752 420 10754
rect 364 9266 420 9268
rect 364 9214 366 9266
rect 366 9214 418 9266
rect 418 9214 420 9266
rect 364 9212 420 9214
rect 364 7726 420 7728
rect 364 7674 366 7726
rect 366 7674 418 7726
rect 418 7674 420 7726
rect 364 7672 420 7674
rect 364 6186 420 6188
rect 364 6134 366 6186
rect 366 6134 418 6186
rect 418 6134 420 6186
rect 364 6132 420 6134
rect 364 4646 420 4648
rect 364 4594 366 4646
rect 366 4594 418 4646
rect 418 4594 420 4646
rect 364 4592 420 4594
rect 364 3106 420 3108
rect 364 3054 366 3106
rect 366 3054 418 3106
rect 418 3054 420 3106
rect 364 3052 420 3054
rect 364 1566 420 1568
rect 364 1514 366 1566
rect 366 1514 418 1566
rect 418 1514 420 1566
rect 364 1512 420 1514
rect 1404 12294 1406 12346
rect 1406 12294 1458 12346
rect 1458 12294 1460 12346
rect 1404 12292 1460 12294
rect 1404 10806 1460 10808
rect 1404 10754 1406 10806
rect 1406 10754 1458 10806
rect 1458 10754 1460 10806
rect 1404 10752 1460 10754
rect 1404 9266 1460 9268
rect 1404 9214 1406 9266
rect 1406 9214 1458 9266
rect 1458 9214 1460 9266
rect 1404 9212 1460 9214
rect 1404 7726 1460 7728
rect 1404 7674 1406 7726
rect 1406 7674 1458 7726
rect 1458 7674 1460 7726
rect 1404 7672 1460 7674
rect 1404 6186 1460 6188
rect 1404 6134 1406 6186
rect 1406 6134 1458 6186
rect 1458 6134 1460 6186
rect 1404 6132 1460 6134
rect 1404 4646 1460 4648
rect 1404 4594 1406 4646
rect 1406 4594 1458 4646
rect 1458 4594 1460 4646
rect 1404 4592 1460 4594
rect 1404 3106 1460 3108
rect 1404 3054 1406 3106
rect 1406 3054 1458 3106
rect 1458 3054 1460 3106
rect 1404 3052 1460 3054
rect 1404 1566 1460 1568
rect 1404 1514 1406 1566
rect 1406 1514 1458 1566
rect 1458 1514 1460 1566
rect 1404 1512 1460 1514
rect 364 26 420 28
rect 364 -26 366 26
rect 366 -26 418 26
rect 418 -26 420 26
rect 364 -28 420 -26
rect 1404 26 1460 28
rect 1404 -26 1406 26
rect 1406 -26 1458 26
rect 1458 -26 1460 26
rect 1404 -28 1460 -26
<< metal3 >>
rect 326 12348 458 12357
rect 326 12292 364 12348
rect 420 12292 458 12348
rect 326 12283 458 12292
rect 1366 12348 1498 12357
rect 1366 12292 1404 12348
rect 1460 12292 1498 12348
rect 1366 12283 1498 12292
rect 326 10808 458 10817
rect 326 10752 364 10808
rect 420 10752 458 10808
rect 326 10743 458 10752
rect 1366 10808 1498 10817
rect 1366 10752 1404 10808
rect 1460 10752 1498 10808
rect 1366 10743 1498 10752
rect 326 9268 458 9277
rect 326 9212 364 9268
rect 420 9212 458 9268
rect 326 9203 458 9212
rect 1366 9268 1498 9277
rect 1366 9212 1404 9268
rect 1460 9212 1498 9268
rect 1366 9203 1498 9212
rect 326 7728 458 7737
rect 326 7672 364 7728
rect 420 7672 458 7728
rect 326 7663 458 7672
rect 1366 7728 1498 7737
rect 1366 7672 1404 7728
rect 1460 7672 1498 7728
rect 1366 7663 1498 7672
rect 326 6188 458 6197
rect 326 6132 364 6188
rect 420 6132 458 6188
rect 326 6123 458 6132
rect 1366 6188 1498 6197
rect 1366 6132 1404 6188
rect 1460 6132 1498 6188
rect 1366 6123 1498 6132
rect 326 4648 458 4657
rect 326 4592 364 4648
rect 420 4592 458 4648
rect 326 4583 458 4592
rect 1366 4648 1498 4657
rect 1366 4592 1404 4648
rect 1460 4592 1498 4648
rect 1366 4583 1498 4592
rect 326 3108 458 3117
rect 326 3052 364 3108
rect 420 3052 458 3108
rect 326 3043 458 3052
rect 1366 3108 1498 3117
rect 1366 3052 1404 3108
rect 1460 3052 1498 3108
rect 1366 3043 1498 3052
rect 326 1568 458 1577
rect 326 1512 364 1568
rect 420 1512 458 1568
rect 326 1503 458 1512
rect 1366 1568 1498 1577
rect 1366 1512 1404 1568
rect 1460 1512 1498 1568
rect 1366 1503 1498 1512
rect 326 28 458 37
rect 326 -28 364 28
rect 420 -28 458 28
rect 326 -37 458 -28
rect 1366 28 1498 37
rect 1366 -28 1404 28
rect 1460 -28 1498 28
rect 1366 -37 1498 -28
use contact_18  contact_18_0
timestamp 1644969367
transform 1 0 1366 0 1 12283
box 0 0 1 1
use contact_17  contact_17_0
timestamp 1644969367
transform 1 0 1400 0 1 12288
box 0 0 1 1
use contact_13  contact_13_0
timestamp 1644969367
transform 1 0 1403 0 1 12297
box 0 0 1 1
use contact_18  contact_18_1
timestamp 1644969367
transform 1 0 326 0 1 12283
box 0 0 1 1
use contact_17  contact_17_1
timestamp 1644969367
transform 1 0 360 0 1 12288
box 0 0 1 1
use contact_13  contact_13_1
timestamp 1644969367
transform 1 0 363 0 1 12297
box 0 0 1 1
use contact_18  contact_18_2
timestamp 1644969367
transform 1 0 1366 0 1 10743
box 0 0 1 1
use contact_17  contact_17_2
timestamp 1644969367
transform 1 0 1400 0 1 10748
box 0 0 1 1
use contact_13  contact_13_2
timestamp 1644969367
transform 1 0 1403 0 1 10757
box 0 0 1 1
use contact_18  contact_18_3
timestamp 1644969367
transform 1 0 326 0 1 10743
box 0 0 1 1
use contact_17  contact_17_3
timestamp 1644969367
transform 1 0 360 0 1 10748
box 0 0 1 1
use contact_13  contact_13_3
timestamp 1644969367
transform 1 0 363 0 1 10757
box 0 0 1 1
use contact_18  contact_18_4
timestamp 1644969367
transform 1 0 1366 0 1 9203
box 0 0 1 1
use contact_17  contact_17_4
timestamp 1644969367
transform 1 0 1400 0 1 9208
box 0 0 1 1
use contact_13  contact_13_4
timestamp 1644969367
transform 1 0 1403 0 1 9217
box 0 0 1 1
use contact_18  contact_18_5
timestamp 1644969367
transform 1 0 326 0 1 9203
box 0 0 1 1
use contact_17  contact_17_5
timestamp 1644969367
transform 1 0 360 0 1 9208
box 0 0 1 1
use contact_13  contact_13_5
timestamp 1644969367
transform 1 0 363 0 1 9217
box 0 0 1 1
use contact_18  contact_18_6
timestamp 1644969367
transform 1 0 1366 0 1 10743
box 0 0 1 1
use contact_17  contact_17_6
timestamp 1644969367
transform 1 0 1400 0 1 10748
box 0 0 1 1
use contact_13  contact_13_6
timestamp 1644969367
transform 1 0 1403 0 1 10757
box 0 0 1 1
use contact_18  contact_18_7
timestamp 1644969367
transform 1 0 326 0 1 10743
box 0 0 1 1
use contact_17  contact_17_7
timestamp 1644969367
transform 1 0 360 0 1 10748
box 0 0 1 1
use contact_13  contact_13_7
timestamp 1644969367
transform 1 0 363 0 1 10757
box 0 0 1 1
use contact_18  contact_18_8
timestamp 1644969367
transform 1 0 1366 0 1 9203
box 0 0 1 1
use contact_17  contact_17_8
timestamp 1644969367
transform 1 0 1400 0 1 9208
box 0 0 1 1
use contact_13  contact_13_8
timestamp 1644969367
transform 1 0 1403 0 1 9217
box 0 0 1 1
use contact_18  contact_18_9
timestamp 1644969367
transform 1 0 326 0 1 9203
box 0 0 1 1
use contact_17  contact_17_9
timestamp 1644969367
transform 1 0 360 0 1 9208
box 0 0 1 1
use contact_13  contact_13_9
timestamp 1644969367
transform 1 0 363 0 1 9217
box 0 0 1 1
use contact_18  contact_18_10
timestamp 1644969367
transform 1 0 1366 0 1 7663
box 0 0 1 1
use contact_17  contact_17_10
timestamp 1644969367
transform 1 0 1400 0 1 7668
box 0 0 1 1
use contact_13  contact_13_10
timestamp 1644969367
transform 1 0 1403 0 1 7677
box 0 0 1 1
use contact_18  contact_18_11
timestamp 1644969367
transform 1 0 326 0 1 7663
box 0 0 1 1
use contact_17  contact_17_11
timestamp 1644969367
transform 1 0 360 0 1 7668
box 0 0 1 1
use contact_13  contact_13_11
timestamp 1644969367
transform 1 0 363 0 1 7677
box 0 0 1 1
use contact_18  contact_18_12
timestamp 1644969367
transform 1 0 1366 0 1 6123
box 0 0 1 1
use contact_17  contact_17_12
timestamp 1644969367
transform 1 0 1400 0 1 6128
box 0 0 1 1
use contact_13  contact_13_12
timestamp 1644969367
transform 1 0 1403 0 1 6137
box 0 0 1 1
use contact_18  contact_18_13
timestamp 1644969367
transform 1 0 326 0 1 6123
box 0 0 1 1
use contact_17  contact_17_13
timestamp 1644969367
transform 1 0 360 0 1 6128
box 0 0 1 1
use contact_13  contact_13_13
timestamp 1644969367
transform 1 0 363 0 1 6137
box 0 0 1 1
use contact_18  contact_18_14
timestamp 1644969367
transform 1 0 1366 0 1 7663
box 0 0 1 1
use contact_17  contact_17_14
timestamp 1644969367
transform 1 0 1400 0 1 7668
box 0 0 1 1
use contact_13  contact_13_14
timestamp 1644969367
transform 1 0 1403 0 1 7677
box 0 0 1 1
use contact_18  contact_18_15
timestamp 1644969367
transform 1 0 326 0 1 7663
box 0 0 1 1
use contact_17  contact_17_15
timestamp 1644969367
transform 1 0 360 0 1 7668
box 0 0 1 1
use contact_13  contact_13_15
timestamp 1644969367
transform 1 0 363 0 1 7677
box 0 0 1 1
use contact_18  contact_18_16
timestamp 1644969367
transform 1 0 1366 0 1 6123
box 0 0 1 1
use contact_17  contact_17_16
timestamp 1644969367
transform 1 0 1400 0 1 6128
box 0 0 1 1
use contact_13  contact_13_16
timestamp 1644969367
transform 1 0 1403 0 1 6137
box 0 0 1 1
use contact_18  contact_18_17
timestamp 1644969367
transform 1 0 326 0 1 6123
box 0 0 1 1
use contact_17  contact_17_17
timestamp 1644969367
transform 1 0 360 0 1 6128
box 0 0 1 1
use contact_13  contact_13_17
timestamp 1644969367
transform 1 0 363 0 1 6137
box 0 0 1 1
use contact_18  contact_18_18
timestamp 1644969367
transform 1 0 1366 0 1 4583
box 0 0 1 1
use contact_17  contact_17_18
timestamp 1644969367
transform 1 0 1400 0 1 4588
box 0 0 1 1
use contact_13  contact_13_18
timestamp 1644969367
transform 1 0 1403 0 1 4597
box 0 0 1 1
use contact_18  contact_18_19
timestamp 1644969367
transform 1 0 326 0 1 4583
box 0 0 1 1
use contact_17  contact_17_19
timestamp 1644969367
transform 1 0 360 0 1 4588
box 0 0 1 1
use contact_13  contact_13_19
timestamp 1644969367
transform 1 0 363 0 1 4597
box 0 0 1 1
use contact_18  contact_18_20
timestamp 1644969367
transform 1 0 1366 0 1 3043
box 0 0 1 1
use contact_17  contact_17_20
timestamp 1644969367
transform 1 0 1400 0 1 3048
box 0 0 1 1
use contact_13  contact_13_20
timestamp 1644969367
transform 1 0 1403 0 1 3057
box 0 0 1 1
use contact_18  contact_18_21
timestamp 1644969367
transform 1 0 326 0 1 3043
box 0 0 1 1
use contact_17  contact_17_21
timestamp 1644969367
transform 1 0 360 0 1 3048
box 0 0 1 1
use contact_13  contact_13_21
timestamp 1644969367
transform 1 0 363 0 1 3057
box 0 0 1 1
use contact_18  contact_18_22
timestamp 1644969367
transform 1 0 1366 0 1 4583
box 0 0 1 1
use contact_17  contact_17_22
timestamp 1644969367
transform 1 0 1400 0 1 4588
box 0 0 1 1
use contact_13  contact_13_22
timestamp 1644969367
transform 1 0 1403 0 1 4597
box 0 0 1 1
use contact_18  contact_18_23
timestamp 1644969367
transform 1 0 326 0 1 4583
box 0 0 1 1
use contact_17  contact_17_23
timestamp 1644969367
transform 1 0 360 0 1 4588
box 0 0 1 1
use contact_13  contact_13_23
timestamp 1644969367
transform 1 0 363 0 1 4597
box 0 0 1 1
use contact_18  contact_18_24
timestamp 1644969367
transform 1 0 1366 0 1 3043
box 0 0 1 1
use contact_17  contact_17_24
timestamp 1644969367
transform 1 0 1400 0 1 3048
box 0 0 1 1
use contact_13  contact_13_24
timestamp 1644969367
transform 1 0 1403 0 1 3057
box 0 0 1 1
use contact_18  contact_18_25
timestamp 1644969367
transform 1 0 326 0 1 3043
box 0 0 1 1
use contact_17  contact_17_25
timestamp 1644969367
transform 1 0 360 0 1 3048
box 0 0 1 1
use contact_13  contact_13_25
timestamp 1644969367
transform 1 0 363 0 1 3057
box 0 0 1 1
use contact_18  contact_18_26
timestamp 1644969367
transform 1 0 1366 0 1 1503
box 0 0 1 1
use contact_17  contact_17_26
timestamp 1644969367
transform 1 0 1400 0 1 1508
box 0 0 1 1
use contact_13  contact_13_26
timestamp 1644969367
transform 1 0 1403 0 1 1517
box 0 0 1 1
use contact_18  contact_18_27
timestamp 1644969367
transform 1 0 326 0 1 1503
box 0 0 1 1
use contact_17  contact_17_27
timestamp 1644969367
transform 1 0 360 0 1 1508
box 0 0 1 1
use contact_13  contact_13_27
timestamp 1644969367
transform 1 0 363 0 1 1517
box 0 0 1 1
use contact_18  contact_18_28
timestamp 1644969367
transform 1 0 1366 0 1 -37
box 0 0 1 1
use contact_17  contact_17_28
timestamp 1644969367
transform 1 0 1400 0 1 -32
box 0 0 1 1
use contact_13  contact_13_28
timestamp 1644969367
transform 1 0 1403 0 1 -23
box 0 0 1 1
use contact_18  contact_18_29
timestamp 1644969367
transform 1 0 326 0 1 -37
box 0 0 1 1
use contact_17  contact_17_29
timestamp 1644969367
transform 1 0 360 0 1 -32
box 0 0 1 1
use contact_13  contact_13_29
timestamp 1644969367
transform 1 0 363 0 1 -23
box 0 0 1 1
use contact_18  contact_18_30
timestamp 1644969367
transform 1 0 1366 0 1 1503
box 0 0 1 1
use contact_17  contact_17_30
timestamp 1644969367
transform 1 0 1400 0 1 1508
box 0 0 1 1
use contact_13  contact_13_30
timestamp 1644969367
transform 1 0 1403 0 1 1517
box 0 0 1 1
use contact_18  contact_18_31
timestamp 1644969367
transform 1 0 326 0 1 1503
box 0 0 1 1
use contact_17  contact_17_31
timestamp 1644969367
transform 1 0 360 0 1 1508
box 0 0 1 1
use contact_13  contact_13_31
timestamp 1644969367
transform 1 0 363 0 1 1517
box 0 0 1 1
use contact_17  contact_17_32
timestamp 1644969367
transform 1 0 1274 0 1 11750
box 0 0 1 1
use contact_17  contact_17_33
timestamp 1644969367
transform 1 0 234 0 1 11750
box 0 0 1 1
use contact_17  contact_17_34
timestamp 1644969367
transform 1 0 1190 0 1 11874
box 0 0 1 1
use contact_17  contact_17_35
timestamp 1644969367
transform 1 0 150 0 1 11874
box 0 0 1 1
use contact_17  contact_17_36
timestamp 1644969367
transform 1 0 1106 0 1 11998
box 0 0 1 1
use contact_17  contact_17_37
timestamp 1644969367
transform 1 0 66 0 1 11998
box 0 0 1 1
use contact_14  contact_14_0
timestamp 1644969367
transform 1 0 1022 0 1 4508
box 0 0 1 1
use contact_13  contact_13_32
timestamp 1644969367
transform 1 0 604 0 1 3785
box 0 0 1 1
use contact_14  contact_14_1
timestamp 1644969367
transform 1 0 938 0 1 2968
box 0 0 1 1
use contact_13  contact_13_33
timestamp 1644969367
transform 1 0 604 0 1 2329
box 0 0 1 1
use contact_14  contact_14_2
timestamp 1644969367
transform 1 0 854 0 1 1428
box 0 0 1 1
use contact_13  contact_13_34
timestamp 1644969367
transform 1 0 604 0 1 705
box 0 0 1 1
use contact_15  contact_15_0
timestamp 1644969367
transform 1 0 1793 0 1 11759
box 0 0 1 1
use contact_14  contact_14_3
timestamp 1644969367
transform 1 0 1274 0 1 11750
box 0 0 1 1
use contact_15  contact_15_1
timestamp 1644969367
transform 1 0 1660 0 1 11883
box 0 0 1 1
use contact_14  contact_14_4
timestamp 1644969367
transform 1 0 1190 0 1 11874
box 0 0 1 1
use contact_13  contact_13_35
timestamp 1644969367
transform 1 0 1527 0 1 12007
box 0 0 1 1
use contact_14  contact_14_5
timestamp 1644969367
transform 1 0 1106 0 1 11998
box 0 0 1 1
use contact_15  contact_15_2
timestamp 1644969367
transform 1 0 1793 0 1 9755
box 0 0 1 1
use contact_14  contact_14_6
timestamp 1644969367
transform 1 0 1274 0 1 9746
box 0 0 1 1
use contact_15  contact_15_3
timestamp 1644969367
transform 1 0 1660 0 1 9631
box 0 0 1 1
use contact_14  contact_14_7
timestamp 1644969367
transform 1 0 1190 0 1 9622
box 0 0 1 1
use contact_13  contact_13_36
timestamp 1644969367
transform 1 0 1527 0 1 9507
box 0 0 1 1
use contact_14  contact_14_8
timestamp 1644969367
transform 1 0 854 0 1 9498
box 0 0 1 1
use contact_15  contact_15_4
timestamp 1644969367
transform 1 0 1793 0 1 8679
box 0 0 1 1
use contact_14  contact_14_9
timestamp 1644969367
transform 1 0 1274 0 1 8670
box 0 0 1 1
use contact_15  contact_15_5
timestamp 1644969367
transform 1 0 1660 0 1 8803
box 0 0 1 1
use contact_14  contact_14_10
timestamp 1644969367
transform 1 0 938 0 1 8794
box 0 0 1 1
use contact_13  contact_13_37
timestamp 1644969367
transform 1 0 1527 0 1 8927
box 0 0 1 1
use contact_14  contact_14_11
timestamp 1644969367
transform 1 0 1106 0 1 8918
box 0 0 1 1
use contact_15  contact_15_6
timestamp 1644969367
transform 1 0 1793 0 1 6675
box 0 0 1 1
use contact_14  contact_14_12
timestamp 1644969367
transform 1 0 1274 0 1 6666
box 0 0 1 1
use contact_15  contact_15_7
timestamp 1644969367
transform 1 0 1660 0 1 6551
box 0 0 1 1
use contact_14  contact_14_13
timestamp 1644969367
transform 1 0 938 0 1 6542
box 0 0 1 1
use contact_13  contact_13_38
timestamp 1644969367
transform 1 0 1527 0 1 6427
box 0 0 1 1
use contact_14  contact_14_14
timestamp 1644969367
transform 1 0 854 0 1 6418
box 0 0 1 1
use contact_15  contact_15_8
timestamp 1644969367
transform 1 0 1793 0 1 5599
box 0 0 1 1
use contact_14  contact_14_15
timestamp 1644969367
transform 1 0 1022 0 1 5590
box 0 0 1 1
use contact_15  contact_15_9
timestamp 1644969367
transform 1 0 1660 0 1 5723
box 0 0 1 1
use contact_14  contact_14_16
timestamp 1644969367
transform 1 0 1190 0 1 5714
box 0 0 1 1
use contact_13  contact_13_39
timestamp 1644969367
transform 1 0 1527 0 1 5847
box 0 0 1 1
use contact_14  contact_14_17
timestamp 1644969367
transform 1 0 1106 0 1 5838
box 0 0 1 1
use contact_15  contact_15_10
timestamp 1644969367
transform 1 0 1793 0 1 3595
box 0 0 1 1
use contact_14  contact_14_18
timestamp 1644969367
transform 1 0 1022 0 1 3586
box 0 0 1 1
use contact_15  contact_15_11
timestamp 1644969367
transform 1 0 1660 0 1 3471
box 0 0 1 1
use contact_14  contact_14_19
timestamp 1644969367
transform 1 0 1190 0 1 3462
box 0 0 1 1
use contact_13  contact_13_40
timestamp 1644969367
transform 1 0 1527 0 1 3347
box 0 0 1 1
use contact_14  contact_14_20
timestamp 1644969367
transform 1 0 854 0 1 3338
box 0 0 1 1
use contact_15  contact_15_12
timestamp 1644969367
transform 1 0 1793 0 1 2519
box 0 0 1 1
use contact_14  contact_14_21
timestamp 1644969367
transform 1 0 1022 0 1 2510
box 0 0 1 1
use contact_15  contact_15_13
timestamp 1644969367
transform 1 0 1660 0 1 2643
box 0 0 1 1
use contact_14  contact_14_22
timestamp 1644969367
transform 1 0 938 0 1 2634
box 0 0 1 1
use contact_13  contact_13_41
timestamp 1644969367
transform 1 0 1527 0 1 2767
box 0 0 1 1
use contact_14  contact_14_23
timestamp 1644969367
transform 1 0 1106 0 1 2758
box 0 0 1 1
use contact_15  contact_15_14
timestamp 1644969367
transform 1 0 1793 0 1 515
box 0 0 1 1
use contact_14  contact_14_24
timestamp 1644969367
transform 1 0 1022 0 1 506
box 0 0 1 1
use contact_15  contact_15_15
timestamp 1644969367
transform 1 0 1660 0 1 391
box 0 0 1 1
use contact_14  contact_14_25
timestamp 1644969367
transform 1 0 938 0 1 382
box 0 0 1 1
use contact_13  contact_13_42
timestamp 1644969367
transform 1 0 1527 0 1 267
box 0 0 1 1
use contact_14  contact_14_26
timestamp 1644969367
transform 1 0 854 0 1 258
box 0 0 1 1
use contact_14  contact_14_27
timestamp 1644969367
transform 1 0 234 0 1 3776
box 0 0 1 1
use contact_13  contact_13_43
timestamp 1644969367
transform 1 0 472 0 1 3785
box 0 0 1 1
use contact_14  contact_14_28
timestamp 1644969367
transform 1 0 150 0 1 2320
box 0 0 1 1
use contact_13  contact_13_44
timestamp 1644969367
transform 1 0 472 0 1 2329
box 0 0 1 1
use contact_14  contact_14_29
timestamp 1644969367
transform 1 0 66 0 1 696
box 0 0 1 1
use contact_13  contact_13_45
timestamp 1644969367
transform 1 0 472 0 1 705
box 0 0 1 1
use and3_dec  and3_dec_0
timestamp 1644969367
transform 1 0 1460 0 -1 12320
box -36 -17 1052 1597
use and3_dec  and3_dec_1
timestamp 1644969367
transform 1 0 1460 0 1 9240
box -36 -17 1052 1597
use and3_dec  and3_dec_2
timestamp 1644969367
transform 1 0 1460 0 -1 9240
box -36 -17 1052 1597
use and3_dec  and3_dec_3
timestamp 1644969367
transform 1 0 1460 0 1 6160
box -36 -17 1052 1597
use and3_dec  and3_dec_4
timestamp 1644969367
transform 1 0 1460 0 -1 6160
box -36 -17 1052 1597
use and3_dec  and3_dec_5
timestamp 1644969367
transform 1 0 1460 0 1 3080
box -36 -17 1052 1597
use and3_dec  and3_dec_6
timestamp 1644969367
transform 1 0 1460 0 -1 3080
box -36 -17 1052 1597
use and3_dec  and3_dec_7
timestamp 1644969367
transform 1 0 1460 0 1 0
box -36 -17 1052 1597
use pinv  pinv_0
timestamp 1644969367
transform 1 0 420 0 1 3080
box -36 -17 404 1597
use pinv  pinv_1
timestamp 1644969367
transform 1 0 420 0 -1 3080
box -36 -17 404 1597
use pinv  pinv_2
timestamp 1644969367
transform 1 0 420 0 1 0
box -36 -17 404 1597
<< labels >>
rlabel metal2 s 72 696 124 760 4 in_0
rlabel metal2 s 156 2320 208 2384 4 in_1
rlabel metal2 s 240 3776 292 3840 4 in_2
rlabel locali s 2304 728 2304 728 4 out_0
rlabel locali s 2304 2352 2304 2352 4 out_1
rlabel locali s 2304 3808 2304 3808 4 out_2
rlabel locali s 2304 5432 2304 5432 4 out_3
rlabel locali s 2304 6888 2304 6888 4 out_4
rlabel locali s 2304 8512 2304 8512 4 out_5
rlabel locali s 2304 9968 2304 9968 4 out_6
rlabel locali s 2304 11592 2304 11592 4 out_7
rlabel metal3 s 1366 7663 1498 7737 4 vdd
rlabel metal3 s 326 10743 458 10817 4 vdd
rlabel metal3 s 392 10780 392 10780 4 vdd
rlabel metal3 s 326 4583 458 4657 4 vdd
rlabel metal3 s 1366 4583 1498 4657 4 vdd
rlabel metal3 s 1366 10743 1498 10817 4 vdd
rlabel metal3 s 1366 1503 1498 1577 4 vdd
rlabel metal3 s 1432 10780 1432 10780 4 vdd
rlabel metal3 s 326 1503 458 1577 4 vdd
rlabel metal3 s 326 7663 458 7737 4 vdd
rlabel metal3 s 326 12283 458 12357 4 gnd
rlabel metal3 s 1366 9203 1498 9277 4 gnd
rlabel metal3 s 326 3043 458 3117 4 gnd
rlabel metal3 s 1366 6123 1498 6197 4 gnd
rlabel metal3 s 1366 -37 1498 37 4 gnd
rlabel metal3 s 326 9203 458 9277 4 gnd
rlabel metal3 s 1366 3043 1498 3117 4 gnd
rlabel metal3 s 326 -37 458 37 4 gnd
rlabel metal3 s 1366 12283 1498 12357 4 gnd
rlabel metal3 s 326 6123 458 6197 4 gnd
<< properties >>
string FIXED_BBOX 1366 -37 1498 0
string GDS_FILE sram_0rw2r1w_32_128_sky130A.gds
string GDS_END 3095176
string GDS_START 3074312
<< end >>
