magic
tech sky130A
magscale 1 2
timestamp 1644949024
<< checkpaint >>
rect -1319 -1316 3089 1598
<< nwell >>
rect -54 226 1824 338
rect -59 58 1829 226
rect -54 -54 1824 58
<< scpmos >>
rect 60 0 90 284
rect 168 0 198 284
rect 276 0 306 284
rect 384 0 414 284
rect 492 0 522 284
rect 600 0 630 284
rect 708 0 738 284
rect 816 0 846 284
rect 924 0 954 284
rect 1032 0 1062 284
rect 1140 0 1170 284
rect 1248 0 1278 284
rect 1356 0 1386 284
rect 1464 0 1494 284
rect 1572 0 1602 284
rect 1680 0 1710 284
<< pdiff >>
rect 0 159 60 284
rect 0 125 8 159
rect 42 125 60 159
rect 0 0 60 125
rect 90 159 168 284
rect 90 125 112 159
rect 146 125 168 159
rect 90 0 168 125
rect 198 159 276 284
rect 198 125 220 159
rect 254 125 276 159
rect 198 0 276 125
rect 306 159 384 284
rect 306 125 328 159
rect 362 125 384 159
rect 306 0 384 125
rect 414 159 492 284
rect 414 125 436 159
rect 470 125 492 159
rect 414 0 492 125
rect 522 159 600 284
rect 522 125 544 159
rect 578 125 600 159
rect 522 0 600 125
rect 630 159 708 284
rect 630 125 652 159
rect 686 125 708 159
rect 630 0 708 125
rect 738 159 816 284
rect 738 125 760 159
rect 794 125 816 159
rect 738 0 816 125
rect 846 159 924 284
rect 846 125 868 159
rect 902 125 924 159
rect 846 0 924 125
rect 954 159 1032 284
rect 954 125 976 159
rect 1010 125 1032 159
rect 954 0 1032 125
rect 1062 159 1140 284
rect 1062 125 1084 159
rect 1118 125 1140 159
rect 1062 0 1140 125
rect 1170 159 1248 284
rect 1170 125 1192 159
rect 1226 125 1248 159
rect 1170 0 1248 125
rect 1278 159 1356 284
rect 1278 125 1300 159
rect 1334 125 1356 159
rect 1278 0 1356 125
rect 1386 159 1464 284
rect 1386 125 1408 159
rect 1442 125 1464 159
rect 1386 0 1464 125
rect 1494 159 1572 284
rect 1494 125 1516 159
rect 1550 125 1572 159
rect 1494 0 1572 125
rect 1602 159 1680 284
rect 1602 125 1624 159
rect 1658 125 1680 159
rect 1602 0 1680 125
rect 1710 159 1770 284
rect 1710 125 1728 159
rect 1762 125 1770 159
rect 1710 0 1770 125
<< pdiffc >>
rect 8 125 42 159
rect 112 125 146 159
rect 220 125 254 159
rect 328 125 362 159
rect 436 125 470 159
rect 544 125 578 159
rect 652 125 686 159
rect 760 125 794 159
rect 868 125 902 159
rect 976 125 1010 159
rect 1084 125 1118 159
rect 1192 125 1226 159
rect 1300 125 1334 159
rect 1408 125 1442 159
rect 1516 125 1550 159
rect 1624 125 1658 159
rect 1728 125 1762 159
<< poly >>
rect 60 284 90 310
rect 168 284 198 310
rect 276 284 306 310
rect 384 284 414 310
rect 492 284 522 310
rect 600 284 630 310
rect 708 284 738 310
rect 816 284 846 310
rect 924 284 954 310
rect 1032 284 1062 310
rect 1140 284 1170 310
rect 1248 284 1278 310
rect 1356 284 1386 310
rect 1464 284 1494 310
rect 1572 284 1602 310
rect 1680 284 1710 310
rect 60 -26 90 0
rect 168 -26 198 0
rect 276 -26 306 0
rect 384 -26 414 0
rect 492 -26 522 0
rect 600 -26 630 0
rect 708 -26 738 0
rect 816 -26 846 0
rect 924 -26 954 0
rect 1032 -26 1062 0
rect 1140 -26 1170 0
rect 1248 -26 1278 0
rect 1356 -26 1386 0
rect 1464 -26 1494 0
rect 1572 -26 1602 0
rect 1680 -26 1710 0
rect 60 -56 1710 -26
<< locali >>
rect 8 159 42 175
rect 8 109 42 125
rect 112 159 146 175
rect 112 75 146 125
rect 220 159 254 175
rect 220 109 254 125
rect 328 159 362 175
rect 328 75 362 125
rect 436 159 470 175
rect 436 109 470 125
rect 544 159 578 175
rect 544 75 578 125
rect 652 159 686 175
rect 652 109 686 125
rect 760 159 794 175
rect 760 75 794 125
rect 868 159 902 175
rect 868 109 902 125
rect 976 159 1010 175
rect 976 75 1010 125
rect 1084 159 1118 175
rect 1084 109 1118 125
rect 1192 159 1226 175
rect 1192 75 1226 125
rect 1300 159 1334 175
rect 1300 109 1334 125
rect 1408 159 1442 175
rect 1408 75 1442 125
rect 1516 159 1550 175
rect 1516 109 1550 125
rect 1624 159 1658 175
rect 1624 75 1658 125
rect 1728 159 1762 175
rect 1728 109 1762 125
rect 112 41 1658 75
use contact_9  contact_9_0
timestamp 1644949024
transform 1 0 1720 0 1 101
box 0 0 2 2
use contact_9  contact_9_1
timestamp 1644949024
transform 1 0 1616 0 1 101
box 0 0 2 2
use contact_9  contact_9_2
timestamp 1644949024
transform 1 0 1508 0 1 101
box 0 0 2 2
use contact_9  contact_9_3
timestamp 1644949024
transform 1 0 1400 0 1 101
box 0 0 2 2
use contact_9  contact_9_4
timestamp 1644949024
transform 1 0 1292 0 1 101
box 0 0 2 2
use contact_9  contact_9_5
timestamp 1644949024
transform 1 0 1184 0 1 101
box 0 0 2 2
use contact_9  contact_9_6
timestamp 1644949024
transform 1 0 1076 0 1 101
box 0 0 2 2
use contact_9  contact_9_7
timestamp 1644949024
transform 1 0 968 0 1 101
box 0 0 2 2
use contact_9  contact_9_8
timestamp 1644949024
transform 1 0 860 0 1 101
box 0 0 2 2
use contact_9  contact_9_9
timestamp 1644949024
transform 1 0 752 0 1 101
box 0 0 2 2
use contact_9  contact_9_10
timestamp 1644949024
transform 1 0 644 0 1 101
box 0 0 2 2
use contact_9  contact_9_11
timestamp 1644949024
transform 1 0 536 0 1 101
box 0 0 2 2
use contact_9  contact_9_12
timestamp 1644949024
transform 1 0 428 0 1 101
box 0 0 2 2
use contact_9  contact_9_13
timestamp 1644949024
transform 1 0 320 0 1 101
box 0 0 2 2
use contact_9  contact_9_14
timestamp 1644949024
transform 1 0 212 0 1 101
box 0 0 2 2
use contact_9  contact_9_15
timestamp 1644949024
transform 1 0 104 0 1 101
box 0 0 2 2
use contact_9  contact_9_16
timestamp 1644949024
transform 1 0 0 0 1 101
box 0 0 2 2
<< labels >>
rlabel mvvaractor s 885 -41 885 -41 4 G
rlabel locali s 1317 142 1317 142 4 S
rlabel locali s 1533 142 1533 142 4 S
rlabel locali s 1101 142 1101 142 4 S
rlabel locali s 237 142 237 142 4 S
rlabel locali s 453 142 453 142 4 S
rlabel locali s 669 142 669 142 4 S
rlabel locali s 885 142 885 142 4 S
rlabel locali s 25 142 25 142 4 S
rlabel locali s 1745 142 1745 142 4 S
rlabel locali s 885 58 885 58 4 D
<< properties >>
string FIXED_BBOX -54 -56 1824 58
string GDS_FILE sram_0rw2r1w_4_16_sky130A.gds
string GDS_END 480558
string GDS_START 476698
<< end >>
