magic
tech sky130A
magscale 1 2
timestamp 1643671299
<< checkpaint >>
rect -1260 -1302 2754 2876
<< nwell >>
rect 0 976 1494 1616
<< pwell >>
rect 240 -42 312 42
rect 554 -42 626 42
rect 868 -42 940 42
rect 1182 -42 1254 42
<< nmos >>
rect 94 230 124 430
rect 190 230 220 430
rect 286 230 316 430
rect 382 230 412 430
rect 478 230 508 430
rect 574 230 604 430
rect 778 230 808 430
rect 874 230 904 430
rect 970 230 1000 430
rect 1074 230 1104 314
rect 1274 230 1304 314
rect 1370 230 1400 314
<< pmos >>
rect 94 1012 124 1096
rect 190 1012 220 1096
rect 286 1012 316 1096
rect 382 1012 412 1096
rect 478 1012 508 1096
rect 574 1012 604 1096
rect 778 1012 808 1096
rect 874 1012 904 1096
rect 970 1012 1000 1096
rect 1074 1012 1104 1282
rect 1274 1012 1304 1282
rect 1370 1012 1400 1282
<< ndiff >>
rect 36 396 94 430
rect 36 362 44 396
rect 78 362 94 396
rect 36 298 94 362
rect 36 264 44 298
rect 78 264 94 298
rect 36 230 94 264
rect 124 230 190 430
rect 220 230 286 430
rect 316 396 382 430
rect 316 362 332 396
rect 366 362 382 396
rect 316 298 382 362
rect 316 264 332 298
rect 366 264 382 298
rect 316 230 382 264
rect 412 230 478 430
rect 508 230 574 430
rect 604 396 662 430
rect 604 362 620 396
rect 654 362 662 396
rect 604 298 662 362
rect 604 264 620 298
rect 654 264 662 298
rect 604 230 662 264
rect 720 396 778 430
rect 720 362 728 396
rect 762 362 778 396
rect 720 298 778 362
rect 720 264 728 298
rect 762 264 778 298
rect 720 230 778 264
rect 808 230 874 430
rect 904 230 970 430
rect 1000 396 1058 430
rect 1000 362 1016 396
rect 1050 362 1058 396
rect 1000 314 1058 362
rect 1000 298 1074 314
rect 1000 264 1016 298
rect 1050 264 1074 298
rect 1000 230 1074 264
rect 1104 288 1162 314
rect 1104 254 1120 288
rect 1154 254 1162 288
rect 1104 230 1162 254
rect 1216 288 1274 314
rect 1216 254 1224 288
rect 1258 254 1274 288
rect 1216 230 1274 254
rect 1304 288 1370 314
rect 1304 254 1320 288
rect 1354 254 1370 288
rect 1304 230 1370 254
rect 1400 288 1458 314
rect 1400 254 1416 288
rect 1450 254 1458 288
rect 1400 230 1458 254
<< pdiff >>
rect 1016 1248 1074 1282
rect 1016 1214 1024 1248
rect 1058 1214 1074 1248
rect 1016 1164 1074 1214
rect 1016 1130 1024 1164
rect 1058 1130 1074 1164
rect 1016 1096 1074 1130
rect 36 1070 94 1096
rect 36 1036 44 1070
rect 78 1036 94 1070
rect 36 1012 94 1036
rect 124 1070 190 1096
rect 124 1036 140 1070
rect 174 1036 190 1070
rect 124 1012 190 1036
rect 220 1070 286 1096
rect 220 1036 236 1070
rect 270 1036 286 1070
rect 220 1012 286 1036
rect 316 1070 382 1096
rect 316 1036 332 1070
rect 366 1036 382 1070
rect 316 1012 382 1036
rect 412 1070 478 1096
rect 412 1036 428 1070
rect 462 1036 478 1070
rect 412 1012 478 1036
rect 508 1070 574 1096
rect 508 1036 524 1070
rect 558 1036 574 1070
rect 508 1012 574 1036
rect 604 1070 662 1096
rect 604 1036 620 1070
rect 654 1036 662 1070
rect 604 1012 662 1036
rect 720 1070 778 1096
rect 720 1036 728 1070
rect 762 1036 778 1070
rect 720 1012 778 1036
rect 808 1070 874 1096
rect 808 1036 824 1070
rect 858 1036 874 1070
rect 808 1012 874 1036
rect 904 1070 970 1096
rect 904 1036 920 1070
rect 954 1036 970 1070
rect 904 1012 970 1036
rect 1000 1080 1074 1096
rect 1000 1046 1024 1080
rect 1058 1046 1074 1080
rect 1000 1012 1074 1046
rect 1104 1248 1162 1282
rect 1104 1214 1120 1248
rect 1154 1214 1162 1248
rect 1104 1164 1162 1214
rect 1104 1130 1120 1164
rect 1154 1130 1162 1164
rect 1104 1080 1162 1130
rect 1104 1046 1120 1080
rect 1154 1046 1162 1080
rect 1104 1012 1162 1046
rect 1216 1248 1274 1282
rect 1216 1214 1224 1248
rect 1258 1214 1274 1248
rect 1216 1164 1274 1214
rect 1216 1130 1224 1164
rect 1258 1130 1274 1164
rect 1216 1080 1274 1130
rect 1216 1046 1224 1080
rect 1258 1046 1274 1080
rect 1216 1012 1274 1046
rect 1304 1248 1370 1282
rect 1304 1214 1320 1248
rect 1354 1214 1370 1248
rect 1304 1164 1370 1214
rect 1304 1130 1320 1164
rect 1354 1130 1370 1164
rect 1304 1080 1370 1130
rect 1304 1046 1320 1080
rect 1354 1046 1370 1080
rect 1304 1012 1370 1046
rect 1400 1248 1458 1282
rect 1400 1214 1416 1248
rect 1450 1214 1458 1248
rect 1400 1164 1458 1214
rect 1400 1130 1416 1164
rect 1450 1130 1458 1164
rect 1400 1080 1458 1130
rect 1400 1046 1416 1080
rect 1450 1046 1458 1080
rect 1400 1012 1458 1046
<< ndiffc >>
rect 44 362 78 396
rect 44 264 78 298
rect 332 362 366 396
rect 332 264 366 298
rect 620 362 654 396
rect 620 264 654 298
rect 728 362 762 396
rect 728 264 762 298
rect 1016 362 1050 396
rect 1016 264 1050 298
rect 1120 254 1154 288
rect 1224 254 1258 288
rect 1320 254 1354 288
rect 1416 254 1450 288
<< pdiffc >>
rect 1024 1214 1058 1248
rect 1024 1130 1058 1164
rect 44 1036 78 1070
rect 140 1036 174 1070
rect 236 1036 270 1070
rect 332 1036 366 1070
rect 428 1036 462 1070
rect 524 1036 558 1070
rect 620 1036 654 1070
rect 728 1036 762 1070
rect 824 1036 858 1070
rect 920 1036 954 1070
rect 1024 1046 1058 1080
rect 1120 1214 1154 1248
rect 1120 1130 1154 1164
rect 1120 1046 1154 1080
rect 1224 1214 1258 1248
rect 1224 1130 1258 1164
rect 1224 1046 1258 1080
rect 1320 1214 1354 1248
rect 1320 1130 1354 1164
rect 1320 1046 1354 1080
rect 1416 1214 1450 1248
rect 1416 1130 1450 1164
rect 1416 1046 1450 1080
<< psubdiff >>
rect 240 17 312 42
rect 240 -17 259 17
rect 293 -17 312 17
rect 240 -42 312 -17
rect 554 17 626 42
rect 554 -17 573 17
rect 607 -17 626 17
rect 554 -42 626 -17
rect 868 17 940 42
rect 868 -17 887 17
rect 921 -17 940 17
rect 868 -42 940 -17
rect 1182 17 1254 42
rect 1182 -17 1201 17
rect 1235 -17 1254 17
rect 1182 -42 1254 -17
<< nsubdiff >>
rect 240 1531 312 1556
rect 240 1497 259 1531
rect 293 1497 312 1531
rect 240 1472 312 1497
rect 554 1531 626 1556
rect 554 1497 573 1531
rect 607 1497 626 1531
rect 554 1472 626 1497
rect 868 1531 940 1556
rect 868 1497 887 1531
rect 921 1497 940 1531
rect 868 1472 940 1497
rect 1182 1531 1254 1556
rect 1182 1497 1201 1531
rect 1235 1497 1254 1531
rect 1182 1472 1254 1497
<< psubdiffcont >>
rect 259 -17 293 17
rect 573 -17 607 17
rect 887 -17 921 17
rect 1201 -17 1235 17
<< nsubdiffcont >>
rect 259 1497 293 1531
rect 573 1497 607 1531
rect 887 1497 921 1531
rect 1201 1497 1235 1531
<< poly >>
rect 1074 1282 1104 1308
rect 1274 1282 1304 1308
rect 1370 1282 1400 1308
rect 94 1096 124 1122
rect 190 1096 220 1122
rect 286 1096 316 1122
rect 382 1096 412 1122
rect 478 1096 508 1122
rect 574 1096 604 1122
rect 778 1096 808 1122
rect 874 1096 904 1122
rect 970 1096 1000 1122
rect 94 978 124 1012
rect 70 962 124 978
rect 70 928 80 962
rect 114 928 124 962
rect 70 912 124 928
rect 190 922 220 1012
rect 94 430 124 912
rect 166 906 220 922
rect 166 872 176 906
rect 210 872 220 906
rect 166 856 220 872
rect 286 866 316 1012
rect 190 430 220 856
rect 262 850 316 866
rect 262 816 272 850
rect 306 816 316 850
rect 262 800 316 816
rect 382 810 412 1012
rect 286 430 316 800
rect 358 794 412 810
rect 358 760 368 794
rect 402 760 412 794
rect 358 744 412 760
rect 478 754 508 1012
rect 382 430 412 744
rect 454 738 508 754
rect 454 704 464 738
rect 498 704 508 738
rect 454 688 508 704
rect 574 698 604 1012
rect 478 430 508 688
rect 550 682 604 698
rect 550 648 560 682
rect 594 648 604 682
rect 550 632 604 648
rect 778 642 808 1012
rect 574 430 604 632
rect 754 626 808 642
rect 754 592 764 626
rect 798 592 808 626
rect 754 576 808 592
rect 874 586 904 1012
rect 778 430 808 576
rect 850 570 904 586
rect 850 536 860 570
rect 894 536 904 570
rect 850 520 904 536
rect 970 530 1000 1012
rect 1074 638 1104 1012
rect 1050 622 1104 638
rect 1050 588 1060 622
rect 1094 588 1104 622
rect 1050 572 1104 588
rect 874 430 904 520
rect 946 514 1000 530
rect 946 480 956 514
rect 990 480 1000 514
rect 946 464 1000 480
rect 970 430 1000 464
rect 1074 314 1104 572
rect 1274 840 1304 1012
rect 1370 978 1400 1012
rect 1346 962 1400 978
rect 1346 928 1356 962
rect 1390 928 1400 962
rect 1346 912 1400 928
rect 1274 824 1328 840
rect 1274 790 1284 824
rect 1318 790 1328 824
rect 1274 774 1328 790
rect 1274 314 1304 774
rect 1370 314 1400 912
rect 94 204 124 230
rect 190 204 220 230
rect 286 204 316 230
rect 382 204 412 230
rect 478 204 508 230
rect 574 204 604 230
rect 778 204 808 230
rect 874 204 904 230
rect 970 204 1000 230
rect 1074 204 1104 230
rect 1274 204 1304 230
rect 1370 204 1400 230
<< polycont >>
rect 80 928 114 962
rect 176 872 210 906
rect 272 816 306 850
rect 368 760 402 794
rect 464 704 498 738
rect 560 648 594 682
rect 764 592 798 626
rect 860 536 894 570
rect 1060 588 1094 622
rect 956 480 990 514
rect 1356 928 1390 962
rect 1284 790 1318 824
<< locali >>
rect 258 1532 294 1548
rect 572 1532 608 1548
rect 886 1532 922 1548
rect 1200 1532 1236 1548
rect 140 1531 1354 1532
rect 140 1497 259 1531
rect 293 1497 573 1531
rect 607 1497 887 1531
rect 921 1497 1201 1531
rect 1235 1497 1354 1531
rect 140 1496 1354 1497
rect 140 1096 174 1496
rect 258 1480 294 1496
rect 332 1096 366 1496
rect 524 1480 608 1496
rect 824 1480 922 1496
rect 524 1096 558 1480
rect 824 1096 858 1480
rect 1024 1282 1058 1496
rect 1200 1480 1236 1496
rect 1320 1282 1354 1496
rect 1016 1248 1064 1282
rect 1016 1214 1024 1248
rect 1058 1214 1064 1248
rect 1016 1164 1064 1214
rect 1016 1130 1024 1164
rect 1058 1130 1064 1164
rect 36 1070 84 1096
rect 36 1036 44 1070
rect 78 1036 84 1070
rect 36 1012 84 1036
rect 134 1070 180 1096
rect 134 1036 140 1070
rect 174 1036 180 1070
rect 134 1012 180 1036
rect 230 1070 276 1096
rect 230 1036 236 1070
rect 270 1036 276 1070
rect 230 1012 276 1036
rect 326 1070 372 1096
rect 326 1036 332 1070
rect 366 1036 372 1070
rect 326 1012 372 1036
rect 422 1070 468 1096
rect 422 1036 428 1070
rect 462 1036 468 1070
rect 422 1012 468 1036
rect 518 1070 564 1096
rect 518 1036 524 1070
rect 558 1036 564 1070
rect 518 1012 564 1036
rect 614 1070 662 1096
rect 614 1036 620 1070
rect 654 1036 662 1070
rect 614 1012 662 1036
rect 720 1070 768 1096
rect 720 1036 728 1070
rect 762 1036 768 1070
rect 720 1012 768 1036
rect 818 1070 864 1096
rect 818 1036 824 1070
rect 858 1036 864 1070
rect 818 1012 864 1036
rect 914 1070 960 1096
rect 914 1036 920 1070
rect 954 1036 960 1070
rect 914 1012 960 1036
rect 1016 1080 1064 1130
rect 1016 1046 1024 1080
rect 1058 1046 1064 1080
rect 1016 1012 1064 1046
rect 1114 1248 1162 1282
rect 1114 1214 1120 1248
rect 1154 1214 1162 1248
rect 1114 1164 1162 1214
rect 1114 1130 1120 1164
rect 1154 1130 1162 1164
rect 1114 1080 1162 1130
rect 1114 1046 1120 1080
rect 1154 1046 1162 1080
rect 1114 1012 1162 1046
rect 80 962 114 978
rect 80 912 114 928
rect 696 934 728 968
rect 176 906 210 922
rect 176 856 210 872
rect 272 850 306 866
rect 272 800 306 816
rect 368 794 402 810
rect 614 776 662 810
rect 368 744 402 760
rect 464 738 498 754
rect 464 688 498 704
rect 560 682 594 698
rect 560 632 594 648
rect 628 598 662 776
rect 44 564 662 598
rect 44 430 78 564
rect 696 530 730 934
rect 926 654 960 1012
rect 764 626 798 642
rect 926 622 1094 654
rect 926 620 1060 622
rect 764 576 798 592
rect 620 496 730 530
rect 860 570 894 586
rect 1060 572 1094 588
rect 1128 608 1162 1012
rect 1216 1248 1264 1282
rect 1216 1214 1224 1248
rect 1258 1214 1264 1248
rect 1216 1164 1264 1214
rect 1216 1130 1224 1164
rect 1258 1130 1264 1164
rect 1216 1080 1264 1130
rect 1216 1046 1224 1080
rect 1258 1046 1264 1080
rect 1216 1012 1264 1046
rect 1314 1248 1360 1282
rect 1314 1214 1320 1248
rect 1354 1214 1360 1248
rect 1314 1164 1360 1214
rect 1314 1130 1320 1164
rect 1354 1130 1360 1164
rect 1314 1080 1360 1130
rect 1314 1046 1320 1080
rect 1354 1046 1360 1080
rect 1314 1012 1360 1046
rect 1410 1248 1458 1282
rect 1410 1214 1416 1248
rect 1450 1214 1458 1248
rect 1410 1164 1458 1214
rect 1410 1130 1416 1164
rect 1450 1130 1458 1164
rect 1410 1080 1458 1130
rect 1410 1046 1416 1080
rect 1450 1046 1458 1080
rect 1410 1012 1458 1046
rect 1216 730 1250 1012
rect 1356 962 1390 978
rect 1356 912 1390 928
rect 1424 876 1458 1012
rect 1284 824 1318 840
rect 1284 774 1318 790
rect 1128 574 1134 608
rect 860 520 894 536
rect 956 514 990 530
rect 620 430 654 496
rect 956 464 990 480
rect 36 396 84 430
rect 36 362 44 396
rect 78 362 84 396
rect 36 298 84 362
rect 36 264 44 298
rect 78 264 84 298
rect 36 230 84 264
rect 326 396 372 430
rect 326 362 332 396
rect 366 362 372 396
rect 326 298 372 362
rect 326 264 332 298
rect 366 264 372 298
rect 326 230 372 264
rect 614 396 662 430
rect 614 362 620 396
rect 654 362 662 396
rect 614 298 662 362
rect 614 264 620 298
rect 654 264 662 298
rect 614 230 662 264
rect 720 396 768 430
rect 720 362 728 396
rect 762 362 768 396
rect 720 298 768 362
rect 720 264 728 298
rect 762 264 768 298
rect 720 230 768 264
rect 1010 396 1058 430
rect 1010 362 1016 396
rect 1050 362 1058 396
rect 1010 298 1058 362
rect 1128 314 1162 574
rect 1010 264 1016 298
rect 1050 264 1058 298
rect 1010 230 1058 264
rect 1114 288 1162 314
rect 1114 254 1120 288
rect 1154 254 1162 288
rect 1114 230 1162 254
rect 1216 314 1250 696
rect 1424 314 1458 842
rect 1216 288 1264 314
rect 1216 254 1224 288
rect 1258 254 1264 288
rect 1216 230 1264 254
rect 1314 288 1360 314
rect 1314 254 1320 288
rect 1354 254 1360 288
rect 1314 230 1360 254
rect 1410 288 1458 314
rect 1410 254 1416 288
rect 1450 254 1458 288
rect 1410 230 1458 254
rect 258 18 294 42
rect 332 18 366 230
rect 572 18 608 42
rect 886 18 922 42
rect 1016 18 1050 230
rect 1200 18 1236 42
rect 1320 18 1354 230
rect 140 17 1354 18
rect 140 -17 259 17
rect 293 -17 573 17
rect 607 -17 887 17
rect 921 -17 1201 17
rect 1235 -17 1354 17
rect 140 -18 1354 -17
rect 258 -42 294 -18
rect 572 -42 608 -18
rect 886 -42 922 -18
rect 1200 -42 1236 -18
<< viali >>
rect 259 1497 293 1531
rect 573 1497 607 1531
rect 887 1497 921 1531
rect 1201 1497 1235 1531
rect 44 1036 78 1070
rect 236 1036 270 1070
rect 428 1036 462 1070
rect 620 1036 654 1070
rect 728 1036 762 1070
rect 920 1036 954 1070
rect 80 928 114 962
rect 728 934 762 968
rect 176 872 210 906
rect 272 816 306 850
rect 368 760 402 794
rect 580 776 614 810
rect 464 704 498 738
rect 560 648 594 682
rect 764 592 798 626
rect 1060 588 1094 622
rect 1356 928 1390 962
rect 1424 842 1458 876
rect 1284 790 1318 824
rect 1216 696 1250 730
rect 1134 574 1168 608
rect 860 536 894 570
rect 956 480 990 514
rect 728 264 762 298
rect 259 -17 293 17
rect 573 -17 607 17
rect 887 -17 921 17
rect 1201 -17 1235 17
<< metal1 >>
rect 0 1531 1494 1544
rect 0 1497 259 1531
rect 293 1497 573 1531
rect 607 1497 887 1531
rect 921 1497 1201 1531
rect 1235 1497 1494 1531
rect 0 1484 1494 1497
rect 38 1070 276 1082
rect 38 1036 44 1070
rect 78 1054 236 1070
rect 78 1036 84 1054
rect 38 1024 84 1036
rect 230 1036 236 1054
rect 270 1036 276 1070
rect 230 1024 276 1036
rect 422 1070 660 1082
rect 422 1036 428 1070
rect 462 1054 620 1070
rect 462 1036 468 1054
rect 422 1024 468 1036
rect 614 1036 620 1054
rect 654 1036 660 1070
rect 614 1024 660 1036
rect 722 1070 960 1082
rect 722 1036 728 1070
rect 762 1054 920 1070
rect 762 1036 768 1054
rect 722 1024 768 1036
rect 914 1036 920 1054
rect 954 1036 960 1070
rect 914 1024 960 1036
rect 248 988 276 1024
rect 72 962 126 976
rect 72 942 80 962
rect 70 928 80 942
rect 114 928 126 962
rect 248 960 506 988
rect 70 914 126 928
rect 168 906 222 920
rect 168 886 176 906
rect 166 872 176 886
rect 210 872 222 906
rect 166 858 222 872
rect 264 850 318 864
rect 264 830 272 850
rect 262 816 272 830
rect 306 816 318 850
rect 262 802 318 816
rect 478 836 506 960
rect 632 980 660 1024
rect 632 974 768 980
rect 632 968 1396 974
rect 632 952 728 968
rect 722 934 728 952
rect 762 962 1396 968
rect 762 946 1356 962
rect 762 934 768 946
rect 722 922 768 934
rect 1350 928 1356 946
rect 1390 928 1396 962
rect 1350 916 1396 928
rect 1418 876 1464 888
rect 1418 842 1424 876
rect 1458 848 1494 876
rect 1458 842 1464 848
rect 478 824 1324 836
rect 1418 830 1464 842
rect 478 810 1284 824
rect 478 808 580 810
rect 360 794 414 808
rect 360 774 368 794
rect 358 760 368 774
rect 402 760 414 794
rect 574 776 580 808
rect 614 808 1284 810
rect 614 776 620 808
rect 1278 790 1284 808
rect 1318 790 1324 824
rect 1278 778 1324 790
rect 574 764 620 776
rect 358 746 414 760
rect 456 738 510 752
rect 456 718 464 738
rect 454 704 464 718
rect 498 704 510 738
rect 454 690 510 704
rect 1210 730 1256 742
rect 1210 696 1216 730
rect 1250 702 1494 730
rect 1250 696 1256 702
rect 552 682 606 696
rect 1210 684 1256 696
rect 552 662 560 682
rect 550 648 560 662
rect 594 648 606 682
rect 550 634 606 648
rect 756 626 810 640
rect 756 606 764 626
rect 754 592 764 606
rect 798 592 810 626
rect 754 578 810 592
rect 1054 622 1100 634
rect 1054 588 1060 622
rect 1094 588 1100 622
rect 852 570 906 584
rect 1054 576 1100 588
rect 852 550 860 570
rect 850 536 860 550
rect 894 536 906 570
rect 850 522 906 536
rect 948 514 1002 528
rect 948 494 956 514
rect 946 480 956 494
rect 990 480 1002 514
rect 946 466 1002 480
rect 1072 310 1100 576
rect 1128 608 1174 620
rect 1128 574 1134 608
rect 1168 580 1494 608
rect 1168 574 1174 580
rect 1128 562 1174 574
rect 722 298 1100 310
rect 722 264 728 298
rect 762 282 1100 298
rect 762 264 768 282
rect 722 252 768 264
rect 0 17 1494 30
rect 0 -17 259 17
rect 293 -17 573 17
rect 607 -17 887 17
rect 921 -17 1201 17
rect 1235 -17 1494 17
rect 0 -30 1494 -17
<< labels >>
rlabel metal1 s 358 964 358 964 4 net3
rlabel mvpsubdiff s 434 316 434 316 4 net4
rlabel mvpsubdiff s 532 314 532 314 4 net5
rlabel metal1 s 652 960 652 960 4 net6
rlabel mvpsubdiff s 252 314 252 314 4 net1
rlabel mvpsubdiff s 158 306 158 306 4 net2
rlabel mvpsubdiff s 932 340 932 340 4 net7
rlabel mvpsubdiff s 840 336 840 336 4 net8
rlabel locali s 950 750 950 750 4 net9
rlabel metal1 s 70 914 126 942 4 A0
port 1 nsew
rlabel metal1 s 166 858 222 886 4 B0
port 2 nsew
rlabel metal1 s 262 802 318 830 4 C0
port 3 nsew
rlabel metal1 s 358 746 414 774 4 A1
port 4 nsew
rlabel metal1 s 454 690 510 718 4 B1
port 5 nsew
rlabel metal1 s 550 634 606 662 4 C1
port 6 nsew
rlabel metal1 s 754 578 810 606 4 A2
port 7 nsew
rlabel metal1 s 850 522 906 550 4 B2
port 8 nsew
rlabel metal1 s 946 466 1002 494 4 C2
port 9 nsew
rlabel metal1 s 1418 848 1494 876 4 OUT1
port 10 nsew
rlabel metal1 s 1210 702 1494 730 4 OUT0
port 11 nsew
rlabel metal1 s 1128 580 1494 608 4 OUT2
port 12 nsew
rlabel metal1 s 0 1484 1494 1544 4 vdd
port 13 nsew
rlabel metal1 s 0 -30 1494 30 4 gnd
port 14 nsew
rlabel metal1 s 98 928 98 928 4 A0
rlabel metal1 s 194 872 194 872 4 B0
rlabel metal1 s 290 816 290 816 4 C0
rlabel metal1 s 386 760 386 760 4 A1
rlabel metal1 s 482 704 482 704 4 B1
rlabel metal1 s 578 648 578 648 4 C1
rlabel metal1 s 782 592 782 592 4 A2
rlabel metal1 s 878 536 878 536 4 B2
rlabel metal1 s 974 480 974 480 4 C2
rlabel metal1 s 1352 716 1352 716 4 OUT0
rlabel metal1 s 1456 862 1456 862 4 OUT1
rlabel metal1 s 1311 594 1311 594 4 OUT2
rlabel metal1 s 747 1514 747 1514 4 vdd
rlabel metal1 s 747 0 747 0 4 gnd
<< properties >>
string FIXED_BBOX 0 0 1494 1514
string GDS_FILE sram_0rw2r1w_16_32_sky130A.gds
string GDS_END 1048788
string GDS_START 1024274
<< end >>
