magic
tech sky130A
magscale 1 2
timestamp 1644969367
<< checkpaint >>
rect -1296 -1277 13008 2155
<< nwell >>
rect -36 402 11748 895
<< locali >>
rect 0 821 11712 855
rect 48 344 114 410
rect 196 360 449 394
rect 564 360 817 394
rect 1025 354 1401 388
rect 1842 354 2417 388
rect 3597 352 4945 386
rect 8285 352 8319 386
rect 0 -17 11712 17
use pinv_10  pinv_10_0
timestamp 1644969367
transform 1 0 4864 0 1 0
box -36 -17 6884 895
use pinv_9  pinv_9_0
timestamp 1644969367
transform 1 0 2336 0 1 0
box -36 -17 2564 895
use pinv_8  pinv_8_0
timestamp 1644969367
transform 1 0 1320 0 1 0
box -36 -17 1052 895
use pinv_7  pinv_7_0
timestamp 1644969367
transform 1 0 736 0 1 0
box -36 -17 620 895
use pinv_6  pinv_6_0
timestamp 1644969367
transform 1 0 368 0 1 0
box -36 -17 404 895
use pinv_6  pinv_6_1
timestamp 1644969367
transform 1 0 0 0 1 0
box -36 -17 404 895
<< labels >>
rlabel locali s 8302 369 8302 369 4 Z
rlabel locali s 81 377 81 377 4 A
rlabel locali s 5856 0 5856 0 4 gnd
rlabel locali s 5856 838 5856 838 4 vdd
<< properties >>
string FIXED_BBOX 0 0 11712 838
string GDS_FILE sram_0rw2r1w_32_128_sky130A.gds
string GDS_END 3305240
string GDS_START 3303638
<< end >>
