magic
tech sky130A
magscale 1 2
timestamp 1644969367
<< checkpaint >>
rect -1260 -1302 7792 99734
<< viali >>
rect 3022 36207 3056 36241
rect 3022 34583 3056 34617
rect 3022 33127 3056 33161
rect 3022 31503 3056 31537
rect 3022 30047 3056 30081
rect 3022 28423 3056 28457
rect 3022 26967 3056 27001
rect 3022 25343 3056 25377
rect 3022 20811 3056 20845
rect 3022 19187 3056 19221
rect 3022 17731 3056 17765
rect 3022 16107 3056 16141
rect 3022 14651 3056 14685
rect 3022 13027 3056 13061
rect 3022 11571 3056 11605
rect 3022 9947 3056 9981
rect 3022 5415 3056 5449
rect 3022 3791 3056 3825
rect 3022 2335 3056 2369
rect 3022 711 3056 745
<< metal1 >>
rect 6434 98406 6440 98458
rect 6492 98406 6498 98458
rect 4688 98024 4694 98076
rect 4746 98064 4752 98076
rect 4746 98036 5946 98064
rect 4746 98024 4752 98036
rect 4184 97938 4190 97990
rect 4242 97978 4248 97990
rect 4242 97950 5850 97978
rect 4242 97938 4248 97950
rect 3428 97852 3434 97904
rect 3486 97892 3492 97904
rect 3486 97864 5754 97892
rect 3486 97852 3492 97864
rect 6086 97824 6452 97852
rect 4688 97766 4694 97818
rect 4746 97806 4752 97818
rect 4746 97778 5550 97806
rect 4746 97766 4752 97778
rect 4184 97680 4190 97732
rect 4242 97720 4248 97732
rect 4242 97692 5454 97720
rect 6168 97702 6452 97730
rect 4242 97680 4248 97692
rect 3344 97594 3350 97646
rect 3402 97634 3408 97646
rect 3402 97606 5358 97634
rect 3402 97594 3408 97606
rect 4688 97508 4694 97560
rect 4746 97548 4752 97560
rect 6376 97556 6452 97584
rect 4746 97520 5262 97548
rect 4746 97508 4752 97520
rect 4184 97422 4190 97474
rect 4242 97462 4248 97474
rect 4242 97434 5166 97462
rect 4242 97422 4248 97434
rect 3260 97336 3266 97388
rect 3318 97376 3324 97388
rect 3318 97348 5070 97376
rect 3318 97336 3324 97348
rect 6434 96868 6440 96920
rect 6492 96868 6498 96920
rect 3344 96400 3350 96452
rect 3402 96440 3408 96452
rect 3402 96412 5070 96440
rect 3402 96400 3408 96412
rect 4100 96314 4106 96366
rect 4158 96354 4164 96366
rect 4158 96326 5166 96354
rect 4158 96314 4164 96326
rect 4688 96228 4694 96280
rect 4746 96268 4752 96280
rect 4746 96240 5262 96268
rect 4746 96228 4752 96240
rect 6376 96204 6452 96232
rect 3428 96142 3434 96194
rect 3486 96182 3492 96194
rect 3486 96154 5358 96182
rect 3486 96142 3492 96154
rect 4100 96056 4106 96108
rect 4158 96096 4164 96108
rect 4158 96068 5454 96096
rect 4158 96056 4164 96068
rect 6168 96058 6452 96086
rect 4688 95970 4694 96022
rect 4746 96010 4752 96022
rect 4746 95982 5550 96010
rect 4746 95970 4752 95982
rect 6086 95936 6452 95964
rect 3512 95884 3518 95936
rect 3570 95924 3576 95936
rect 3570 95896 5754 95924
rect 3570 95884 3576 95896
rect 4100 95798 4106 95850
rect 4158 95838 4164 95850
rect 4158 95810 5850 95838
rect 4158 95798 4164 95810
rect 4688 95712 4694 95764
rect 4746 95752 4752 95764
rect 4746 95724 5946 95752
rect 4746 95712 4752 95724
rect 6434 95330 6440 95382
rect 6492 95330 6498 95382
rect 4688 94948 4694 95000
rect 4746 94988 4752 95000
rect 4746 94960 5946 94988
rect 4746 94948 4752 94960
rect 4100 94862 4106 94914
rect 4158 94902 4164 94914
rect 4158 94874 5850 94902
rect 4158 94862 4164 94874
rect 3260 94776 3266 94828
rect 3318 94816 3324 94828
rect 3318 94788 5754 94816
rect 3318 94776 3324 94788
rect 6086 94748 6452 94776
rect 4688 94690 4694 94742
rect 4746 94730 4752 94742
rect 4746 94702 5550 94730
rect 4746 94690 4752 94702
rect 4016 94604 4022 94656
rect 4074 94644 4080 94656
rect 4074 94616 5454 94644
rect 6168 94626 6452 94654
rect 4074 94604 4080 94616
rect 3512 94518 3518 94570
rect 3570 94558 3576 94570
rect 3570 94530 5358 94558
rect 3570 94518 3576 94530
rect 4688 94432 4694 94484
rect 4746 94472 4752 94484
rect 6376 94480 6452 94508
rect 4746 94444 5262 94472
rect 4746 94432 4752 94444
rect 4016 94346 4022 94398
rect 4074 94386 4080 94398
rect 4074 94358 5166 94386
rect 4074 94346 4080 94358
rect 3428 94260 3434 94312
rect 3486 94300 3492 94312
rect 3486 94272 5070 94300
rect 3486 94260 3492 94272
rect 6434 93792 6440 93844
rect 6492 93792 6498 93844
rect 3512 93324 3518 93376
rect 3570 93364 3576 93376
rect 3570 93336 5070 93364
rect 3570 93324 3576 93336
rect 3932 93238 3938 93290
rect 3990 93278 3996 93290
rect 3990 93250 5166 93278
rect 3990 93238 3996 93250
rect 4688 93152 4694 93204
rect 4746 93192 4752 93204
rect 4746 93164 5262 93192
rect 4746 93152 4752 93164
rect 6376 93128 6452 93156
rect 3260 93066 3266 93118
rect 3318 93106 3324 93118
rect 3318 93078 5358 93106
rect 3318 93066 3324 93078
rect 4016 92980 4022 93032
rect 4074 93020 4080 93032
rect 4074 92992 5454 93020
rect 4074 92980 4080 92992
rect 6168 92982 6452 93010
rect 4688 92894 4694 92946
rect 4746 92934 4752 92946
rect 4746 92906 5550 92934
rect 4746 92894 4752 92906
rect 6086 92860 6452 92888
rect 3344 92808 3350 92860
rect 3402 92848 3408 92860
rect 3402 92820 5754 92848
rect 3402 92808 3408 92820
rect 4016 92722 4022 92774
rect 4074 92762 4080 92774
rect 4074 92734 5850 92762
rect 4074 92722 4080 92734
rect 4688 92636 4694 92688
rect 4746 92676 4752 92688
rect 4746 92648 5946 92676
rect 4746 92636 4752 92648
rect 6434 92254 6440 92306
rect 6492 92254 6498 92306
rect 4688 91872 4694 91924
rect 4746 91912 4752 91924
rect 4746 91884 5946 91912
rect 4746 91872 4752 91884
rect 3932 91786 3938 91838
rect 3990 91826 3996 91838
rect 3990 91798 5850 91826
rect 3990 91786 3996 91798
rect 3428 91700 3434 91752
rect 3486 91740 3492 91752
rect 3486 91712 5754 91740
rect 3486 91700 3492 91712
rect 6086 91672 6452 91700
rect 4688 91614 4694 91666
rect 4746 91654 4752 91666
rect 4746 91626 5550 91654
rect 4746 91614 4752 91626
rect 3932 91528 3938 91580
rect 3990 91568 3996 91580
rect 3990 91540 5454 91568
rect 6168 91550 6452 91578
rect 3990 91528 3996 91540
rect 3344 91442 3350 91494
rect 3402 91482 3408 91494
rect 3402 91454 5358 91482
rect 3402 91442 3408 91454
rect 4688 91356 4694 91408
rect 4746 91396 4752 91408
rect 6376 91404 6452 91432
rect 4746 91368 5262 91396
rect 4746 91356 4752 91368
rect 3932 91270 3938 91322
rect 3990 91310 3996 91322
rect 3990 91282 5166 91310
rect 3990 91270 3996 91282
rect 3260 91184 3266 91236
rect 3318 91224 3324 91236
rect 3318 91196 5070 91224
rect 3318 91184 3324 91196
rect 6434 90716 6440 90768
rect 6492 90716 6498 90768
rect 3344 90248 3350 90300
rect 3402 90288 3408 90300
rect 3402 90260 5070 90288
rect 3402 90248 3408 90260
rect 3848 90162 3854 90214
rect 3906 90202 3912 90214
rect 3906 90174 5166 90202
rect 3906 90162 3912 90174
rect 4688 90076 4694 90128
rect 4746 90116 4752 90128
rect 4746 90088 5262 90116
rect 4746 90076 4752 90088
rect 6376 90052 6452 90080
rect 3428 89990 3434 90042
rect 3486 90030 3492 90042
rect 3486 90002 5358 90030
rect 3486 89990 3492 90002
rect 3848 89904 3854 89956
rect 3906 89944 3912 89956
rect 3906 89916 5454 89944
rect 3906 89904 3912 89916
rect 6168 89906 6452 89934
rect 4688 89818 4694 89870
rect 4746 89858 4752 89870
rect 4746 89830 5550 89858
rect 4746 89818 4752 89830
rect 6086 89784 6452 89812
rect 3512 89732 3518 89784
rect 3570 89772 3576 89784
rect 3570 89744 5754 89772
rect 3570 89732 3576 89744
rect 3848 89646 3854 89698
rect 3906 89686 3912 89698
rect 3906 89658 5850 89686
rect 3906 89646 3912 89658
rect 4688 89560 4694 89612
rect 4746 89600 4752 89612
rect 4746 89572 5946 89600
rect 4746 89560 4752 89572
rect 6434 89178 6440 89230
rect 6492 89178 6498 89230
rect 4688 88796 4694 88848
rect 4746 88836 4752 88848
rect 4746 88808 5946 88836
rect 4746 88796 4752 88808
rect 3848 88710 3854 88762
rect 3906 88750 3912 88762
rect 3906 88722 5850 88750
rect 3906 88710 3912 88722
rect 3260 88624 3266 88676
rect 3318 88664 3324 88676
rect 3318 88636 5754 88664
rect 3318 88624 3324 88636
rect 6086 88596 6452 88624
rect 4688 88538 4694 88590
rect 4746 88578 4752 88590
rect 4746 88550 5550 88578
rect 4746 88538 4752 88550
rect 3764 88452 3770 88504
rect 3822 88492 3828 88504
rect 3822 88464 5454 88492
rect 6168 88474 6452 88502
rect 3822 88452 3828 88464
rect 3512 88366 3518 88418
rect 3570 88406 3576 88418
rect 3570 88378 5358 88406
rect 3570 88366 3576 88378
rect 4688 88280 4694 88332
rect 4746 88320 4752 88332
rect 6376 88328 6452 88356
rect 4746 88292 5262 88320
rect 4746 88280 4752 88292
rect 3764 88194 3770 88246
rect 3822 88234 3828 88246
rect 3822 88206 5166 88234
rect 3822 88194 3828 88206
rect 3428 88108 3434 88160
rect 3486 88148 3492 88160
rect 3486 88120 5070 88148
rect 3486 88108 3492 88120
rect 6434 87640 6440 87692
rect 6492 87640 6498 87692
rect 3512 87172 3518 87224
rect 3570 87212 3576 87224
rect 3570 87184 5070 87212
rect 3570 87172 3576 87184
rect 3680 87086 3686 87138
rect 3738 87126 3744 87138
rect 3738 87098 5166 87126
rect 3738 87086 3744 87098
rect 4688 87000 4694 87052
rect 4746 87040 4752 87052
rect 4746 87012 5262 87040
rect 4746 87000 4752 87012
rect 6376 86976 6452 87004
rect 3260 86914 3266 86966
rect 3318 86954 3324 86966
rect 3318 86926 5358 86954
rect 3318 86914 3324 86926
rect 3764 86828 3770 86880
rect 3822 86868 3828 86880
rect 3822 86840 5454 86868
rect 3822 86828 3828 86840
rect 6168 86830 6452 86858
rect 4688 86742 4694 86794
rect 4746 86782 4752 86794
rect 4746 86754 5550 86782
rect 4746 86742 4752 86754
rect 6086 86708 6452 86736
rect 3344 86656 3350 86708
rect 3402 86696 3408 86708
rect 3402 86668 5754 86696
rect 3402 86656 3408 86668
rect 3764 86570 3770 86622
rect 3822 86610 3828 86622
rect 3822 86582 5850 86610
rect 3822 86570 3828 86582
rect 4688 86484 4694 86536
rect 4746 86524 4752 86536
rect 4746 86496 5946 86524
rect 4746 86484 4752 86496
rect 6434 86102 6440 86154
rect 6492 86102 6498 86154
rect 4688 85720 4694 85772
rect 4746 85760 4752 85772
rect 4746 85732 5946 85760
rect 4746 85720 4752 85732
rect 3680 85634 3686 85686
rect 3738 85674 3744 85686
rect 3738 85646 5850 85674
rect 3738 85634 3744 85646
rect 3428 85548 3434 85600
rect 3486 85588 3492 85600
rect 3486 85560 5754 85588
rect 3486 85548 3492 85560
rect 6086 85520 6452 85548
rect 4688 85462 4694 85514
rect 4746 85502 4752 85514
rect 4746 85474 5550 85502
rect 4746 85462 4752 85474
rect 3680 85376 3686 85428
rect 3738 85416 3744 85428
rect 3738 85388 5454 85416
rect 6168 85398 6452 85426
rect 3738 85376 3744 85388
rect 3344 85290 3350 85342
rect 3402 85330 3408 85342
rect 3402 85302 5358 85330
rect 3402 85290 3408 85302
rect 4688 85204 4694 85256
rect 4746 85244 4752 85256
rect 6376 85252 6452 85280
rect 4746 85216 5262 85244
rect 4746 85204 4752 85216
rect 3680 85118 3686 85170
rect 3738 85158 3744 85170
rect 3738 85130 5166 85158
rect 3738 85118 3744 85130
rect 3260 85032 3266 85084
rect 3318 85072 3324 85084
rect 3318 85044 5070 85072
rect 3318 85032 3324 85044
rect 6434 84564 6440 84616
rect 6492 84564 6498 84616
rect 3344 84096 3350 84148
rect 3402 84136 3408 84148
rect 3402 84108 5070 84136
rect 3402 84096 3408 84108
rect 3596 84010 3602 84062
rect 3654 84050 3660 84062
rect 3654 84022 5166 84050
rect 3654 84010 3660 84022
rect 4688 83924 4694 83976
rect 4746 83964 4752 83976
rect 4746 83936 5262 83964
rect 4746 83924 4752 83936
rect 6376 83900 6452 83928
rect 3428 83838 3434 83890
rect 3486 83878 3492 83890
rect 3486 83850 5358 83878
rect 3486 83838 3492 83850
rect 3596 83752 3602 83804
rect 3654 83792 3660 83804
rect 3654 83764 5454 83792
rect 3654 83752 3660 83764
rect 6168 83754 6452 83782
rect 4688 83666 4694 83718
rect 4746 83706 4752 83718
rect 4746 83678 5550 83706
rect 4746 83666 4752 83678
rect 6086 83632 6452 83660
rect 3512 83580 3518 83632
rect 3570 83620 3576 83632
rect 3570 83592 5754 83620
rect 3570 83580 3576 83592
rect 3596 83494 3602 83546
rect 3654 83534 3660 83546
rect 3654 83506 5850 83534
rect 3654 83494 3660 83506
rect 4688 83408 4694 83460
rect 4746 83448 4752 83460
rect 4746 83420 5946 83448
rect 4746 83408 4752 83420
rect 6434 83026 6440 83078
rect 6492 83026 6498 83078
rect 4688 82644 4694 82696
rect 4746 82684 4752 82696
rect 4746 82656 5946 82684
rect 4746 82644 4752 82656
rect 3596 82558 3602 82610
rect 3654 82598 3660 82610
rect 3654 82570 5850 82598
rect 3654 82558 3660 82570
rect 3260 82472 3266 82524
rect 3318 82512 3324 82524
rect 3318 82484 5754 82512
rect 3318 82472 3324 82484
rect 6086 82444 6452 82472
rect 4604 82386 4610 82438
rect 4662 82426 4668 82438
rect 4662 82398 5550 82426
rect 4662 82386 4668 82398
rect 4184 82300 4190 82352
rect 4242 82340 4248 82352
rect 4242 82312 5454 82340
rect 6168 82322 6452 82350
rect 4242 82300 4248 82312
rect 3512 82214 3518 82266
rect 3570 82254 3576 82266
rect 3570 82226 5358 82254
rect 3570 82214 3576 82226
rect 4604 82128 4610 82180
rect 4662 82168 4668 82180
rect 6376 82176 6452 82204
rect 4662 82140 5262 82168
rect 4662 82128 4668 82140
rect 4184 82042 4190 82094
rect 4242 82082 4248 82094
rect 4242 82054 5166 82082
rect 4242 82042 4248 82054
rect 3428 81956 3434 82008
rect 3486 81996 3492 82008
rect 3486 81968 5070 81996
rect 3486 81956 3492 81968
rect 6434 81488 6440 81540
rect 6492 81488 6498 81540
rect 3512 81020 3518 81072
rect 3570 81060 3576 81072
rect 3570 81032 5070 81060
rect 3570 81020 3576 81032
rect 4100 80934 4106 80986
rect 4158 80974 4164 80986
rect 4158 80946 5166 80974
rect 4158 80934 4164 80946
rect 4604 80848 4610 80900
rect 4662 80888 4668 80900
rect 4662 80860 5262 80888
rect 4662 80848 4668 80860
rect 6376 80824 6452 80852
rect 3260 80762 3266 80814
rect 3318 80802 3324 80814
rect 3318 80774 5358 80802
rect 3318 80762 3324 80774
rect 4184 80676 4190 80728
rect 4242 80716 4248 80728
rect 4242 80688 5454 80716
rect 4242 80676 4248 80688
rect 6168 80678 6452 80706
rect 4604 80590 4610 80642
rect 4662 80630 4668 80642
rect 4662 80602 5550 80630
rect 4662 80590 4668 80602
rect 6086 80556 6452 80584
rect 3344 80504 3350 80556
rect 3402 80544 3408 80556
rect 3402 80516 5754 80544
rect 3402 80504 3408 80516
rect 4184 80418 4190 80470
rect 4242 80458 4248 80470
rect 4242 80430 5850 80458
rect 4242 80418 4248 80430
rect 4604 80332 4610 80384
rect 4662 80372 4668 80384
rect 4662 80344 5946 80372
rect 4662 80332 4668 80344
rect 6434 79950 6440 80002
rect 6492 79950 6498 80002
rect 4604 79568 4610 79620
rect 4662 79608 4668 79620
rect 4662 79580 5946 79608
rect 4662 79568 4668 79580
rect 4100 79482 4106 79534
rect 4158 79522 4164 79534
rect 4158 79494 5850 79522
rect 4158 79482 4164 79494
rect 3428 79396 3434 79448
rect 3486 79436 3492 79448
rect 3486 79408 5754 79436
rect 3486 79396 3492 79408
rect 6086 79368 6452 79396
rect 4604 79310 4610 79362
rect 4662 79350 4668 79362
rect 4662 79322 5550 79350
rect 4662 79310 4668 79322
rect 4100 79224 4106 79276
rect 4158 79264 4164 79276
rect 4158 79236 5454 79264
rect 6168 79246 6452 79274
rect 4158 79224 4164 79236
rect 3344 79138 3350 79190
rect 3402 79178 3408 79190
rect 3402 79150 5358 79178
rect 3402 79138 3408 79150
rect 4604 79052 4610 79104
rect 4662 79092 4668 79104
rect 6376 79100 6452 79128
rect 4662 79064 5262 79092
rect 4662 79052 4668 79064
rect 4100 78966 4106 79018
rect 4158 79006 4164 79018
rect 4158 78978 5166 79006
rect 4158 78966 4164 78978
rect 3260 78880 3266 78932
rect 3318 78920 3324 78932
rect 3318 78892 5070 78920
rect 3318 78880 3324 78892
rect 6434 78412 6440 78464
rect 6492 78412 6498 78464
rect 3344 77944 3350 77996
rect 3402 77984 3408 77996
rect 3402 77956 5070 77984
rect 3402 77944 3408 77956
rect 4016 77858 4022 77910
rect 4074 77898 4080 77910
rect 4074 77870 5166 77898
rect 4074 77858 4080 77870
rect 4604 77772 4610 77824
rect 4662 77812 4668 77824
rect 4662 77784 5262 77812
rect 4662 77772 4668 77784
rect 6376 77748 6452 77776
rect 3428 77686 3434 77738
rect 3486 77726 3492 77738
rect 3486 77698 5358 77726
rect 3486 77686 3492 77698
rect 4016 77600 4022 77652
rect 4074 77640 4080 77652
rect 4074 77612 5454 77640
rect 4074 77600 4080 77612
rect 6168 77602 6452 77630
rect 4604 77514 4610 77566
rect 4662 77554 4668 77566
rect 4662 77526 5550 77554
rect 4662 77514 4668 77526
rect 6086 77480 6452 77508
rect 3512 77428 3518 77480
rect 3570 77468 3576 77480
rect 3570 77440 5754 77468
rect 3570 77428 3576 77440
rect 4016 77342 4022 77394
rect 4074 77382 4080 77394
rect 4074 77354 5850 77382
rect 4074 77342 4080 77354
rect 4604 77256 4610 77308
rect 4662 77296 4668 77308
rect 4662 77268 5946 77296
rect 4662 77256 4668 77268
rect 6434 76874 6440 76926
rect 6492 76874 6498 76926
rect 4604 76492 4610 76544
rect 4662 76532 4668 76544
rect 4662 76504 5946 76532
rect 4662 76492 4668 76504
rect 4016 76406 4022 76458
rect 4074 76446 4080 76458
rect 4074 76418 5850 76446
rect 4074 76406 4080 76418
rect 3260 76320 3266 76372
rect 3318 76360 3324 76372
rect 3318 76332 5754 76360
rect 3318 76320 3324 76332
rect 6086 76292 6452 76320
rect 4604 76234 4610 76286
rect 4662 76274 4668 76286
rect 4662 76246 5550 76274
rect 4662 76234 4668 76246
rect 3932 76148 3938 76200
rect 3990 76188 3996 76200
rect 3990 76160 5454 76188
rect 6168 76170 6452 76198
rect 3990 76148 3996 76160
rect 3512 76062 3518 76114
rect 3570 76102 3576 76114
rect 3570 76074 5358 76102
rect 3570 76062 3576 76074
rect 4604 75976 4610 76028
rect 4662 76016 4668 76028
rect 6376 76024 6452 76052
rect 4662 75988 5262 76016
rect 4662 75976 4668 75988
rect 3932 75890 3938 75942
rect 3990 75930 3996 75942
rect 3990 75902 5166 75930
rect 3990 75890 3996 75902
rect 3428 75804 3434 75856
rect 3486 75844 3492 75856
rect 3486 75816 5070 75844
rect 3486 75804 3492 75816
rect 6434 75336 6440 75388
rect 6492 75336 6498 75388
rect 3512 74868 3518 74920
rect 3570 74908 3576 74920
rect 3570 74880 5070 74908
rect 3570 74868 3576 74880
rect 3848 74782 3854 74834
rect 3906 74822 3912 74834
rect 3906 74794 5166 74822
rect 3906 74782 3912 74794
rect 4604 74696 4610 74748
rect 4662 74736 4668 74748
rect 4662 74708 5262 74736
rect 4662 74696 4668 74708
rect 6376 74672 6452 74700
rect 3260 74610 3266 74662
rect 3318 74650 3324 74662
rect 3318 74622 5358 74650
rect 3318 74610 3324 74622
rect 3932 74524 3938 74576
rect 3990 74564 3996 74576
rect 3990 74536 5454 74564
rect 3990 74524 3996 74536
rect 6168 74526 6452 74554
rect 4604 74438 4610 74490
rect 4662 74478 4668 74490
rect 4662 74450 5550 74478
rect 4662 74438 4668 74450
rect 6086 74404 6452 74432
rect 3344 74352 3350 74404
rect 3402 74392 3408 74404
rect 3402 74364 5754 74392
rect 3402 74352 3408 74364
rect 3932 74266 3938 74318
rect 3990 74306 3996 74318
rect 3990 74278 5850 74306
rect 3990 74266 3996 74278
rect 4604 74180 4610 74232
rect 4662 74220 4668 74232
rect 4662 74192 5946 74220
rect 4662 74180 4668 74192
rect 6434 73798 6440 73850
rect 6492 73798 6498 73850
rect 4604 73416 4610 73468
rect 4662 73456 4668 73468
rect 4662 73428 5946 73456
rect 4662 73416 4668 73428
rect 3848 73330 3854 73382
rect 3906 73370 3912 73382
rect 3906 73342 5850 73370
rect 3906 73330 3912 73342
rect 3428 73244 3434 73296
rect 3486 73284 3492 73296
rect 3486 73256 5754 73284
rect 3486 73244 3492 73256
rect 6086 73216 6452 73244
rect 4604 73158 4610 73210
rect 4662 73198 4668 73210
rect 4662 73170 5550 73198
rect 4662 73158 4668 73170
rect 3848 73072 3854 73124
rect 3906 73112 3912 73124
rect 3906 73084 5454 73112
rect 6168 73094 6452 73122
rect 3906 73072 3912 73084
rect 3344 72986 3350 73038
rect 3402 73026 3408 73038
rect 3402 72998 5358 73026
rect 3402 72986 3408 72998
rect 4604 72900 4610 72952
rect 4662 72940 4668 72952
rect 6376 72948 6452 72976
rect 4662 72912 5262 72940
rect 4662 72900 4668 72912
rect 3848 72814 3854 72866
rect 3906 72854 3912 72866
rect 3906 72826 5166 72854
rect 3906 72814 3912 72826
rect 3260 72728 3266 72780
rect 3318 72768 3324 72780
rect 3318 72740 5070 72768
rect 3318 72728 3324 72740
rect 6434 72260 6440 72312
rect 6492 72260 6498 72312
rect 3344 71792 3350 71844
rect 3402 71832 3408 71844
rect 3402 71804 5070 71832
rect 3402 71792 3408 71804
rect 3764 71706 3770 71758
rect 3822 71746 3828 71758
rect 3822 71718 5166 71746
rect 3822 71706 3828 71718
rect 4604 71620 4610 71672
rect 4662 71660 4668 71672
rect 4662 71632 5262 71660
rect 4662 71620 4668 71632
rect 6376 71596 6452 71624
rect 3428 71534 3434 71586
rect 3486 71574 3492 71586
rect 3486 71546 5358 71574
rect 3486 71534 3492 71546
rect 3764 71448 3770 71500
rect 3822 71488 3828 71500
rect 3822 71460 5454 71488
rect 3822 71448 3828 71460
rect 6168 71450 6452 71478
rect 4604 71362 4610 71414
rect 4662 71402 4668 71414
rect 4662 71374 5550 71402
rect 4662 71362 4668 71374
rect 6086 71328 6452 71356
rect 3512 71276 3518 71328
rect 3570 71316 3576 71328
rect 3570 71288 5754 71316
rect 3570 71276 3576 71288
rect 3764 71190 3770 71242
rect 3822 71230 3828 71242
rect 3822 71202 5850 71230
rect 3822 71190 3828 71202
rect 4604 71104 4610 71156
rect 4662 71144 4668 71156
rect 4662 71116 5946 71144
rect 4662 71104 4668 71116
rect 6434 70722 6440 70774
rect 6492 70722 6498 70774
rect 4604 70340 4610 70392
rect 4662 70380 4668 70392
rect 4662 70352 5946 70380
rect 4662 70340 4668 70352
rect 3764 70254 3770 70306
rect 3822 70294 3828 70306
rect 3822 70266 5850 70294
rect 3822 70254 3828 70266
rect 3260 70168 3266 70220
rect 3318 70208 3324 70220
rect 3318 70180 5754 70208
rect 3318 70168 3324 70180
rect 6086 70140 6452 70168
rect 4604 70082 4610 70134
rect 4662 70122 4668 70134
rect 4662 70094 5550 70122
rect 4662 70082 4668 70094
rect 3680 69996 3686 70048
rect 3738 70036 3744 70048
rect 3738 70008 5454 70036
rect 6168 70018 6452 70046
rect 3738 69996 3744 70008
rect 3512 69910 3518 69962
rect 3570 69950 3576 69962
rect 3570 69922 5358 69950
rect 3570 69910 3576 69922
rect 4604 69824 4610 69876
rect 4662 69864 4668 69876
rect 6376 69872 6452 69900
rect 4662 69836 5262 69864
rect 4662 69824 4668 69836
rect 3680 69738 3686 69790
rect 3738 69778 3744 69790
rect 3738 69750 5166 69778
rect 3738 69738 3744 69750
rect 3428 69652 3434 69704
rect 3486 69692 3492 69704
rect 3486 69664 5070 69692
rect 3486 69652 3492 69664
rect 6434 69184 6440 69236
rect 6492 69184 6498 69236
rect 3512 68716 3518 68768
rect 3570 68756 3576 68768
rect 3570 68728 5070 68756
rect 3570 68716 3576 68728
rect 3596 68630 3602 68682
rect 3654 68670 3660 68682
rect 3654 68642 5166 68670
rect 3654 68630 3660 68642
rect 4604 68544 4610 68596
rect 4662 68584 4668 68596
rect 4662 68556 5262 68584
rect 4662 68544 4668 68556
rect 6376 68520 6452 68548
rect 3260 68458 3266 68510
rect 3318 68498 3324 68510
rect 3318 68470 5358 68498
rect 3318 68458 3324 68470
rect 3680 68372 3686 68424
rect 3738 68412 3744 68424
rect 3738 68384 5454 68412
rect 3738 68372 3744 68384
rect 6168 68374 6452 68402
rect 4604 68286 4610 68338
rect 4662 68326 4668 68338
rect 4662 68298 5550 68326
rect 4662 68286 4668 68298
rect 6086 68252 6452 68280
rect 3344 68200 3350 68252
rect 3402 68240 3408 68252
rect 3402 68212 5754 68240
rect 3402 68200 3408 68212
rect 3680 68114 3686 68166
rect 3738 68154 3744 68166
rect 3738 68126 5850 68154
rect 3738 68114 3744 68126
rect 4604 68028 4610 68080
rect 4662 68068 4668 68080
rect 4662 68040 5946 68068
rect 4662 68028 4668 68040
rect 6434 67646 6440 67698
rect 6492 67646 6498 67698
rect 4604 67264 4610 67316
rect 4662 67304 4668 67316
rect 4662 67276 5946 67304
rect 4662 67264 4668 67276
rect 3596 67178 3602 67230
rect 3654 67218 3660 67230
rect 3654 67190 5850 67218
rect 3654 67178 3660 67190
rect 3428 67092 3434 67144
rect 3486 67132 3492 67144
rect 3486 67104 5754 67132
rect 3486 67092 3492 67104
rect 6086 67064 6452 67092
rect 4604 67006 4610 67058
rect 4662 67046 4668 67058
rect 4662 67018 5550 67046
rect 4662 67006 4668 67018
rect 3596 66920 3602 66972
rect 3654 66960 3660 66972
rect 3654 66932 5454 66960
rect 6168 66942 6452 66970
rect 3654 66920 3660 66932
rect 3344 66834 3350 66886
rect 3402 66874 3408 66886
rect 3402 66846 5358 66874
rect 3402 66834 3408 66846
rect 4604 66748 4610 66800
rect 4662 66788 4668 66800
rect 6376 66796 6452 66824
rect 4662 66760 5262 66788
rect 4662 66748 4668 66760
rect 3596 66662 3602 66714
rect 3654 66702 3660 66714
rect 3654 66674 5166 66702
rect 3654 66662 3660 66674
rect 3260 66576 3266 66628
rect 3318 66616 3324 66628
rect 3318 66588 5070 66616
rect 3318 66576 3324 66588
rect 6434 66108 6440 66160
rect 6492 66108 6498 66160
rect 3344 65640 3350 65692
rect 3402 65680 3408 65692
rect 3402 65652 5070 65680
rect 3402 65640 3408 65652
rect 4184 65554 4190 65606
rect 4242 65594 4248 65606
rect 4242 65566 5166 65594
rect 4242 65554 4248 65566
rect 4520 65468 4526 65520
rect 4578 65508 4584 65520
rect 4578 65480 5262 65508
rect 4578 65468 4584 65480
rect 6376 65444 6452 65472
rect 3428 65382 3434 65434
rect 3486 65422 3492 65434
rect 3486 65394 5358 65422
rect 3486 65382 3492 65394
rect 4184 65296 4190 65348
rect 4242 65336 4248 65348
rect 4242 65308 5454 65336
rect 4242 65296 4248 65308
rect 6168 65298 6452 65326
rect 4520 65210 4526 65262
rect 4578 65250 4584 65262
rect 4578 65222 5550 65250
rect 4578 65210 4584 65222
rect 6086 65176 6452 65204
rect 3512 65124 3518 65176
rect 3570 65164 3576 65176
rect 3570 65136 5754 65164
rect 3570 65124 3576 65136
rect 4184 65038 4190 65090
rect 4242 65078 4248 65090
rect 4242 65050 5850 65078
rect 4242 65038 4248 65050
rect 4520 64952 4526 65004
rect 4578 64992 4584 65004
rect 4578 64964 5946 64992
rect 4578 64952 4584 64964
rect 6434 64570 6440 64622
rect 6492 64570 6498 64622
rect 4520 64188 4526 64240
rect 4578 64228 4584 64240
rect 4578 64200 5946 64228
rect 4578 64188 4584 64200
rect 4184 64102 4190 64154
rect 4242 64142 4248 64154
rect 4242 64114 5850 64142
rect 4242 64102 4248 64114
rect 3260 64016 3266 64068
rect 3318 64056 3324 64068
rect 3318 64028 5754 64056
rect 3318 64016 3324 64028
rect 6086 63988 6452 64016
rect 4520 63930 4526 63982
rect 4578 63970 4584 63982
rect 4578 63942 5550 63970
rect 4578 63930 4584 63942
rect 4100 63844 4106 63896
rect 4158 63884 4164 63896
rect 4158 63856 5454 63884
rect 6168 63866 6452 63894
rect 4158 63844 4164 63856
rect 3512 63758 3518 63810
rect 3570 63798 3576 63810
rect 3570 63770 5358 63798
rect 3570 63758 3576 63770
rect 4520 63672 4526 63724
rect 4578 63712 4584 63724
rect 6376 63720 6452 63748
rect 4578 63684 5262 63712
rect 4578 63672 4584 63684
rect 4100 63586 4106 63638
rect 4158 63626 4164 63638
rect 4158 63598 5166 63626
rect 4158 63586 4164 63598
rect 3428 63500 3434 63552
rect 3486 63540 3492 63552
rect 3486 63512 5070 63540
rect 3486 63500 3492 63512
rect 6434 63032 6440 63084
rect 6492 63032 6498 63084
rect 3512 62564 3518 62616
rect 3570 62604 3576 62616
rect 3570 62576 5070 62604
rect 3570 62564 3576 62576
rect 4016 62478 4022 62530
rect 4074 62518 4080 62530
rect 4074 62490 5166 62518
rect 4074 62478 4080 62490
rect 4520 62392 4526 62444
rect 4578 62432 4584 62444
rect 4578 62404 5262 62432
rect 4578 62392 4584 62404
rect 6376 62368 6452 62396
rect 3260 62306 3266 62358
rect 3318 62346 3324 62358
rect 3318 62318 5358 62346
rect 3318 62306 3324 62318
rect 4100 62220 4106 62272
rect 4158 62260 4164 62272
rect 4158 62232 5454 62260
rect 4158 62220 4164 62232
rect 6168 62222 6452 62250
rect 4520 62134 4526 62186
rect 4578 62174 4584 62186
rect 4578 62146 5550 62174
rect 4578 62134 4584 62146
rect 6086 62100 6452 62128
rect 3344 62048 3350 62100
rect 3402 62088 3408 62100
rect 3402 62060 5754 62088
rect 3402 62048 3408 62060
rect 4100 61962 4106 62014
rect 4158 62002 4164 62014
rect 4158 61974 5850 62002
rect 4158 61962 4164 61974
rect 4520 61876 4526 61928
rect 4578 61916 4584 61928
rect 4578 61888 5946 61916
rect 4578 61876 4584 61888
rect 6434 61494 6440 61546
rect 6492 61494 6498 61546
rect 4520 61112 4526 61164
rect 4578 61152 4584 61164
rect 4578 61124 5946 61152
rect 4578 61112 4584 61124
rect 4016 61026 4022 61078
rect 4074 61066 4080 61078
rect 4074 61038 5850 61066
rect 4074 61026 4080 61038
rect 3428 60940 3434 60992
rect 3486 60980 3492 60992
rect 3486 60952 5754 60980
rect 3486 60940 3492 60952
rect 6086 60912 6452 60940
rect 4520 60854 4526 60906
rect 4578 60894 4584 60906
rect 4578 60866 5550 60894
rect 4578 60854 4584 60866
rect 4016 60768 4022 60820
rect 4074 60808 4080 60820
rect 4074 60780 5454 60808
rect 6168 60790 6452 60818
rect 4074 60768 4080 60780
rect 3344 60682 3350 60734
rect 3402 60722 3408 60734
rect 3402 60694 5358 60722
rect 3402 60682 3408 60694
rect 4520 60596 4526 60648
rect 4578 60636 4584 60648
rect 6376 60644 6452 60672
rect 4578 60608 5262 60636
rect 4578 60596 4584 60608
rect 4016 60510 4022 60562
rect 4074 60550 4080 60562
rect 4074 60522 5166 60550
rect 4074 60510 4080 60522
rect 3260 60424 3266 60476
rect 3318 60464 3324 60476
rect 3318 60436 5070 60464
rect 3318 60424 3324 60436
rect 6434 59956 6440 60008
rect 6492 59956 6498 60008
rect 3344 59488 3350 59540
rect 3402 59528 3408 59540
rect 3402 59500 5070 59528
rect 3402 59488 3408 59500
rect 3932 59402 3938 59454
rect 3990 59442 3996 59454
rect 3990 59414 5166 59442
rect 3990 59402 3996 59414
rect 4520 59316 4526 59368
rect 4578 59356 4584 59368
rect 4578 59328 5262 59356
rect 4578 59316 4584 59328
rect 6376 59292 6452 59320
rect 3428 59230 3434 59282
rect 3486 59270 3492 59282
rect 3486 59242 5358 59270
rect 3486 59230 3492 59242
rect 3932 59144 3938 59196
rect 3990 59184 3996 59196
rect 3990 59156 5454 59184
rect 3990 59144 3996 59156
rect 6168 59146 6452 59174
rect 4520 59058 4526 59110
rect 4578 59098 4584 59110
rect 4578 59070 5550 59098
rect 4578 59058 4584 59070
rect 6086 59024 6452 59052
rect 3512 58972 3518 59024
rect 3570 59012 3576 59024
rect 3570 58984 5754 59012
rect 3570 58972 3576 58984
rect 3932 58886 3938 58938
rect 3990 58926 3996 58938
rect 3990 58898 5850 58926
rect 3990 58886 3996 58898
rect 4520 58800 4526 58852
rect 4578 58840 4584 58852
rect 4578 58812 5946 58840
rect 4578 58800 4584 58812
rect 6434 58418 6440 58470
rect 6492 58418 6498 58470
rect 4520 58036 4526 58088
rect 4578 58076 4584 58088
rect 4578 58048 5946 58076
rect 4578 58036 4584 58048
rect 3932 57950 3938 58002
rect 3990 57990 3996 58002
rect 3990 57962 5850 57990
rect 3990 57950 3996 57962
rect 3260 57864 3266 57916
rect 3318 57904 3324 57916
rect 3318 57876 5754 57904
rect 3318 57864 3324 57876
rect 6086 57836 6452 57864
rect 4520 57778 4526 57830
rect 4578 57818 4584 57830
rect 4578 57790 5550 57818
rect 4578 57778 4584 57790
rect 3848 57692 3854 57744
rect 3906 57732 3912 57744
rect 3906 57704 5454 57732
rect 6168 57714 6452 57742
rect 3906 57692 3912 57704
rect 3512 57606 3518 57658
rect 3570 57646 3576 57658
rect 3570 57618 5358 57646
rect 3570 57606 3576 57618
rect 4520 57520 4526 57572
rect 4578 57560 4584 57572
rect 6376 57568 6452 57596
rect 4578 57532 5262 57560
rect 4578 57520 4584 57532
rect 3848 57434 3854 57486
rect 3906 57474 3912 57486
rect 3906 57446 5166 57474
rect 3906 57434 3912 57446
rect 3428 57348 3434 57400
rect 3486 57388 3492 57400
rect 3486 57360 5070 57388
rect 3486 57348 3492 57360
rect 6434 56880 6440 56932
rect 6492 56880 6498 56932
rect 3512 56412 3518 56464
rect 3570 56452 3576 56464
rect 3570 56424 5070 56452
rect 3570 56412 3576 56424
rect 3764 56326 3770 56378
rect 3822 56366 3828 56378
rect 3822 56338 5166 56366
rect 3822 56326 3828 56338
rect 4520 56240 4526 56292
rect 4578 56280 4584 56292
rect 4578 56252 5262 56280
rect 4578 56240 4584 56252
rect 6376 56216 6452 56244
rect 3260 56154 3266 56206
rect 3318 56194 3324 56206
rect 3318 56166 5358 56194
rect 3318 56154 3324 56166
rect 3848 56068 3854 56120
rect 3906 56108 3912 56120
rect 3906 56080 5454 56108
rect 3906 56068 3912 56080
rect 6168 56070 6452 56098
rect 4520 55982 4526 56034
rect 4578 56022 4584 56034
rect 4578 55994 5550 56022
rect 4578 55982 4584 55994
rect 6086 55948 6452 55976
rect 3344 55896 3350 55948
rect 3402 55936 3408 55948
rect 3402 55908 5754 55936
rect 3402 55896 3408 55908
rect 3848 55810 3854 55862
rect 3906 55850 3912 55862
rect 3906 55822 5850 55850
rect 3906 55810 3912 55822
rect 4520 55724 4526 55776
rect 4578 55764 4584 55776
rect 4578 55736 5946 55764
rect 4578 55724 4584 55736
rect 6434 55342 6440 55394
rect 6492 55342 6498 55394
rect 4520 54960 4526 55012
rect 4578 55000 4584 55012
rect 4578 54972 5946 55000
rect 4578 54960 4584 54972
rect 3764 54874 3770 54926
rect 3822 54914 3828 54926
rect 3822 54886 5850 54914
rect 3822 54874 3828 54886
rect 3428 54788 3434 54840
rect 3486 54828 3492 54840
rect 3486 54800 5754 54828
rect 3486 54788 3492 54800
rect 6086 54760 6452 54788
rect 4520 54702 4526 54754
rect 4578 54742 4584 54754
rect 4578 54714 5550 54742
rect 4578 54702 4584 54714
rect 3764 54616 3770 54668
rect 3822 54656 3828 54668
rect 3822 54628 5454 54656
rect 6168 54638 6452 54666
rect 3822 54616 3828 54628
rect 3344 54530 3350 54582
rect 3402 54570 3408 54582
rect 3402 54542 5358 54570
rect 3402 54530 3408 54542
rect 4520 54444 4526 54496
rect 4578 54484 4584 54496
rect 6376 54492 6452 54520
rect 4578 54456 5262 54484
rect 4578 54444 4584 54456
rect 3764 54358 3770 54410
rect 3822 54398 3828 54410
rect 3822 54370 5166 54398
rect 3822 54358 3828 54370
rect 3260 54272 3266 54324
rect 3318 54312 3324 54324
rect 3318 54284 5070 54312
rect 3318 54272 3324 54284
rect 6434 53804 6440 53856
rect 6492 53804 6498 53856
rect 3344 53336 3350 53388
rect 3402 53376 3408 53388
rect 3402 53348 5070 53376
rect 3402 53336 3408 53348
rect 3680 53250 3686 53302
rect 3738 53290 3744 53302
rect 3738 53262 5166 53290
rect 3738 53250 3744 53262
rect 4520 53164 4526 53216
rect 4578 53204 4584 53216
rect 4578 53176 5262 53204
rect 4578 53164 4584 53176
rect 6376 53140 6452 53168
rect 3428 53078 3434 53130
rect 3486 53118 3492 53130
rect 3486 53090 5358 53118
rect 3486 53078 3492 53090
rect 3680 52992 3686 53044
rect 3738 53032 3744 53044
rect 3738 53004 5454 53032
rect 3738 52992 3744 53004
rect 6168 52994 6452 53022
rect 4520 52906 4526 52958
rect 4578 52946 4584 52958
rect 4578 52918 5550 52946
rect 4578 52906 4584 52918
rect 6086 52872 6452 52900
rect 3512 52820 3518 52872
rect 3570 52860 3576 52872
rect 3570 52832 5754 52860
rect 3570 52820 3576 52832
rect 3680 52734 3686 52786
rect 3738 52774 3744 52786
rect 3738 52746 5850 52774
rect 3738 52734 3744 52746
rect 4520 52648 4526 52700
rect 4578 52688 4584 52700
rect 4578 52660 5946 52688
rect 4578 52648 4584 52660
rect 6434 52266 6440 52318
rect 6492 52266 6498 52318
rect 4520 51884 4526 51936
rect 4578 51924 4584 51936
rect 4578 51896 5946 51924
rect 4578 51884 4584 51896
rect 3680 51798 3686 51850
rect 3738 51838 3744 51850
rect 3738 51810 5850 51838
rect 3738 51798 3744 51810
rect 3260 51712 3266 51764
rect 3318 51752 3324 51764
rect 3318 51724 5754 51752
rect 3318 51712 3324 51724
rect 6086 51684 6452 51712
rect 4520 51626 4526 51678
rect 4578 51666 4584 51678
rect 4578 51638 5550 51666
rect 4578 51626 4584 51638
rect 3596 51540 3602 51592
rect 3654 51580 3660 51592
rect 3654 51552 5454 51580
rect 6168 51562 6452 51590
rect 3654 51540 3660 51552
rect 3512 51454 3518 51506
rect 3570 51494 3576 51506
rect 3570 51466 5358 51494
rect 3570 51454 3576 51466
rect 4520 51368 4526 51420
rect 4578 51408 4584 51420
rect 6376 51416 6452 51444
rect 4578 51380 5262 51408
rect 4578 51368 4584 51380
rect 3596 51282 3602 51334
rect 3654 51322 3660 51334
rect 3654 51294 5166 51322
rect 3654 51282 3660 51294
rect 3428 51196 3434 51248
rect 3486 51236 3492 51248
rect 3486 51208 5070 51236
rect 3486 51196 3492 51208
rect 6434 50728 6440 50780
rect 6492 50728 6498 50780
rect 3512 50260 3518 50312
rect 3570 50300 3576 50312
rect 3570 50272 5070 50300
rect 3570 50260 3576 50272
rect 4184 50174 4190 50226
rect 4242 50214 4248 50226
rect 4242 50186 5166 50214
rect 4242 50174 4248 50186
rect 4436 50088 4442 50140
rect 4494 50128 4500 50140
rect 4494 50100 5262 50128
rect 4494 50088 4500 50100
rect 6376 50064 6452 50092
rect 3260 50002 3266 50054
rect 3318 50042 3324 50054
rect 3318 50014 5358 50042
rect 3318 50002 3324 50014
rect 3596 49916 3602 49968
rect 3654 49956 3660 49968
rect 3654 49928 5454 49956
rect 3654 49916 3660 49928
rect 6168 49918 6452 49946
rect 4520 49830 4526 49882
rect 4578 49870 4584 49882
rect 4578 49842 5550 49870
rect 4578 49830 4584 49842
rect 6086 49796 6452 49824
rect 3344 49744 3350 49796
rect 3402 49784 3408 49796
rect 3402 49756 5754 49784
rect 3402 49744 3408 49756
rect 3596 49658 3602 49710
rect 3654 49698 3660 49710
rect 3654 49670 5850 49698
rect 3654 49658 3660 49670
rect 4520 49572 4526 49624
rect 4578 49612 4584 49624
rect 4578 49584 5946 49612
rect 4578 49572 4584 49584
rect 6434 49190 6440 49242
rect 6492 49190 6498 49242
rect 4436 48808 4442 48860
rect 4494 48848 4500 48860
rect 4494 48820 5946 48848
rect 4494 48808 4500 48820
rect 4184 48722 4190 48774
rect 4242 48762 4248 48774
rect 4242 48734 5850 48762
rect 4242 48722 4248 48734
rect 3428 48636 3434 48688
rect 3486 48676 3492 48688
rect 3486 48648 5754 48676
rect 3486 48636 3492 48648
rect 6086 48608 6452 48636
rect 4436 48550 4442 48602
rect 4494 48590 4500 48602
rect 4494 48562 5550 48590
rect 4494 48550 4500 48562
rect 4184 48464 4190 48516
rect 4242 48504 4248 48516
rect 4242 48476 5454 48504
rect 6168 48486 6452 48514
rect 4242 48464 4248 48476
rect 3344 48378 3350 48430
rect 3402 48418 3408 48430
rect 3402 48390 5358 48418
rect 3402 48378 3408 48390
rect 4436 48292 4442 48344
rect 4494 48332 4500 48344
rect 6376 48340 6452 48368
rect 4494 48304 5262 48332
rect 4494 48292 4500 48304
rect 4184 48206 4190 48258
rect 4242 48246 4248 48258
rect 4242 48218 5166 48246
rect 4242 48206 4248 48218
rect 3260 48120 3266 48172
rect 3318 48160 3324 48172
rect 3318 48132 5070 48160
rect 3318 48120 3324 48132
rect 6434 47652 6440 47704
rect 6492 47652 6498 47704
rect 3344 47184 3350 47236
rect 3402 47224 3408 47236
rect 3402 47196 5070 47224
rect 3402 47184 3408 47196
rect 4100 47098 4106 47150
rect 4158 47138 4164 47150
rect 4158 47110 5166 47138
rect 4158 47098 4164 47110
rect 4436 47012 4442 47064
rect 4494 47052 4500 47064
rect 4494 47024 5262 47052
rect 4494 47012 4500 47024
rect 6376 46988 6452 47016
rect 3428 46926 3434 46978
rect 3486 46966 3492 46978
rect 3486 46938 5358 46966
rect 3486 46926 3492 46938
rect 4100 46840 4106 46892
rect 4158 46880 4164 46892
rect 4158 46852 5454 46880
rect 4158 46840 4164 46852
rect 6168 46842 6452 46870
rect 4436 46754 4442 46806
rect 4494 46794 4500 46806
rect 4494 46766 5550 46794
rect 4494 46754 4500 46766
rect 6086 46720 6452 46748
rect 3512 46668 3518 46720
rect 3570 46708 3576 46720
rect 3570 46680 5754 46708
rect 3570 46668 3576 46680
rect 4100 46582 4106 46634
rect 4158 46622 4164 46634
rect 4158 46594 5850 46622
rect 4158 46582 4164 46594
rect 4436 46496 4442 46548
rect 4494 46536 4500 46548
rect 4494 46508 5946 46536
rect 4494 46496 4500 46508
rect 6434 46114 6440 46166
rect 6492 46114 6498 46166
rect 4436 45732 4442 45784
rect 4494 45772 4500 45784
rect 4494 45744 5946 45772
rect 4494 45732 4500 45744
rect 4100 45646 4106 45698
rect 4158 45686 4164 45698
rect 4158 45658 5850 45686
rect 4158 45646 4164 45658
rect 3260 45560 3266 45612
rect 3318 45600 3324 45612
rect 3318 45572 5754 45600
rect 3318 45560 3324 45572
rect 6086 45532 6452 45560
rect 4436 45474 4442 45526
rect 4494 45514 4500 45526
rect 4494 45486 5550 45514
rect 4494 45474 4500 45486
rect 4016 45388 4022 45440
rect 4074 45428 4080 45440
rect 4074 45400 5454 45428
rect 6168 45410 6452 45438
rect 4074 45388 4080 45400
rect 3512 45302 3518 45354
rect 3570 45342 3576 45354
rect 3570 45314 5358 45342
rect 3570 45302 3576 45314
rect 4436 45216 4442 45268
rect 4494 45256 4500 45268
rect 6376 45264 6452 45292
rect 4494 45228 5262 45256
rect 4494 45216 4500 45228
rect 4016 45130 4022 45182
rect 4074 45170 4080 45182
rect 4074 45142 5166 45170
rect 4074 45130 4080 45142
rect 3428 45044 3434 45096
rect 3486 45084 3492 45096
rect 3486 45056 5070 45084
rect 3486 45044 3492 45056
rect 6434 44576 6440 44628
rect 6492 44576 6498 44628
rect 3512 44108 3518 44160
rect 3570 44148 3576 44160
rect 3570 44120 5070 44148
rect 3570 44108 3576 44120
rect 3932 44022 3938 44074
rect 3990 44062 3996 44074
rect 3990 44034 5166 44062
rect 3990 44022 3996 44034
rect 4436 43936 4442 43988
rect 4494 43976 4500 43988
rect 4494 43948 5262 43976
rect 4494 43936 4500 43948
rect 6376 43912 6452 43940
rect 3260 43850 3266 43902
rect 3318 43890 3324 43902
rect 3318 43862 5358 43890
rect 3318 43850 3324 43862
rect 4016 43764 4022 43816
rect 4074 43804 4080 43816
rect 4074 43776 5454 43804
rect 4074 43764 4080 43776
rect 6168 43766 6452 43794
rect 4436 43678 4442 43730
rect 4494 43718 4500 43730
rect 4494 43690 5550 43718
rect 4494 43678 4500 43690
rect 6086 43644 6452 43672
rect 3344 43592 3350 43644
rect 3402 43632 3408 43644
rect 3402 43604 5754 43632
rect 3402 43592 3408 43604
rect 4016 43506 4022 43558
rect 4074 43546 4080 43558
rect 4074 43518 5850 43546
rect 4074 43506 4080 43518
rect 4436 43420 4442 43472
rect 4494 43460 4500 43472
rect 4494 43432 5946 43460
rect 4494 43420 4500 43432
rect 6434 43038 6440 43090
rect 6492 43038 6498 43090
rect 4436 42656 4442 42708
rect 4494 42696 4500 42708
rect 4494 42668 5946 42696
rect 4494 42656 4500 42668
rect 3932 42570 3938 42622
rect 3990 42610 3996 42622
rect 3990 42582 5850 42610
rect 3990 42570 3996 42582
rect 3428 42484 3434 42536
rect 3486 42524 3492 42536
rect 3486 42496 5754 42524
rect 3486 42484 3492 42496
rect 6086 42456 6452 42484
rect 4436 42398 4442 42450
rect 4494 42438 4500 42450
rect 4494 42410 5550 42438
rect 4494 42398 4500 42410
rect 3932 42312 3938 42364
rect 3990 42352 3996 42364
rect 3990 42324 5454 42352
rect 6168 42334 6452 42362
rect 3990 42312 3996 42324
rect 3344 42226 3350 42278
rect 3402 42266 3408 42278
rect 3402 42238 5358 42266
rect 3402 42226 3408 42238
rect 4436 42140 4442 42192
rect 4494 42180 4500 42192
rect 6376 42188 6452 42216
rect 4494 42152 5262 42180
rect 4494 42140 4500 42152
rect 3932 42054 3938 42106
rect 3990 42094 3996 42106
rect 3990 42066 5166 42094
rect 3990 42054 3996 42066
rect 3260 41968 3266 42020
rect 3318 42008 3324 42020
rect 3318 41980 5070 42008
rect 3318 41968 3324 41980
rect 6434 41500 6440 41552
rect 6492 41500 6498 41552
rect 3344 41032 3350 41084
rect 3402 41072 3408 41084
rect 3402 41044 5070 41072
rect 3402 41032 3408 41044
rect 3848 40946 3854 40998
rect 3906 40986 3912 40998
rect 3906 40958 5166 40986
rect 3906 40946 3912 40958
rect 4436 40860 4442 40912
rect 4494 40900 4500 40912
rect 4494 40872 5262 40900
rect 4494 40860 4500 40872
rect 6376 40836 6452 40864
rect 3428 40774 3434 40826
rect 3486 40814 3492 40826
rect 3486 40786 5358 40814
rect 3486 40774 3492 40786
rect 3848 40688 3854 40740
rect 3906 40728 3912 40740
rect 3906 40700 5454 40728
rect 3906 40688 3912 40700
rect 6168 40690 6452 40718
rect 4436 40602 4442 40654
rect 4494 40642 4500 40654
rect 4494 40614 5550 40642
rect 4494 40602 4500 40614
rect 6086 40568 6452 40596
rect 3512 40516 3518 40568
rect 3570 40556 3576 40568
rect 3570 40528 5754 40556
rect 3570 40516 3576 40528
rect 3848 40430 3854 40482
rect 3906 40470 3912 40482
rect 3906 40442 5850 40470
rect 3906 40430 3912 40442
rect 4436 40344 4442 40396
rect 4494 40384 4500 40396
rect 4494 40356 5946 40384
rect 4494 40344 4500 40356
rect 6434 39962 6440 40014
rect 6492 39962 6498 40014
rect 4436 39580 4442 39632
rect 4494 39620 4500 39632
rect 4494 39592 5946 39620
rect 4494 39580 4500 39592
rect 3848 39494 3854 39546
rect 3906 39534 3912 39546
rect 3906 39506 5850 39534
rect 3906 39494 3912 39506
rect 3260 39408 3266 39460
rect 3318 39448 3324 39460
rect 3318 39420 5754 39448
rect 3318 39408 3324 39420
rect 6086 39380 6452 39408
rect 4436 39322 4442 39374
rect 4494 39362 4500 39374
rect 4494 39334 5550 39362
rect 4494 39322 4500 39334
rect 3764 39236 3770 39288
rect 3822 39276 3828 39288
rect 3822 39248 5454 39276
rect 6168 39258 6452 39286
rect 3822 39236 3828 39248
rect 3512 39150 3518 39202
rect 3570 39190 3576 39202
rect 3570 39162 5358 39190
rect 3570 39150 3576 39162
rect 4436 39064 4442 39116
rect 4494 39104 4500 39116
rect 6376 39112 6452 39140
rect 4494 39076 5262 39104
rect 4494 39064 4500 39076
rect 3764 38978 3770 39030
rect 3822 39018 3828 39030
rect 3822 38990 5166 39018
rect 3822 38978 3828 38990
rect 3428 38892 3434 38944
rect 3486 38932 3492 38944
rect 3486 38904 5070 38932
rect 3486 38892 3492 38904
rect 6434 38424 6440 38476
rect 6492 38424 6498 38476
rect 3512 37956 3518 38008
rect 3570 37996 3576 38008
rect 3570 37968 5070 37996
rect 3570 37956 3576 37968
rect 3680 37870 3686 37922
rect 3738 37910 3744 37922
rect 3738 37882 5166 37910
rect 3738 37870 3744 37882
rect 4436 37784 4442 37836
rect 4494 37824 4500 37836
rect 4494 37796 5262 37824
rect 4494 37784 4500 37796
rect 6376 37760 6452 37788
rect 3260 37698 3266 37750
rect 3318 37738 3324 37750
rect 3318 37710 5358 37738
rect 3318 37698 3324 37710
rect 3764 37612 3770 37664
rect 3822 37652 3828 37664
rect 3822 37624 5454 37652
rect 3822 37612 3828 37624
rect 6168 37614 6452 37642
rect 4436 37526 4442 37578
rect 4494 37566 4500 37578
rect 4494 37538 5550 37566
rect 4494 37526 4500 37538
rect 6086 37492 6452 37520
rect 3344 37440 3350 37492
rect 3402 37480 3408 37492
rect 3402 37452 5754 37480
rect 3402 37440 3408 37452
rect 3764 37354 3770 37406
rect 3822 37394 3828 37406
rect 3822 37366 5850 37394
rect 3822 37354 3828 37366
rect 4436 37268 4442 37320
rect 4494 37308 4500 37320
rect 4494 37280 5946 37308
rect 4494 37268 4500 37280
rect 6434 36886 6440 36938
rect 6492 36886 6498 36938
rect 4436 36504 4442 36556
rect 4494 36544 4500 36556
rect 4494 36516 5946 36544
rect 4494 36504 4500 36516
rect 3680 36418 3686 36470
rect 3738 36458 3744 36470
rect 3738 36430 5850 36458
rect 3738 36418 3744 36430
rect 3428 36332 3434 36384
rect 3486 36372 3492 36384
rect 3486 36344 5754 36372
rect 3486 36332 3492 36344
rect 6086 36304 6452 36332
rect 3007 36198 3013 36250
rect 3065 36198 3071 36250
rect 4436 36246 4442 36298
rect 4494 36286 4500 36298
rect 4494 36258 5550 36286
rect 4494 36246 4500 36258
rect 3680 36160 3686 36212
rect 3738 36200 3744 36212
rect 3738 36172 5454 36200
rect 6168 36182 6452 36210
rect 3738 36160 3744 36172
rect 3344 36074 3350 36126
rect 3402 36114 3408 36126
rect 3402 36086 5358 36114
rect 3402 36074 3408 36086
rect 4436 35988 4442 36040
rect 4494 36028 4500 36040
rect 6376 36036 6452 36064
rect 4494 36000 5262 36028
rect 4494 35988 4500 36000
rect 3680 35902 3686 35954
rect 3738 35942 3744 35954
rect 3738 35914 5166 35942
rect 3738 35902 3744 35914
rect 3260 35816 3266 35868
rect 3318 35856 3324 35868
rect 3318 35828 5070 35856
rect 3318 35816 3324 35828
rect 6434 35348 6440 35400
rect 6492 35348 6498 35400
rect 3344 34880 3350 34932
rect 3402 34920 3408 34932
rect 3402 34892 5070 34920
rect 3402 34880 3408 34892
rect 3596 34794 3602 34846
rect 3654 34834 3660 34846
rect 3654 34806 5166 34834
rect 3654 34794 3660 34806
rect 4436 34708 4442 34760
rect 4494 34748 4500 34760
rect 4494 34720 5262 34748
rect 4494 34708 4500 34720
rect 6376 34684 6452 34712
rect 3007 34574 3013 34626
rect 3065 34574 3071 34626
rect 3428 34622 3434 34674
rect 3486 34662 3492 34674
rect 3486 34634 5358 34662
rect 3486 34622 3492 34634
rect 3596 34536 3602 34588
rect 3654 34576 3660 34588
rect 3654 34548 5454 34576
rect 3654 34536 3660 34548
rect 6168 34538 6452 34566
rect 4436 34450 4442 34502
rect 4494 34490 4500 34502
rect 4494 34462 5550 34490
rect 4494 34450 4500 34462
rect 6086 34416 6452 34444
rect 3512 34364 3518 34416
rect 3570 34404 3576 34416
rect 3570 34376 5754 34404
rect 3570 34364 3576 34376
rect 3596 34278 3602 34330
rect 3654 34318 3660 34330
rect 3654 34290 5850 34318
rect 3654 34278 3660 34290
rect 4436 34192 4442 34244
rect 4494 34232 4500 34244
rect 4494 34204 5946 34232
rect 4494 34192 4500 34204
rect 6434 33810 6440 33862
rect 6492 33810 6498 33862
rect 4436 33428 4442 33480
rect 4494 33468 4500 33480
rect 4494 33440 5946 33468
rect 4494 33428 4500 33440
rect 3596 33342 3602 33394
rect 3654 33382 3660 33394
rect 3654 33354 5850 33382
rect 3654 33342 3660 33354
rect 3260 33256 3266 33308
rect 3318 33296 3324 33308
rect 3318 33268 5754 33296
rect 3318 33256 3324 33268
rect 6086 33228 6452 33256
rect 4352 33170 4358 33222
rect 4410 33210 4416 33222
rect 4410 33182 5550 33210
rect 4410 33170 4416 33182
rect 3007 33118 3013 33170
rect 3065 33118 3071 33170
rect 4184 33084 4190 33136
rect 4242 33124 4248 33136
rect 4242 33096 5454 33124
rect 6168 33106 6452 33134
rect 4242 33084 4248 33096
rect 3512 32998 3518 33050
rect 3570 33038 3576 33050
rect 3570 33010 5358 33038
rect 3570 32998 3576 33010
rect 4352 32912 4358 32964
rect 4410 32952 4416 32964
rect 6376 32960 6452 32988
rect 4410 32924 5262 32952
rect 4410 32912 4416 32924
rect 4184 32826 4190 32878
rect 4242 32866 4248 32878
rect 4242 32838 5166 32866
rect 4242 32826 4248 32838
rect 3428 32740 3434 32792
rect 3486 32780 3492 32792
rect 3486 32752 5070 32780
rect 3486 32740 3492 32752
rect 6434 32272 6440 32324
rect 6492 32272 6498 32324
rect 3512 31804 3518 31856
rect 3570 31844 3576 31856
rect 3570 31816 5070 31844
rect 3570 31804 3576 31816
rect 4100 31718 4106 31770
rect 4158 31758 4164 31770
rect 4158 31730 5166 31758
rect 4158 31718 4164 31730
rect 4352 31632 4358 31684
rect 4410 31672 4416 31684
rect 4410 31644 5262 31672
rect 4410 31632 4416 31644
rect 6376 31608 6452 31636
rect 3260 31546 3266 31598
rect 3318 31586 3324 31598
rect 3318 31558 5358 31586
rect 3318 31546 3324 31558
rect 3007 31494 3013 31546
rect 3065 31494 3071 31546
rect 4184 31460 4190 31512
rect 4242 31500 4248 31512
rect 4242 31472 5454 31500
rect 4242 31460 4248 31472
rect 6168 31462 6452 31490
rect 4352 31374 4358 31426
rect 4410 31414 4416 31426
rect 4410 31386 5550 31414
rect 4410 31374 4416 31386
rect 6086 31340 6452 31368
rect 3344 31288 3350 31340
rect 3402 31328 3408 31340
rect 3402 31300 5754 31328
rect 3402 31288 3408 31300
rect 4184 31202 4190 31254
rect 4242 31242 4248 31254
rect 4242 31214 5850 31242
rect 4242 31202 4248 31214
rect 4352 31116 4358 31168
rect 4410 31156 4416 31168
rect 4410 31128 5946 31156
rect 4410 31116 4416 31128
rect 6434 30734 6440 30786
rect 6492 30734 6498 30786
rect 4352 30352 4358 30404
rect 4410 30392 4416 30404
rect 4410 30364 5946 30392
rect 4410 30352 4416 30364
rect 4100 30266 4106 30318
rect 4158 30306 4164 30318
rect 4158 30278 5850 30306
rect 4158 30266 4164 30278
rect 3428 30180 3434 30232
rect 3486 30220 3492 30232
rect 3486 30192 5754 30220
rect 3486 30180 3492 30192
rect 6086 30152 6452 30180
rect 4352 30094 4358 30146
rect 4410 30134 4416 30146
rect 4410 30106 5550 30134
rect 4410 30094 4416 30106
rect 3007 30038 3013 30090
rect 3065 30038 3071 30090
rect 4100 30008 4106 30060
rect 4158 30048 4164 30060
rect 4158 30020 5454 30048
rect 6168 30030 6452 30058
rect 4158 30008 4164 30020
rect 3344 29922 3350 29974
rect 3402 29962 3408 29974
rect 3402 29934 5358 29962
rect 3402 29922 3408 29934
rect 4352 29836 4358 29888
rect 4410 29876 4416 29888
rect 6376 29884 6452 29912
rect 4410 29848 5262 29876
rect 4410 29836 4416 29848
rect 4100 29750 4106 29802
rect 4158 29790 4164 29802
rect 4158 29762 5166 29790
rect 4158 29750 4164 29762
rect 3260 29664 3266 29716
rect 3318 29704 3324 29716
rect 3318 29676 5070 29704
rect 3318 29664 3324 29676
rect 6434 29196 6440 29248
rect 6492 29196 6498 29248
rect 3344 28728 3350 28780
rect 3402 28768 3408 28780
rect 3402 28740 5070 28768
rect 3402 28728 3408 28740
rect 4016 28642 4022 28694
rect 4074 28682 4080 28694
rect 4074 28654 5166 28682
rect 4074 28642 4080 28654
rect 4352 28556 4358 28608
rect 4410 28596 4416 28608
rect 4410 28568 5262 28596
rect 4410 28556 4416 28568
rect 6376 28532 6452 28560
rect 3428 28470 3434 28522
rect 3486 28510 3492 28522
rect 3486 28482 5358 28510
rect 3486 28470 3492 28482
rect 588 28414 594 28466
rect 646 28454 652 28466
rect 952 28454 958 28466
rect 646 28426 958 28454
rect 646 28414 652 28426
rect 952 28414 958 28426
rect 1010 28414 1016 28466
rect 3007 28414 3013 28466
rect 3065 28414 3071 28466
rect 4016 28384 4022 28436
rect 4074 28424 4080 28436
rect 4074 28396 5454 28424
rect 4074 28384 4080 28396
rect 6168 28386 6452 28414
rect 4352 28298 4358 28350
rect 4410 28338 4416 28350
rect 4410 28310 5550 28338
rect 4410 28298 4416 28310
rect 6086 28264 6452 28292
rect 3512 28212 3518 28264
rect 3570 28252 3576 28264
rect 3570 28224 5754 28252
rect 3570 28212 3576 28224
rect 4016 28126 4022 28178
rect 4074 28166 4080 28178
rect 4074 28138 5850 28166
rect 4074 28126 4080 28138
rect 4352 28040 4358 28092
rect 4410 28080 4416 28092
rect 4410 28052 5946 28080
rect 4410 28040 4416 28052
rect 6434 27658 6440 27710
rect 6492 27658 6498 27710
rect 4352 27276 4358 27328
rect 4410 27316 4416 27328
rect 4410 27288 5946 27316
rect 4410 27276 4416 27288
rect 4016 27190 4022 27242
rect 4074 27230 4080 27242
rect 4074 27202 5850 27230
rect 4074 27190 4080 27202
rect 3260 27104 3266 27156
rect 3318 27144 3324 27156
rect 3318 27116 5754 27144
rect 3318 27104 3324 27116
rect 6086 27076 6452 27104
rect 4352 27018 4358 27070
rect 4410 27058 4416 27070
rect 4410 27030 5550 27058
rect 4410 27018 4416 27030
rect 504 26958 510 27010
rect 562 26998 568 27010
rect 868 26998 874 27010
rect 562 26970 874 26998
rect 562 26958 568 26970
rect 868 26958 874 26970
rect 926 26958 932 27010
rect 3007 26958 3013 27010
rect 3065 26958 3071 27010
rect 3932 26932 3938 26984
rect 3990 26972 3996 26984
rect 3990 26944 5454 26972
rect 6168 26954 6452 26982
rect 3990 26932 3996 26944
rect 3512 26846 3518 26898
rect 3570 26886 3576 26898
rect 3570 26858 5358 26886
rect 3570 26846 3576 26858
rect 4352 26760 4358 26812
rect 4410 26800 4416 26812
rect 6376 26808 6452 26836
rect 4410 26772 5262 26800
rect 4410 26760 4416 26772
rect 3932 26674 3938 26726
rect 3990 26714 3996 26726
rect 3990 26686 5166 26714
rect 3990 26674 3996 26686
rect 3428 26588 3434 26640
rect 3486 26628 3492 26640
rect 3486 26600 5070 26628
rect 3486 26588 3492 26600
rect 6434 26120 6440 26172
rect 6492 26120 6498 26172
rect 3512 25652 3518 25704
rect 3570 25692 3576 25704
rect 3570 25664 5070 25692
rect 3570 25652 3576 25664
rect 3848 25566 3854 25618
rect 3906 25606 3912 25618
rect 3906 25578 5166 25606
rect 3906 25566 3912 25578
rect 4352 25480 4358 25532
rect 4410 25520 4416 25532
rect 4410 25492 5262 25520
rect 4410 25480 4416 25492
rect 6376 25456 6452 25484
rect 3260 25394 3266 25446
rect 3318 25434 3324 25446
rect 3318 25406 5358 25434
rect 3318 25394 3324 25406
rect 420 25334 426 25386
rect 478 25374 484 25386
rect 784 25374 790 25386
rect 478 25346 790 25374
rect 478 25334 484 25346
rect 784 25334 790 25346
rect 842 25334 848 25386
rect 3007 25334 3013 25386
rect 3065 25334 3071 25386
rect 3932 25308 3938 25360
rect 3990 25348 3996 25360
rect 3990 25320 5454 25348
rect 3990 25308 3996 25320
rect 6168 25310 6452 25338
rect 4352 25222 4358 25274
rect 4410 25262 4416 25274
rect 4410 25234 5550 25262
rect 4410 25222 4416 25234
rect 6086 25188 6452 25216
rect 3344 25136 3350 25188
rect 3402 25176 3408 25188
rect 3402 25148 5754 25176
rect 3402 25136 3408 25148
rect 3932 25050 3938 25102
rect 3990 25090 3996 25102
rect 3990 25062 5850 25090
rect 3990 25050 3996 25062
rect 4352 24964 4358 25016
rect 4410 25004 4416 25016
rect 4410 24976 5946 25004
rect 4410 24964 4416 24976
rect 6434 24582 6440 24634
rect 6492 24582 6498 24634
rect 4352 24200 4358 24252
rect 4410 24240 4416 24252
rect 4410 24212 5946 24240
rect 4410 24200 4416 24212
rect 3848 24114 3854 24166
rect 3906 24154 3912 24166
rect 3906 24126 5850 24154
rect 3906 24114 3912 24126
rect 3428 24028 3434 24080
rect 3486 24068 3492 24080
rect 3486 24040 5754 24068
rect 3486 24028 3492 24040
rect 6086 24000 6452 24028
rect 4352 23942 4358 23994
rect 4410 23982 4416 23994
rect 4410 23954 5550 23982
rect 4410 23942 4416 23954
rect 3848 23856 3854 23908
rect 3906 23896 3912 23908
rect 3906 23868 5454 23896
rect 6168 23878 6452 23906
rect 3906 23856 3912 23868
rect 3344 23770 3350 23822
rect 3402 23810 3408 23822
rect 3402 23782 5358 23810
rect 3402 23770 3408 23782
rect 4352 23684 4358 23736
rect 4410 23724 4416 23736
rect 6376 23732 6452 23760
rect 4410 23696 5262 23724
rect 4410 23684 4416 23696
rect 3848 23598 3854 23650
rect 3906 23638 3912 23650
rect 3906 23610 5166 23638
rect 3906 23598 3912 23610
rect 3260 23512 3266 23564
rect 3318 23552 3324 23564
rect 3318 23524 5070 23552
rect 3318 23512 3324 23524
rect 6434 23044 6440 23096
rect 6492 23044 6498 23096
rect 3344 22576 3350 22628
rect 3402 22616 3408 22628
rect 3402 22588 5070 22616
rect 3402 22576 3408 22588
rect 3764 22490 3770 22542
rect 3822 22530 3828 22542
rect 3822 22502 5166 22530
rect 3822 22490 3828 22502
rect 4352 22404 4358 22456
rect 4410 22444 4416 22456
rect 4410 22416 5262 22444
rect 4410 22404 4416 22416
rect 6376 22380 6452 22408
rect 3428 22318 3434 22370
rect 3486 22358 3492 22370
rect 3486 22330 5358 22358
rect 3486 22318 3492 22330
rect 3764 22232 3770 22284
rect 3822 22272 3828 22284
rect 3822 22244 5454 22272
rect 3822 22232 3828 22244
rect 6168 22234 6452 22262
rect 4352 22146 4358 22198
rect 4410 22186 4416 22198
rect 4410 22158 5550 22186
rect 4410 22146 4416 22158
rect 6086 22112 6452 22140
rect 3512 22060 3518 22112
rect 3570 22100 3576 22112
rect 3570 22072 5754 22100
rect 3570 22060 3576 22072
rect 3764 21974 3770 22026
rect 3822 22014 3828 22026
rect 3822 21986 5850 22014
rect 3822 21974 3828 21986
rect 4352 21888 4358 21940
rect 4410 21928 4416 21940
rect 4410 21900 5946 21928
rect 4410 21888 4416 21900
rect 6434 21506 6440 21558
rect 6492 21506 6498 21558
rect 4352 21124 4358 21176
rect 4410 21164 4416 21176
rect 4410 21136 5946 21164
rect 4410 21124 4416 21136
rect 3764 21038 3770 21090
rect 3822 21078 3828 21090
rect 3822 21050 5850 21078
rect 3822 21038 3828 21050
rect 3260 20952 3266 21004
rect 3318 20992 3324 21004
rect 3318 20964 5754 20992
rect 3318 20952 3324 20964
rect 6086 20924 6452 20952
rect 4352 20866 4358 20918
rect 4410 20906 4416 20918
rect 4410 20878 5550 20906
rect 4410 20866 4416 20878
rect 3007 20802 3013 20854
rect 3065 20802 3071 20854
rect 3680 20780 3686 20832
rect 3738 20820 3744 20832
rect 3738 20792 5454 20820
rect 6168 20802 6452 20830
rect 3738 20780 3744 20792
rect 3512 20694 3518 20746
rect 3570 20734 3576 20746
rect 3570 20706 5358 20734
rect 3570 20694 3576 20706
rect 4352 20608 4358 20660
rect 4410 20648 4416 20660
rect 6376 20656 6452 20684
rect 4410 20620 5262 20648
rect 4410 20608 4416 20620
rect 3680 20522 3686 20574
rect 3738 20562 3744 20574
rect 3738 20534 5166 20562
rect 3738 20522 3744 20534
rect 3428 20436 3434 20488
rect 3486 20476 3492 20488
rect 3486 20448 5070 20476
rect 3486 20436 3492 20448
rect 6434 19968 6440 20020
rect 6492 19968 6498 20020
rect 3512 19500 3518 19552
rect 3570 19540 3576 19552
rect 3570 19512 5070 19540
rect 3570 19500 3576 19512
rect 3596 19414 3602 19466
rect 3654 19454 3660 19466
rect 3654 19426 5166 19454
rect 3654 19414 3660 19426
rect 4352 19328 4358 19380
rect 4410 19368 4416 19380
rect 4410 19340 5262 19368
rect 4410 19328 4416 19340
rect 6376 19304 6452 19332
rect 3260 19242 3266 19294
rect 3318 19282 3324 19294
rect 3318 19254 5358 19282
rect 3318 19242 3324 19254
rect 3007 19178 3013 19230
rect 3065 19178 3071 19230
rect 3680 19156 3686 19208
rect 3738 19196 3744 19208
rect 3738 19168 5454 19196
rect 3738 19156 3744 19168
rect 6168 19158 6452 19186
rect 4352 19070 4358 19122
rect 4410 19110 4416 19122
rect 4410 19082 5550 19110
rect 4410 19070 4416 19082
rect 6086 19036 6452 19064
rect 3344 18984 3350 19036
rect 3402 19024 3408 19036
rect 3402 18996 5754 19024
rect 3402 18984 3408 18996
rect 3680 18898 3686 18950
rect 3738 18938 3744 18950
rect 3738 18910 5850 18938
rect 3738 18898 3744 18910
rect 4352 18812 4358 18864
rect 4410 18852 4416 18864
rect 4410 18824 5946 18852
rect 4410 18812 4416 18824
rect 6434 18430 6440 18482
rect 6492 18430 6498 18482
rect 4352 18048 4358 18100
rect 4410 18088 4416 18100
rect 4410 18060 5946 18088
rect 4410 18048 4416 18060
rect 3596 17962 3602 18014
rect 3654 18002 3660 18014
rect 3654 17974 5850 18002
rect 3654 17962 3660 17974
rect 3428 17876 3434 17928
rect 3486 17916 3492 17928
rect 3486 17888 5754 17916
rect 3486 17876 3492 17888
rect 6086 17848 6452 17876
rect 4352 17790 4358 17842
rect 4410 17830 4416 17842
rect 4410 17802 5550 17830
rect 4410 17790 4416 17802
rect 3007 17722 3013 17774
rect 3065 17722 3071 17774
rect 3596 17704 3602 17756
rect 3654 17744 3660 17756
rect 3654 17716 5454 17744
rect 6168 17726 6452 17754
rect 3654 17704 3660 17716
rect 3344 17618 3350 17670
rect 3402 17658 3408 17670
rect 3402 17630 5358 17658
rect 3402 17618 3408 17630
rect 4352 17532 4358 17584
rect 4410 17572 4416 17584
rect 6376 17580 6452 17608
rect 4410 17544 5262 17572
rect 4410 17532 4416 17544
rect 3596 17446 3602 17498
rect 3654 17486 3660 17498
rect 3654 17458 5166 17486
rect 3654 17446 3660 17458
rect 3260 17360 3266 17412
rect 3318 17400 3324 17412
rect 3318 17372 5070 17400
rect 3318 17360 3324 17372
rect 6434 16892 6440 16944
rect 6492 16892 6498 16944
rect 3344 16424 3350 16476
rect 3402 16464 3408 16476
rect 3402 16436 5070 16464
rect 3402 16424 3408 16436
rect 4184 16338 4190 16390
rect 4242 16378 4248 16390
rect 4242 16350 5166 16378
rect 4242 16338 4248 16350
rect 4268 16252 4274 16304
rect 4326 16292 4332 16304
rect 4326 16264 5262 16292
rect 4326 16252 4332 16264
rect 6376 16228 6452 16256
rect 3428 16166 3434 16218
rect 3486 16206 3492 16218
rect 3486 16178 5358 16206
rect 3486 16166 3492 16178
rect 3007 16098 3013 16150
rect 3065 16098 3071 16150
rect 4184 16080 4190 16132
rect 4242 16120 4248 16132
rect 4242 16092 5454 16120
rect 4242 16080 4248 16092
rect 6168 16082 6452 16110
rect 4268 15994 4274 16046
rect 4326 16034 4332 16046
rect 4326 16006 5550 16034
rect 4326 15994 4332 16006
rect 6086 15960 6452 15988
rect 3512 15908 3518 15960
rect 3570 15948 3576 15960
rect 3570 15920 5754 15948
rect 3570 15908 3576 15920
rect 4184 15822 4190 15874
rect 4242 15862 4248 15874
rect 4242 15834 5850 15862
rect 4242 15822 4248 15834
rect 4268 15736 4274 15788
rect 4326 15776 4332 15788
rect 4326 15748 5946 15776
rect 4326 15736 4332 15748
rect 6434 15354 6440 15406
rect 6492 15354 6498 15406
rect 4268 14972 4274 15024
rect 4326 15012 4332 15024
rect 4326 14984 5946 15012
rect 4326 14972 4332 14984
rect 4184 14886 4190 14938
rect 4242 14926 4248 14938
rect 4242 14898 5850 14926
rect 4242 14886 4248 14898
rect 3260 14800 3266 14852
rect 3318 14840 3324 14852
rect 3318 14812 5754 14840
rect 3318 14800 3324 14812
rect 6086 14772 6452 14800
rect 4268 14714 4274 14766
rect 4326 14754 4332 14766
rect 4326 14726 5550 14754
rect 4326 14714 4332 14726
rect 3007 14642 3013 14694
rect 3065 14642 3071 14694
rect 4100 14628 4106 14680
rect 4158 14668 4164 14680
rect 4158 14640 5454 14668
rect 6168 14650 6452 14678
rect 4158 14628 4164 14640
rect 3512 14542 3518 14594
rect 3570 14582 3576 14594
rect 3570 14554 5358 14582
rect 3570 14542 3576 14554
rect 4268 14456 4274 14508
rect 4326 14496 4332 14508
rect 6376 14504 6452 14532
rect 4326 14468 5262 14496
rect 4326 14456 4332 14468
rect 4100 14370 4106 14422
rect 4158 14410 4164 14422
rect 4158 14382 5166 14410
rect 4158 14370 4164 14382
rect 3428 14284 3434 14336
rect 3486 14324 3492 14336
rect 3486 14296 5070 14324
rect 3486 14284 3492 14296
rect 6434 13816 6440 13868
rect 6492 13816 6498 13868
rect 3512 13348 3518 13400
rect 3570 13388 3576 13400
rect 3570 13360 5070 13388
rect 3570 13348 3576 13360
rect 4016 13262 4022 13314
rect 4074 13302 4080 13314
rect 4074 13274 5166 13302
rect 4074 13262 4080 13274
rect 4268 13176 4274 13228
rect 4326 13216 4332 13228
rect 4326 13188 5262 13216
rect 4326 13176 4332 13188
rect 6376 13152 6452 13180
rect 3260 13090 3266 13142
rect 3318 13130 3324 13142
rect 3318 13102 5358 13130
rect 3318 13090 3324 13102
rect 336 13018 342 13070
rect 394 13058 400 13070
rect 952 13058 958 13070
rect 394 13030 958 13058
rect 394 13018 400 13030
rect 952 13018 958 13030
rect 1010 13018 1016 13070
rect 3007 13018 3013 13070
rect 3065 13018 3071 13070
rect 4100 13004 4106 13056
rect 4158 13044 4164 13056
rect 4158 13016 5454 13044
rect 4158 13004 4164 13016
rect 6168 13006 6452 13034
rect 4268 12918 4274 12970
rect 4326 12958 4332 12970
rect 4326 12930 5550 12958
rect 4326 12918 4332 12930
rect 6086 12884 6452 12912
rect 3344 12832 3350 12884
rect 3402 12872 3408 12884
rect 3402 12844 5754 12872
rect 3402 12832 3408 12844
rect 4100 12746 4106 12798
rect 4158 12786 4164 12798
rect 4158 12758 5850 12786
rect 4158 12746 4164 12758
rect 4268 12660 4274 12712
rect 4326 12700 4332 12712
rect 4326 12672 5946 12700
rect 4326 12660 4332 12672
rect 6434 12278 6440 12330
rect 6492 12278 6498 12330
rect 4268 11896 4274 11948
rect 4326 11936 4332 11948
rect 4326 11908 5946 11936
rect 4326 11896 4332 11908
rect 4016 11810 4022 11862
rect 4074 11850 4080 11862
rect 4074 11822 5850 11850
rect 4074 11810 4080 11822
rect 3428 11724 3434 11776
rect 3486 11764 3492 11776
rect 3486 11736 5754 11764
rect 3486 11724 3492 11736
rect 6086 11696 6452 11724
rect 4268 11638 4274 11690
rect 4326 11678 4332 11690
rect 4326 11650 5550 11678
rect 4326 11638 4332 11650
rect 252 11562 258 11614
rect 310 11602 316 11614
rect 868 11602 874 11614
rect 310 11574 874 11602
rect 310 11562 316 11574
rect 868 11562 874 11574
rect 926 11562 932 11614
rect 3007 11562 3013 11614
rect 3065 11562 3071 11614
rect 4016 11552 4022 11604
rect 4074 11592 4080 11604
rect 4074 11564 5454 11592
rect 6168 11574 6452 11602
rect 4074 11552 4080 11564
rect 3344 11466 3350 11518
rect 3402 11506 3408 11518
rect 3402 11478 5358 11506
rect 3402 11466 3408 11478
rect 4268 11380 4274 11432
rect 4326 11420 4332 11432
rect 6376 11428 6452 11456
rect 4326 11392 5262 11420
rect 4326 11380 4332 11392
rect 4016 11294 4022 11346
rect 4074 11334 4080 11346
rect 4074 11306 5166 11334
rect 4074 11294 4080 11306
rect 3260 11208 3266 11260
rect 3318 11248 3324 11260
rect 3318 11220 5070 11248
rect 3318 11208 3324 11220
rect 6434 10740 6440 10792
rect 6492 10740 6498 10792
rect 3344 10272 3350 10324
rect 3402 10312 3408 10324
rect 3402 10284 5070 10312
rect 3402 10272 3408 10284
rect 3932 10186 3938 10238
rect 3990 10226 3996 10238
rect 3990 10198 5166 10226
rect 3990 10186 3996 10198
rect 4268 10100 4274 10152
rect 4326 10140 4332 10152
rect 4326 10112 5262 10140
rect 4326 10100 4332 10112
rect 6376 10076 6452 10104
rect 3428 10014 3434 10066
rect 3486 10054 3492 10066
rect 3486 10026 5358 10054
rect 3486 10014 3492 10026
rect 168 9938 174 9990
rect 226 9978 232 9990
rect 784 9978 790 9990
rect 226 9950 790 9978
rect 226 9938 232 9950
rect 784 9938 790 9950
rect 842 9938 848 9990
rect 3007 9938 3013 9990
rect 3065 9938 3071 9990
rect 3932 9928 3938 9980
rect 3990 9968 3996 9980
rect 3990 9940 5454 9968
rect 3990 9928 3996 9940
rect 6168 9930 6452 9958
rect 4268 9842 4274 9894
rect 4326 9882 4332 9894
rect 4326 9854 5550 9882
rect 4326 9842 4332 9854
rect 6086 9808 6452 9836
rect 3512 9756 3518 9808
rect 3570 9796 3576 9808
rect 3570 9768 5754 9796
rect 3570 9756 3576 9768
rect 3932 9670 3938 9722
rect 3990 9710 3996 9722
rect 3990 9682 5850 9710
rect 3990 9670 3996 9682
rect 4268 9584 4274 9636
rect 4326 9624 4332 9636
rect 4326 9596 5946 9624
rect 4326 9584 4332 9596
rect 6434 9202 6440 9254
rect 6492 9202 6498 9254
rect 4268 8820 4274 8872
rect 4326 8860 4332 8872
rect 4326 8832 5946 8860
rect 4326 8820 4332 8832
rect 3932 8734 3938 8786
rect 3990 8774 3996 8786
rect 3990 8746 5850 8774
rect 3990 8734 3996 8746
rect 3260 8648 3266 8700
rect 3318 8688 3324 8700
rect 3318 8660 5754 8688
rect 3318 8648 3324 8660
rect 6086 8620 6452 8648
rect 4268 8562 4274 8614
rect 4326 8602 4332 8614
rect 4326 8574 5550 8602
rect 4326 8562 4332 8574
rect 3848 8476 3854 8528
rect 3906 8516 3912 8528
rect 3906 8488 5454 8516
rect 6168 8498 6452 8526
rect 3906 8476 3912 8488
rect 3512 8390 3518 8442
rect 3570 8430 3576 8442
rect 3570 8402 5358 8430
rect 3570 8390 3576 8402
rect 4268 8304 4274 8356
rect 4326 8344 4332 8356
rect 6376 8352 6452 8380
rect 4326 8316 5262 8344
rect 4326 8304 4332 8316
rect 3848 8218 3854 8270
rect 3906 8258 3912 8270
rect 3906 8230 5166 8258
rect 3906 8218 3912 8230
rect 3428 8132 3434 8184
rect 3486 8172 3492 8184
rect 3486 8144 5070 8172
rect 3486 8132 3492 8144
rect 6434 7664 6440 7716
rect 6492 7664 6498 7716
rect 3512 7196 3518 7248
rect 3570 7236 3576 7248
rect 3570 7208 5070 7236
rect 3570 7196 3576 7208
rect 3764 7110 3770 7162
rect 3822 7150 3828 7162
rect 3822 7122 5166 7150
rect 3822 7110 3828 7122
rect 4268 7024 4274 7076
rect 4326 7064 4332 7076
rect 4326 7036 5262 7064
rect 4326 7024 4332 7036
rect 6376 7000 6452 7028
rect 3260 6938 3266 6990
rect 3318 6978 3324 6990
rect 3318 6950 5358 6978
rect 3318 6938 3324 6950
rect 3848 6852 3854 6904
rect 3906 6892 3912 6904
rect 3906 6864 5454 6892
rect 3906 6852 3912 6864
rect 6168 6854 6452 6882
rect 4268 6766 4274 6818
rect 4326 6806 4332 6818
rect 4326 6778 5550 6806
rect 4326 6766 4332 6778
rect 6086 6732 6452 6760
rect 3344 6680 3350 6732
rect 3402 6720 3408 6732
rect 3402 6692 5754 6720
rect 3402 6680 3408 6692
rect 3848 6594 3854 6646
rect 3906 6634 3912 6646
rect 3906 6606 5850 6634
rect 3906 6594 3912 6606
rect 4268 6508 4274 6560
rect 4326 6548 4332 6560
rect 4326 6520 5946 6548
rect 4326 6508 4332 6520
rect 6434 6126 6440 6178
rect 6492 6126 6498 6178
rect 4268 5744 4274 5796
rect 4326 5784 4332 5796
rect 4326 5756 5946 5784
rect 4326 5744 4332 5756
rect 3764 5658 3770 5710
rect 3822 5698 3828 5710
rect 3822 5670 5850 5698
rect 3822 5658 3828 5670
rect 3428 5572 3434 5624
rect 3486 5612 3492 5624
rect 3486 5584 5754 5612
rect 3486 5572 3492 5584
rect 6086 5544 6452 5572
rect 4268 5486 4274 5538
rect 4326 5526 4332 5538
rect 4326 5498 5550 5526
rect 4326 5486 4332 5498
rect 3007 5406 3013 5458
rect 3065 5406 3071 5458
rect 3764 5400 3770 5452
rect 3822 5440 3828 5452
rect 3822 5412 5454 5440
rect 6168 5422 6452 5450
rect 3822 5400 3828 5412
rect 3344 5314 3350 5366
rect 3402 5354 3408 5366
rect 3402 5326 5358 5354
rect 3402 5314 3408 5326
rect 4268 5228 4274 5280
rect 4326 5268 4332 5280
rect 6376 5276 6452 5304
rect 4326 5240 5262 5268
rect 4326 5228 4332 5240
rect 3764 5142 3770 5194
rect 3822 5182 3828 5194
rect 3822 5154 5166 5182
rect 3822 5142 3828 5154
rect 3260 5056 3266 5108
rect 3318 5096 3324 5108
rect 3318 5068 5070 5096
rect 3318 5056 3324 5068
rect 6434 4588 6440 4640
rect 6492 4588 6498 4640
rect 3344 4120 3350 4172
rect 3402 4160 3408 4172
rect 3402 4132 5070 4160
rect 3402 4120 3408 4132
rect 3680 4034 3686 4086
rect 3738 4074 3744 4086
rect 3738 4046 5166 4074
rect 3738 4034 3744 4046
rect 4268 3948 4274 4000
rect 4326 3988 4332 4000
rect 4326 3960 5262 3988
rect 4326 3948 4332 3960
rect 6376 3924 6452 3952
rect 3428 3862 3434 3914
rect 3486 3902 3492 3914
rect 3486 3874 5358 3902
rect 3486 3862 3492 3874
rect 3007 3782 3013 3834
rect 3065 3782 3071 3834
rect 3680 3776 3686 3828
rect 3738 3816 3744 3828
rect 3738 3788 5454 3816
rect 3738 3776 3744 3788
rect 6168 3778 6452 3806
rect 4268 3690 4274 3742
rect 4326 3730 4332 3742
rect 4326 3702 5550 3730
rect 4326 3690 4332 3702
rect 6086 3656 6452 3684
rect 3512 3604 3518 3656
rect 3570 3644 3576 3656
rect 3570 3616 5754 3644
rect 3570 3604 3576 3616
rect 3680 3518 3686 3570
rect 3738 3558 3744 3570
rect 3738 3530 5850 3558
rect 3738 3518 3744 3530
rect 4268 3432 4274 3484
rect 4326 3472 4332 3484
rect 4326 3444 5946 3472
rect 4326 3432 4332 3444
rect 6434 3050 6440 3102
rect 6492 3050 6498 3102
rect 4268 2668 4274 2720
rect 4326 2708 4332 2720
rect 4326 2680 5946 2708
rect 4326 2668 4332 2680
rect 3680 2582 3686 2634
rect 3738 2622 3744 2634
rect 3738 2594 5850 2622
rect 3738 2582 3744 2594
rect 3260 2496 3266 2548
rect 3318 2536 3324 2548
rect 3318 2508 5754 2536
rect 3318 2496 3324 2508
rect 6086 2468 6452 2496
rect 4268 2410 4274 2462
rect 4326 2450 4332 2462
rect 4326 2422 5550 2450
rect 4326 2410 4332 2422
rect 84 2326 90 2378
rect 142 2366 148 2378
rect 1300 2366 1306 2378
rect 142 2338 1306 2366
rect 142 2326 148 2338
rect 1300 2326 1306 2338
rect 1358 2326 1364 2378
rect 3007 2326 3013 2378
rect 3065 2326 3071 2378
rect 3596 2324 3602 2376
rect 3654 2364 3660 2376
rect 3654 2336 5454 2364
rect 6168 2346 6452 2374
rect 3654 2324 3660 2336
rect 3512 2238 3518 2290
rect 3570 2278 3576 2290
rect 3570 2250 5358 2278
rect 3570 2238 3576 2250
rect 4268 2152 4274 2204
rect 4326 2192 4332 2204
rect 6376 2200 6452 2228
rect 4326 2164 5262 2192
rect 4326 2152 4332 2164
rect 3596 2066 3602 2118
rect 3654 2106 3660 2118
rect 3654 2078 5166 2106
rect 3654 2066 3660 2078
rect 3428 1980 3434 2032
rect 3486 2020 3492 2032
rect 3486 1992 5070 2020
rect 3486 1980 3492 1992
rect 6434 1512 6440 1564
rect 6492 1512 6498 1564
rect 6376 848 6452 876
rect 3260 786 3266 838
rect 3318 826 3324 838
rect 3318 798 5358 826
rect 3318 786 3324 798
rect 0 702 6 754
rect 58 742 64 754
rect 1216 742 1222 754
rect 58 714 1222 742
rect 58 702 64 714
rect 1216 702 1222 714
rect 1274 702 1280 754
rect 3007 702 3013 754
rect 3065 702 3071 754
rect 3596 700 3602 752
rect 3654 740 3660 752
rect 3654 712 5454 740
rect 3654 700 3660 712
rect 6168 702 6452 730
rect 4268 614 4274 666
rect 4326 654 4332 666
rect 4326 626 5550 654
rect 4326 614 4332 626
rect 6086 580 6452 608
rect 3344 528 3350 580
rect 3402 568 3408 580
rect 3402 540 5754 568
rect 3402 528 3408 540
rect 3596 442 3602 494
rect 3654 482 3660 494
rect 3654 454 5850 482
rect 3654 442 3660 454
rect 4268 356 4274 408
rect 4326 396 4332 408
rect 4326 368 5946 396
rect 4326 356 4332 368
rect 6434 -26 6440 26
rect 6492 -26 6498 26
<< via1 >>
rect 6440 98406 6492 98458
rect 4694 98024 4746 98076
rect 4190 97938 4242 97990
rect 3434 97852 3486 97904
rect 4694 97766 4746 97818
rect 4190 97680 4242 97732
rect 3350 97594 3402 97646
rect 4694 97508 4746 97560
rect 4190 97422 4242 97474
rect 3266 97336 3318 97388
rect 6440 96868 6492 96920
rect 3350 96400 3402 96452
rect 4106 96314 4158 96366
rect 4694 96228 4746 96280
rect 3434 96142 3486 96194
rect 4106 96056 4158 96108
rect 4694 95970 4746 96022
rect 3518 95884 3570 95936
rect 4106 95798 4158 95850
rect 4694 95712 4746 95764
rect 6440 95330 6492 95382
rect 4694 94948 4746 95000
rect 4106 94862 4158 94914
rect 3266 94776 3318 94828
rect 4694 94690 4746 94742
rect 4022 94604 4074 94656
rect 3518 94518 3570 94570
rect 4694 94432 4746 94484
rect 4022 94346 4074 94398
rect 3434 94260 3486 94312
rect 6440 93792 6492 93844
rect 3518 93324 3570 93376
rect 3938 93238 3990 93290
rect 4694 93152 4746 93204
rect 3266 93066 3318 93118
rect 4022 92980 4074 93032
rect 4694 92894 4746 92946
rect 3350 92808 3402 92860
rect 4022 92722 4074 92774
rect 4694 92636 4746 92688
rect 6440 92254 6492 92306
rect 4694 91872 4746 91924
rect 3938 91786 3990 91838
rect 3434 91700 3486 91752
rect 4694 91614 4746 91666
rect 3938 91528 3990 91580
rect 3350 91442 3402 91494
rect 4694 91356 4746 91408
rect 3938 91270 3990 91322
rect 3266 91184 3318 91236
rect 6440 90716 6492 90768
rect 3350 90248 3402 90300
rect 3854 90162 3906 90214
rect 4694 90076 4746 90128
rect 3434 89990 3486 90042
rect 3854 89904 3906 89956
rect 4694 89818 4746 89870
rect 3518 89732 3570 89784
rect 3854 89646 3906 89698
rect 4694 89560 4746 89612
rect 6440 89178 6492 89230
rect 4694 88796 4746 88848
rect 3854 88710 3906 88762
rect 3266 88624 3318 88676
rect 4694 88538 4746 88590
rect 3770 88452 3822 88504
rect 3518 88366 3570 88418
rect 4694 88280 4746 88332
rect 3770 88194 3822 88246
rect 3434 88108 3486 88160
rect 6440 87640 6492 87692
rect 3518 87172 3570 87224
rect 3686 87086 3738 87138
rect 4694 87000 4746 87052
rect 3266 86914 3318 86966
rect 3770 86828 3822 86880
rect 4694 86742 4746 86794
rect 3350 86656 3402 86708
rect 3770 86570 3822 86622
rect 4694 86484 4746 86536
rect 6440 86102 6492 86154
rect 4694 85720 4746 85772
rect 3686 85634 3738 85686
rect 3434 85548 3486 85600
rect 4694 85462 4746 85514
rect 3686 85376 3738 85428
rect 3350 85290 3402 85342
rect 4694 85204 4746 85256
rect 3686 85118 3738 85170
rect 3266 85032 3318 85084
rect 6440 84564 6492 84616
rect 3350 84096 3402 84148
rect 3602 84010 3654 84062
rect 4694 83924 4746 83976
rect 3434 83838 3486 83890
rect 3602 83752 3654 83804
rect 4694 83666 4746 83718
rect 3518 83580 3570 83632
rect 3602 83494 3654 83546
rect 4694 83408 4746 83460
rect 6440 83026 6492 83078
rect 4694 82644 4746 82696
rect 3602 82558 3654 82610
rect 3266 82472 3318 82524
rect 4610 82386 4662 82438
rect 4190 82300 4242 82352
rect 3518 82214 3570 82266
rect 4610 82128 4662 82180
rect 4190 82042 4242 82094
rect 3434 81956 3486 82008
rect 6440 81488 6492 81540
rect 3518 81020 3570 81072
rect 4106 80934 4158 80986
rect 4610 80848 4662 80900
rect 3266 80762 3318 80814
rect 4190 80676 4242 80728
rect 4610 80590 4662 80642
rect 3350 80504 3402 80556
rect 4190 80418 4242 80470
rect 4610 80332 4662 80384
rect 6440 79950 6492 80002
rect 4610 79568 4662 79620
rect 4106 79482 4158 79534
rect 3434 79396 3486 79448
rect 4610 79310 4662 79362
rect 4106 79224 4158 79276
rect 3350 79138 3402 79190
rect 4610 79052 4662 79104
rect 4106 78966 4158 79018
rect 3266 78880 3318 78932
rect 6440 78412 6492 78464
rect 3350 77944 3402 77996
rect 4022 77858 4074 77910
rect 4610 77772 4662 77824
rect 3434 77686 3486 77738
rect 4022 77600 4074 77652
rect 4610 77514 4662 77566
rect 3518 77428 3570 77480
rect 4022 77342 4074 77394
rect 4610 77256 4662 77308
rect 6440 76874 6492 76926
rect 4610 76492 4662 76544
rect 4022 76406 4074 76458
rect 3266 76320 3318 76372
rect 4610 76234 4662 76286
rect 3938 76148 3990 76200
rect 3518 76062 3570 76114
rect 4610 75976 4662 76028
rect 3938 75890 3990 75942
rect 3434 75804 3486 75856
rect 6440 75336 6492 75388
rect 3518 74868 3570 74920
rect 3854 74782 3906 74834
rect 4610 74696 4662 74748
rect 3266 74610 3318 74662
rect 3938 74524 3990 74576
rect 4610 74438 4662 74490
rect 3350 74352 3402 74404
rect 3938 74266 3990 74318
rect 4610 74180 4662 74232
rect 6440 73798 6492 73850
rect 4610 73416 4662 73468
rect 3854 73330 3906 73382
rect 3434 73244 3486 73296
rect 4610 73158 4662 73210
rect 3854 73072 3906 73124
rect 3350 72986 3402 73038
rect 4610 72900 4662 72952
rect 3854 72814 3906 72866
rect 3266 72728 3318 72780
rect 6440 72260 6492 72312
rect 3350 71792 3402 71844
rect 3770 71706 3822 71758
rect 4610 71620 4662 71672
rect 3434 71534 3486 71586
rect 3770 71448 3822 71500
rect 4610 71362 4662 71414
rect 3518 71276 3570 71328
rect 3770 71190 3822 71242
rect 4610 71104 4662 71156
rect 6440 70722 6492 70774
rect 4610 70340 4662 70392
rect 3770 70254 3822 70306
rect 3266 70168 3318 70220
rect 4610 70082 4662 70134
rect 3686 69996 3738 70048
rect 3518 69910 3570 69962
rect 4610 69824 4662 69876
rect 3686 69738 3738 69790
rect 3434 69652 3486 69704
rect 6440 69184 6492 69236
rect 3518 68716 3570 68768
rect 3602 68630 3654 68682
rect 4610 68544 4662 68596
rect 3266 68458 3318 68510
rect 3686 68372 3738 68424
rect 4610 68286 4662 68338
rect 3350 68200 3402 68252
rect 3686 68114 3738 68166
rect 4610 68028 4662 68080
rect 6440 67646 6492 67698
rect 4610 67264 4662 67316
rect 3602 67178 3654 67230
rect 3434 67092 3486 67144
rect 4610 67006 4662 67058
rect 3602 66920 3654 66972
rect 3350 66834 3402 66886
rect 4610 66748 4662 66800
rect 3602 66662 3654 66714
rect 3266 66576 3318 66628
rect 6440 66108 6492 66160
rect 3350 65640 3402 65692
rect 4190 65554 4242 65606
rect 4526 65468 4578 65520
rect 3434 65382 3486 65434
rect 4190 65296 4242 65348
rect 4526 65210 4578 65262
rect 3518 65124 3570 65176
rect 4190 65038 4242 65090
rect 4526 64952 4578 65004
rect 6440 64570 6492 64622
rect 4526 64188 4578 64240
rect 4190 64102 4242 64154
rect 3266 64016 3318 64068
rect 4526 63930 4578 63982
rect 4106 63844 4158 63896
rect 3518 63758 3570 63810
rect 4526 63672 4578 63724
rect 4106 63586 4158 63638
rect 3434 63500 3486 63552
rect 6440 63032 6492 63084
rect 3518 62564 3570 62616
rect 4022 62478 4074 62530
rect 4526 62392 4578 62444
rect 3266 62306 3318 62358
rect 4106 62220 4158 62272
rect 4526 62134 4578 62186
rect 3350 62048 3402 62100
rect 4106 61962 4158 62014
rect 4526 61876 4578 61928
rect 6440 61494 6492 61546
rect 4526 61112 4578 61164
rect 4022 61026 4074 61078
rect 3434 60940 3486 60992
rect 4526 60854 4578 60906
rect 4022 60768 4074 60820
rect 3350 60682 3402 60734
rect 4526 60596 4578 60648
rect 4022 60510 4074 60562
rect 3266 60424 3318 60476
rect 6440 59956 6492 60008
rect 3350 59488 3402 59540
rect 3938 59402 3990 59454
rect 4526 59316 4578 59368
rect 3434 59230 3486 59282
rect 3938 59144 3990 59196
rect 4526 59058 4578 59110
rect 3518 58972 3570 59024
rect 3938 58886 3990 58938
rect 4526 58800 4578 58852
rect 6440 58418 6492 58470
rect 4526 58036 4578 58088
rect 3938 57950 3990 58002
rect 3266 57864 3318 57916
rect 4526 57778 4578 57830
rect 3854 57692 3906 57744
rect 3518 57606 3570 57658
rect 4526 57520 4578 57572
rect 3854 57434 3906 57486
rect 3434 57348 3486 57400
rect 6440 56880 6492 56932
rect 3518 56412 3570 56464
rect 3770 56326 3822 56378
rect 4526 56240 4578 56292
rect 3266 56154 3318 56206
rect 3854 56068 3906 56120
rect 4526 55982 4578 56034
rect 3350 55896 3402 55948
rect 3854 55810 3906 55862
rect 4526 55724 4578 55776
rect 6440 55342 6492 55394
rect 4526 54960 4578 55012
rect 3770 54874 3822 54926
rect 3434 54788 3486 54840
rect 4526 54702 4578 54754
rect 3770 54616 3822 54668
rect 3350 54530 3402 54582
rect 4526 54444 4578 54496
rect 3770 54358 3822 54410
rect 3266 54272 3318 54324
rect 6440 53804 6492 53856
rect 3350 53336 3402 53388
rect 3686 53250 3738 53302
rect 4526 53164 4578 53216
rect 3434 53078 3486 53130
rect 3686 52992 3738 53044
rect 4526 52906 4578 52958
rect 3518 52820 3570 52872
rect 3686 52734 3738 52786
rect 4526 52648 4578 52700
rect 6440 52266 6492 52318
rect 4526 51884 4578 51936
rect 3686 51798 3738 51850
rect 3266 51712 3318 51764
rect 4526 51626 4578 51678
rect 3602 51540 3654 51592
rect 3518 51454 3570 51506
rect 4526 51368 4578 51420
rect 3602 51282 3654 51334
rect 3434 51196 3486 51248
rect 6440 50728 6492 50780
rect 3518 50260 3570 50312
rect 4190 50174 4242 50226
rect 4442 50088 4494 50140
rect 3266 50002 3318 50054
rect 3602 49916 3654 49968
rect 4526 49830 4578 49882
rect 3350 49744 3402 49796
rect 3602 49658 3654 49710
rect 4526 49572 4578 49624
rect 6440 49190 6492 49242
rect 4442 48808 4494 48860
rect 4190 48722 4242 48774
rect 3434 48636 3486 48688
rect 4442 48550 4494 48602
rect 4190 48464 4242 48516
rect 3350 48378 3402 48430
rect 4442 48292 4494 48344
rect 4190 48206 4242 48258
rect 3266 48120 3318 48172
rect 6440 47652 6492 47704
rect 3350 47184 3402 47236
rect 4106 47098 4158 47150
rect 4442 47012 4494 47064
rect 3434 46926 3486 46978
rect 4106 46840 4158 46892
rect 4442 46754 4494 46806
rect 3518 46668 3570 46720
rect 4106 46582 4158 46634
rect 4442 46496 4494 46548
rect 6440 46114 6492 46166
rect 4442 45732 4494 45784
rect 4106 45646 4158 45698
rect 3266 45560 3318 45612
rect 4442 45474 4494 45526
rect 4022 45388 4074 45440
rect 3518 45302 3570 45354
rect 4442 45216 4494 45268
rect 4022 45130 4074 45182
rect 3434 45044 3486 45096
rect 6440 44576 6492 44628
rect 3518 44108 3570 44160
rect 3938 44022 3990 44074
rect 4442 43936 4494 43988
rect 3266 43850 3318 43902
rect 4022 43764 4074 43816
rect 4442 43678 4494 43730
rect 3350 43592 3402 43644
rect 4022 43506 4074 43558
rect 4442 43420 4494 43472
rect 6440 43038 6492 43090
rect 4442 42656 4494 42708
rect 3938 42570 3990 42622
rect 3434 42484 3486 42536
rect 4442 42398 4494 42450
rect 3938 42312 3990 42364
rect 3350 42226 3402 42278
rect 4442 42140 4494 42192
rect 3938 42054 3990 42106
rect 3266 41968 3318 42020
rect 6440 41500 6492 41552
rect 3350 41032 3402 41084
rect 3854 40946 3906 40998
rect 4442 40860 4494 40912
rect 3434 40774 3486 40826
rect 3854 40688 3906 40740
rect 4442 40602 4494 40654
rect 3518 40516 3570 40568
rect 3854 40430 3906 40482
rect 4442 40344 4494 40396
rect 6440 39962 6492 40014
rect 4442 39580 4494 39632
rect 3854 39494 3906 39546
rect 3266 39408 3318 39460
rect 4442 39322 4494 39374
rect 3770 39236 3822 39288
rect 3518 39150 3570 39202
rect 4442 39064 4494 39116
rect 3770 38978 3822 39030
rect 3434 38892 3486 38944
rect 6440 38424 6492 38476
rect 3518 37956 3570 38008
rect 3686 37870 3738 37922
rect 4442 37784 4494 37836
rect 3266 37698 3318 37750
rect 3770 37612 3822 37664
rect 4442 37526 4494 37578
rect 3350 37440 3402 37492
rect 3770 37354 3822 37406
rect 4442 37268 4494 37320
rect 6440 36886 6492 36938
rect 4442 36504 4494 36556
rect 3686 36418 3738 36470
rect 3434 36332 3486 36384
rect 3013 36241 3065 36250
rect 3013 36207 3022 36241
rect 3022 36207 3056 36241
rect 3056 36207 3065 36241
rect 3013 36198 3065 36207
rect 4442 36246 4494 36298
rect 3686 36160 3738 36212
rect 3350 36074 3402 36126
rect 4442 35988 4494 36040
rect 3686 35902 3738 35954
rect 3266 35816 3318 35868
rect 6440 35348 6492 35400
rect 3350 34880 3402 34932
rect 3602 34794 3654 34846
rect 4442 34708 4494 34760
rect 3013 34617 3065 34626
rect 3013 34583 3022 34617
rect 3022 34583 3056 34617
rect 3056 34583 3065 34617
rect 3013 34574 3065 34583
rect 3434 34622 3486 34674
rect 3602 34536 3654 34588
rect 4442 34450 4494 34502
rect 3518 34364 3570 34416
rect 3602 34278 3654 34330
rect 4442 34192 4494 34244
rect 6440 33810 6492 33862
rect 4442 33428 4494 33480
rect 3602 33342 3654 33394
rect 3266 33256 3318 33308
rect 4358 33170 4410 33222
rect 3013 33161 3065 33170
rect 3013 33127 3022 33161
rect 3022 33127 3056 33161
rect 3056 33127 3065 33161
rect 3013 33118 3065 33127
rect 4190 33084 4242 33136
rect 3518 32998 3570 33050
rect 4358 32912 4410 32964
rect 4190 32826 4242 32878
rect 3434 32740 3486 32792
rect 6440 32272 6492 32324
rect 3518 31804 3570 31856
rect 4106 31718 4158 31770
rect 4358 31632 4410 31684
rect 3266 31546 3318 31598
rect 3013 31537 3065 31546
rect 3013 31503 3022 31537
rect 3022 31503 3056 31537
rect 3056 31503 3065 31537
rect 3013 31494 3065 31503
rect 4190 31460 4242 31512
rect 4358 31374 4410 31426
rect 3350 31288 3402 31340
rect 4190 31202 4242 31254
rect 4358 31116 4410 31168
rect 6440 30734 6492 30786
rect 4358 30352 4410 30404
rect 4106 30266 4158 30318
rect 3434 30180 3486 30232
rect 4358 30094 4410 30146
rect 3013 30081 3065 30090
rect 3013 30047 3022 30081
rect 3022 30047 3056 30081
rect 3056 30047 3065 30081
rect 3013 30038 3065 30047
rect 4106 30008 4158 30060
rect 3350 29922 3402 29974
rect 4358 29836 4410 29888
rect 4106 29750 4158 29802
rect 3266 29664 3318 29716
rect 6440 29196 6492 29248
rect 3350 28728 3402 28780
rect 4022 28642 4074 28694
rect 4358 28556 4410 28608
rect 3434 28470 3486 28522
rect 594 28414 646 28466
rect 958 28414 1010 28466
rect 3013 28457 3065 28466
rect 3013 28423 3022 28457
rect 3022 28423 3056 28457
rect 3056 28423 3065 28457
rect 3013 28414 3065 28423
rect 4022 28384 4074 28436
rect 4358 28298 4410 28350
rect 3518 28212 3570 28264
rect 4022 28126 4074 28178
rect 4358 28040 4410 28092
rect 6440 27658 6492 27710
rect 4358 27276 4410 27328
rect 4022 27190 4074 27242
rect 3266 27104 3318 27156
rect 4358 27018 4410 27070
rect 510 26958 562 27010
rect 874 26958 926 27010
rect 3013 27001 3065 27010
rect 3013 26967 3022 27001
rect 3022 26967 3056 27001
rect 3056 26967 3065 27001
rect 3013 26958 3065 26967
rect 3938 26932 3990 26984
rect 3518 26846 3570 26898
rect 4358 26760 4410 26812
rect 3938 26674 3990 26726
rect 3434 26588 3486 26640
rect 6440 26120 6492 26172
rect 3518 25652 3570 25704
rect 3854 25566 3906 25618
rect 4358 25480 4410 25532
rect 3266 25394 3318 25446
rect 426 25334 478 25386
rect 790 25334 842 25386
rect 3013 25377 3065 25386
rect 3013 25343 3022 25377
rect 3022 25343 3056 25377
rect 3056 25343 3065 25377
rect 3013 25334 3065 25343
rect 3938 25308 3990 25360
rect 4358 25222 4410 25274
rect 3350 25136 3402 25188
rect 3938 25050 3990 25102
rect 4358 24964 4410 25016
rect 6440 24582 6492 24634
rect 4358 24200 4410 24252
rect 3854 24114 3906 24166
rect 3434 24028 3486 24080
rect 4358 23942 4410 23994
rect 3854 23856 3906 23908
rect 3350 23770 3402 23822
rect 4358 23684 4410 23736
rect 3854 23598 3906 23650
rect 3266 23512 3318 23564
rect 6440 23044 6492 23096
rect 3350 22576 3402 22628
rect 3770 22490 3822 22542
rect 4358 22404 4410 22456
rect 3434 22318 3486 22370
rect 3770 22232 3822 22284
rect 4358 22146 4410 22198
rect 3518 22060 3570 22112
rect 3770 21974 3822 22026
rect 4358 21888 4410 21940
rect 6440 21506 6492 21558
rect 4358 21124 4410 21176
rect 3770 21038 3822 21090
rect 3266 20952 3318 21004
rect 4358 20866 4410 20918
rect 3013 20845 3065 20854
rect 3013 20811 3022 20845
rect 3022 20811 3056 20845
rect 3056 20811 3065 20845
rect 3013 20802 3065 20811
rect 3686 20780 3738 20832
rect 3518 20694 3570 20746
rect 4358 20608 4410 20660
rect 3686 20522 3738 20574
rect 3434 20436 3486 20488
rect 6440 19968 6492 20020
rect 3518 19500 3570 19552
rect 3602 19414 3654 19466
rect 4358 19328 4410 19380
rect 3266 19242 3318 19294
rect 3013 19221 3065 19230
rect 3013 19187 3022 19221
rect 3022 19187 3056 19221
rect 3056 19187 3065 19221
rect 3013 19178 3065 19187
rect 3686 19156 3738 19208
rect 4358 19070 4410 19122
rect 3350 18984 3402 19036
rect 3686 18898 3738 18950
rect 4358 18812 4410 18864
rect 6440 18430 6492 18482
rect 4358 18048 4410 18100
rect 3602 17962 3654 18014
rect 3434 17876 3486 17928
rect 4358 17790 4410 17842
rect 3013 17765 3065 17774
rect 3013 17731 3022 17765
rect 3022 17731 3056 17765
rect 3056 17731 3065 17765
rect 3013 17722 3065 17731
rect 3602 17704 3654 17756
rect 3350 17618 3402 17670
rect 4358 17532 4410 17584
rect 3602 17446 3654 17498
rect 3266 17360 3318 17412
rect 6440 16892 6492 16944
rect 3350 16424 3402 16476
rect 4190 16338 4242 16390
rect 4274 16252 4326 16304
rect 3434 16166 3486 16218
rect 3013 16141 3065 16150
rect 3013 16107 3022 16141
rect 3022 16107 3056 16141
rect 3056 16107 3065 16141
rect 3013 16098 3065 16107
rect 4190 16080 4242 16132
rect 4274 15994 4326 16046
rect 3518 15908 3570 15960
rect 4190 15822 4242 15874
rect 4274 15736 4326 15788
rect 6440 15354 6492 15406
rect 4274 14972 4326 15024
rect 4190 14886 4242 14938
rect 3266 14800 3318 14852
rect 4274 14714 4326 14766
rect 3013 14685 3065 14694
rect 3013 14651 3022 14685
rect 3022 14651 3056 14685
rect 3056 14651 3065 14685
rect 3013 14642 3065 14651
rect 4106 14628 4158 14680
rect 3518 14542 3570 14594
rect 4274 14456 4326 14508
rect 4106 14370 4158 14422
rect 3434 14284 3486 14336
rect 6440 13816 6492 13868
rect 3518 13348 3570 13400
rect 4022 13262 4074 13314
rect 4274 13176 4326 13228
rect 3266 13090 3318 13142
rect 342 13018 394 13070
rect 958 13018 1010 13070
rect 3013 13061 3065 13070
rect 3013 13027 3022 13061
rect 3022 13027 3056 13061
rect 3056 13027 3065 13061
rect 3013 13018 3065 13027
rect 4106 13004 4158 13056
rect 4274 12918 4326 12970
rect 3350 12832 3402 12884
rect 4106 12746 4158 12798
rect 4274 12660 4326 12712
rect 6440 12278 6492 12330
rect 4274 11896 4326 11948
rect 4022 11810 4074 11862
rect 3434 11724 3486 11776
rect 4274 11638 4326 11690
rect 258 11562 310 11614
rect 874 11562 926 11614
rect 3013 11605 3065 11614
rect 3013 11571 3022 11605
rect 3022 11571 3056 11605
rect 3056 11571 3065 11605
rect 3013 11562 3065 11571
rect 4022 11552 4074 11604
rect 3350 11466 3402 11518
rect 4274 11380 4326 11432
rect 4022 11294 4074 11346
rect 3266 11208 3318 11260
rect 6440 10740 6492 10792
rect 3350 10272 3402 10324
rect 3938 10186 3990 10238
rect 4274 10100 4326 10152
rect 3434 10014 3486 10066
rect 174 9938 226 9990
rect 790 9938 842 9990
rect 3013 9981 3065 9990
rect 3013 9947 3022 9981
rect 3022 9947 3056 9981
rect 3056 9947 3065 9981
rect 3013 9938 3065 9947
rect 3938 9928 3990 9980
rect 4274 9842 4326 9894
rect 3518 9756 3570 9808
rect 3938 9670 3990 9722
rect 4274 9584 4326 9636
rect 6440 9202 6492 9254
rect 4274 8820 4326 8872
rect 3938 8734 3990 8786
rect 3266 8648 3318 8700
rect 4274 8562 4326 8614
rect 3854 8476 3906 8528
rect 3518 8390 3570 8442
rect 4274 8304 4326 8356
rect 3854 8218 3906 8270
rect 3434 8132 3486 8184
rect 6440 7664 6492 7716
rect 3518 7196 3570 7248
rect 3770 7110 3822 7162
rect 4274 7024 4326 7076
rect 3266 6938 3318 6990
rect 3854 6852 3906 6904
rect 4274 6766 4326 6818
rect 3350 6680 3402 6732
rect 3854 6594 3906 6646
rect 4274 6508 4326 6560
rect 6440 6126 6492 6178
rect 4274 5744 4326 5796
rect 3770 5658 3822 5710
rect 3434 5572 3486 5624
rect 4274 5486 4326 5538
rect 3013 5449 3065 5458
rect 3013 5415 3022 5449
rect 3022 5415 3056 5449
rect 3056 5415 3065 5449
rect 3013 5406 3065 5415
rect 3770 5400 3822 5452
rect 3350 5314 3402 5366
rect 4274 5228 4326 5280
rect 3770 5142 3822 5194
rect 3266 5056 3318 5108
rect 6440 4588 6492 4640
rect 3350 4120 3402 4172
rect 3686 4034 3738 4086
rect 4274 3948 4326 4000
rect 3434 3862 3486 3914
rect 3013 3825 3065 3834
rect 3013 3791 3022 3825
rect 3022 3791 3056 3825
rect 3056 3791 3065 3825
rect 3013 3782 3065 3791
rect 3686 3776 3738 3828
rect 4274 3690 4326 3742
rect 3518 3604 3570 3656
rect 3686 3518 3738 3570
rect 4274 3432 4326 3484
rect 6440 3050 6492 3102
rect 4274 2668 4326 2720
rect 3686 2582 3738 2634
rect 3266 2496 3318 2548
rect 4274 2410 4326 2462
rect 90 2326 142 2378
rect 1306 2326 1358 2378
rect 3013 2369 3065 2378
rect 3013 2335 3022 2369
rect 3022 2335 3056 2369
rect 3056 2335 3065 2369
rect 3013 2326 3065 2335
rect 3602 2324 3654 2376
rect 3518 2238 3570 2290
rect 4274 2152 4326 2204
rect 3602 2066 3654 2118
rect 3434 1980 3486 2032
rect 6440 1512 6492 1564
rect 3266 786 3318 838
rect 6 702 58 754
rect 1222 702 1274 754
rect 3013 745 3065 754
rect 3013 711 3022 745
rect 3022 711 3056 745
rect 3056 711 3065 745
rect 3013 702 3065 711
rect 3602 700 3654 752
rect 4274 614 4326 666
rect 3350 528 3402 580
rect 3602 442 3654 494
rect 4274 356 4326 408
rect 6440 -26 6492 26
<< metal2 >>
rect 6438 98460 6494 98469
rect 3278 97394 3306 98460
rect 3362 97652 3390 98460
rect 3446 97910 3474 98460
rect 3434 97904 3486 97910
rect 3434 97846 3486 97852
rect 3350 97646 3402 97652
rect 3350 97588 3402 97594
rect 3266 97388 3318 97394
rect 3266 97330 3318 97336
rect 3278 94834 3306 97330
rect 3362 96458 3390 97588
rect 3350 96452 3402 96458
rect 3350 96394 3402 96400
rect 3266 94828 3318 94834
rect 3266 94770 3318 94776
rect 3278 93124 3306 94770
rect 3266 93118 3318 93124
rect 3266 93060 3318 93066
rect 3278 91242 3306 93060
rect 3362 92866 3390 96394
rect 3446 96200 3474 97846
rect 3434 96194 3486 96200
rect 3434 96136 3486 96142
rect 3446 94318 3474 96136
rect 3530 95942 3558 98460
rect 3518 95936 3570 95942
rect 3518 95878 3570 95884
rect 3530 94576 3558 95878
rect 3518 94570 3570 94576
rect 3518 94512 3570 94518
rect 3434 94312 3486 94318
rect 3434 94254 3486 94260
rect 3350 92860 3402 92866
rect 3350 92802 3402 92808
rect 3362 91500 3390 92802
rect 3446 91758 3474 94254
rect 3530 93382 3558 94512
rect 3518 93376 3570 93382
rect 3518 93318 3570 93324
rect 3434 91752 3486 91758
rect 3434 91694 3486 91700
rect 3350 91494 3402 91500
rect 3350 91436 3402 91442
rect 3266 91236 3318 91242
rect 3266 91178 3318 91184
rect 3278 88682 3306 91178
rect 3362 90306 3390 91436
rect 3350 90300 3402 90306
rect 3350 90242 3402 90248
rect 3266 88676 3318 88682
rect 3266 88618 3318 88624
rect 3278 86972 3306 88618
rect 3266 86966 3318 86972
rect 3266 86908 3318 86914
rect 3278 85090 3306 86908
rect 3362 86714 3390 90242
rect 3446 90048 3474 91694
rect 3434 90042 3486 90048
rect 3434 89984 3486 89990
rect 3446 88166 3474 89984
rect 3530 89790 3558 93318
rect 3518 89784 3570 89790
rect 3518 89726 3570 89732
rect 3530 88424 3558 89726
rect 3518 88418 3570 88424
rect 3518 88360 3570 88366
rect 3434 88160 3486 88166
rect 3434 88102 3486 88108
rect 3350 86708 3402 86714
rect 3350 86650 3402 86656
rect 3362 85348 3390 86650
rect 3446 85606 3474 88102
rect 3530 87230 3558 88360
rect 3518 87224 3570 87230
rect 3518 87166 3570 87172
rect 3434 85600 3486 85606
rect 3434 85542 3486 85548
rect 3350 85342 3402 85348
rect 3350 85284 3402 85290
rect 3266 85084 3318 85090
rect 3266 85026 3318 85032
rect 3278 82530 3306 85026
rect 3362 84154 3390 85284
rect 3350 84148 3402 84154
rect 3350 84090 3402 84096
rect 3266 82524 3318 82530
rect 3266 82466 3318 82472
rect 3278 80820 3306 82466
rect 3266 80814 3318 80820
rect 3266 80756 3318 80762
rect 3278 78938 3306 80756
rect 3362 80562 3390 84090
rect 3446 83896 3474 85542
rect 3434 83890 3486 83896
rect 3434 83832 3486 83838
rect 3446 82014 3474 83832
rect 3530 83638 3558 87166
rect 3614 84068 3642 98460
rect 3698 87144 3726 98460
rect 3782 88510 3810 98460
rect 3866 90220 3894 98460
rect 3950 93296 3978 98460
rect 4034 94662 4062 98460
rect 4118 96372 4146 98460
rect 4202 97996 4230 98460
rect 4190 97990 4242 97996
rect 4190 97932 4242 97938
rect 4202 97738 4230 97932
rect 4190 97732 4242 97738
rect 4190 97674 4242 97680
rect 4202 97480 4230 97674
rect 4190 97474 4242 97480
rect 4190 97416 4242 97422
rect 4106 96366 4158 96372
rect 4106 96308 4158 96314
rect 4118 96114 4146 96308
rect 4106 96108 4158 96114
rect 4106 96050 4158 96056
rect 4118 95856 4146 96050
rect 4106 95850 4158 95856
rect 4106 95792 4158 95798
rect 4118 94920 4146 95792
rect 4106 94914 4158 94920
rect 4106 94856 4158 94862
rect 4022 94656 4074 94662
rect 4022 94598 4074 94604
rect 4034 94404 4062 94598
rect 4022 94398 4074 94404
rect 4022 94340 4074 94346
rect 3938 93290 3990 93296
rect 3938 93232 3990 93238
rect 3950 91844 3978 93232
rect 4034 93038 4062 94340
rect 4022 93032 4074 93038
rect 4022 92974 4074 92980
rect 4034 92780 4062 92974
rect 4022 92774 4074 92780
rect 4022 92716 4074 92722
rect 3938 91838 3990 91844
rect 3938 91780 3990 91786
rect 3950 91586 3978 91780
rect 3938 91580 3990 91586
rect 3938 91522 3990 91528
rect 3950 91328 3978 91522
rect 3938 91322 3990 91328
rect 3938 91264 3990 91270
rect 3854 90214 3906 90220
rect 3854 90156 3906 90162
rect 3866 89962 3894 90156
rect 3854 89956 3906 89962
rect 3854 89898 3906 89904
rect 3866 89704 3894 89898
rect 3854 89698 3906 89704
rect 3854 89640 3906 89646
rect 3866 88768 3894 89640
rect 3854 88762 3906 88768
rect 3854 88704 3906 88710
rect 3770 88504 3822 88510
rect 3770 88446 3822 88452
rect 3782 88252 3810 88446
rect 3770 88246 3822 88252
rect 3770 88188 3822 88194
rect 3686 87138 3738 87144
rect 3686 87080 3738 87086
rect 3698 85692 3726 87080
rect 3782 86886 3810 88188
rect 3770 86880 3822 86886
rect 3770 86822 3822 86828
rect 3782 86628 3810 86822
rect 3770 86622 3822 86628
rect 3770 86564 3822 86570
rect 3686 85686 3738 85692
rect 3686 85628 3738 85634
rect 3698 85434 3726 85628
rect 3686 85428 3738 85434
rect 3686 85370 3738 85376
rect 3698 85176 3726 85370
rect 3686 85170 3738 85176
rect 3686 85112 3738 85118
rect 3602 84062 3654 84068
rect 3602 84004 3654 84010
rect 3614 83810 3642 84004
rect 3602 83804 3654 83810
rect 3602 83746 3654 83752
rect 3518 83632 3570 83638
rect 3518 83574 3570 83580
rect 3530 82272 3558 83574
rect 3614 83552 3642 83746
rect 3602 83546 3654 83552
rect 3602 83488 3654 83494
rect 3614 82616 3642 83488
rect 3602 82610 3654 82616
rect 3602 82552 3654 82558
rect 3518 82266 3570 82272
rect 3518 82208 3570 82214
rect 3434 82008 3486 82014
rect 3434 81950 3486 81956
rect 3350 80556 3402 80562
rect 3350 80498 3402 80504
rect 3362 79196 3390 80498
rect 3446 79454 3474 81950
rect 3530 81078 3558 82208
rect 3518 81072 3570 81078
rect 3518 81014 3570 81020
rect 3434 79448 3486 79454
rect 3434 79390 3486 79396
rect 3350 79190 3402 79196
rect 3350 79132 3402 79138
rect 3266 78932 3318 78938
rect 3266 78874 3318 78880
rect 3278 76378 3306 78874
rect 3362 78002 3390 79132
rect 3350 77996 3402 78002
rect 3350 77938 3402 77944
rect 3266 76372 3318 76378
rect 3266 76314 3318 76320
rect 3278 74668 3306 76314
rect 3266 74662 3318 74668
rect 3266 74604 3318 74610
rect 3278 72786 3306 74604
rect 3362 74410 3390 77938
rect 3446 77744 3474 79390
rect 3434 77738 3486 77744
rect 3434 77680 3486 77686
rect 3446 75862 3474 77680
rect 3530 77486 3558 81014
rect 3518 77480 3570 77486
rect 3518 77422 3570 77428
rect 3530 76120 3558 77422
rect 3518 76114 3570 76120
rect 3518 76056 3570 76062
rect 3434 75856 3486 75862
rect 3434 75798 3486 75804
rect 3350 74404 3402 74410
rect 3350 74346 3402 74352
rect 3362 73044 3390 74346
rect 3446 73302 3474 75798
rect 3530 74926 3558 76056
rect 3518 74920 3570 74926
rect 3518 74862 3570 74868
rect 3434 73296 3486 73302
rect 3434 73238 3486 73244
rect 3350 73038 3402 73044
rect 3350 72980 3402 72986
rect 3266 72780 3318 72786
rect 3266 72722 3318 72728
rect 3278 70226 3306 72722
rect 3362 71850 3390 72980
rect 3350 71844 3402 71850
rect 3350 71786 3402 71792
rect 3266 70220 3318 70226
rect 3266 70162 3318 70168
rect 3278 68516 3306 70162
rect 3266 68510 3318 68516
rect 3266 68452 3318 68458
rect 3278 66634 3306 68452
rect 3362 68258 3390 71786
rect 3446 71592 3474 73238
rect 3434 71586 3486 71592
rect 3434 71528 3486 71534
rect 3446 69710 3474 71528
rect 3530 71334 3558 74862
rect 3518 71328 3570 71334
rect 3518 71270 3570 71276
rect 3530 69968 3558 71270
rect 3518 69962 3570 69968
rect 3518 69904 3570 69910
rect 3434 69704 3486 69710
rect 3434 69646 3486 69652
rect 3350 68252 3402 68258
rect 3350 68194 3402 68200
rect 3362 66892 3390 68194
rect 3446 67150 3474 69646
rect 3530 68774 3558 69904
rect 3518 68768 3570 68774
rect 3518 68710 3570 68716
rect 3434 67144 3486 67150
rect 3434 67086 3486 67092
rect 3350 66886 3402 66892
rect 3350 66828 3402 66834
rect 3266 66628 3318 66634
rect 3266 66570 3318 66576
rect 3278 64074 3306 66570
rect 3362 65698 3390 66828
rect 3350 65692 3402 65698
rect 3350 65634 3402 65640
rect 3266 64068 3318 64074
rect 3266 64010 3318 64016
rect 3278 62364 3306 64010
rect 3266 62358 3318 62364
rect 3266 62300 3318 62306
rect 3278 60482 3306 62300
rect 3362 62106 3390 65634
rect 3446 65440 3474 67086
rect 3434 65434 3486 65440
rect 3434 65376 3486 65382
rect 3446 63558 3474 65376
rect 3530 65182 3558 68710
rect 3614 68688 3642 82552
rect 3698 70054 3726 85112
rect 3782 71764 3810 86564
rect 3866 74840 3894 88704
rect 3950 76206 3978 91264
rect 4034 77916 4062 92716
rect 4118 80992 4146 94856
rect 4202 82358 4230 97416
rect 4190 82352 4242 82358
rect 4190 82294 4242 82300
rect 4202 82100 4230 82294
rect 4190 82094 4242 82100
rect 4190 82036 4242 82042
rect 4106 80986 4158 80992
rect 4106 80928 4158 80934
rect 4118 79540 4146 80928
rect 4202 80734 4230 82036
rect 4190 80728 4242 80734
rect 4190 80670 4242 80676
rect 4202 80476 4230 80670
rect 4190 80470 4242 80476
rect 4190 80412 4242 80418
rect 4106 79534 4158 79540
rect 4106 79476 4158 79482
rect 4118 79282 4146 79476
rect 4106 79276 4158 79282
rect 4106 79218 4158 79224
rect 4118 79024 4146 79218
rect 4106 79018 4158 79024
rect 4106 78960 4158 78966
rect 4022 77910 4074 77916
rect 4022 77852 4074 77858
rect 4034 77658 4062 77852
rect 4022 77652 4074 77658
rect 4022 77594 4074 77600
rect 4034 77400 4062 77594
rect 4022 77394 4074 77400
rect 4022 77336 4074 77342
rect 4034 76464 4062 77336
rect 4022 76458 4074 76464
rect 4022 76400 4074 76406
rect 3938 76200 3990 76206
rect 3938 76142 3990 76148
rect 3950 75948 3978 76142
rect 3938 75942 3990 75948
rect 3938 75884 3990 75890
rect 3854 74834 3906 74840
rect 3854 74776 3906 74782
rect 3866 73388 3894 74776
rect 3950 74582 3978 75884
rect 3938 74576 3990 74582
rect 3938 74518 3990 74524
rect 3950 74324 3978 74518
rect 3938 74318 3990 74324
rect 3938 74260 3990 74266
rect 3854 73382 3906 73388
rect 3854 73324 3906 73330
rect 3866 73130 3894 73324
rect 3854 73124 3906 73130
rect 3854 73066 3906 73072
rect 3866 72872 3894 73066
rect 3854 72866 3906 72872
rect 3854 72808 3906 72814
rect 3770 71758 3822 71764
rect 3770 71700 3822 71706
rect 3782 71506 3810 71700
rect 3770 71500 3822 71506
rect 3770 71442 3822 71448
rect 3782 71248 3810 71442
rect 3770 71242 3822 71248
rect 3770 71184 3822 71190
rect 3782 70312 3810 71184
rect 3770 70306 3822 70312
rect 3770 70248 3822 70254
rect 3686 70048 3738 70054
rect 3686 69990 3738 69996
rect 3698 69796 3726 69990
rect 3686 69790 3738 69796
rect 3686 69732 3738 69738
rect 3602 68682 3654 68688
rect 3602 68624 3654 68630
rect 3614 67236 3642 68624
rect 3698 68430 3726 69732
rect 3686 68424 3738 68430
rect 3686 68366 3738 68372
rect 3698 68172 3726 68366
rect 3686 68166 3738 68172
rect 3686 68108 3738 68114
rect 3602 67230 3654 67236
rect 3602 67172 3654 67178
rect 3614 66978 3642 67172
rect 3602 66972 3654 66978
rect 3602 66914 3654 66920
rect 3614 66720 3642 66914
rect 3602 66714 3654 66720
rect 3602 66656 3654 66662
rect 3518 65176 3570 65182
rect 3518 65118 3570 65124
rect 3530 63816 3558 65118
rect 3518 63810 3570 63816
rect 3518 63752 3570 63758
rect 3434 63552 3486 63558
rect 3434 63494 3486 63500
rect 3350 62100 3402 62106
rect 3350 62042 3402 62048
rect 3362 60740 3390 62042
rect 3446 60998 3474 63494
rect 3530 62622 3558 63752
rect 3518 62616 3570 62622
rect 3518 62558 3570 62564
rect 3434 60992 3486 60998
rect 3434 60934 3486 60940
rect 3350 60734 3402 60740
rect 3350 60676 3402 60682
rect 3266 60476 3318 60482
rect 3266 60418 3318 60424
rect 3278 57922 3306 60418
rect 3362 59546 3390 60676
rect 3350 59540 3402 59546
rect 3350 59482 3402 59488
rect 3266 57916 3318 57922
rect 3266 57858 3318 57864
rect 3278 56212 3306 57858
rect 3266 56206 3318 56212
rect 3266 56148 3318 56154
rect 3278 54330 3306 56148
rect 3362 55954 3390 59482
rect 3446 59288 3474 60934
rect 3434 59282 3486 59288
rect 3434 59224 3486 59230
rect 3446 57406 3474 59224
rect 3530 59030 3558 62558
rect 3518 59024 3570 59030
rect 3518 58966 3570 58972
rect 3530 57664 3558 58966
rect 3518 57658 3570 57664
rect 3518 57600 3570 57606
rect 3434 57400 3486 57406
rect 3434 57342 3486 57348
rect 3350 55948 3402 55954
rect 3350 55890 3402 55896
rect 3362 54588 3390 55890
rect 3446 54846 3474 57342
rect 3530 56470 3558 57600
rect 3518 56464 3570 56470
rect 3518 56406 3570 56412
rect 3434 54840 3486 54846
rect 3434 54782 3486 54788
rect 3350 54582 3402 54588
rect 3350 54524 3402 54530
rect 3266 54324 3318 54330
rect 3266 54266 3318 54272
rect 3278 51770 3306 54266
rect 3362 53394 3390 54524
rect 3350 53388 3402 53394
rect 3350 53330 3402 53336
rect 3266 51764 3318 51770
rect 3266 51706 3318 51712
rect 3278 50060 3306 51706
rect 3266 50054 3318 50060
rect 3266 49996 3318 50002
rect 3278 48178 3306 49996
rect 3362 49802 3390 53330
rect 3446 53136 3474 54782
rect 3434 53130 3486 53136
rect 3434 53072 3486 53078
rect 3446 51254 3474 53072
rect 3530 52878 3558 56406
rect 3518 52872 3570 52878
rect 3518 52814 3570 52820
rect 3530 51512 3558 52814
rect 3614 51598 3642 66656
rect 3698 53308 3726 68108
rect 3782 56384 3810 70248
rect 3866 57750 3894 72808
rect 3950 59460 3978 74260
rect 4034 62536 4062 76400
rect 4118 63902 4146 78960
rect 4202 65612 4230 80412
rect 4190 65606 4242 65612
rect 4190 65548 4242 65554
rect 4202 65354 4230 65548
rect 4190 65348 4242 65354
rect 4190 65290 4242 65296
rect 4202 65096 4230 65290
rect 4190 65090 4242 65096
rect 4190 65032 4242 65038
rect 4202 64160 4230 65032
rect 4190 64154 4242 64160
rect 4190 64096 4242 64102
rect 4106 63896 4158 63902
rect 4106 63838 4158 63844
rect 4118 63644 4146 63838
rect 4106 63638 4158 63644
rect 4106 63580 4158 63586
rect 4022 62530 4074 62536
rect 4022 62472 4074 62478
rect 4034 61084 4062 62472
rect 4118 62278 4146 63580
rect 4106 62272 4158 62278
rect 4106 62214 4158 62220
rect 4118 62020 4146 62214
rect 4106 62014 4158 62020
rect 4106 61956 4158 61962
rect 4022 61078 4074 61084
rect 4022 61020 4074 61026
rect 4034 60826 4062 61020
rect 4022 60820 4074 60826
rect 4022 60762 4074 60768
rect 4034 60568 4062 60762
rect 4022 60562 4074 60568
rect 4022 60504 4074 60510
rect 3938 59454 3990 59460
rect 3938 59396 3990 59402
rect 3950 59202 3978 59396
rect 3938 59196 3990 59202
rect 3938 59138 3990 59144
rect 3950 58944 3978 59138
rect 3938 58938 3990 58944
rect 3938 58880 3990 58886
rect 3950 58008 3978 58880
rect 3938 58002 3990 58008
rect 3938 57944 3990 57950
rect 3854 57744 3906 57750
rect 3854 57686 3906 57692
rect 3866 57492 3894 57686
rect 3854 57486 3906 57492
rect 3854 57428 3906 57434
rect 3770 56378 3822 56384
rect 3770 56320 3822 56326
rect 3782 54932 3810 56320
rect 3866 56126 3894 57428
rect 3854 56120 3906 56126
rect 3854 56062 3906 56068
rect 3866 55868 3894 56062
rect 3854 55862 3906 55868
rect 3854 55804 3906 55810
rect 3770 54926 3822 54932
rect 3770 54868 3822 54874
rect 3782 54674 3810 54868
rect 3770 54668 3822 54674
rect 3770 54610 3822 54616
rect 3782 54416 3810 54610
rect 3770 54410 3822 54416
rect 3770 54352 3822 54358
rect 3686 53302 3738 53308
rect 3686 53244 3738 53250
rect 3698 53050 3726 53244
rect 3686 53044 3738 53050
rect 3686 52986 3738 52992
rect 3698 52792 3726 52986
rect 3686 52786 3738 52792
rect 3686 52728 3738 52734
rect 3698 51856 3726 52728
rect 3686 51850 3738 51856
rect 3686 51792 3738 51798
rect 3602 51592 3654 51598
rect 3602 51534 3654 51540
rect 3518 51506 3570 51512
rect 3518 51448 3570 51454
rect 3434 51248 3486 51254
rect 3434 51190 3486 51196
rect 3350 49796 3402 49802
rect 3350 49738 3402 49744
rect 3362 48436 3390 49738
rect 3446 48694 3474 51190
rect 3530 50318 3558 51448
rect 3614 51340 3642 51534
rect 3602 51334 3654 51340
rect 3602 51276 3654 51282
rect 3518 50312 3570 50318
rect 3518 50254 3570 50260
rect 3434 48688 3486 48694
rect 3434 48630 3486 48636
rect 3350 48430 3402 48436
rect 3350 48372 3402 48378
rect 3266 48172 3318 48178
rect 3266 48114 3318 48120
rect 3278 45618 3306 48114
rect 3362 47242 3390 48372
rect 3350 47236 3402 47242
rect 3350 47178 3402 47184
rect 3266 45612 3318 45618
rect 3266 45554 3318 45560
rect 3278 43908 3306 45554
rect 3266 43902 3318 43908
rect 3266 43844 3318 43850
rect 3278 42026 3306 43844
rect 3362 43650 3390 47178
rect 3446 46984 3474 48630
rect 3434 46978 3486 46984
rect 3434 46920 3486 46926
rect 3446 45102 3474 46920
rect 3530 46726 3558 50254
rect 3614 49974 3642 51276
rect 3602 49968 3654 49974
rect 3602 49910 3654 49916
rect 3614 49716 3642 49910
rect 3602 49710 3654 49716
rect 3602 49652 3654 49658
rect 3518 46720 3570 46726
rect 3518 46662 3570 46668
rect 3530 45360 3558 46662
rect 3518 45354 3570 45360
rect 3518 45296 3570 45302
rect 3434 45096 3486 45102
rect 3434 45038 3486 45044
rect 3350 43644 3402 43650
rect 3350 43586 3402 43592
rect 3362 42284 3390 43586
rect 3446 42542 3474 45038
rect 3530 44166 3558 45296
rect 3518 44160 3570 44166
rect 3518 44102 3570 44108
rect 3434 42536 3486 42542
rect 3434 42478 3486 42484
rect 3350 42278 3402 42284
rect 3350 42220 3402 42226
rect 3266 42020 3318 42026
rect 3266 41962 3318 41968
rect 3278 39466 3306 41962
rect 3362 41090 3390 42220
rect 3350 41084 3402 41090
rect 3350 41026 3402 41032
rect 3266 39460 3318 39466
rect 3266 39402 3318 39408
rect 3278 37756 3306 39402
rect 3266 37750 3318 37756
rect 3266 37692 3318 37698
rect 18 760 46 36952
rect 102 2384 130 36952
rect 186 9996 214 36952
rect 270 11620 298 36952
rect 354 13076 382 36952
rect 438 25392 466 36952
rect 522 27016 550 36952
rect 606 28472 634 36952
rect 3011 36252 3067 36261
rect 3011 36187 3067 36196
rect 3278 35874 3306 37692
rect 3362 37498 3390 41026
rect 3446 40832 3474 42478
rect 3434 40826 3486 40832
rect 3434 40768 3486 40774
rect 3446 38950 3474 40768
rect 3530 40574 3558 44102
rect 3518 40568 3570 40574
rect 3518 40510 3570 40516
rect 3530 39208 3558 40510
rect 3518 39202 3570 39208
rect 3518 39144 3570 39150
rect 3434 38944 3486 38950
rect 3434 38886 3486 38892
rect 3350 37492 3402 37498
rect 3350 37434 3402 37440
rect 3362 36132 3390 37434
rect 3446 36390 3474 38886
rect 3530 38014 3558 39144
rect 3518 38008 3570 38014
rect 3518 37950 3570 37956
rect 3434 36384 3486 36390
rect 3434 36326 3486 36332
rect 3350 36126 3402 36132
rect 3350 36068 3402 36074
rect 3266 35868 3318 35874
rect 3266 35810 3318 35816
rect 3011 34628 3067 34637
rect 3011 34563 3067 34572
rect 3278 33314 3306 35810
rect 3362 34938 3390 36068
rect 3350 34932 3402 34938
rect 3350 34874 3402 34880
rect 3266 33308 3318 33314
rect 3266 33250 3318 33256
rect 3011 33172 3067 33181
rect 3011 33107 3067 33116
rect 3278 31604 3306 33250
rect 3266 31598 3318 31604
rect 3011 31548 3067 31557
rect 3266 31540 3318 31546
rect 3011 31483 3067 31492
rect 3011 30092 3067 30101
rect 3011 30027 3067 30036
rect 3278 29722 3306 31540
rect 3362 31346 3390 34874
rect 3446 34680 3474 36326
rect 3434 34674 3486 34680
rect 3434 34616 3486 34622
rect 3446 32798 3474 34616
rect 3530 34422 3558 37950
rect 3614 34852 3642 49652
rect 3698 37928 3726 51792
rect 3782 39294 3810 54352
rect 3866 41004 3894 55804
rect 3950 44080 3978 57944
rect 4034 45446 4062 60504
rect 4118 47156 4146 61956
rect 4202 50232 4230 64096
rect 4190 50226 4242 50232
rect 4190 50168 4242 50174
rect 4202 48780 4230 50168
rect 4190 48774 4242 48780
rect 4190 48716 4242 48722
rect 4202 48522 4230 48716
rect 4190 48516 4242 48522
rect 4190 48458 4242 48464
rect 4202 48264 4230 48458
rect 4190 48258 4242 48264
rect 4190 48200 4242 48206
rect 4106 47150 4158 47156
rect 4106 47092 4158 47098
rect 4118 46898 4146 47092
rect 4106 46892 4158 46898
rect 4106 46834 4158 46840
rect 4118 46640 4146 46834
rect 4106 46634 4158 46640
rect 4106 46576 4158 46582
rect 4118 45704 4146 46576
rect 4106 45698 4158 45704
rect 4106 45640 4158 45646
rect 4022 45440 4074 45446
rect 4022 45382 4074 45388
rect 4034 45188 4062 45382
rect 4022 45182 4074 45188
rect 4022 45124 4074 45130
rect 3938 44074 3990 44080
rect 3938 44016 3990 44022
rect 3950 42628 3978 44016
rect 4034 43822 4062 45124
rect 4022 43816 4074 43822
rect 4022 43758 4074 43764
rect 4034 43564 4062 43758
rect 4022 43558 4074 43564
rect 4022 43500 4074 43506
rect 3938 42622 3990 42628
rect 3938 42564 3990 42570
rect 3950 42370 3978 42564
rect 3938 42364 3990 42370
rect 3938 42306 3990 42312
rect 3950 42112 3978 42306
rect 3938 42106 3990 42112
rect 3938 42048 3990 42054
rect 3854 40998 3906 41004
rect 3854 40940 3906 40946
rect 3866 40746 3894 40940
rect 3854 40740 3906 40746
rect 3854 40682 3906 40688
rect 3866 40488 3894 40682
rect 3854 40482 3906 40488
rect 3854 40424 3906 40430
rect 3866 39552 3894 40424
rect 3854 39546 3906 39552
rect 3854 39488 3906 39494
rect 3770 39288 3822 39294
rect 3770 39230 3822 39236
rect 3782 39036 3810 39230
rect 3770 39030 3822 39036
rect 3770 38972 3822 38978
rect 3686 37922 3738 37928
rect 3686 37864 3738 37870
rect 3698 36476 3726 37864
rect 3782 37670 3810 38972
rect 3770 37664 3822 37670
rect 3770 37606 3822 37612
rect 3782 37412 3810 37606
rect 3770 37406 3822 37412
rect 3770 37348 3822 37354
rect 3686 36470 3738 36476
rect 3686 36412 3738 36418
rect 3698 36218 3726 36412
rect 3686 36212 3738 36218
rect 3686 36154 3738 36160
rect 3698 35960 3726 36154
rect 3686 35954 3738 35960
rect 3686 35896 3738 35902
rect 3602 34846 3654 34852
rect 3602 34788 3654 34794
rect 3614 34594 3642 34788
rect 3602 34588 3654 34594
rect 3602 34530 3654 34536
rect 3518 34416 3570 34422
rect 3518 34358 3570 34364
rect 3530 33056 3558 34358
rect 3614 34336 3642 34530
rect 3602 34330 3654 34336
rect 3602 34272 3654 34278
rect 3614 33400 3642 34272
rect 3602 33394 3654 33400
rect 3602 33336 3654 33342
rect 3518 33050 3570 33056
rect 3518 32992 3570 32998
rect 3434 32792 3486 32798
rect 3434 32734 3486 32740
rect 3350 31340 3402 31346
rect 3350 31282 3402 31288
rect 3362 29980 3390 31282
rect 3446 30238 3474 32734
rect 3530 31862 3558 32992
rect 3518 31856 3570 31862
rect 3518 31798 3570 31804
rect 3434 30232 3486 30238
rect 3434 30174 3486 30180
rect 3350 29974 3402 29980
rect 3350 29916 3402 29922
rect 3266 29716 3318 29722
rect 3266 29658 3318 29664
rect 594 28466 646 28472
rect 594 28408 646 28414
rect 958 28466 1010 28472
rect 958 28408 1010 28414
rect 3011 28468 3067 28477
rect 510 27010 562 27016
rect 510 26952 562 26958
rect 426 25386 478 25392
rect 426 25328 478 25334
rect 342 13070 394 13076
rect 342 13012 394 13018
rect 258 11614 310 11620
rect 258 11556 310 11562
rect 174 9990 226 9996
rect 174 9932 226 9938
rect 90 2378 142 2384
rect 90 2320 142 2326
rect 6 754 58 760
rect 6 696 58 702
rect 18 0 46 696
rect 102 0 130 2320
rect 186 0 214 9932
rect 270 0 298 11556
rect 354 0 382 13012
rect 438 0 466 25328
rect 522 0 550 26952
rect 606 0 634 28408
rect 3011 28403 3067 28412
rect 3278 27162 3306 29658
rect 3362 28786 3390 29916
rect 3350 28780 3402 28786
rect 3350 28722 3402 28728
rect 3266 27156 3318 27162
rect 3266 27098 3318 27104
rect 874 27010 926 27016
rect 874 26952 926 26958
rect 3011 27012 3067 27021
rect 3011 26947 3067 26956
rect 3278 25452 3306 27098
rect 3266 25446 3318 25452
rect 790 25386 842 25392
rect 790 25328 842 25334
rect 3011 25388 3067 25397
rect 3266 25388 3318 25394
rect 3011 25323 3067 25332
rect 3278 23570 3306 25388
rect 3362 25194 3390 28722
rect 3446 28528 3474 30174
rect 3434 28522 3486 28528
rect 3434 28464 3486 28470
rect 3446 26646 3474 28464
rect 3530 28270 3558 31798
rect 3518 28264 3570 28270
rect 3518 28206 3570 28212
rect 3530 26904 3558 28206
rect 3518 26898 3570 26904
rect 3518 26840 3570 26846
rect 3434 26640 3486 26646
rect 3434 26582 3486 26588
rect 3350 25188 3402 25194
rect 3350 25130 3402 25136
rect 3362 23828 3390 25130
rect 3446 24086 3474 26582
rect 3530 25710 3558 26840
rect 3518 25704 3570 25710
rect 3518 25646 3570 25652
rect 3434 24080 3486 24086
rect 3434 24022 3486 24028
rect 3350 23822 3402 23828
rect 3350 23764 3402 23770
rect 3266 23564 3318 23570
rect 3266 23506 3318 23512
rect 3278 21010 3306 23506
rect 3362 22634 3390 23764
rect 3350 22628 3402 22634
rect 3350 22570 3402 22576
rect 3266 21004 3318 21010
rect 3266 20946 3318 20952
rect 3011 20856 3067 20865
rect 3011 20791 3067 20800
rect 3278 19300 3306 20946
rect 3266 19294 3318 19300
rect 3011 19232 3067 19241
rect 3266 19236 3318 19242
rect 3011 19167 3067 19176
rect 3011 17776 3067 17785
rect 3011 17711 3067 17720
rect 3278 17418 3306 19236
rect 3362 19042 3390 22570
rect 3446 22376 3474 24022
rect 3434 22370 3486 22376
rect 3434 22312 3486 22318
rect 3446 20494 3474 22312
rect 3530 22118 3558 25646
rect 3518 22112 3570 22118
rect 3518 22054 3570 22060
rect 3530 20752 3558 22054
rect 3518 20746 3570 20752
rect 3518 20688 3570 20694
rect 3434 20488 3486 20494
rect 3434 20430 3486 20436
rect 3350 19036 3402 19042
rect 3350 18978 3402 18984
rect 3362 17676 3390 18978
rect 3446 17934 3474 20430
rect 3530 19558 3558 20688
rect 3518 19552 3570 19558
rect 3518 19494 3570 19500
rect 3434 17928 3486 17934
rect 3434 17870 3486 17876
rect 3350 17670 3402 17676
rect 3350 17612 3402 17618
rect 3266 17412 3318 17418
rect 3266 17354 3318 17360
rect 3011 16152 3067 16161
rect 3011 16087 3067 16096
rect 3278 14858 3306 17354
rect 3362 16482 3390 17612
rect 3350 16476 3402 16482
rect 3350 16418 3402 16424
rect 3266 14852 3318 14858
rect 3266 14794 3318 14800
rect 3011 14696 3067 14705
rect 3011 14631 3067 14640
rect 3278 13148 3306 14794
rect 3266 13142 3318 13148
rect 3266 13084 3318 13090
rect 958 13070 1010 13076
rect 958 13012 1010 13018
rect 3011 13072 3067 13081
rect 3011 13007 3067 13016
rect 874 11614 926 11620
rect 874 11556 926 11562
rect 3011 11616 3067 11625
rect 3011 11551 3067 11560
rect 3278 11266 3306 13084
rect 3362 12890 3390 16418
rect 3446 16224 3474 17870
rect 3434 16218 3486 16224
rect 3434 16160 3486 16166
rect 3446 14342 3474 16160
rect 3530 15966 3558 19494
rect 3614 19472 3642 33336
rect 3698 20838 3726 35896
rect 3782 22548 3810 37348
rect 3866 25624 3894 39488
rect 3950 26990 3978 42048
rect 4034 28700 4062 43500
rect 4118 31776 4146 45640
rect 4202 33142 4230 48200
rect 4190 33136 4242 33142
rect 4190 33078 4242 33084
rect 4202 32884 4230 33078
rect 4190 32878 4242 32884
rect 4190 32820 4242 32826
rect 4106 31770 4158 31776
rect 4106 31712 4158 31718
rect 4118 30324 4146 31712
rect 4202 31518 4230 32820
rect 4190 31512 4242 31518
rect 4190 31454 4242 31460
rect 4202 31260 4230 31454
rect 4190 31254 4242 31260
rect 4190 31196 4242 31202
rect 4106 30318 4158 30324
rect 4106 30260 4158 30266
rect 4118 30066 4146 30260
rect 4106 30060 4158 30066
rect 4106 30002 4158 30008
rect 4118 29808 4146 30002
rect 4106 29802 4158 29808
rect 4106 29744 4158 29750
rect 4022 28694 4074 28700
rect 4022 28636 4074 28642
rect 4034 28442 4062 28636
rect 4022 28436 4074 28442
rect 4022 28378 4074 28384
rect 4034 28184 4062 28378
rect 4022 28178 4074 28184
rect 4022 28120 4074 28126
rect 4034 27248 4062 28120
rect 4022 27242 4074 27248
rect 4022 27184 4074 27190
rect 3938 26984 3990 26990
rect 3938 26926 3990 26932
rect 3950 26732 3978 26926
rect 3938 26726 3990 26732
rect 3938 26668 3990 26674
rect 3854 25618 3906 25624
rect 3854 25560 3906 25566
rect 3866 24172 3894 25560
rect 3950 25366 3978 26668
rect 3938 25360 3990 25366
rect 3938 25302 3990 25308
rect 3950 25108 3978 25302
rect 3938 25102 3990 25108
rect 3938 25044 3990 25050
rect 3854 24166 3906 24172
rect 3854 24108 3906 24114
rect 3866 23914 3894 24108
rect 3854 23908 3906 23914
rect 3854 23850 3906 23856
rect 3866 23656 3894 23850
rect 3854 23650 3906 23656
rect 3854 23592 3906 23598
rect 3770 22542 3822 22548
rect 3770 22484 3822 22490
rect 3782 22290 3810 22484
rect 3770 22284 3822 22290
rect 3770 22226 3822 22232
rect 3782 22032 3810 22226
rect 3770 22026 3822 22032
rect 3770 21968 3822 21974
rect 3782 21096 3810 21968
rect 3770 21090 3822 21096
rect 3770 21032 3822 21038
rect 3686 20832 3738 20838
rect 3686 20774 3738 20780
rect 3698 20580 3726 20774
rect 3686 20574 3738 20580
rect 3686 20516 3738 20522
rect 3602 19466 3654 19472
rect 3602 19408 3654 19414
rect 3614 18020 3642 19408
rect 3698 19214 3726 20516
rect 3686 19208 3738 19214
rect 3686 19150 3738 19156
rect 3698 18956 3726 19150
rect 3686 18950 3738 18956
rect 3686 18892 3738 18898
rect 3602 18014 3654 18020
rect 3602 17956 3654 17962
rect 3614 17762 3642 17956
rect 3602 17756 3654 17762
rect 3602 17698 3654 17704
rect 3614 17504 3642 17698
rect 3602 17498 3654 17504
rect 3602 17440 3654 17446
rect 3518 15960 3570 15966
rect 3518 15902 3570 15908
rect 3530 14600 3558 15902
rect 3518 14594 3570 14600
rect 3518 14536 3570 14542
rect 3434 14336 3486 14342
rect 3434 14278 3486 14284
rect 3350 12884 3402 12890
rect 3350 12826 3402 12832
rect 3362 11524 3390 12826
rect 3446 11782 3474 14278
rect 3530 13406 3558 14536
rect 3518 13400 3570 13406
rect 3518 13342 3570 13348
rect 3434 11776 3486 11782
rect 3434 11718 3486 11724
rect 3350 11518 3402 11524
rect 3350 11460 3402 11466
rect 3266 11260 3318 11266
rect 3266 11202 3318 11208
rect 790 9990 842 9996
rect 790 9932 842 9938
rect 3011 9992 3067 10001
rect 3011 9927 3067 9936
rect 3278 8706 3306 11202
rect 3362 10330 3390 11460
rect 3350 10324 3402 10330
rect 3350 10266 3402 10272
rect 3266 8700 3318 8706
rect 3266 8642 3318 8648
rect 3278 6996 3306 8642
rect 3266 6990 3318 6996
rect 3266 6932 3318 6938
rect 3011 5460 3067 5469
rect 3011 5395 3067 5404
rect 3278 5114 3306 6932
rect 3362 6738 3390 10266
rect 3446 10072 3474 11718
rect 3434 10066 3486 10072
rect 3434 10008 3486 10014
rect 3446 8190 3474 10008
rect 3530 9814 3558 13342
rect 3518 9808 3570 9814
rect 3518 9750 3570 9756
rect 3530 8448 3558 9750
rect 3614 9273 3642 17440
rect 3698 10813 3726 18892
rect 3782 12353 3810 21032
rect 3866 13893 3894 23592
rect 3950 15433 3978 25044
rect 4034 16973 4062 27184
rect 4118 18513 4146 29744
rect 4202 20053 4230 31196
rect 4286 24669 4314 98460
rect 4370 33228 4398 98460
rect 4454 50146 4482 98460
rect 4538 65526 4566 98460
rect 4622 82444 4650 98460
rect 4706 98082 4734 98460
rect 4694 98076 4746 98082
rect 4694 98018 4746 98024
rect 4706 97824 4734 98018
rect 4694 97818 4746 97824
rect 4694 97760 4746 97766
rect 4706 97566 4734 97760
rect 4694 97560 4746 97566
rect 4694 97502 4746 97508
rect 4706 96286 4734 97502
rect 4694 96280 4746 96286
rect 4694 96222 4746 96228
rect 4706 96028 4734 96222
rect 4694 96022 4746 96028
rect 4694 95964 4746 95970
rect 4706 95770 4734 95964
rect 4694 95764 4746 95770
rect 4694 95706 4746 95712
rect 4706 95006 4734 95706
rect 4694 95000 4746 95006
rect 4694 94942 4746 94948
rect 4706 94748 4734 94942
rect 4694 94742 4746 94748
rect 4694 94684 4746 94690
rect 4706 94490 4734 94684
rect 4694 94484 4746 94490
rect 4694 94426 4746 94432
rect 4706 93210 4734 94426
rect 4694 93204 4746 93210
rect 4694 93146 4746 93152
rect 4706 92952 4734 93146
rect 4694 92946 4746 92952
rect 4694 92888 4746 92894
rect 4706 92694 4734 92888
rect 4694 92688 4746 92694
rect 4694 92630 4746 92636
rect 4706 91930 4734 92630
rect 4694 91924 4746 91930
rect 4694 91866 4746 91872
rect 4706 91672 4734 91866
rect 4694 91666 4746 91672
rect 4694 91608 4746 91614
rect 4706 91414 4734 91608
rect 4694 91408 4746 91414
rect 4694 91350 4746 91356
rect 4706 90134 4734 91350
rect 4694 90128 4746 90134
rect 4694 90070 4746 90076
rect 4706 89876 4734 90070
rect 4694 89870 4746 89876
rect 4694 89812 4746 89818
rect 4706 89618 4734 89812
rect 4694 89612 4746 89618
rect 4694 89554 4746 89560
rect 4706 88854 4734 89554
rect 4694 88848 4746 88854
rect 4694 88790 4746 88796
rect 4706 88596 4734 88790
rect 4694 88590 4746 88596
rect 4694 88532 4746 88538
rect 4706 88338 4734 88532
rect 4694 88332 4746 88338
rect 4694 88274 4746 88280
rect 4706 87058 4734 88274
rect 4694 87052 4746 87058
rect 4694 86994 4746 87000
rect 4706 86800 4734 86994
rect 4694 86794 4746 86800
rect 4694 86736 4746 86742
rect 4706 86542 4734 86736
rect 4694 86536 4746 86542
rect 4694 86478 4746 86484
rect 4706 85778 4734 86478
rect 4694 85772 4746 85778
rect 4694 85714 4746 85720
rect 4706 85520 4734 85714
rect 4694 85514 4746 85520
rect 4694 85456 4746 85462
rect 4706 85262 4734 85456
rect 4694 85256 4746 85262
rect 4694 85198 4746 85204
rect 4706 83982 4734 85198
rect 4694 83976 4746 83982
rect 4694 83918 4746 83924
rect 4706 83724 4734 83918
rect 4694 83718 4746 83724
rect 4694 83660 4746 83666
rect 4706 83466 4734 83660
rect 4694 83460 4746 83466
rect 4694 83402 4746 83408
rect 4706 82702 4734 83402
rect 4694 82696 4746 82702
rect 4694 82638 4746 82644
rect 4610 82438 4662 82444
rect 4610 82380 4662 82386
rect 4622 82186 4650 82380
rect 4610 82180 4662 82186
rect 4610 82122 4662 82128
rect 4622 80906 4650 82122
rect 4610 80900 4662 80906
rect 4610 80842 4662 80848
rect 4622 80648 4650 80842
rect 4610 80642 4662 80648
rect 4610 80584 4662 80590
rect 4622 80390 4650 80584
rect 4610 80384 4662 80390
rect 4610 80326 4662 80332
rect 4622 79626 4650 80326
rect 4610 79620 4662 79626
rect 4610 79562 4662 79568
rect 4622 79368 4650 79562
rect 4610 79362 4662 79368
rect 4610 79304 4662 79310
rect 4622 79110 4650 79304
rect 4610 79104 4662 79110
rect 4610 79046 4662 79052
rect 4622 77830 4650 79046
rect 4610 77824 4662 77830
rect 4610 77766 4662 77772
rect 4622 77572 4650 77766
rect 4610 77566 4662 77572
rect 4610 77508 4662 77514
rect 4622 77314 4650 77508
rect 4610 77308 4662 77314
rect 4610 77250 4662 77256
rect 4622 76550 4650 77250
rect 4610 76544 4662 76550
rect 4610 76486 4662 76492
rect 4622 76292 4650 76486
rect 4610 76286 4662 76292
rect 4610 76228 4662 76234
rect 4622 76034 4650 76228
rect 4610 76028 4662 76034
rect 4610 75970 4662 75976
rect 4622 74754 4650 75970
rect 4610 74748 4662 74754
rect 4610 74690 4662 74696
rect 4622 74496 4650 74690
rect 4610 74490 4662 74496
rect 4610 74432 4662 74438
rect 4622 74238 4650 74432
rect 4610 74232 4662 74238
rect 4610 74174 4662 74180
rect 4622 73474 4650 74174
rect 4610 73468 4662 73474
rect 4610 73410 4662 73416
rect 4622 73216 4650 73410
rect 4610 73210 4662 73216
rect 4610 73152 4662 73158
rect 4622 72958 4650 73152
rect 4610 72952 4662 72958
rect 4610 72894 4662 72900
rect 4622 71678 4650 72894
rect 4610 71672 4662 71678
rect 4610 71614 4662 71620
rect 4622 71420 4650 71614
rect 4610 71414 4662 71420
rect 4610 71356 4662 71362
rect 4622 71162 4650 71356
rect 4610 71156 4662 71162
rect 4610 71098 4662 71104
rect 4622 70398 4650 71098
rect 4610 70392 4662 70398
rect 4610 70334 4662 70340
rect 4622 70140 4650 70334
rect 4610 70134 4662 70140
rect 4610 70076 4662 70082
rect 4622 69882 4650 70076
rect 4610 69876 4662 69882
rect 4610 69818 4662 69824
rect 4622 68602 4650 69818
rect 4610 68596 4662 68602
rect 4610 68538 4662 68544
rect 4622 68344 4650 68538
rect 4610 68338 4662 68344
rect 4610 68280 4662 68286
rect 4622 68086 4650 68280
rect 4610 68080 4662 68086
rect 4610 68022 4662 68028
rect 4622 67322 4650 68022
rect 4610 67316 4662 67322
rect 4610 67258 4662 67264
rect 4622 67064 4650 67258
rect 4610 67058 4662 67064
rect 4610 67000 4662 67006
rect 4622 66806 4650 67000
rect 4610 66800 4662 66806
rect 4610 66742 4662 66748
rect 4526 65520 4578 65526
rect 4526 65462 4578 65468
rect 4538 65268 4566 65462
rect 4526 65262 4578 65268
rect 4526 65204 4578 65210
rect 4538 65010 4566 65204
rect 4526 65004 4578 65010
rect 4526 64946 4578 64952
rect 4538 64246 4566 64946
rect 4526 64240 4578 64246
rect 4526 64182 4578 64188
rect 4538 63988 4566 64182
rect 4526 63982 4578 63988
rect 4526 63924 4578 63930
rect 4538 63730 4566 63924
rect 4526 63724 4578 63730
rect 4526 63666 4578 63672
rect 4538 62450 4566 63666
rect 4526 62444 4578 62450
rect 4526 62386 4578 62392
rect 4538 62192 4566 62386
rect 4526 62186 4578 62192
rect 4526 62128 4578 62134
rect 4538 61934 4566 62128
rect 4526 61928 4578 61934
rect 4526 61870 4578 61876
rect 4538 61170 4566 61870
rect 4526 61164 4578 61170
rect 4526 61106 4578 61112
rect 4538 60912 4566 61106
rect 4526 60906 4578 60912
rect 4526 60848 4578 60854
rect 4538 60654 4566 60848
rect 4526 60648 4578 60654
rect 4526 60590 4578 60596
rect 4538 59374 4566 60590
rect 4526 59368 4578 59374
rect 4526 59310 4578 59316
rect 4538 59116 4566 59310
rect 4526 59110 4578 59116
rect 4526 59052 4578 59058
rect 4538 58858 4566 59052
rect 4526 58852 4578 58858
rect 4526 58794 4578 58800
rect 4538 58094 4566 58794
rect 4526 58088 4578 58094
rect 4526 58030 4578 58036
rect 4538 57836 4566 58030
rect 4526 57830 4578 57836
rect 4526 57772 4578 57778
rect 4538 57578 4566 57772
rect 4526 57572 4578 57578
rect 4526 57514 4578 57520
rect 4538 56298 4566 57514
rect 4526 56292 4578 56298
rect 4526 56234 4578 56240
rect 4538 56040 4566 56234
rect 4526 56034 4578 56040
rect 4526 55976 4578 55982
rect 4538 55782 4566 55976
rect 4526 55776 4578 55782
rect 4526 55718 4578 55724
rect 4538 55018 4566 55718
rect 4526 55012 4578 55018
rect 4526 54954 4578 54960
rect 4538 54760 4566 54954
rect 4526 54754 4578 54760
rect 4526 54696 4578 54702
rect 4538 54502 4566 54696
rect 4526 54496 4578 54502
rect 4526 54438 4578 54444
rect 4538 53222 4566 54438
rect 4526 53216 4578 53222
rect 4526 53158 4578 53164
rect 4538 52964 4566 53158
rect 4526 52958 4578 52964
rect 4526 52900 4578 52906
rect 4538 52706 4566 52900
rect 4526 52700 4578 52706
rect 4526 52642 4578 52648
rect 4538 51942 4566 52642
rect 4526 51936 4578 51942
rect 4526 51878 4578 51884
rect 4538 51684 4566 51878
rect 4526 51678 4578 51684
rect 4526 51620 4578 51626
rect 4538 51426 4566 51620
rect 4526 51420 4578 51426
rect 4526 51362 4578 51368
rect 4442 50140 4494 50146
rect 4442 50082 4494 50088
rect 4454 48866 4482 50082
rect 4538 49888 4566 51362
rect 4526 49882 4578 49888
rect 4526 49824 4578 49830
rect 4538 49630 4566 49824
rect 4526 49624 4578 49630
rect 4526 49566 4578 49572
rect 4442 48860 4494 48866
rect 4442 48802 4494 48808
rect 4454 48608 4482 48802
rect 4442 48602 4494 48608
rect 4442 48544 4494 48550
rect 4454 48350 4482 48544
rect 4442 48344 4494 48350
rect 4442 48286 4494 48292
rect 4454 47070 4482 48286
rect 4442 47064 4494 47070
rect 4442 47006 4494 47012
rect 4454 46812 4482 47006
rect 4442 46806 4494 46812
rect 4442 46748 4494 46754
rect 4454 46554 4482 46748
rect 4442 46548 4494 46554
rect 4442 46490 4494 46496
rect 4454 45790 4482 46490
rect 4442 45784 4494 45790
rect 4442 45726 4494 45732
rect 4454 45532 4482 45726
rect 4442 45526 4494 45532
rect 4442 45468 4494 45474
rect 4454 45274 4482 45468
rect 4442 45268 4494 45274
rect 4442 45210 4494 45216
rect 4454 43994 4482 45210
rect 4442 43988 4494 43994
rect 4442 43930 4494 43936
rect 4454 43736 4482 43930
rect 4442 43730 4494 43736
rect 4442 43672 4494 43678
rect 4454 43478 4482 43672
rect 4442 43472 4494 43478
rect 4442 43414 4494 43420
rect 4454 42714 4482 43414
rect 4442 42708 4494 42714
rect 4442 42650 4494 42656
rect 4454 42456 4482 42650
rect 4442 42450 4494 42456
rect 4442 42392 4494 42398
rect 4454 42198 4482 42392
rect 4442 42192 4494 42198
rect 4442 42134 4494 42140
rect 4454 40918 4482 42134
rect 4442 40912 4494 40918
rect 4442 40854 4494 40860
rect 4454 40660 4482 40854
rect 4442 40654 4494 40660
rect 4442 40596 4494 40602
rect 4454 40402 4482 40596
rect 4442 40396 4494 40402
rect 4442 40338 4494 40344
rect 4454 39638 4482 40338
rect 4442 39632 4494 39638
rect 4442 39574 4494 39580
rect 4454 39380 4482 39574
rect 4442 39374 4494 39380
rect 4442 39316 4494 39322
rect 4454 39122 4482 39316
rect 4442 39116 4494 39122
rect 4442 39058 4494 39064
rect 4454 37842 4482 39058
rect 4442 37836 4494 37842
rect 4442 37778 4494 37784
rect 4454 37584 4482 37778
rect 4442 37578 4494 37584
rect 4442 37520 4494 37526
rect 4454 37326 4482 37520
rect 4442 37320 4494 37326
rect 4442 37262 4494 37268
rect 4454 36562 4482 37262
rect 4442 36556 4494 36562
rect 4442 36498 4494 36504
rect 4454 36304 4482 36498
rect 4442 36298 4494 36304
rect 4442 36240 4494 36246
rect 4454 36046 4482 36240
rect 4442 36040 4494 36046
rect 4442 35982 4494 35988
rect 4454 34766 4482 35982
rect 4442 34760 4494 34766
rect 4442 34702 4494 34708
rect 4454 34508 4482 34702
rect 4442 34502 4494 34508
rect 4442 34444 4494 34450
rect 4454 34250 4482 34444
rect 4442 34244 4494 34250
rect 4442 34186 4494 34192
rect 4454 33486 4482 34186
rect 4442 33480 4494 33486
rect 4442 33422 4494 33428
rect 4358 33222 4410 33228
rect 4358 33164 4410 33170
rect 4370 32970 4398 33164
rect 4358 32964 4410 32970
rect 4358 32906 4410 32912
rect 4370 31690 4398 32906
rect 4358 31684 4410 31690
rect 4358 31626 4410 31632
rect 4370 31432 4398 31626
rect 4358 31426 4410 31432
rect 4358 31368 4410 31374
rect 4370 31174 4398 31368
rect 4358 31168 4410 31174
rect 4358 31110 4410 31116
rect 4370 30410 4398 31110
rect 4358 30404 4410 30410
rect 4358 30346 4410 30352
rect 4370 30152 4398 30346
rect 4358 30146 4410 30152
rect 4358 30088 4410 30094
rect 4370 29894 4398 30088
rect 4358 29888 4410 29894
rect 4358 29830 4410 29836
rect 4370 28614 4398 29830
rect 4358 28608 4410 28614
rect 4358 28550 4410 28556
rect 4370 28356 4398 28550
rect 4358 28350 4410 28356
rect 4358 28292 4410 28298
rect 4370 28098 4398 28292
rect 4358 28092 4410 28098
rect 4358 28034 4410 28040
rect 4370 27334 4398 28034
rect 4454 27749 4482 33422
rect 4538 29289 4566 49566
rect 4622 30829 4650 66742
rect 4706 32369 4734 82638
rect 4790 33909 4818 98460
rect 4874 35449 4902 98460
rect 6438 98395 6494 98404
rect 6438 96922 6494 96931
rect 6438 96857 6494 96866
rect 6438 95384 6494 95393
rect 6438 95319 6494 95328
rect 6438 93846 6494 93855
rect 6438 93781 6494 93790
rect 6438 92308 6494 92317
rect 6438 92243 6494 92252
rect 6438 90770 6494 90779
rect 6438 90705 6494 90714
rect 6438 89232 6494 89241
rect 6438 89167 6494 89176
rect 6438 87694 6494 87703
rect 6438 87629 6494 87638
rect 6438 86156 6494 86165
rect 6438 86091 6494 86100
rect 6438 84618 6494 84627
rect 6438 84553 6494 84562
rect 6438 83080 6494 83089
rect 6438 83015 6494 83024
rect 6438 81542 6494 81551
rect 6438 81477 6494 81486
rect 6438 80004 6494 80013
rect 6438 79939 6494 79948
rect 6438 78466 6494 78475
rect 6438 78401 6494 78410
rect 6438 76928 6494 76937
rect 6438 76863 6494 76872
rect 6438 75390 6494 75399
rect 6438 75325 6494 75334
rect 6438 73852 6494 73861
rect 6438 73787 6494 73796
rect 6438 72314 6494 72323
rect 6438 72249 6494 72258
rect 6438 70776 6494 70785
rect 6438 70711 6494 70720
rect 6438 69238 6494 69247
rect 6438 69173 6494 69182
rect 6438 67700 6494 67709
rect 6438 67635 6494 67644
rect 6438 66162 6494 66171
rect 6438 66097 6494 66106
rect 6438 64624 6494 64633
rect 6438 64559 6494 64568
rect 6438 63086 6494 63095
rect 6438 63021 6494 63030
rect 6438 61548 6494 61557
rect 6438 61483 6494 61492
rect 6438 60010 6494 60019
rect 6438 59945 6494 59954
rect 6438 58472 6494 58481
rect 6438 58407 6494 58416
rect 6438 56934 6494 56943
rect 6438 56869 6494 56878
rect 6438 55396 6494 55405
rect 6438 55331 6494 55340
rect 6438 53858 6494 53867
rect 6438 53793 6494 53802
rect 6438 52320 6494 52329
rect 6438 52255 6494 52264
rect 6438 50782 6494 50791
rect 6438 50717 6494 50726
rect 6438 49244 6494 49253
rect 6438 49179 6494 49188
rect 6438 47706 6494 47715
rect 6438 47641 6494 47650
rect 6438 46168 6494 46177
rect 6438 46103 6494 46112
rect 6438 44630 6494 44639
rect 6438 44565 6494 44574
rect 6438 43092 6494 43101
rect 6438 43027 6494 43036
rect 6438 41554 6494 41563
rect 6438 41489 6494 41498
rect 6438 40016 6494 40025
rect 6438 39951 6494 39960
rect 6438 38478 6494 38487
rect 6438 38413 6494 38422
rect 6438 36940 6494 36949
rect 6438 36875 6494 36884
rect 4860 35440 4916 35449
rect 4860 35375 4916 35384
rect 6438 35402 6494 35411
rect 4776 33900 4832 33909
rect 4776 33835 4832 33844
rect 4692 32360 4748 32369
rect 4692 32295 4748 32304
rect 4608 30820 4664 30829
rect 4608 30755 4664 30764
rect 4524 29280 4580 29289
rect 4524 29215 4580 29224
rect 4440 27740 4496 27749
rect 4440 27675 4496 27684
rect 4358 27328 4410 27334
rect 4358 27270 4410 27276
rect 4370 27076 4398 27270
rect 4358 27070 4410 27076
rect 4358 27012 4410 27018
rect 4370 26818 4398 27012
rect 4358 26812 4410 26818
rect 4358 26754 4410 26760
rect 4370 26209 4398 26754
rect 4356 26200 4412 26209
rect 4356 26135 4412 26144
rect 4370 25538 4398 26135
rect 4358 25532 4410 25538
rect 4358 25474 4410 25480
rect 4370 25280 4398 25474
rect 4358 25274 4410 25280
rect 4358 25216 4410 25222
rect 4370 25022 4398 25216
rect 4358 25016 4410 25022
rect 4358 24958 4410 24964
rect 4272 24660 4328 24669
rect 4272 24595 4328 24604
rect 4188 20044 4244 20053
rect 4188 19979 4244 19988
rect 4104 18504 4160 18513
rect 4104 18439 4160 18448
rect 4020 16964 4076 16973
rect 4020 16899 4076 16908
rect 3936 15424 3992 15433
rect 3936 15359 3992 15368
rect 3852 13884 3908 13893
rect 3852 13819 3908 13828
rect 3768 12344 3824 12353
rect 3768 12279 3824 12288
rect 3684 10804 3740 10813
rect 3684 10739 3740 10748
rect 3600 9264 3656 9273
rect 3600 9199 3656 9208
rect 3518 8442 3570 8448
rect 3518 8384 3570 8390
rect 3434 8184 3486 8190
rect 3434 8126 3486 8132
rect 3350 6732 3402 6738
rect 3350 6674 3402 6680
rect 3362 5372 3390 6674
rect 3446 5630 3474 8126
rect 3530 7254 3558 8384
rect 3518 7248 3570 7254
rect 3518 7190 3570 7196
rect 3434 5624 3486 5630
rect 3434 5566 3486 5572
rect 3350 5366 3402 5372
rect 3350 5308 3402 5314
rect 3266 5108 3318 5114
rect 3266 5050 3318 5056
rect 3011 3836 3067 3845
rect 3011 3771 3067 3780
rect 3278 2554 3306 5050
rect 3362 4178 3390 5308
rect 3350 4172 3402 4178
rect 3350 4114 3402 4120
rect 3266 2548 3318 2554
rect 3266 2490 3318 2496
rect 1306 2378 1358 2384
rect 1306 2320 1358 2326
rect 3011 2380 3067 2389
rect 3011 2315 3067 2324
rect 3278 844 3306 2490
rect 3362 1577 3390 4114
rect 3446 3920 3474 5566
rect 3530 4657 3558 7190
rect 3516 4648 3572 4657
rect 3516 4583 3572 4592
rect 3434 3914 3486 3920
rect 3434 3856 3486 3862
rect 3446 3117 3474 3856
rect 3530 3662 3558 4583
rect 3518 3656 3570 3662
rect 3518 3598 3570 3604
rect 3432 3108 3488 3117
rect 3432 3043 3488 3052
rect 3446 2038 3474 3043
rect 3530 2296 3558 3598
rect 3614 2382 3642 9199
rect 3698 4092 3726 10739
rect 3782 7168 3810 12279
rect 3866 8534 3894 13819
rect 3950 10244 3978 15359
rect 4034 13320 4062 16899
rect 4118 14686 4146 18439
rect 4202 16396 4230 19979
rect 4190 16390 4242 16396
rect 4190 16332 4242 16338
rect 4202 16138 4230 16332
rect 4286 16310 4314 24595
rect 4370 24258 4398 24958
rect 4358 24252 4410 24258
rect 4358 24194 4410 24200
rect 4370 24000 4398 24194
rect 4358 23994 4410 24000
rect 4358 23936 4410 23942
rect 4370 23742 4398 23936
rect 4358 23736 4410 23742
rect 4358 23678 4410 23684
rect 4370 22462 4398 23678
rect 4358 22456 4410 22462
rect 4358 22398 4410 22404
rect 4370 22204 4398 22398
rect 4358 22198 4410 22204
rect 4358 22140 4410 22146
rect 4370 21946 4398 22140
rect 4358 21940 4410 21946
rect 4358 21882 4410 21888
rect 4370 21182 4398 21882
rect 4358 21176 4410 21182
rect 4358 21118 4410 21124
rect 4370 20924 4398 21118
rect 4358 20918 4410 20924
rect 4358 20860 4410 20866
rect 4370 20666 4398 20860
rect 4358 20660 4410 20666
rect 4358 20602 4410 20608
rect 4370 19386 4398 20602
rect 4358 19380 4410 19386
rect 4358 19322 4410 19328
rect 4370 19128 4398 19322
rect 4358 19122 4410 19128
rect 4358 19064 4410 19070
rect 4370 18870 4398 19064
rect 4358 18864 4410 18870
rect 4358 18806 4410 18812
rect 4370 18106 4398 18806
rect 4358 18100 4410 18106
rect 4358 18042 4410 18048
rect 4370 17848 4398 18042
rect 4358 17842 4410 17848
rect 4358 17784 4410 17790
rect 4370 17590 4398 17784
rect 4358 17584 4410 17590
rect 4358 17526 4410 17532
rect 4274 16304 4326 16310
rect 4274 16246 4326 16252
rect 4190 16132 4242 16138
rect 4190 16074 4242 16080
rect 4202 15880 4230 16074
rect 4286 16052 4314 16246
rect 4274 16046 4326 16052
rect 4274 15988 4326 15994
rect 4190 15874 4242 15880
rect 4190 15816 4242 15822
rect 4202 14944 4230 15816
rect 4286 15794 4314 15988
rect 4274 15788 4326 15794
rect 4274 15730 4326 15736
rect 4286 15030 4314 15730
rect 4274 15024 4326 15030
rect 4274 14966 4326 14972
rect 4190 14938 4242 14944
rect 4190 14880 4242 14886
rect 4106 14680 4158 14686
rect 4106 14622 4158 14628
rect 4118 14428 4146 14622
rect 4106 14422 4158 14428
rect 4106 14364 4158 14370
rect 4022 13314 4074 13320
rect 4022 13256 4074 13262
rect 4034 11868 4062 13256
rect 4118 13062 4146 14364
rect 4106 13056 4158 13062
rect 4106 12998 4158 13004
rect 4118 12804 4146 12998
rect 4106 12798 4158 12804
rect 4106 12740 4158 12746
rect 4022 11862 4074 11868
rect 4022 11804 4074 11810
rect 4034 11610 4062 11804
rect 4022 11604 4074 11610
rect 4022 11546 4074 11552
rect 4034 11352 4062 11546
rect 4022 11346 4074 11352
rect 4022 11288 4074 11294
rect 3938 10238 3990 10244
rect 3938 10180 3990 10186
rect 3950 9986 3978 10180
rect 3938 9980 3990 9986
rect 3938 9922 3990 9928
rect 3950 9728 3978 9922
rect 3938 9722 3990 9728
rect 3938 9664 3990 9670
rect 3950 8792 3978 9664
rect 3938 8786 3990 8792
rect 3938 8728 3990 8734
rect 3854 8528 3906 8534
rect 3854 8470 3906 8476
rect 3866 8276 3894 8470
rect 3854 8270 3906 8276
rect 3854 8212 3906 8218
rect 3770 7162 3822 7168
rect 3770 7104 3822 7110
rect 3782 5716 3810 7104
rect 3866 6910 3894 8212
rect 3854 6904 3906 6910
rect 3854 6846 3906 6852
rect 3866 6652 3894 6846
rect 3854 6646 3906 6652
rect 3854 6588 3906 6594
rect 3770 5710 3822 5716
rect 3770 5652 3822 5658
rect 3782 5458 3810 5652
rect 3770 5452 3822 5458
rect 3770 5394 3822 5400
rect 3782 5200 3810 5394
rect 3770 5194 3822 5200
rect 3770 5136 3822 5142
rect 3686 4086 3738 4092
rect 3686 4028 3738 4034
rect 3698 3834 3726 4028
rect 3686 3828 3738 3834
rect 3686 3770 3738 3776
rect 3698 3576 3726 3770
rect 3686 3570 3738 3576
rect 3686 3512 3738 3518
rect 3698 2640 3726 3512
rect 3686 2634 3738 2640
rect 3686 2576 3738 2582
rect 3602 2376 3654 2382
rect 3602 2318 3654 2324
rect 3518 2290 3570 2296
rect 3518 2232 3570 2238
rect 3434 2032 3486 2038
rect 3434 1974 3486 1980
rect 3348 1568 3404 1577
rect 3348 1503 3404 1512
rect 3266 838 3318 844
rect 3266 780 3318 786
rect 1222 754 1274 760
rect 1222 696 1274 702
rect 3011 756 3067 765
rect 3011 691 3067 700
rect 3278 37 3306 780
rect 3362 586 3390 1503
rect 3350 580 3402 586
rect 3350 522 3402 528
rect 3264 28 3320 37
rect 3362 0 3390 522
rect 3446 0 3474 1974
rect 3530 0 3558 2232
rect 3614 2124 3642 2318
rect 3602 2118 3654 2124
rect 3602 2060 3654 2066
rect 3614 758 3642 2060
rect 3602 752 3654 758
rect 3602 694 3654 700
rect 3614 500 3642 694
rect 3602 494 3654 500
rect 3602 436 3654 442
rect 3614 0 3642 436
rect 3698 0 3726 2576
rect 3782 0 3810 5136
rect 3866 0 3894 6588
rect 3950 0 3978 8728
rect 4034 0 4062 11288
rect 4118 0 4146 12740
rect 4202 0 4230 14880
rect 4286 14772 4314 14966
rect 4274 14766 4326 14772
rect 4274 14708 4326 14714
rect 4286 14514 4314 14708
rect 4274 14508 4326 14514
rect 4274 14450 4326 14456
rect 4286 13234 4314 14450
rect 4274 13228 4326 13234
rect 4274 13170 4326 13176
rect 4286 12976 4314 13170
rect 4274 12970 4326 12976
rect 4274 12912 4326 12918
rect 4286 12718 4314 12912
rect 4274 12712 4326 12718
rect 4274 12654 4326 12660
rect 4286 11954 4314 12654
rect 4274 11948 4326 11954
rect 4274 11890 4326 11896
rect 4286 11696 4314 11890
rect 4274 11690 4326 11696
rect 4274 11632 4326 11638
rect 4286 11438 4314 11632
rect 4274 11432 4326 11438
rect 4274 11374 4326 11380
rect 4286 10158 4314 11374
rect 4274 10152 4326 10158
rect 4274 10094 4326 10100
rect 4286 9900 4314 10094
rect 4274 9894 4326 9900
rect 4274 9836 4326 9842
rect 4286 9642 4314 9836
rect 4274 9636 4326 9642
rect 4274 9578 4326 9584
rect 4286 8878 4314 9578
rect 4274 8872 4326 8878
rect 4274 8814 4326 8820
rect 4286 8620 4314 8814
rect 4274 8614 4326 8620
rect 4274 8556 4326 8562
rect 4286 8362 4314 8556
rect 4274 8356 4326 8362
rect 4274 8298 4326 8304
rect 4286 7082 4314 8298
rect 4274 7076 4326 7082
rect 4274 7018 4326 7024
rect 4286 6824 4314 7018
rect 4274 6818 4326 6824
rect 4274 6760 4326 6766
rect 4286 6566 4314 6760
rect 4274 6560 4326 6566
rect 4274 6502 4326 6508
rect 4286 5802 4314 6502
rect 4274 5796 4326 5802
rect 4274 5738 4326 5744
rect 4286 5544 4314 5738
rect 4274 5538 4326 5544
rect 4274 5480 4326 5486
rect 4286 5286 4314 5480
rect 4274 5280 4326 5286
rect 4274 5222 4326 5228
rect 4286 4006 4314 5222
rect 4274 4000 4326 4006
rect 4274 3942 4326 3948
rect 4286 3748 4314 3942
rect 4274 3742 4326 3748
rect 4274 3684 4326 3690
rect 4286 3490 4314 3684
rect 4274 3484 4326 3490
rect 4274 3426 4326 3432
rect 4286 2726 4314 3426
rect 4274 2720 4326 2726
rect 4274 2662 4326 2668
rect 4286 2468 4314 2662
rect 4274 2462 4326 2468
rect 4274 2404 4326 2410
rect 4286 2210 4314 2404
rect 4274 2204 4326 2210
rect 4274 2146 4326 2152
rect 4286 672 4314 2146
rect 4274 666 4326 672
rect 4274 608 4326 614
rect 4286 414 4314 608
rect 4274 408 4326 414
rect 4274 350 4326 356
rect 4286 0 4314 350
rect 4370 0 4398 17526
rect 4454 0 4482 27675
rect 4538 0 4566 29215
rect 4622 0 4650 30755
rect 4706 0 4734 32295
rect 4790 0 4818 33835
rect 4874 0 4902 35375
rect 6438 35337 6494 35346
rect 6438 33864 6494 33873
rect 6438 33799 6494 33808
rect 6438 32326 6494 32335
rect 6438 32261 6494 32270
rect 6438 30788 6494 30797
rect 6438 30723 6494 30732
rect 6438 29250 6494 29259
rect 6438 29185 6494 29194
rect 6438 27712 6494 27721
rect 6438 27647 6494 27656
rect 6438 26174 6494 26183
rect 6438 26109 6494 26118
rect 6438 24636 6494 24645
rect 6438 24571 6494 24580
rect 6438 23098 6494 23107
rect 6438 23033 6494 23042
rect 6438 21560 6494 21569
rect 6438 21495 6494 21504
rect 6438 20022 6494 20031
rect 6438 19957 6494 19966
rect 6438 18484 6494 18493
rect 6438 18419 6494 18428
rect 6438 16946 6494 16955
rect 6438 16881 6494 16890
rect 6438 15408 6494 15417
rect 6438 15343 6494 15352
rect 6438 13870 6494 13879
rect 6438 13805 6494 13814
rect 6438 12332 6494 12341
rect 6438 12267 6494 12276
rect 6438 10794 6494 10803
rect 6438 10729 6494 10738
rect 6438 9256 6494 9265
rect 6438 9191 6494 9200
rect 6438 7718 6494 7727
rect 6438 7653 6494 7662
rect 6438 6180 6494 6189
rect 6438 6115 6494 6124
rect 6438 4642 6494 4651
rect 6438 4577 6494 4586
rect 6438 3104 6494 3113
rect 6438 3039 6494 3048
rect 6438 1566 6494 1575
rect 6438 1501 6494 1510
rect 6438 28 6494 37
rect 3264 -37 3320 -28
rect 6438 -37 6494 -28
<< via2 >>
rect 3011 36250 3067 36252
rect 3011 36198 3013 36250
rect 3013 36198 3065 36250
rect 3065 36198 3067 36250
rect 3011 36196 3067 36198
rect 3011 34626 3067 34628
rect 3011 34574 3013 34626
rect 3013 34574 3065 34626
rect 3065 34574 3067 34626
rect 3011 34572 3067 34574
rect 3011 33170 3067 33172
rect 3011 33118 3013 33170
rect 3013 33118 3065 33170
rect 3065 33118 3067 33170
rect 3011 33116 3067 33118
rect 3011 31546 3067 31548
rect 3011 31494 3013 31546
rect 3013 31494 3065 31546
rect 3065 31494 3067 31546
rect 3011 31492 3067 31494
rect 3011 30090 3067 30092
rect 3011 30038 3013 30090
rect 3013 30038 3065 30090
rect 3065 30038 3067 30090
rect 3011 30036 3067 30038
rect 3011 28466 3067 28468
rect 3011 28414 3013 28466
rect 3013 28414 3065 28466
rect 3065 28414 3067 28466
rect 3011 28412 3067 28414
rect 3011 27010 3067 27012
rect 3011 26958 3013 27010
rect 3013 26958 3065 27010
rect 3065 26958 3067 27010
rect 3011 26956 3067 26958
rect 3011 25386 3067 25388
rect 3011 25334 3013 25386
rect 3013 25334 3065 25386
rect 3065 25334 3067 25386
rect 3011 25332 3067 25334
rect 3011 20854 3067 20856
rect 3011 20802 3013 20854
rect 3013 20802 3065 20854
rect 3065 20802 3067 20854
rect 3011 20800 3067 20802
rect 3011 19230 3067 19232
rect 3011 19178 3013 19230
rect 3013 19178 3065 19230
rect 3065 19178 3067 19230
rect 3011 19176 3067 19178
rect 3011 17774 3067 17776
rect 3011 17722 3013 17774
rect 3013 17722 3065 17774
rect 3065 17722 3067 17774
rect 3011 17720 3067 17722
rect 3011 16150 3067 16152
rect 3011 16098 3013 16150
rect 3013 16098 3065 16150
rect 3065 16098 3067 16150
rect 3011 16096 3067 16098
rect 3011 14694 3067 14696
rect 3011 14642 3013 14694
rect 3013 14642 3065 14694
rect 3065 14642 3067 14694
rect 3011 14640 3067 14642
rect 3011 13070 3067 13072
rect 3011 13018 3013 13070
rect 3013 13018 3065 13070
rect 3065 13018 3067 13070
rect 3011 13016 3067 13018
rect 3011 11614 3067 11616
rect 3011 11562 3013 11614
rect 3013 11562 3065 11614
rect 3065 11562 3067 11614
rect 3011 11560 3067 11562
rect 3011 9990 3067 9992
rect 3011 9938 3013 9990
rect 3013 9938 3065 9990
rect 3065 9938 3067 9990
rect 3011 9936 3067 9938
rect 3011 5458 3067 5460
rect 3011 5406 3013 5458
rect 3013 5406 3065 5458
rect 3065 5406 3067 5458
rect 3011 5404 3067 5406
rect 6438 98458 6494 98460
rect 6438 98406 6440 98458
rect 6440 98406 6492 98458
rect 6492 98406 6494 98458
rect 6438 98404 6494 98406
rect 6438 96920 6494 96922
rect 6438 96868 6440 96920
rect 6440 96868 6492 96920
rect 6492 96868 6494 96920
rect 6438 96866 6494 96868
rect 6438 95382 6494 95384
rect 6438 95330 6440 95382
rect 6440 95330 6492 95382
rect 6492 95330 6494 95382
rect 6438 95328 6494 95330
rect 6438 93844 6494 93846
rect 6438 93792 6440 93844
rect 6440 93792 6492 93844
rect 6492 93792 6494 93844
rect 6438 93790 6494 93792
rect 6438 92306 6494 92308
rect 6438 92254 6440 92306
rect 6440 92254 6492 92306
rect 6492 92254 6494 92306
rect 6438 92252 6494 92254
rect 6438 90768 6494 90770
rect 6438 90716 6440 90768
rect 6440 90716 6492 90768
rect 6492 90716 6494 90768
rect 6438 90714 6494 90716
rect 6438 89230 6494 89232
rect 6438 89178 6440 89230
rect 6440 89178 6492 89230
rect 6492 89178 6494 89230
rect 6438 89176 6494 89178
rect 6438 87692 6494 87694
rect 6438 87640 6440 87692
rect 6440 87640 6492 87692
rect 6492 87640 6494 87692
rect 6438 87638 6494 87640
rect 6438 86154 6494 86156
rect 6438 86102 6440 86154
rect 6440 86102 6492 86154
rect 6492 86102 6494 86154
rect 6438 86100 6494 86102
rect 6438 84616 6494 84618
rect 6438 84564 6440 84616
rect 6440 84564 6492 84616
rect 6492 84564 6494 84616
rect 6438 84562 6494 84564
rect 6438 83078 6494 83080
rect 6438 83026 6440 83078
rect 6440 83026 6492 83078
rect 6492 83026 6494 83078
rect 6438 83024 6494 83026
rect 6438 81540 6494 81542
rect 6438 81488 6440 81540
rect 6440 81488 6492 81540
rect 6492 81488 6494 81540
rect 6438 81486 6494 81488
rect 6438 80002 6494 80004
rect 6438 79950 6440 80002
rect 6440 79950 6492 80002
rect 6492 79950 6494 80002
rect 6438 79948 6494 79950
rect 6438 78464 6494 78466
rect 6438 78412 6440 78464
rect 6440 78412 6492 78464
rect 6492 78412 6494 78464
rect 6438 78410 6494 78412
rect 6438 76926 6494 76928
rect 6438 76874 6440 76926
rect 6440 76874 6492 76926
rect 6492 76874 6494 76926
rect 6438 76872 6494 76874
rect 6438 75388 6494 75390
rect 6438 75336 6440 75388
rect 6440 75336 6492 75388
rect 6492 75336 6494 75388
rect 6438 75334 6494 75336
rect 6438 73850 6494 73852
rect 6438 73798 6440 73850
rect 6440 73798 6492 73850
rect 6492 73798 6494 73850
rect 6438 73796 6494 73798
rect 6438 72312 6494 72314
rect 6438 72260 6440 72312
rect 6440 72260 6492 72312
rect 6492 72260 6494 72312
rect 6438 72258 6494 72260
rect 6438 70774 6494 70776
rect 6438 70722 6440 70774
rect 6440 70722 6492 70774
rect 6492 70722 6494 70774
rect 6438 70720 6494 70722
rect 6438 69236 6494 69238
rect 6438 69184 6440 69236
rect 6440 69184 6492 69236
rect 6492 69184 6494 69236
rect 6438 69182 6494 69184
rect 6438 67698 6494 67700
rect 6438 67646 6440 67698
rect 6440 67646 6492 67698
rect 6492 67646 6494 67698
rect 6438 67644 6494 67646
rect 6438 66160 6494 66162
rect 6438 66108 6440 66160
rect 6440 66108 6492 66160
rect 6492 66108 6494 66160
rect 6438 66106 6494 66108
rect 6438 64622 6494 64624
rect 6438 64570 6440 64622
rect 6440 64570 6492 64622
rect 6492 64570 6494 64622
rect 6438 64568 6494 64570
rect 6438 63084 6494 63086
rect 6438 63032 6440 63084
rect 6440 63032 6492 63084
rect 6492 63032 6494 63084
rect 6438 63030 6494 63032
rect 6438 61546 6494 61548
rect 6438 61494 6440 61546
rect 6440 61494 6492 61546
rect 6492 61494 6494 61546
rect 6438 61492 6494 61494
rect 6438 60008 6494 60010
rect 6438 59956 6440 60008
rect 6440 59956 6492 60008
rect 6492 59956 6494 60008
rect 6438 59954 6494 59956
rect 6438 58470 6494 58472
rect 6438 58418 6440 58470
rect 6440 58418 6492 58470
rect 6492 58418 6494 58470
rect 6438 58416 6494 58418
rect 6438 56932 6494 56934
rect 6438 56880 6440 56932
rect 6440 56880 6492 56932
rect 6492 56880 6494 56932
rect 6438 56878 6494 56880
rect 6438 55394 6494 55396
rect 6438 55342 6440 55394
rect 6440 55342 6492 55394
rect 6492 55342 6494 55394
rect 6438 55340 6494 55342
rect 6438 53856 6494 53858
rect 6438 53804 6440 53856
rect 6440 53804 6492 53856
rect 6492 53804 6494 53856
rect 6438 53802 6494 53804
rect 6438 52318 6494 52320
rect 6438 52266 6440 52318
rect 6440 52266 6492 52318
rect 6492 52266 6494 52318
rect 6438 52264 6494 52266
rect 6438 50780 6494 50782
rect 6438 50728 6440 50780
rect 6440 50728 6492 50780
rect 6492 50728 6494 50780
rect 6438 50726 6494 50728
rect 6438 49242 6494 49244
rect 6438 49190 6440 49242
rect 6440 49190 6492 49242
rect 6492 49190 6494 49242
rect 6438 49188 6494 49190
rect 6438 47704 6494 47706
rect 6438 47652 6440 47704
rect 6440 47652 6492 47704
rect 6492 47652 6494 47704
rect 6438 47650 6494 47652
rect 6438 46166 6494 46168
rect 6438 46114 6440 46166
rect 6440 46114 6492 46166
rect 6492 46114 6494 46166
rect 6438 46112 6494 46114
rect 6438 44628 6494 44630
rect 6438 44576 6440 44628
rect 6440 44576 6492 44628
rect 6492 44576 6494 44628
rect 6438 44574 6494 44576
rect 6438 43090 6494 43092
rect 6438 43038 6440 43090
rect 6440 43038 6492 43090
rect 6492 43038 6494 43090
rect 6438 43036 6494 43038
rect 6438 41552 6494 41554
rect 6438 41500 6440 41552
rect 6440 41500 6492 41552
rect 6492 41500 6494 41552
rect 6438 41498 6494 41500
rect 6438 40014 6494 40016
rect 6438 39962 6440 40014
rect 6440 39962 6492 40014
rect 6492 39962 6494 40014
rect 6438 39960 6494 39962
rect 6438 38476 6494 38478
rect 6438 38424 6440 38476
rect 6440 38424 6492 38476
rect 6492 38424 6494 38476
rect 6438 38422 6494 38424
rect 6438 36938 6494 36940
rect 6438 36886 6440 36938
rect 6440 36886 6492 36938
rect 6492 36886 6494 36938
rect 6438 36884 6494 36886
rect 4860 35384 4916 35440
rect 6438 35400 6494 35402
rect 4776 33844 4832 33900
rect 4692 32304 4748 32360
rect 4608 30764 4664 30820
rect 4524 29224 4580 29280
rect 4440 27684 4496 27740
rect 4356 26144 4412 26200
rect 4272 24604 4328 24660
rect 4188 19988 4244 20044
rect 4104 18448 4160 18504
rect 4020 16908 4076 16964
rect 3936 15368 3992 15424
rect 3852 13828 3908 13884
rect 3768 12288 3824 12344
rect 3684 10748 3740 10804
rect 3600 9208 3656 9264
rect 3011 3834 3067 3836
rect 3011 3782 3013 3834
rect 3013 3782 3065 3834
rect 3065 3782 3067 3834
rect 3011 3780 3067 3782
rect 3011 2378 3067 2380
rect 3011 2326 3013 2378
rect 3013 2326 3065 2378
rect 3065 2326 3067 2378
rect 3011 2324 3067 2326
rect 3516 4592 3572 4648
rect 3432 3052 3488 3108
rect 3348 1512 3404 1568
rect 3011 754 3067 756
rect 3011 702 3013 754
rect 3013 702 3065 754
rect 3065 702 3067 754
rect 3011 700 3067 702
rect 3264 -28 3320 28
rect 6438 35348 6440 35400
rect 6440 35348 6492 35400
rect 6492 35348 6494 35400
rect 6438 35346 6494 35348
rect 6438 33862 6494 33864
rect 6438 33810 6440 33862
rect 6440 33810 6492 33862
rect 6492 33810 6494 33862
rect 6438 33808 6494 33810
rect 6438 32324 6494 32326
rect 6438 32272 6440 32324
rect 6440 32272 6492 32324
rect 6492 32272 6494 32324
rect 6438 32270 6494 32272
rect 6438 30786 6494 30788
rect 6438 30734 6440 30786
rect 6440 30734 6492 30786
rect 6492 30734 6494 30786
rect 6438 30732 6494 30734
rect 6438 29248 6494 29250
rect 6438 29196 6440 29248
rect 6440 29196 6492 29248
rect 6492 29196 6494 29248
rect 6438 29194 6494 29196
rect 6438 27710 6494 27712
rect 6438 27658 6440 27710
rect 6440 27658 6492 27710
rect 6492 27658 6494 27710
rect 6438 27656 6494 27658
rect 6438 26172 6494 26174
rect 6438 26120 6440 26172
rect 6440 26120 6492 26172
rect 6492 26120 6494 26172
rect 6438 26118 6494 26120
rect 6438 24634 6494 24636
rect 6438 24582 6440 24634
rect 6440 24582 6492 24634
rect 6492 24582 6494 24634
rect 6438 24580 6494 24582
rect 6438 23096 6494 23098
rect 6438 23044 6440 23096
rect 6440 23044 6492 23096
rect 6492 23044 6494 23096
rect 6438 23042 6494 23044
rect 6438 21558 6494 21560
rect 6438 21506 6440 21558
rect 6440 21506 6492 21558
rect 6492 21506 6494 21558
rect 6438 21504 6494 21506
rect 6438 20020 6494 20022
rect 6438 19968 6440 20020
rect 6440 19968 6492 20020
rect 6492 19968 6494 20020
rect 6438 19966 6494 19968
rect 6438 18482 6494 18484
rect 6438 18430 6440 18482
rect 6440 18430 6492 18482
rect 6492 18430 6494 18482
rect 6438 18428 6494 18430
rect 6438 16944 6494 16946
rect 6438 16892 6440 16944
rect 6440 16892 6492 16944
rect 6492 16892 6494 16944
rect 6438 16890 6494 16892
rect 6438 15406 6494 15408
rect 6438 15354 6440 15406
rect 6440 15354 6492 15406
rect 6492 15354 6494 15406
rect 6438 15352 6494 15354
rect 6438 13868 6494 13870
rect 6438 13816 6440 13868
rect 6440 13816 6492 13868
rect 6492 13816 6494 13868
rect 6438 13814 6494 13816
rect 6438 12330 6494 12332
rect 6438 12278 6440 12330
rect 6440 12278 6492 12330
rect 6492 12278 6494 12330
rect 6438 12276 6494 12278
rect 6438 10792 6494 10794
rect 6438 10740 6440 10792
rect 6440 10740 6492 10792
rect 6492 10740 6494 10792
rect 6438 10738 6494 10740
rect 6438 9254 6494 9256
rect 6438 9202 6440 9254
rect 6440 9202 6492 9254
rect 6492 9202 6494 9254
rect 6438 9200 6494 9202
rect 6438 7716 6494 7718
rect 6438 7664 6440 7716
rect 6440 7664 6492 7716
rect 6492 7664 6494 7716
rect 6438 7662 6494 7664
rect 6438 6178 6494 6180
rect 6438 6126 6440 6178
rect 6440 6126 6492 6178
rect 6492 6126 6494 6178
rect 6438 6124 6494 6126
rect 6438 4640 6494 4642
rect 6438 4588 6440 4640
rect 6440 4588 6492 4640
rect 6492 4588 6494 4640
rect 6438 4586 6494 4588
rect 6438 3102 6494 3104
rect 6438 3050 6440 3102
rect 6440 3050 6492 3102
rect 6492 3050 6494 3102
rect 6438 3048 6494 3050
rect 6438 1564 6494 1566
rect 6438 1512 6440 1564
rect 6440 1512 6492 1564
rect 6492 1512 6494 1564
rect 6438 1510 6494 1512
rect 6438 26 6494 28
rect 6438 -26 6440 26
rect 6440 -26 6492 26
rect 6492 -26 6494 26
rect 6438 -28 6494 -26
<< metal3 >>
rect 6400 98460 6532 98469
rect 6400 98404 6438 98460
rect 6494 98404 6532 98460
rect 6400 98395 6532 98404
rect 6400 96922 6532 96931
rect 6400 96866 6438 96922
rect 6494 96866 6532 96922
rect 6400 96857 6532 96866
rect 6400 95384 6532 95393
rect 6400 95328 6438 95384
rect 6494 95328 6532 95384
rect 6400 95319 6532 95328
rect 6400 93846 6532 93855
rect 6400 93790 6438 93846
rect 6494 93790 6532 93846
rect 6400 93781 6532 93790
rect 6400 92308 6532 92317
rect 6400 92252 6438 92308
rect 6494 92252 6532 92308
rect 6400 92243 6532 92252
rect 6400 90770 6532 90779
rect 6400 90714 6438 90770
rect 6494 90714 6532 90770
rect 6400 90705 6532 90714
rect 6400 89232 6532 89241
rect 6400 89176 6438 89232
rect 6494 89176 6532 89232
rect 6400 89167 6532 89176
rect 6400 87694 6532 87703
rect 6400 87638 6438 87694
rect 6494 87638 6532 87694
rect 6400 87629 6532 87638
rect 6400 86156 6532 86165
rect 6400 86100 6438 86156
rect 6494 86100 6532 86156
rect 6400 86091 6532 86100
rect 6400 84618 6532 84627
rect 6400 84562 6438 84618
rect 6494 84562 6532 84618
rect 6400 84553 6532 84562
rect 6400 83080 6532 83089
rect 6400 83024 6438 83080
rect 6494 83024 6532 83080
rect 6400 83015 6532 83024
rect 6400 81542 6532 81551
rect 6400 81486 6438 81542
rect 6494 81486 6532 81542
rect 6400 81477 6532 81486
rect 6400 80004 6532 80013
rect 6400 79948 6438 80004
rect 6494 79948 6532 80004
rect 6400 79939 6532 79948
rect 6400 78466 6532 78475
rect 6400 78410 6438 78466
rect 6494 78410 6532 78466
rect 6400 78401 6532 78410
rect 6400 76928 6532 76937
rect 6400 76872 6438 76928
rect 6494 76872 6532 76928
rect 6400 76863 6532 76872
rect 6400 75390 6532 75399
rect 6400 75334 6438 75390
rect 6494 75334 6532 75390
rect 6400 75325 6532 75334
rect 6400 73852 6532 73861
rect 6400 73796 6438 73852
rect 6494 73796 6532 73852
rect 6400 73787 6532 73796
rect 6400 72314 6532 72323
rect 6400 72258 6438 72314
rect 6494 72258 6532 72314
rect 6400 72249 6532 72258
rect 6400 70776 6532 70785
rect 6400 70720 6438 70776
rect 6494 70720 6532 70776
rect 6400 70711 6532 70720
rect 6400 69238 6532 69247
rect 6400 69182 6438 69238
rect 6494 69182 6532 69238
rect 6400 69173 6532 69182
rect 6400 67700 6532 67709
rect 6400 67644 6438 67700
rect 6494 67644 6532 67700
rect 6400 67635 6532 67644
rect 6400 66162 6532 66171
rect 6400 66106 6438 66162
rect 6494 66106 6532 66162
rect 6400 66097 6532 66106
rect 6400 64624 6532 64633
rect 6400 64568 6438 64624
rect 6494 64568 6532 64624
rect 6400 64559 6532 64568
rect 6400 63086 6532 63095
rect 6400 63030 6438 63086
rect 6494 63030 6532 63086
rect 6400 63021 6532 63030
rect 6400 61548 6532 61557
rect 6400 61492 6438 61548
rect 6494 61492 6532 61548
rect 6400 61483 6532 61492
rect 6400 60010 6532 60019
rect 6400 59954 6438 60010
rect 6494 59954 6532 60010
rect 6400 59945 6532 59954
rect 6400 58472 6532 58481
rect 6400 58416 6438 58472
rect 6494 58416 6532 58472
rect 6400 58407 6532 58416
rect 6400 56934 6532 56943
rect 6400 56878 6438 56934
rect 6494 56878 6532 56934
rect 6400 56869 6532 56878
rect 6400 55396 6532 55405
rect 6400 55340 6438 55396
rect 6494 55340 6532 55396
rect 6400 55331 6532 55340
rect 6400 53858 6532 53867
rect 6400 53802 6438 53858
rect 6494 53802 6532 53858
rect 6400 53793 6532 53802
rect 6400 52320 6532 52329
rect 6400 52264 6438 52320
rect 6494 52264 6532 52320
rect 6400 52255 6532 52264
rect 6400 50782 6532 50791
rect 6400 50726 6438 50782
rect 6494 50726 6532 50782
rect 6400 50717 6532 50726
rect 6400 49244 6532 49253
rect 6400 49188 6438 49244
rect 6494 49188 6532 49244
rect 6400 49179 6532 49188
rect 6400 47706 6532 47715
rect 6400 47650 6438 47706
rect 6494 47650 6532 47706
rect 6400 47641 6532 47650
rect 6400 46168 6532 46177
rect 6400 46112 6438 46168
rect 6494 46112 6532 46168
rect 6400 46103 6532 46112
rect 6400 44630 6532 44639
rect 6400 44574 6438 44630
rect 6494 44574 6532 44630
rect 6400 44565 6532 44574
rect 6400 43092 6532 43101
rect 6400 43036 6438 43092
rect 6494 43036 6532 43092
rect 6400 43027 6532 43036
rect 6400 41554 6532 41563
rect 6400 41498 6438 41554
rect 6494 41498 6532 41554
rect 6400 41489 6532 41498
rect 6400 40016 6532 40025
rect 6400 39960 6438 40016
rect 6494 39960 6532 40016
rect 6400 39951 6532 39960
rect 6400 38478 6532 38487
rect 6400 38422 6438 38478
rect 6494 38422 6532 38478
rect 6400 38413 6532 38422
rect 1044 36915 1176 36989
rect 2084 36915 2216 36989
rect 6400 36940 6532 36949
rect 6400 36884 6438 36940
rect 6494 36884 6532 36940
rect 6400 36875 6532 36884
rect 2973 36252 3105 36257
rect 2973 36196 3011 36252
rect 3067 36196 3105 36252
rect 2973 36191 3105 36196
rect 1044 35375 1176 35449
rect 2084 35375 2216 35449
rect 3009 35442 3069 36191
rect 4822 35442 4954 35445
rect 3009 35440 4954 35442
rect 3009 35384 4860 35440
rect 4916 35384 4954 35440
rect 3009 35382 4954 35384
rect 4822 35379 4954 35382
rect 6400 35402 6532 35411
rect 6400 35346 6438 35402
rect 6494 35346 6532 35402
rect 6400 35337 6532 35346
rect 2973 34628 3105 34633
rect 2973 34572 3011 34628
rect 3067 34572 3105 34628
rect 2973 34567 3105 34572
rect 1044 33835 1176 33909
rect 2084 33835 2216 33909
rect 3009 33902 3069 34567
rect 4738 33902 4870 33905
rect 3009 33900 4870 33902
rect 3009 33844 4776 33900
rect 4832 33844 4870 33900
rect 3009 33842 4870 33844
rect 4738 33839 4870 33842
rect 6400 33864 6532 33873
rect 6400 33808 6438 33864
rect 6494 33808 6532 33864
rect 6400 33799 6532 33808
rect 2973 33172 3105 33177
rect 2973 33116 3011 33172
rect 3067 33116 3105 33172
rect 2973 33111 3105 33116
rect 1044 32295 1176 32369
rect 2084 32295 2216 32369
rect 3009 32362 3069 33111
rect 4654 32362 4786 32365
rect 3009 32360 4786 32362
rect 3009 32304 4692 32360
rect 4748 32304 4786 32360
rect 3009 32302 4786 32304
rect 4654 32299 4786 32302
rect 6400 32326 6532 32335
rect 6400 32270 6438 32326
rect 6494 32270 6532 32326
rect 6400 32261 6532 32270
rect 2973 31548 3105 31553
rect 2973 31492 3011 31548
rect 3067 31492 3105 31548
rect 2973 31487 3105 31492
rect 1044 30755 1176 30829
rect 2084 30755 2216 30829
rect 3009 30822 3069 31487
rect 4570 30822 4702 30825
rect 3009 30820 4702 30822
rect 3009 30764 4608 30820
rect 4664 30764 4702 30820
rect 3009 30762 4702 30764
rect 4570 30759 4702 30762
rect 6400 30788 6532 30797
rect 6400 30732 6438 30788
rect 6494 30732 6532 30788
rect 6400 30723 6532 30732
rect 2973 30092 3105 30097
rect 2973 30036 3011 30092
rect 3067 30036 3105 30092
rect 2973 30031 3105 30036
rect 1044 29215 1176 29289
rect 2084 29215 2216 29289
rect 3009 29282 3069 30031
rect 4486 29282 4618 29285
rect 3009 29280 4618 29282
rect 3009 29224 4524 29280
rect 4580 29224 4618 29280
rect 3009 29222 4618 29224
rect 4486 29219 4618 29222
rect 6400 29250 6532 29259
rect 6400 29194 6438 29250
rect 6494 29194 6532 29250
rect 6400 29185 6532 29194
rect 2973 28468 3105 28473
rect 2973 28412 3011 28468
rect 3067 28412 3105 28468
rect 2973 28407 3105 28412
rect 1044 27675 1176 27749
rect 2084 27675 2216 27749
rect 3009 27742 3069 28407
rect 4402 27742 4534 27745
rect 3009 27740 4534 27742
rect 3009 27684 4440 27740
rect 4496 27684 4534 27740
rect 3009 27682 4534 27684
rect 4402 27679 4534 27682
rect 6400 27712 6532 27721
rect 6400 27656 6438 27712
rect 6494 27656 6532 27712
rect 6400 27647 6532 27656
rect 2973 27012 3105 27017
rect 2973 26956 3011 27012
rect 3067 26956 3105 27012
rect 2973 26951 3105 26956
rect 1044 26135 1176 26209
rect 2084 26135 2216 26209
rect 3009 26202 3069 26951
rect 4318 26202 4450 26205
rect 3009 26200 4450 26202
rect 3009 26144 4356 26200
rect 4412 26144 4450 26200
rect 3009 26142 4450 26144
rect 4318 26139 4450 26142
rect 6400 26174 6532 26183
rect 6400 26118 6438 26174
rect 6494 26118 6532 26174
rect 6400 26109 6532 26118
rect 2973 25388 3105 25393
rect 2973 25332 3011 25388
rect 3067 25332 3105 25388
rect 2973 25327 3105 25332
rect 1044 24595 1176 24669
rect 2084 24595 2216 24669
rect 3009 24662 3069 25327
rect 4234 24662 4366 24665
rect 3009 24660 4366 24662
rect 3009 24604 4272 24660
rect 4328 24604 4366 24660
rect 3009 24602 4366 24604
rect 4234 24599 4366 24602
rect 6400 24636 6532 24645
rect 6400 24580 6438 24636
rect 6494 24580 6532 24636
rect 6400 24571 6532 24580
rect 6400 23098 6532 23107
rect 6400 23042 6438 23098
rect 6494 23042 6532 23098
rect 6400 23033 6532 23042
rect 1044 21519 1176 21593
rect 2084 21519 2216 21593
rect 6400 21560 6532 21569
rect 6400 21504 6438 21560
rect 6494 21504 6532 21560
rect 6400 21495 6532 21504
rect 2973 20856 3105 20861
rect 2973 20800 3011 20856
rect 3067 20800 3105 20856
rect 2973 20795 3105 20800
rect 1044 19979 1176 20053
rect 2084 19979 2216 20053
rect 3009 20046 3069 20795
rect 4150 20046 4282 20049
rect 3009 20044 4282 20046
rect 3009 19988 4188 20044
rect 4244 19988 4282 20044
rect 3009 19986 4282 19988
rect 4150 19983 4282 19986
rect 6400 20022 6532 20031
rect 6400 19966 6438 20022
rect 6494 19966 6532 20022
rect 6400 19957 6532 19966
rect 2973 19232 3105 19237
rect 2973 19176 3011 19232
rect 3067 19176 3105 19232
rect 2973 19171 3105 19176
rect 1044 18439 1176 18513
rect 2084 18439 2216 18513
rect 3009 18506 3069 19171
rect 4066 18506 4198 18509
rect 3009 18504 4198 18506
rect 3009 18448 4104 18504
rect 4160 18448 4198 18504
rect 3009 18446 4198 18448
rect 4066 18443 4198 18446
rect 6400 18484 6532 18493
rect 6400 18428 6438 18484
rect 6494 18428 6532 18484
rect 6400 18419 6532 18428
rect 2973 17776 3105 17781
rect 2973 17720 3011 17776
rect 3067 17720 3105 17776
rect 2973 17715 3105 17720
rect 1044 16899 1176 16973
rect 2084 16899 2216 16973
rect 3009 16966 3069 17715
rect 3982 16966 4114 16969
rect 3009 16964 4114 16966
rect 3009 16908 4020 16964
rect 4076 16908 4114 16964
rect 3009 16906 4114 16908
rect 3982 16903 4114 16906
rect 6400 16946 6532 16955
rect 6400 16890 6438 16946
rect 6494 16890 6532 16946
rect 6400 16881 6532 16890
rect 2973 16152 3105 16157
rect 2973 16096 3011 16152
rect 3067 16096 3105 16152
rect 2973 16091 3105 16096
rect 1044 15359 1176 15433
rect 2084 15359 2216 15433
rect 3009 15426 3069 16091
rect 3898 15426 4030 15429
rect 3009 15424 4030 15426
rect 3009 15368 3936 15424
rect 3992 15368 4030 15424
rect 3009 15366 4030 15368
rect 3898 15363 4030 15366
rect 6400 15408 6532 15417
rect 6400 15352 6438 15408
rect 6494 15352 6532 15408
rect 6400 15343 6532 15352
rect 2973 14696 3105 14701
rect 2973 14640 3011 14696
rect 3067 14640 3105 14696
rect 2973 14635 3105 14640
rect 1044 13819 1176 13893
rect 2084 13819 2216 13893
rect 3009 13886 3069 14635
rect 3814 13886 3946 13889
rect 3009 13884 3946 13886
rect 3009 13828 3852 13884
rect 3908 13828 3946 13884
rect 3009 13826 3946 13828
rect 3814 13823 3946 13826
rect 6400 13870 6532 13879
rect 6400 13814 6438 13870
rect 6494 13814 6532 13870
rect 6400 13805 6532 13814
rect 2973 13072 3105 13077
rect 2973 13016 3011 13072
rect 3067 13016 3105 13072
rect 2973 13011 3105 13016
rect 1044 12279 1176 12353
rect 2084 12279 2216 12353
rect 3009 12346 3069 13011
rect 3730 12346 3862 12349
rect 3009 12344 3862 12346
rect 3009 12288 3768 12344
rect 3824 12288 3862 12344
rect 3009 12286 3862 12288
rect 3730 12283 3862 12286
rect 6400 12332 6532 12341
rect 6400 12276 6438 12332
rect 6494 12276 6532 12332
rect 6400 12267 6532 12276
rect 2973 11616 3105 11621
rect 2973 11560 3011 11616
rect 3067 11560 3105 11616
rect 2973 11555 3105 11560
rect 1044 10739 1176 10813
rect 2084 10739 2216 10813
rect 3009 10806 3069 11555
rect 3646 10806 3778 10809
rect 3009 10804 3778 10806
rect 3009 10748 3684 10804
rect 3740 10748 3778 10804
rect 3009 10746 3778 10748
rect 3646 10743 3778 10746
rect 6400 10794 6532 10803
rect 6400 10738 6438 10794
rect 6494 10738 6532 10794
rect 6400 10729 6532 10738
rect 2973 9992 3105 9997
rect 2973 9936 3011 9992
rect 3067 9936 3105 9992
rect 2973 9931 3105 9936
rect 1044 9199 1176 9273
rect 2084 9199 2216 9273
rect 3009 9266 3069 9931
rect 3562 9266 3694 9269
rect 3009 9264 3694 9266
rect 3009 9208 3600 9264
rect 3656 9208 3694 9264
rect 3009 9206 3694 9208
rect 3562 9203 3694 9206
rect 6400 9256 6532 9265
rect 6400 9200 6438 9256
rect 6494 9200 6532 9256
rect 6400 9191 6532 9200
rect 6400 7718 6532 7727
rect 6400 7662 6438 7718
rect 6494 7662 6532 7718
rect 6400 7653 6532 7662
rect 1392 6123 1524 6197
rect 2264 6123 2396 6197
rect 6400 6180 6532 6189
rect 6400 6124 6438 6180
rect 6494 6124 6532 6180
rect 6400 6115 6532 6124
rect 2973 5460 3105 5465
rect 2973 5404 3011 5460
rect 3067 5404 3105 5460
rect 2973 5399 3105 5404
rect 1392 4583 1524 4657
rect 2264 4583 2396 4657
rect 3009 4650 3069 5399
rect 3478 4650 3610 4653
rect 3009 4648 3610 4650
rect 3009 4592 3516 4648
rect 3572 4592 3610 4648
rect 3009 4590 3610 4592
rect 3478 4587 3610 4590
rect 6400 4642 6532 4651
rect 6400 4586 6438 4642
rect 6494 4586 6532 4642
rect 6400 4577 6532 4586
rect 2973 3836 3105 3841
rect 2973 3780 3011 3836
rect 3067 3780 3105 3836
rect 2973 3775 3105 3780
rect 1392 3043 1524 3117
rect 2264 3043 2396 3117
rect 3009 3110 3069 3775
rect 3394 3110 3526 3113
rect 3009 3108 3526 3110
rect 3009 3052 3432 3108
rect 3488 3052 3526 3108
rect 3009 3050 3526 3052
rect 3394 3047 3526 3050
rect 6400 3104 6532 3113
rect 6400 3048 6438 3104
rect 6494 3048 6532 3104
rect 6400 3039 6532 3048
rect 2973 2380 3105 2385
rect 2973 2324 3011 2380
rect 3067 2324 3105 2380
rect 2973 2319 3105 2324
rect 1392 1503 1524 1577
rect 2264 1503 2396 1577
rect 3009 1570 3069 2319
rect 3310 1570 3442 1573
rect 3009 1568 3442 1570
rect 3009 1512 3348 1568
rect 3404 1512 3442 1568
rect 3009 1510 3442 1512
rect 3310 1507 3442 1510
rect 6400 1566 6532 1575
rect 6400 1510 6438 1566
rect 6494 1510 6532 1566
rect 6400 1501 6532 1510
rect 2973 756 3105 761
rect 2973 700 3011 756
rect 3067 700 3105 756
rect 2973 695 3105 700
rect 1392 -37 1524 37
rect 2264 -37 2396 37
rect 3009 30 3069 695
rect 3226 30 3358 33
rect 3009 28 3358 30
rect 3009 -28 3264 28
rect 3320 -28 3358 28
rect 3009 -30 3358 -28
rect 3226 -33 3358 -30
rect 6400 28 6532 37
rect 6400 -28 6438 28
rect 6494 -28 6532 28
rect 6400 -37 6532 -28
use contact_18  contact_18_0
timestamp 1644969367
transform 1 0 6400 0 1 98395
box 0 0 1 1
use contact_17  contact_17_0
timestamp 1644969367
transform 1 0 6434 0 1 98400
box 0 0 1 1
use contact_18  contact_18_1
timestamp 1644969367
transform 1 0 6400 0 1 96857
box 0 0 1 1
use contact_17  contact_17_1
timestamp 1644969367
transform 1 0 6434 0 1 96862
box 0 0 1 1
use contact_18  contact_18_2
timestamp 1644969367
transform 1 0 6400 0 1 95319
box 0 0 1 1
use contact_17  contact_17_2
timestamp 1644969367
transform 1 0 6434 0 1 95324
box 0 0 1 1
use contact_18  contact_18_3
timestamp 1644969367
transform 1 0 6400 0 1 96857
box 0 0 1 1
use contact_17  contact_17_3
timestamp 1644969367
transform 1 0 6434 0 1 96862
box 0 0 1 1
use contact_18  contact_18_4
timestamp 1644969367
transform 1 0 6400 0 1 95319
box 0 0 1 1
use contact_17  contact_17_4
timestamp 1644969367
transform 1 0 6434 0 1 95324
box 0 0 1 1
use contact_18  contact_18_5
timestamp 1644969367
transform 1 0 6400 0 1 93781
box 0 0 1 1
use contact_17  contact_17_5
timestamp 1644969367
transform 1 0 6434 0 1 93786
box 0 0 1 1
use contact_18  contact_18_6
timestamp 1644969367
transform 1 0 6400 0 1 92243
box 0 0 1 1
use contact_17  contact_17_6
timestamp 1644969367
transform 1 0 6434 0 1 92248
box 0 0 1 1
use contact_18  contact_18_7
timestamp 1644969367
transform 1 0 6400 0 1 93781
box 0 0 1 1
use contact_17  contact_17_7
timestamp 1644969367
transform 1 0 6434 0 1 93786
box 0 0 1 1
use contact_18  contact_18_8
timestamp 1644969367
transform 1 0 6400 0 1 92243
box 0 0 1 1
use contact_17  contact_17_8
timestamp 1644969367
transform 1 0 6434 0 1 92248
box 0 0 1 1
use contact_18  contact_18_9
timestamp 1644969367
transform 1 0 6400 0 1 90705
box 0 0 1 1
use contact_17  contact_17_9
timestamp 1644969367
transform 1 0 6434 0 1 90710
box 0 0 1 1
use contact_18  contact_18_10
timestamp 1644969367
transform 1 0 6400 0 1 89167
box 0 0 1 1
use contact_17  contact_17_10
timestamp 1644969367
transform 1 0 6434 0 1 89172
box 0 0 1 1
use contact_18  contact_18_11
timestamp 1644969367
transform 1 0 6400 0 1 90705
box 0 0 1 1
use contact_17  contact_17_11
timestamp 1644969367
transform 1 0 6434 0 1 90710
box 0 0 1 1
use contact_18  contact_18_12
timestamp 1644969367
transform 1 0 6400 0 1 89167
box 0 0 1 1
use contact_17  contact_17_12
timestamp 1644969367
transform 1 0 6434 0 1 89172
box 0 0 1 1
use contact_18  contact_18_13
timestamp 1644969367
transform 1 0 6400 0 1 87629
box 0 0 1 1
use contact_17  contact_17_13
timestamp 1644969367
transform 1 0 6434 0 1 87634
box 0 0 1 1
use contact_18  contact_18_14
timestamp 1644969367
transform 1 0 6400 0 1 86091
box 0 0 1 1
use contact_17  contact_17_14
timestamp 1644969367
transform 1 0 6434 0 1 86096
box 0 0 1 1
use contact_18  contact_18_15
timestamp 1644969367
transform 1 0 6400 0 1 87629
box 0 0 1 1
use contact_17  contact_17_15
timestamp 1644969367
transform 1 0 6434 0 1 87634
box 0 0 1 1
use contact_18  contact_18_16
timestamp 1644969367
transform 1 0 6400 0 1 86091
box 0 0 1 1
use contact_17  contact_17_16
timestamp 1644969367
transform 1 0 6434 0 1 86096
box 0 0 1 1
use contact_18  contact_18_17
timestamp 1644969367
transform 1 0 6400 0 1 84553
box 0 0 1 1
use contact_17  contact_17_17
timestamp 1644969367
transform 1 0 6434 0 1 84558
box 0 0 1 1
use contact_18  contact_18_18
timestamp 1644969367
transform 1 0 6400 0 1 83015
box 0 0 1 1
use contact_17  contact_17_18
timestamp 1644969367
transform 1 0 6434 0 1 83020
box 0 0 1 1
use contact_18  contact_18_19
timestamp 1644969367
transform 1 0 6400 0 1 84553
box 0 0 1 1
use contact_17  contact_17_19
timestamp 1644969367
transform 1 0 6434 0 1 84558
box 0 0 1 1
use contact_18  contact_18_20
timestamp 1644969367
transform 1 0 6400 0 1 83015
box 0 0 1 1
use contact_17  contact_17_20
timestamp 1644969367
transform 1 0 6434 0 1 83020
box 0 0 1 1
use contact_18  contact_18_21
timestamp 1644969367
transform 1 0 6400 0 1 81477
box 0 0 1 1
use contact_17  contact_17_21
timestamp 1644969367
transform 1 0 6434 0 1 81482
box 0 0 1 1
use contact_18  contact_18_22
timestamp 1644969367
transform 1 0 6400 0 1 79939
box 0 0 1 1
use contact_17  contact_17_22
timestamp 1644969367
transform 1 0 6434 0 1 79944
box 0 0 1 1
use contact_18  contact_18_23
timestamp 1644969367
transform 1 0 6400 0 1 81477
box 0 0 1 1
use contact_17  contact_17_23
timestamp 1644969367
transform 1 0 6434 0 1 81482
box 0 0 1 1
use contact_18  contact_18_24
timestamp 1644969367
transform 1 0 6400 0 1 79939
box 0 0 1 1
use contact_17  contact_17_24
timestamp 1644969367
transform 1 0 6434 0 1 79944
box 0 0 1 1
use contact_18  contact_18_25
timestamp 1644969367
transform 1 0 6400 0 1 78401
box 0 0 1 1
use contact_17  contact_17_25
timestamp 1644969367
transform 1 0 6434 0 1 78406
box 0 0 1 1
use contact_18  contact_18_26
timestamp 1644969367
transform 1 0 6400 0 1 76863
box 0 0 1 1
use contact_17  contact_17_26
timestamp 1644969367
transform 1 0 6434 0 1 76868
box 0 0 1 1
use contact_18  contact_18_27
timestamp 1644969367
transform 1 0 6400 0 1 78401
box 0 0 1 1
use contact_17  contact_17_27
timestamp 1644969367
transform 1 0 6434 0 1 78406
box 0 0 1 1
use contact_18  contact_18_28
timestamp 1644969367
transform 1 0 6400 0 1 76863
box 0 0 1 1
use contact_17  contact_17_28
timestamp 1644969367
transform 1 0 6434 0 1 76868
box 0 0 1 1
use contact_18  contact_18_29
timestamp 1644969367
transform 1 0 6400 0 1 75325
box 0 0 1 1
use contact_17  contact_17_29
timestamp 1644969367
transform 1 0 6434 0 1 75330
box 0 0 1 1
use contact_18  contact_18_30
timestamp 1644969367
transform 1 0 6400 0 1 73787
box 0 0 1 1
use contact_17  contact_17_30
timestamp 1644969367
transform 1 0 6434 0 1 73792
box 0 0 1 1
use contact_18  contact_18_31
timestamp 1644969367
transform 1 0 6400 0 1 75325
box 0 0 1 1
use contact_17  contact_17_31
timestamp 1644969367
transform 1 0 6434 0 1 75330
box 0 0 1 1
use contact_18  contact_18_32
timestamp 1644969367
transform 1 0 6400 0 1 73787
box 0 0 1 1
use contact_17  contact_17_32
timestamp 1644969367
transform 1 0 6434 0 1 73792
box 0 0 1 1
use contact_18  contact_18_33
timestamp 1644969367
transform 1 0 6400 0 1 72249
box 0 0 1 1
use contact_17  contact_17_33
timestamp 1644969367
transform 1 0 6434 0 1 72254
box 0 0 1 1
use contact_18  contact_18_34
timestamp 1644969367
transform 1 0 6400 0 1 70711
box 0 0 1 1
use contact_17  contact_17_34
timestamp 1644969367
transform 1 0 6434 0 1 70716
box 0 0 1 1
use contact_18  contact_18_35
timestamp 1644969367
transform 1 0 6400 0 1 72249
box 0 0 1 1
use contact_17  contact_17_35
timestamp 1644969367
transform 1 0 6434 0 1 72254
box 0 0 1 1
use contact_18  contact_18_36
timestamp 1644969367
transform 1 0 6400 0 1 70711
box 0 0 1 1
use contact_17  contact_17_36
timestamp 1644969367
transform 1 0 6434 0 1 70716
box 0 0 1 1
use contact_18  contact_18_37
timestamp 1644969367
transform 1 0 6400 0 1 69173
box 0 0 1 1
use contact_17  contact_17_37
timestamp 1644969367
transform 1 0 6434 0 1 69178
box 0 0 1 1
use contact_18  contact_18_38
timestamp 1644969367
transform 1 0 6400 0 1 67635
box 0 0 1 1
use contact_17  contact_17_38
timestamp 1644969367
transform 1 0 6434 0 1 67640
box 0 0 1 1
use contact_18  contact_18_39
timestamp 1644969367
transform 1 0 6400 0 1 69173
box 0 0 1 1
use contact_17  contact_17_39
timestamp 1644969367
transform 1 0 6434 0 1 69178
box 0 0 1 1
use contact_18  contact_18_40
timestamp 1644969367
transform 1 0 6400 0 1 67635
box 0 0 1 1
use contact_17  contact_17_40
timestamp 1644969367
transform 1 0 6434 0 1 67640
box 0 0 1 1
use contact_18  contact_18_41
timestamp 1644969367
transform 1 0 6400 0 1 66097
box 0 0 1 1
use contact_17  contact_17_41
timestamp 1644969367
transform 1 0 6434 0 1 66102
box 0 0 1 1
use contact_18  contact_18_42
timestamp 1644969367
transform 1 0 6400 0 1 64559
box 0 0 1 1
use contact_17  contact_17_42
timestamp 1644969367
transform 1 0 6434 0 1 64564
box 0 0 1 1
use contact_18  contact_18_43
timestamp 1644969367
transform 1 0 6400 0 1 66097
box 0 0 1 1
use contact_17  contact_17_43
timestamp 1644969367
transform 1 0 6434 0 1 66102
box 0 0 1 1
use contact_18  contact_18_44
timestamp 1644969367
transform 1 0 6400 0 1 64559
box 0 0 1 1
use contact_17  contact_17_44
timestamp 1644969367
transform 1 0 6434 0 1 64564
box 0 0 1 1
use contact_18  contact_18_45
timestamp 1644969367
transform 1 0 6400 0 1 63021
box 0 0 1 1
use contact_17  contact_17_45
timestamp 1644969367
transform 1 0 6434 0 1 63026
box 0 0 1 1
use contact_18  contact_18_46
timestamp 1644969367
transform 1 0 6400 0 1 61483
box 0 0 1 1
use contact_17  contact_17_46
timestamp 1644969367
transform 1 0 6434 0 1 61488
box 0 0 1 1
use contact_18  contact_18_47
timestamp 1644969367
transform 1 0 6400 0 1 63021
box 0 0 1 1
use contact_17  contact_17_47
timestamp 1644969367
transform 1 0 6434 0 1 63026
box 0 0 1 1
use contact_18  contact_18_48
timestamp 1644969367
transform 1 0 6400 0 1 61483
box 0 0 1 1
use contact_17  contact_17_48
timestamp 1644969367
transform 1 0 6434 0 1 61488
box 0 0 1 1
use contact_18  contact_18_49
timestamp 1644969367
transform 1 0 6400 0 1 59945
box 0 0 1 1
use contact_17  contact_17_49
timestamp 1644969367
transform 1 0 6434 0 1 59950
box 0 0 1 1
use contact_18  contact_18_50
timestamp 1644969367
transform 1 0 6400 0 1 58407
box 0 0 1 1
use contact_17  contact_17_50
timestamp 1644969367
transform 1 0 6434 0 1 58412
box 0 0 1 1
use contact_18  contact_18_51
timestamp 1644969367
transform 1 0 6400 0 1 59945
box 0 0 1 1
use contact_17  contact_17_51
timestamp 1644969367
transform 1 0 6434 0 1 59950
box 0 0 1 1
use contact_18  contact_18_52
timestamp 1644969367
transform 1 0 6400 0 1 58407
box 0 0 1 1
use contact_17  contact_17_52
timestamp 1644969367
transform 1 0 6434 0 1 58412
box 0 0 1 1
use contact_18  contact_18_53
timestamp 1644969367
transform 1 0 6400 0 1 56869
box 0 0 1 1
use contact_17  contact_17_53
timestamp 1644969367
transform 1 0 6434 0 1 56874
box 0 0 1 1
use contact_18  contact_18_54
timestamp 1644969367
transform 1 0 6400 0 1 55331
box 0 0 1 1
use contact_17  contact_17_54
timestamp 1644969367
transform 1 0 6434 0 1 55336
box 0 0 1 1
use contact_18  contact_18_55
timestamp 1644969367
transform 1 0 6400 0 1 56869
box 0 0 1 1
use contact_17  contact_17_55
timestamp 1644969367
transform 1 0 6434 0 1 56874
box 0 0 1 1
use contact_18  contact_18_56
timestamp 1644969367
transform 1 0 6400 0 1 55331
box 0 0 1 1
use contact_17  contact_17_56
timestamp 1644969367
transform 1 0 6434 0 1 55336
box 0 0 1 1
use contact_18  contact_18_57
timestamp 1644969367
transform 1 0 6400 0 1 53793
box 0 0 1 1
use contact_17  contact_17_57
timestamp 1644969367
transform 1 0 6434 0 1 53798
box 0 0 1 1
use contact_18  contact_18_58
timestamp 1644969367
transform 1 0 6400 0 1 52255
box 0 0 1 1
use contact_17  contact_17_58
timestamp 1644969367
transform 1 0 6434 0 1 52260
box 0 0 1 1
use contact_18  contact_18_59
timestamp 1644969367
transform 1 0 6400 0 1 53793
box 0 0 1 1
use contact_17  contact_17_59
timestamp 1644969367
transform 1 0 6434 0 1 53798
box 0 0 1 1
use contact_18  contact_18_60
timestamp 1644969367
transform 1 0 6400 0 1 52255
box 0 0 1 1
use contact_17  contact_17_60
timestamp 1644969367
transform 1 0 6434 0 1 52260
box 0 0 1 1
use contact_18  contact_18_61
timestamp 1644969367
transform 1 0 6400 0 1 50717
box 0 0 1 1
use contact_17  contact_17_61
timestamp 1644969367
transform 1 0 6434 0 1 50722
box 0 0 1 1
use contact_18  contact_18_62
timestamp 1644969367
transform 1 0 6400 0 1 49179
box 0 0 1 1
use contact_17  contact_17_62
timestamp 1644969367
transform 1 0 6434 0 1 49184
box 0 0 1 1
use contact_18  contact_18_63
timestamp 1644969367
transform 1 0 6400 0 1 50717
box 0 0 1 1
use contact_17  contact_17_63
timestamp 1644969367
transform 1 0 6434 0 1 50722
box 0 0 1 1
use contact_18  contact_18_64
timestamp 1644969367
transform 1 0 6400 0 1 49179
box 0 0 1 1
use contact_17  contact_17_64
timestamp 1644969367
transform 1 0 6434 0 1 49184
box 0 0 1 1
use contact_18  contact_18_65
timestamp 1644969367
transform 1 0 6400 0 1 47641
box 0 0 1 1
use contact_17  contact_17_65
timestamp 1644969367
transform 1 0 6434 0 1 47646
box 0 0 1 1
use contact_18  contact_18_66
timestamp 1644969367
transform 1 0 6400 0 1 46103
box 0 0 1 1
use contact_17  contact_17_66
timestamp 1644969367
transform 1 0 6434 0 1 46108
box 0 0 1 1
use contact_18  contact_18_67
timestamp 1644969367
transform 1 0 6400 0 1 47641
box 0 0 1 1
use contact_17  contact_17_67
timestamp 1644969367
transform 1 0 6434 0 1 47646
box 0 0 1 1
use contact_18  contact_18_68
timestamp 1644969367
transform 1 0 6400 0 1 46103
box 0 0 1 1
use contact_17  contact_17_68
timestamp 1644969367
transform 1 0 6434 0 1 46108
box 0 0 1 1
use contact_18  contact_18_69
timestamp 1644969367
transform 1 0 6400 0 1 44565
box 0 0 1 1
use contact_17  contact_17_69
timestamp 1644969367
transform 1 0 6434 0 1 44570
box 0 0 1 1
use contact_18  contact_18_70
timestamp 1644969367
transform 1 0 6400 0 1 43027
box 0 0 1 1
use contact_17  contact_17_70
timestamp 1644969367
transform 1 0 6434 0 1 43032
box 0 0 1 1
use contact_18  contact_18_71
timestamp 1644969367
transform 1 0 6400 0 1 44565
box 0 0 1 1
use contact_17  contact_17_71
timestamp 1644969367
transform 1 0 6434 0 1 44570
box 0 0 1 1
use contact_18  contact_18_72
timestamp 1644969367
transform 1 0 6400 0 1 43027
box 0 0 1 1
use contact_17  contact_17_72
timestamp 1644969367
transform 1 0 6434 0 1 43032
box 0 0 1 1
use contact_18  contact_18_73
timestamp 1644969367
transform 1 0 6400 0 1 41489
box 0 0 1 1
use contact_17  contact_17_73
timestamp 1644969367
transform 1 0 6434 0 1 41494
box 0 0 1 1
use contact_18  contact_18_74
timestamp 1644969367
transform 1 0 6400 0 1 39951
box 0 0 1 1
use contact_17  contact_17_74
timestamp 1644969367
transform 1 0 6434 0 1 39956
box 0 0 1 1
use contact_18  contact_18_75
timestamp 1644969367
transform 1 0 6400 0 1 41489
box 0 0 1 1
use contact_17  contact_17_75
timestamp 1644969367
transform 1 0 6434 0 1 41494
box 0 0 1 1
use contact_18  contact_18_76
timestamp 1644969367
transform 1 0 6400 0 1 39951
box 0 0 1 1
use contact_17  contact_17_76
timestamp 1644969367
transform 1 0 6434 0 1 39956
box 0 0 1 1
use contact_18  contact_18_77
timestamp 1644969367
transform 1 0 6400 0 1 38413
box 0 0 1 1
use contact_17  contact_17_77
timestamp 1644969367
transform 1 0 6434 0 1 38418
box 0 0 1 1
use contact_18  contact_18_78
timestamp 1644969367
transform 1 0 6400 0 1 36875
box 0 0 1 1
use contact_17  contact_17_78
timestamp 1644969367
transform 1 0 6434 0 1 36880
box 0 0 1 1
use contact_18  contact_18_79
timestamp 1644969367
transform 1 0 6400 0 1 38413
box 0 0 1 1
use contact_17  contact_17_79
timestamp 1644969367
transform 1 0 6434 0 1 38418
box 0 0 1 1
use contact_18  contact_18_80
timestamp 1644969367
transform 1 0 6400 0 1 36875
box 0 0 1 1
use contact_17  contact_17_80
timestamp 1644969367
transform 1 0 6434 0 1 36880
box 0 0 1 1
use contact_18  contact_18_81
timestamp 1644969367
transform 1 0 6400 0 1 35337
box 0 0 1 1
use contact_17  contact_17_81
timestamp 1644969367
transform 1 0 6434 0 1 35342
box 0 0 1 1
use contact_18  contact_18_82
timestamp 1644969367
transform 1 0 6400 0 1 33799
box 0 0 1 1
use contact_17  contact_17_82
timestamp 1644969367
transform 1 0 6434 0 1 33804
box 0 0 1 1
use contact_18  contact_18_83
timestamp 1644969367
transform 1 0 6400 0 1 35337
box 0 0 1 1
use contact_17  contact_17_83
timestamp 1644969367
transform 1 0 6434 0 1 35342
box 0 0 1 1
use contact_18  contact_18_84
timestamp 1644969367
transform 1 0 6400 0 1 33799
box 0 0 1 1
use contact_17  contact_17_84
timestamp 1644969367
transform 1 0 6434 0 1 33804
box 0 0 1 1
use contact_18  contact_18_85
timestamp 1644969367
transform 1 0 6400 0 1 32261
box 0 0 1 1
use contact_17  contact_17_85
timestamp 1644969367
transform 1 0 6434 0 1 32266
box 0 0 1 1
use contact_18  contact_18_86
timestamp 1644969367
transform 1 0 6400 0 1 30723
box 0 0 1 1
use contact_17  contact_17_86
timestamp 1644969367
transform 1 0 6434 0 1 30728
box 0 0 1 1
use contact_18  contact_18_87
timestamp 1644969367
transform 1 0 6400 0 1 32261
box 0 0 1 1
use contact_17  contact_17_87
timestamp 1644969367
transform 1 0 6434 0 1 32266
box 0 0 1 1
use contact_18  contact_18_88
timestamp 1644969367
transform 1 0 6400 0 1 30723
box 0 0 1 1
use contact_17  contact_17_88
timestamp 1644969367
transform 1 0 6434 0 1 30728
box 0 0 1 1
use contact_18  contact_18_89
timestamp 1644969367
transform 1 0 6400 0 1 29185
box 0 0 1 1
use contact_17  contact_17_89
timestamp 1644969367
transform 1 0 6434 0 1 29190
box 0 0 1 1
use contact_18  contact_18_90
timestamp 1644969367
transform 1 0 6400 0 1 27647
box 0 0 1 1
use contact_17  contact_17_90
timestamp 1644969367
transform 1 0 6434 0 1 27652
box 0 0 1 1
use contact_18  contact_18_91
timestamp 1644969367
transform 1 0 6400 0 1 29185
box 0 0 1 1
use contact_17  contact_17_91
timestamp 1644969367
transform 1 0 6434 0 1 29190
box 0 0 1 1
use contact_18  contact_18_92
timestamp 1644969367
transform 1 0 6400 0 1 27647
box 0 0 1 1
use contact_17  contact_17_92
timestamp 1644969367
transform 1 0 6434 0 1 27652
box 0 0 1 1
use contact_18  contact_18_93
timestamp 1644969367
transform 1 0 6400 0 1 26109
box 0 0 1 1
use contact_17  contact_17_93
timestamp 1644969367
transform 1 0 6434 0 1 26114
box 0 0 1 1
use contact_18  contact_18_94
timestamp 1644969367
transform 1 0 6400 0 1 24571
box 0 0 1 1
use contact_17  contact_17_94
timestamp 1644969367
transform 1 0 6434 0 1 24576
box 0 0 1 1
use contact_18  contact_18_95
timestamp 1644969367
transform 1 0 6400 0 1 26109
box 0 0 1 1
use contact_17  contact_17_95
timestamp 1644969367
transform 1 0 6434 0 1 26114
box 0 0 1 1
use contact_18  contact_18_96
timestamp 1644969367
transform 1 0 6400 0 1 24571
box 0 0 1 1
use contact_17  contact_17_96
timestamp 1644969367
transform 1 0 6434 0 1 24576
box 0 0 1 1
use contact_18  contact_18_97
timestamp 1644969367
transform 1 0 6400 0 1 23033
box 0 0 1 1
use contact_17  contact_17_97
timestamp 1644969367
transform 1 0 6434 0 1 23038
box 0 0 1 1
use contact_18  contact_18_98
timestamp 1644969367
transform 1 0 6400 0 1 21495
box 0 0 1 1
use contact_17  contact_17_98
timestamp 1644969367
transform 1 0 6434 0 1 21500
box 0 0 1 1
use contact_18  contact_18_99
timestamp 1644969367
transform 1 0 6400 0 1 23033
box 0 0 1 1
use contact_17  contact_17_99
timestamp 1644969367
transform 1 0 6434 0 1 23038
box 0 0 1 1
use contact_18  contact_18_100
timestamp 1644969367
transform 1 0 6400 0 1 21495
box 0 0 1 1
use contact_17  contact_17_100
timestamp 1644969367
transform 1 0 6434 0 1 21500
box 0 0 1 1
use contact_18  contact_18_101
timestamp 1644969367
transform 1 0 6400 0 1 19957
box 0 0 1 1
use contact_17  contact_17_101
timestamp 1644969367
transform 1 0 6434 0 1 19962
box 0 0 1 1
use contact_18  contact_18_102
timestamp 1644969367
transform 1 0 6400 0 1 18419
box 0 0 1 1
use contact_17  contact_17_102
timestamp 1644969367
transform 1 0 6434 0 1 18424
box 0 0 1 1
use contact_18  contact_18_103
timestamp 1644969367
transform 1 0 6400 0 1 19957
box 0 0 1 1
use contact_17  contact_17_103
timestamp 1644969367
transform 1 0 6434 0 1 19962
box 0 0 1 1
use contact_18  contact_18_104
timestamp 1644969367
transform 1 0 6400 0 1 18419
box 0 0 1 1
use contact_17  contact_17_104
timestamp 1644969367
transform 1 0 6434 0 1 18424
box 0 0 1 1
use contact_18  contact_18_105
timestamp 1644969367
transform 1 0 6400 0 1 16881
box 0 0 1 1
use contact_17  contact_17_105
timestamp 1644969367
transform 1 0 6434 0 1 16886
box 0 0 1 1
use contact_18  contact_18_106
timestamp 1644969367
transform 1 0 6400 0 1 15343
box 0 0 1 1
use contact_17  contact_17_106
timestamp 1644969367
transform 1 0 6434 0 1 15348
box 0 0 1 1
use contact_18  contact_18_107
timestamp 1644969367
transform 1 0 6400 0 1 16881
box 0 0 1 1
use contact_17  contact_17_107
timestamp 1644969367
transform 1 0 6434 0 1 16886
box 0 0 1 1
use contact_18  contact_18_108
timestamp 1644969367
transform 1 0 6400 0 1 15343
box 0 0 1 1
use contact_17  contact_17_108
timestamp 1644969367
transform 1 0 6434 0 1 15348
box 0 0 1 1
use contact_18  contact_18_109
timestamp 1644969367
transform 1 0 6400 0 1 13805
box 0 0 1 1
use contact_17  contact_17_109
timestamp 1644969367
transform 1 0 6434 0 1 13810
box 0 0 1 1
use contact_18  contact_18_110
timestamp 1644969367
transform 1 0 6400 0 1 12267
box 0 0 1 1
use contact_17  contact_17_110
timestamp 1644969367
transform 1 0 6434 0 1 12272
box 0 0 1 1
use contact_18  contact_18_111
timestamp 1644969367
transform 1 0 6400 0 1 13805
box 0 0 1 1
use contact_17  contact_17_111
timestamp 1644969367
transform 1 0 6434 0 1 13810
box 0 0 1 1
use contact_18  contact_18_112
timestamp 1644969367
transform 1 0 6400 0 1 12267
box 0 0 1 1
use contact_17  contact_17_112
timestamp 1644969367
transform 1 0 6434 0 1 12272
box 0 0 1 1
use contact_18  contact_18_113
timestamp 1644969367
transform 1 0 6400 0 1 10729
box 0 0 1 1
use contact_17  contact_17_113
timestamp 1644969367
transform 1 0 6434 0 1 10734
box 0 0 1 1
use contact_18  contact_18_114
timestamp 1644969367
transform 1 0 6400 0 1 9191
box 0 0 1 1
use contact_17  contact_17_114
timestamp 1644969367
transform 1 0 6434 0 1 9196
box 0 0 1 1
use contact_18  contact_18_115
timestamp 1644969367
transform 1 0 6400 0 1 10729
box 0 0 1 1
use contact_17  contact_17_115
timestamp 1644969367
transform 1 0 6434 0 1 10734
box 0 0 1 1
use contact_18  contact_18_116
timestamp 1644969367
transform 1 0 6400 0 1 9191
box 0 0 1 1
use contact_17  contact_17_116
timestamp 1644969367
transform 1 0 6434 0 1 9196
box 0 0 1 1
use contact_18  contact_18_117
timestamp 1644969367
transform 1 0 6400 0 1 7653
box 0 0 1 1
use contact_17  contact_17_117
timestamp 1644969367
transform 1 0 6434 0 1 7658
box 0 0 1 1
use contact_18  contact_18_118
timestamp 1644969367
transform 1 0 6400 0 1 6115
box 0 0 1 1
use contact_17  contact_17_118
timestamp 1644969367
transform 1 0 6434 0 1 6120
box 0 0 1 1
use contact_18  contact_18_119
timestamp 1644969367
transform 1 0 6400 0 1 7653
box 0 0 1 1
use contact_17  contact_17_119
timestamp 1644969367
transform 1 0 6434 0 1 7658
box 0 0 1 1
use contact_18  contact_18_120
timestamp 1644969367
transform 1 0 6400 0 1 6115
box 0 0 1 1
use contact_17  contact_17_120
timestamp 1644969367
transform 1 0 6434 0 1 6120
box 0 0 1 1
use contact_18  contact_18_121
timestamp 1644969367
transform 1 0 6400 0 1 4577
box 0 0 1 1
use contact_17  contact_17_121
timestamp 1644969367
transform 1 0 6434 0 1 4582
box 0 0 1 1
use contact_18  contact_18_122
timestamp 1644969367
transform 1 0 6400 0 1 3039
box 0 0 1 1
use contact_17  contact_17_122
timestamp 1644969367
transform 1 0 6434 0 1 3044
box 0 0 1 1
use contact_18  contact_18_123
timestamp 1644969367
transform 1 0 6400 0 1 4577
box 0 0 1 1
use contact_17  contact_17_123
timestamp 1644969367
transform 1 0 6434 0 1 4582
box 0 0 1 1
use contact_18  contact_18_124
timestamp 1644969367
transform 1 0 6400 0 1 3039
box 0 0 1 1
use contact_17  contact_17_124
timestamp 1644969367
transform 1 0 6434 0 1 3044
box 0 0 1 1
use contact_18  contact_18_125
timestamp 1644969367
transform 1 0 6400 0 1 1501
box 0 0 1 1
use contact_17  contact_17_125
timestamp 1644969367
transform 1 0 6434 0 1 1506
box 0 0 1 1
use contact_18  contact_18_126
timestamp 1644969367
transform 1 0 6400 0 1 -37
box 0 0 1 1
use contact_17  contact_17_126
timestamp 1644969367
transform 1 0 6434 0 1 -32
box 0 0 1 1
use contact_18  contact_18_127
timestamp 1644969367
transform 1 0 6400 0 1 1501
box 0 0 1 1
use contact_17  contact_17_127
timestamp 1644969367
transform 1 0 6434 0 1 1506
box 0 0 1 1
use contact_20  contact_20_0
timestamp 1644969367
transform 1 0 4822 0 1 35375
box 0 0 1 1
use contact_18  contact_18_128
timestamp 1644969367
transform 1 0 2973 0 1 36187
box 0 0 1 1
use contact_17  contact_17_128
timestamp 1644969367
transform 1 0 3007 0 1 36192
box 0 0 1 1
use contact_13  contact_13_0
timestamp 1644969367
transform 1 0 3010 0 1 36201
box 0 0 1 1
use contact_20  contact_20_1
timestamp 1644969367
transform 1 0 4738 0 1 33835
box 0 0 1 1
use contact_18  contact_18_129
timestamp 1644969367
transform 1 0 2973 0 1 34563
box 0 0 1 1
use contact_17  contact_17_129
timestamp 1644969367
transform 1 0 3007 0 1 34568
box 0 0 1 1
use contact_13  contact_13_1
timestamp 1644969367
transform 1 0 3010 0 1 34577
box 0 0 1 1
use contact_20  contact_20_2
timestamp 1644969367
transform 1 0 4654 0 1 32295
box 0 0 1 1
use contact_18  contact_18_130
timestamp 1644969367
transform 1 0 2973 0 1 33107
box 0 0 1 1
use contact_17  contact_17_130
timestamp 1644969367
transform 1 0 3007 0 1 33112
box 0 0 1 1
use contact_13  contact_13_2
timestamp 1644969367
transform 1 0 3010 0 1 33121
box 0 0 1 1
use contact_20  contact_20_3
timestamp 1644969367
transform 1 0 4570 0 1 30755
box 0 0 1 1
use contact_18  contact_18_131
timestamp 1644969367
transform 1 0 2973 0 1 31483
box 0 0 1 1
use contact_17  contact_17_131
timestamp 1644969367
transform 1 0 3007 0 1 31488
box 0 0 1 1
use contact_13  contact_13_3
timestamp 1644969367
transform 1 0 3010 0 1 31497
box 0 0 1 1
use contact_20  contact_20_4
timestamp 1644969367
transform 1 0 4486 0 1 29215
box 0 0 1 1
use contact_18  contact_18_132
timestamp 1644969367
transform 1 0 2973 0 1 30027
box 0 0 1 1
use contact_17  contact_17_132
timestamp 1644969367
transform 1 0 3007 0 1 30032
box 0 0 1 1
use contact_13  contact_13_4
timestamp 1644969367
transform 1 0 3010 0 1 30041
box 0 0 1 1
use contact_20  contact_20_5
timestamp 1644969367
transform 1 0 4402 0 1 27675
box 0 0 1 1
use contact_18  contact_18_133
timestamp 1644969367
transform 1 0 2973 0 1 28403
box 0 0 1 1
use contact_17  contact_17_133
timestamp 1644969367
transform 1 0 3007 0 1 28408
box 0 0 1 1
use contact_13  contact_13_5
timestamp 1644969367
transform 1 0 3010 0 1 28417
box 0 0 1 1
use contact_20  contact_20_6
timestamp 1644969367
transform 1 0 4318 0 1 26135
box 0 0 1 1
use contact_18  contact_18_134
timestamp 1644969367
transform 1 0 2973 0 1 26947
box 0 0 1 1
use contact_17  contact_17_134
timestamp 1644969367
transform 1 0 3007 0 1 26952
box 0 0 1 1
use contact_13  contact_13_6
timestamp 1644969367
transform 1 0 3010 0 1 26961
box 0 0 1 1
use contact_20  contact_20_7
timestamp 1644969367
transform 1 0 4234 0 1 24595
box 0 0 1 1
use contact_18  contact_18_135
timestamp 1644969367
transform 1 0 2973 0 1 25323
box 0 0 1 1
use contact_17  contact_17_135
timestamp 1644969367
transform 1 0 3007 0 1 25328
box 0 0 1 1
use contact_13  contact_13_7
timestamp 1644969367
transform 1 0 3010 0 1 25337
box 0 0 1 1
use contact_20  contact_20_8
timestamp 1644969367
transform 1 0 4150 0 1 19979
box 0 0 1 1
use contact_18  contact_18_136
timestamp 1644969367
transform 1 0 2973 0 1 20791
box 0 0 1 1
use contact_17  contact_17_136
timestamp 1644969367
transform 1 0 3007 0 1 20796
box 0 0 1 1
use contact_13  contact_13_8
timestamp 1644969367
transform 1 0 3010 0 1 20805
box 0 0 1 1
use contact_20  contact_20_9
timestamp 1644969367
transform 1 0 4066 0 1 18439
box 0 0 1 1
use contact_18  contact_18_137
timestamp 1644969367
transform 1 0 2973 0 1 19167
box 0 0 1 1
use contact_17  contact_17_137
timestamp 1644969367
transform 1 0 3007 0 1 19172
box 0 0 1 1
use contact_13  contact_13_9
timestamp 1644969367
transform 1 0 3010 0 1 19181
box 0 0 1 1
use contact_20  contact_20_10
timestamp 1644969367
transform 1 0 3982 0 1 16899
box 0 0 1 1
use contact_18  contact_18_138
timestamp 1644969367
transform 1 0 2973 0 1 17711
box 0 0 1 1
use contact_17  contact_17_138
timestamp 1644969367
transform 1 0 3007 0 1 17716
box 0 0 1 1
use contact_13  contact_13_10
timestamp 1644969367
transform 1 0 3010 0 1 17725
box 0 0 1 1
use contact_20  contact_20_11
timestamp 1644969367
transform 1 0 3898 0 1 15359
box 0 0 1 1
use contact_18  contact_18_139
timestamp 1644969367
transform 1 0 2973 0 1 16087
box 0 0 1 1
use contact_17  contact_17_139
timestamp 1644969367
transform 1 0 3007 0 1 16092
box 0 0 1 1
use contact_13  contact_13_11
timestamp 1644969367
transform 1 0 3010 0 1 16101
box 0 0 1 1
use contact_20  contact_20_12
timestamp 1644969367
transform 1 0 3814 0 1 13819
box 0 0 1 1
use contact_18  contact_18_140
timestamp 1644969367
transform 1 0 2973 0 1 14631
box 0 0 1 1
use contact_17  contact_17_140
timestamp 1644969367
transform 1 0 3007 0 1 14636
box 0 0 1 1
use contact_13  contact_13_12
timestamp 1644969367
transform 1 0 3010 0 1 14645
box 0 0 1 1
use contact_20  contact_20_13
timestamp 1644969367
transform 1 0 3730 0 1 12279
box 0 0 1 1
use contact_18  contact_18_141
timestamp 1644969367
transform 1 0 2973 0 1 13007
box 0 0 1 1
use contact_17  contact_17_141
timestamp 1644969367
transform 1 0 3007 0 1 13012
box 0 0 1 1
use contact_13  contact_13_13
timestamp 1644969367
transform 1 0 3010 0 1 13021
box 0 0 1 1
use contact_20  contact_20_14
timestamp 1644969367
transform 1 0 3646 0 1 10739
box 0 0 1 1
use contact_18  contact_18_142
timestamp 1644969367
transform 1 0 2973 0 1 11551
box 0 0 1 1
use contact_17  contact_17_142
timestamp 1644969367
transform 1 0 3007 0 1 11556
box 0 0 1 1
use contact_13  contact_13_14
timestamp 1644969367
transform 1 0 3010 0 1 11565
box 0 0 1 1
use contact_20  contact_20_15
timestamp 1644969367
transform 1 0 3562 0 1 9199
box 0 0 1 1
use contact_18  contact_18_143
timestamp 1644969367
transform 1 0 2973 0 1 9927
box 0 0 1 1
use contact_17  contact_17_143
timestamp 1644969367
transform 1 0 3007 0 1 9932
box 0 0 1 1
use contact_13  contact_13_15
timestamp 1644969367
transform 1 0 3010 0 1 9941
box 0 0 1 1
use contact_20  contact_20_16
timestamp 1644969367
transform 1 0 3478 0 1 4583
box 0 0 1 1
use contact_18  contact_18_144
timestamp 1644969367
transform 1 0 2973 0 1 5395
box 0 0 1 1
use contact_17  contact_17_144
timestamp 1644969367
transform 1 0 3007 0 1 5400
box 0 0 1 1
use contact_13  contact_13_16
timestamp 1644969367
transform 1 0 3010 0 1 5409
box 0 0 1 1
use contact_20  contact_20_17
timestamp 1644969367
transform 1 0 3394 0 1 3043
box 0 0 1 1
use contact_18  contact_18_145
timestamp 1644969367
transform 1 0 2973 0 1 3771
box 0 0 1 1
use contact_17  contact_17_145
timestamp 1644969367
transform 1 0 3007 0 1 3776
box 0 0 1 1
use contact_13  contact_13_17
timestamp 1644969367
transform 1 0 3010 0 1 3785
box 0 0 1 1
use contact_20  contact_20_18
timestamp 1644969367
transform 1 0 3310 0 1 1503
box 0 0 1 1
use contact_18  contact_18_146
timestamp 1644969367
transform 1 0 2973 0 1 2315
box 0 0 1 1
use contact_17  contact_17_146
timestamp 1644969367
transform 1 0 3007 0 1 2320
box 0 0 1 1
use contact_13  contact_13_18
timestamp 1644969367
transform 1 0 3010 0 1 2329
box 0 0 1 1
use contact_20  contact_20_19
timestamp 1644969367
transform 1 0 3226 0 1 -37
box 0 0 1 1
use contact_18  contact_18_147
timestamp 1644969367
transform 1 0 2973 0 1 691
box 0 0 1 1
use contact_17  contact_17_147
timestamp 1644969367
transform 1 0 3007 0 1 696
box 0 0 1 1
use contact_13  contact_13_19
timestamp 1644969367
transform 1 0 3010 0 1 705
box 0 0 1 1
use contact_14  contact_14_0
timestamp 1644969367
transform 1 0 4688 0 1 98018
box 0 0 1 1
use contact_14  contact_14_1
timestamp 1644969367
transform 1 0 4184 0 1 97932
box 0 0 1 1
use contact_14  contact_14_2
timestamp 1644969367
transform 1 0 3428 0 1 97846
box 0 0 1 1
use contact_14  contact_14_3
timestamp 1644969367
transform 1 0 4688 0 1 97760
box 0 0 1 1
use contact_14  contact_14_4
timestamp 1644969367
transform 1 0 4184 0 1 97674
box 0 0 1 1
use contact_14  contact_14_5
timestamp 1644969367
transform 1 0 3344 0 1 97588
box 0 0 1 1
use contact_14  contact_14_6
timestamp 1644969367
transform 1 0 4688 0 1 97502
box 0 0 1 1
use contact_14  contact_14_7
timestamp 1644969367
transform 1 0 4184 0 1 97416
box 0 0 1 1
use contact_14  contact_14_8
timestamp 1644969367
transform 1 0 3260 0 1 97330
box 0 0 1 1
use contact_14  contact_14_9
timestamp 1644969367
transform 1 0 4688 0 1 95706
box 0 0 1 1
use contact_14  contact_14_10
timestamp 1644969367
transform 1 0 4100 0 1 95792
box 0 0 1 1
use contact_14  contact_14_11
timestamp 1644969367
transform 1 0 3512 0 1 95878
box 0 0 1 1
use contact_14  contact_14_12
timestamp 1644969367
transform 1 0 4688 0 1 95964
box 0 0 1 1
use contact_14  contact_14_13
timestamp 1644969367
transform 1 0 4100 0 1 96050
box 0 0 1 1
use contact_14  contact_14_14
timestamp 1644969367
transform 1 0 3428 0 1 96136
box 0 0 1 1
use contact_14  contact_14_15
timestamp 1644969367
transform 1 0 4688 0 1 96222
box 0 0 1 1
use contact_14  contact_14_16
timestamp 1644969367
transform 1 0 4100 0 1 96308
box 0 0 1 1
use contact_14  contact_14_17
timestamp 1644969367
transform 1 0 3344 0 1 96394
box 0 0 1 1
use contact_14  contact_14_18
timestamp 1644969367
transform 1 0 4688 0 1 94942
box 0 0 1 1
use contact_14  contact_14_19
timestamp 1644969367
transform 1 0 4100 0 1 94856
box 0 0 1 1
use contact_14  contact_14_20
timestamp 1644969367
transform 1 0 3260 0 1 94770
box 0 0 1 1
use contact_14  contact_14_21
timestamp 1644969367
transform 1 0 4688 0 1 94684
box 0 0 1 1
use contact_14  contact_14_22
timestamp 1644969367
transform 1 0 4016 0 1 94598
box 0 0 1 1
use contact_14  contact_14_23
timestamp 1644969367
transform 1 0 3512 0 1 94512
box 0 0 1 1
use contact_14  contact_14_24
timestamp 1644969367
transform 1 0 4688 0 1 94426
box 0 0 1 1
use contact_14  contact_14_25
timestamp 1644969367
transform 1 0 4016 0 1 94340
box 0 0 1 1
use contact_14  contact_14_26
timestamp 1644969367
transform 1 0 3428 0 1 94254
box 0 0 1 1
use contact_14  contact_14_27
timestamp 1644969367
transform 1 0 4688 0 1 92630
box 0 0 1 1
use contact_14  contact_14_28
timestamp 1644969367
transform 1 0 4016 0 1 92716
box 0 0 1 1
use contact_14  contact_14_29
timestamp 1644969367
transform 1 0 3344 0 1 92802
box 0 0 1 1
use contact_14  contact_14_30
timestamp 1644969367
transform 1 0 4688 0 1 92888
box 0 0 1 1
use contact_14  contact_14_31
timestamp 1644969367
transform 1 0 4016 0 1 92974
box 0 0 1 1
use contact_14  contact_14_32
timestamp 1644969367
transform 1 0 3260 0 1 93060
box 0 0 1 1
use contact_14  contact_14_33
timestamp 1644969367
transform 1 0 4688 0 1 93146
box 0 0 1 1
use contact_14  contact_14_34
timestamp 1644969367
transform 1 0 3932 0 1 93232
box 0 0 1 1
use contact_14  contact_14_35
timestamp 1644969367
transform 1 0 3512 0 1 93318
box 0 0 1 1
use contact_14  contact_14_36
timestamp 1644969367
transform 1 0 4688 0 1 91866
box 0 0 1 1
use contact_14  contact_14_37
timestamp 1644969367
transform 1 0 3932 0 1 91780
box 0 0 1 1
use contact_14  contact_14_38
timestamp 1644969367
transform 1 0 3428 0 1 91694
box 0 0 1 1
use contact_14  contact_14_39
timestamp 1644969367
transform 1 0 4688 0 1 91608
box 0 0 1 1
use contact_14  contact_14_40
timestamp 1644969367
transform 1 0 3932 0 1 91522
box 0 0 1 1
use contact_14  contact_14_41
timestamp 1644969367
transform 1 0 3344 0 1 91436
box 0 0 1 1
use contact_14  contact_14_42
timestamp 1644969367
transform 1 0 4688 0 1 91350
box 0 0 1 1
use contact_14  contact_14_43
timestamp 1644969367
transform 1 0 3932 0 1 91264
box 0 0 1 1
use contact_14  contact_14_44
timestamp 1644969367
transform 1 0 3260 0 1 91178
box 0 0 1 1
use contact_14  contact_14_45
timestamp 1644969367
transform 1 0 4688 0 1 89554
box 0 0 1 1
use contact_14  contact_14_46
timestamp 1644969367
transform 1 0 3848 0 1 89640
box 0 0 1 1
use contact_14  contact_14_47
timestamp 1644969367
transform 1 0 3512 0 1 89726
box 0 0 1 1
use contact_14  contact_14_48
timestamp 1644969367
transform 1 0 4688 0 1 89812
box 0 0 1 1
use contact_14  contact_14_49
timestamp 1644969367
transform 1 0 3848 0 1 89898
box 0 0 1 1
use contact_14  contact_14_50
timestamp 1644969367
transform 1 0 3428 0 1 89984
box 0 0 1 1
use contact_14  contact_14_51
timestamp 1644969367
transform 1 0 4688 0 1 90070
box 0 0 1 1
use contact_14  contact_14_52
timestamp 1644969367
transform 1 0 3848 0 1 90156
box 0 0 1 1
use contact_14  contact_14_53
timestamp 1644969367
transform 1 0 3344 0 1 90242
box 0 0 1 1
use contact_14  contact_14_54
timestamp 1644969367
transform 1 0 4688 0 1 88790
box 0 0 1 1
use contact_14  contact_14_55
timestamp 1644969367
transform 1 0 3848 0 1 88704
box 0 0 1 1
use contact_14  contact_14_56
timestamp 1644969367
transform 1 0 3260 0 1 88618
box 0 0 1 1
use contact_14  contact_14_57
timestamp 1644969367
transform 1 0 4688 0 1 88532
box 0 0 1 1
use contact_14  contact_14_58
timestamp 1644969367
transform 1 0 3764 0 1 88446
box 0 0 1 1
use contact_14  contact_14_59
timestamp 1644969367
transform 1 0 3512 0 1 88360
box 0 0 1 1
use contact_14  contact_14_60
timestamp 1644969367
transform 1 0 4688 0 1 88274
box 0 0 1 1
use contact_14  contact_14_61
timestamp 1644969367
transform 1 0 3764 0 1 88188
box 0 0 1 1
use contact_14  contact_14_62
timestamp 1644969367
transform 1 0 3428 0 1 88102
box 0 0 1 1
use contact_14  contact_14_63
timestamp 1644969367
transform 1 0 4688 0 1 86478
box 0 0 1 1
use contact_14  contact_14_64
timestamp 1644969367
transform 1 0 3764 0 1 86564
box 0 0 1 1
use contact_14  contact_14_65
timestamp 1644969367
transform 1 0 3344 0 1 86650
box 0 0 1 1
use contact_14  contact_14_66
timestamp 1644969367
transform 1 0 4688 0 1 86736
box 0 0 1 1
use contact_14  contact_14_67
timestamp 1644969367
transform 1 0 3764 0 1 86822
box 0 0 1 1
use contact_14  contact_14_68
timestamp 1644969367
transform 1 0 3260 0 1 86908
box 0 0 1 1
use contact_14  contact_14_69
timestamp 1644969367
transform 1 0 4688 0 1 86994
box 0 0 1 1
use contact_14  contact_14_70
timestamp 1644969367
transform 1 0 3680 0 1 87080
box 0 0 1 1
use contact_14  contact_14_71
timestamp 1644969367
transform 1 0 3512 0 1 87166
box 0 0 1 1
use contact_14  contact_14_72
timestamp 1644969367
transform 1 0 4688 0 1 85714
box 0 0 1 1
use contact_14  contact_14_73
timestamp 1644969367
transform 1 0 3680 0 1 85628
box 0 0 1 1
use contact_14  contact_14_74
timestamp 1644969367
transform 1 0 3428 0 1 85542
box 0 0 1 1
use contact_14  contact_14_75
timestamp 1644969367
transform 1 0 4688 0 1 85456
box 0 0 1 1
use contact_14  contact_14_76
timestamp 1644969367
transform 1 0 3680 0 1 85370
box 0 0 1 1
use contact_14  contact_14_77
timestamp 1644969367
transform 1 0 3344 0 1 85284
box 0 0 1 1
use contact_14  contact_14_78
timestamp 1644969367
transform 1 0 4688 0 1 85198
box 0 0 1 1
use contact_14  contact_14_79
timestamp 1644969367
transform 1 0 3680 0 1 85112
box 0 0 1 1
use contact_14  contact_14_80
timestamp 1644969367
transform 1 0 3260 0 1 85026
box 0 0 1 1
use contact_14  contact_14_81
timestamp 1644969367
transform 1 0 4688 0 1 83402
box 0 0 1 1
use contact_14  contact_14_82
timestamp 1644969367
transform 1 0 3596 0 1 83488
box 0 0 1 1
use contact_14  contact_14_83
timestamp 1644969367
transform 1 0 3512 0 1 83574
box 0 0 1 1
use contact_14  contact_14_84
timestamp 1644969367
transform 1 0 4688 0 1 83660
box 0 0 1 1
use contact_14  contact_14_85
timestamp 1644969367
transform 1 0 3596 0 1 83746
box 0 0 1 1
use contact_14  contact_14_86
timestamp 1644969367
transform 1 0 3428 0 1 83832
box 0 0 1 1
use contact_14  contact_14_87
timestamp 1644969367
transform 1 0 4688 0 1 83918
box 0 0 1 1
use contact_14  contact_14_88
timestamp 1644969367
transform 1 0 3596 0 1 84004
box 0 0 1 1
use contact_14  contact_14_89
timestamp 1644969367
transform 1 0 3344 0 1 84090
box 0 0 1 1
use contact_14  contact_14_90
timestamp 1644969367
transform 1 0 4688 0 1 82638
box 0 0 1 1
use contact_14  contact_14_91
timestamp 1644969367
transform 1 0 3596 0 1 82552
box 0 0 1 1
use contact_14  contact_14_92
timestamp 1644969367
transform 1 0 3260 0 1 82466
box 0 0 1 1
use contact_14  contact_14_93
timestamp 1644969367
transform 1 0 4604 0 1 82380
box 0 0 1 1
use contact_14  contact_14_94
timestamp 1644969367
transform 1 0 4184 0 1 82294
box 0 0 1 1
use contact_14  contact_14_95
timestamp 1644969367
transform 1 0 3512 0 1 82208
box 0 0 1 1
use contact_14  contact_14_96
timestamp 1644969367
transform 1 0 4604 0 1 82122
box 0 0 1 1
use contact_14  contact_14_97
timestamp 1644969367
transform 1 0 4184 0 1 82036
box 0 0 1 1
use contact_14  contact_14_98
timestamp 1644969367
transform 1 0 3428 0 1 81950
box 0 0 1 1
use contact_14  contact_14_99
timestamp 1644969367
transform 1 0 4604 0 1 80326
box 0 0 1 1
use contact_14  contact_14_100
timestamp 1644969367
transform 1 0 4184 0 1 80412
box 0 0 1 1
use contact_14  contact_14_101
timestamp 1644969367
transform 1 0 3344 0 1 80498
box 0 0 1 1
use contact_14  contact_14_102
timestamp 1644969367
transform 1 0 4604 0 1 80584
box 0 0 1 1
use contact_14  contact_14_103
timestamp 1644969367
transform 1 0 4184 0 1 80670
box 0 0 1 1
use contact_14  contact_14_104
timestamp 1644969367
transform 1 0 3260 0 1 80756
box 0 0 1 1
use contact_14  contact_14_105
timestamp 1644969367
transform 1 0 4604 0 1 80842
box 0 0 1 1
use contact_14  contact_14_106
timestamp 1644969367
transform 1 0 4100 0 1 80928
box 0 0 1 1
use contact_14  contact_14_107
timestamp 1644969367
transform 1 0 3512 0 1 81014
box 0 0 1 1
use contact_14  contact_14_108
timestamp 1644969367
transform 1 0 4604 0 1 79562
box 0 0 1 1
use contact_14  contact_14_109
timestamp 1644969367
transform 1 0 4100 0 1 79476
box 0 0 1 1
use contact_14  contact_14_110
timestamp 1644969367
transform 1 0 3428 0 1 79390
box 0 0 1 1
use contact_14  contact_14_111
timestamp 1644969367
transform 1 0 4604 0 1 79304
box 0 0 1 1
use contact_14  contact_14_112
timestamp 1644969367
transform 1 0 4100 0 1 79218
box 0 0 1 1
use contact_14  contact_14_113
timestamp 1644969367
transform 1 0 3344 0 1 79132
box 0 0 1 1
use contact_14  contact_14_114
timestamp 1644969367
transform 1 0 4604 0 1 79046
box 0 0 1 1
use contact_14  contact_14_115
timestamp 1644969367
transform 1 0 4100 0 1 78960
box 0 0 1 1
use contact_14  contact_14_116
timestamp 1644969367
transform 1 0 3260 0 1 78874
box 0 0 1 1
use contact_14  contact_14_117
timestamp 1644969367
transform 1 0 4604 0 1 77250
box 0 0 1 1
use contact_14  contact_14_118
timestamp 1644969367
transform 1 0 4016 0 1 77336
box 0 0 1 1
use contact_14  contact_14_119
timestamp 1644969367
transform 1 0 3512 0 1 77422
box 0 0 1 1
use contact_14  contact_14_120
timestamp 1644969367
transform 1 0 4604 0 1 77508
box 0 0 1 1
use contact_14  contact_14_121
timestamp 1644969367
transform 1 0 4016 0 1 77594
box 0 0 1 1
use contact_14  contact_14_122
timestamp 1644969367
transform 1 0 3428 0 1 77680
box 0 0 1 1
use contact_14  contact_14_123
timestamp 1644969367
transform 1 0 4604 0 1 77766
box 0 0 1 1
use contact_14  contact_14_124
timestamp 1644969367
transform 1 0 4016 0 1 77852
box 0 0 1 1
use contact_14  contact_14_125
timestamp 1644969367
transform 1 0 3344 0 1 77938
box 0 0 1 1
use contact_14  contact_14_126
timestamp 1644969367
transform 1 0 4604 0 1 76486
box 0 0 1 1
use contact_14  contact_14_127
timestamp 1644969367
transform 1 0 4016 0 1 76400
box 0 0 1 1
use contact_14  contact_14_128
timestamp 1644969367
transform 1 0 3260 0 1 76314
box 0 0 1 1
use contact_14  contact_14_129
timestamp 1644969367
transform 1 0 4604 0 1 76228
box 0 0 1 1
use contact_14  contact_14_130
timestamp 1644969367
transform 1 0 3932 0 1 76142
box 0 0 1 1
use contact_14  contact_14_131
timestamp 1644969367
transform 1 0 3512 0 1 76056
box 0 0 1 1
use contact_14  contact_14_132
timestamp 1644969367
transform 1 0 4604 0 1 75970
box 0 0 1 1
use contact_14  contact_14_133
timestamp 1644969367
transform 1 0 3932 0 1 75884
box 0 0 1 1
use contact_14  contact_14_134
timestamp 1644969367
transform 1 0 3428 0 1 75798
box 0 0 1 1
use contact_14  contact_14_135
timestamp 1644969367
transform 1 0 4604 0 1 74174
box 0 0 1 1
use contact_14  contact_14_136
timestamp 1644969367
transform 1 0 3932 0 1 74260
box 0 0 1 1
use contact_14  contact_14_137
timestamp 1644969367
transform 1 0 3344 0 1 74346
box 0 0 1 1
use contact_14  contact_14_138
timestamp 1644969367
transform 1 0 4604 0 1 74432
box 0 0 1 1
use contact_14  contact_14_139
timestamp 1644969367
transform 1 0 3932 0 1 74518
box 0 0 1 1
use contact_14  contact_14_140
timestamp 1644969367
transform 1 0 3260 0 1 74604
box 0 0 1 1
use contact_14  contact_14_141
timestamp 1644969367
transform 1 0 4604 0 1 74690
box 0 0 1 1
use contact_14  contact_14_142
timestamp 1644969367
transform 1 0 3848 0 1 74776
box 0 0 1 1
use contact_14  contact_14_143
timestamp 1644969367
transform 1 0 3512 0 1 74862
box 0 0 1 1
use contact_14  contact_14_144
timestamp 1644969367
transform 1 0 4604 0 1 73410
box 0 0 1 1
use contact_14  contact_14_145
timestamp 1644969367
transform 1 0 3848 0 1 73324
box 0 0 1 1
use contact_14  contact_14_146
timestamp 1644969367
transform 1 0 3428 0 1 73238
box 0 0 1 1
use contact_14  contact_14_147
timestamp 1644969367
transform 1 0 4604 0 1 73152
box 0 0 1 1
use contact_14  contact_14_148
timestamp 1644969367
transform 1 0 3848 0 1 73066
box 0 0 1 1
use contact_14  contact_14_149
timestamp 1644969367
transform 1 0 3344 0 1 72980
box 0 0 1 1
use contact_14  contact_14_150
timestamp 1644969367
transform 1 0 4604 0 1 72894
box 0 0 1 1
use contact_14  contact_14_151
timestamp 1644969367
transform 1 0 3848 0 1 72808
box 0 0 1 1
use contact_14  contact_14_152
timestamp 1644969367
transform 1 0 3260 0 1 72722
box 0 0 1 1
use contact_14  contact_14_153
timestamp 1644969367
transform 1 0 4604 0 1 71098
box 0 0 1 1
use contact_14  contact_14_154
timestamp 1644969367
transform 1 0 3764 0 1 71184
box 0 0 1 1
use contact_14  contact_14_155
timestamp 1644969367
transform 1 0 3512 0 1 71270
box 0 0 1 1
use contact_14  contact_14_156
timestamp 1644969367
transform 1 0 4604 0 1 71356
box 0 0 1 1
use contact_14  contact_14_157
timestamp 1644969367
transform 1 0 3764 0 1 71442
box 0 0 1 1
use contact_14  contact_14_158
timestamp 1644969367
transform 1 0 3428 0 1 71528
box 0 0 1 1
use contact_14  contact_14_159
timestamp 1644969367
transform 1 0 4604 0 1 71614
box 0 0 1 1
use contact_14  contact_14_160
timestamp 1644969367
transform 1 0 3764 0 1 71700
box 0 0 1 1
use contact_14  contact_14_161
timestamp 1644969367
transform 1 0 3344 0 1 71786
box 0 0 1 1
use contact_14  contact_14_162
timestamp 1644969367
transform 1 0 4604 0 1 70334
box 0 0 1 1
use contact_14  contact_14_163
timestamp 1644969367
transform 1 0 3764 0 1 70248
box 0 0 1 1
use contact_14  contact_14_164
timestamp 1644969367
transform 1 0 3260 0 1 70162
box 0 0 1 1
use contact_14  contact_14_165
timestamp 1644969367
transform 1 0 4604 0 1 70076
box 0 0 1 1
use contact_14  contact_14_166
timestamp 1644969367
transform 1 0 3680 0 1 69990
box 0 0 1 1
use contact_14  contact_14_167
timestamp 1644969367
transform 1 0 3512 0 1 69904
box 0 0 1 1
use contact_14  contact_14_168
timestamp 1644969367
transform 1 0 4604 0 1 69818
box 0 0 1 1
use contact_14  contact_14_169
timestamp 1644969367
transform 1 0 3680 0 1 69732
box 0 0 1 1
use contact_14  contact_14_170
timestamp 1644969367
transform 1 0 3428 0 1 69646
box 0 0 1 1
use contact_14  contact_14_171
timestamp 1644969367
transform 1 0 4604 0 1 68022
box 0 0 1 1
use contact_14  contact_14_172
timestamp 1644969367
transform 1 0 3680 0 1 68108
box 0 0 1 1
use contact_14  contact_14_173
timestamp 1644969367
transform 1 0 3344 0 1 68194
box 0 0 1 1
use contact_14  contact_14_174
timestamp 1644969367
transform 1 0 4604 0 1 68280
box 0 0 1 1
use contact_14  contact_14_175
timestamp 1644969367
transform 1 0 3680 0 1 68366
box 0 0 1 1
use contact_14  contact_14_176
timestamp 1644969367
transform 1 0 3260 0 1 68452
box 0 0 1 1
use contact_14  contact_14_177
timestamp 1644969367
transform 1 0 4604 0 1 68538
box 0 0 1 1
use contact_14  contact_14_178
timestamp 1644969367
transform 1 0 3596 0 1 68624
box 0 0 1 1
use contact_14  contact_14_179
timestamp 1644969367
transform 1 0 3512 0 1 68710
box 0 0 1 1
use contact_14  contact_14_180
timestamp 1644969367
transform 1 0 4604 0 1 67258
box 0 0 1 1
use contact_14  contact_14_181
timestamp 1644969367
transform 1 0 3596 0 1 67172
box 0 0 1 1
use contact_14  contact_14_182
timestamp 1644969367
transform 1 0 3428 0 1 67086
box 0 0 1 1
use contact_14  contact_14_183
timestamp 1644969367
transform 1 0 4604 0 1 67000
box 0 0 1 1
use contact_14  contact_14_184
timestamp 1644969367
transform 1 0 3596 0 1 66914
box 0 0 1 1
use contact_14  contact_14_185
timestamp 1644969367
transform 1 0 3344 0 1 66828
box 0 0 1 1
use contact_14  contact_14_186
timestamp 1644969367
transform 1 0 4604 0 1 66742
box 0 0 1 1
use contact_14  contact_14_187
timestamp 1644969367
transform 1 0 3596 0 1 66656
box 0 0 1 1
use contact_14  contact_14_188
timestamp 1644969367
transform 1 0 3260 0 1 66570
box 0 0 1 1
use contact_14  contact_14_189
timestamp 1644969367
transform 1 0 4520 0 1 64946
box 0 0 1 1
use contact_14  contact_14_190
timestamp 1644969367
transform 1 0 4184 0 1 65032
box 0 0 1 1
use contact_14  contact_14_191
timestamp 1644969367
transform 1 0 3512 0 1 65118
box 0 0 1 1
use contact_14  contact_14_192
timestamp 1644969367
transform 1 0 4520 0 1 65204
box 0 0 1 1
use contact_14  contact_14_193
timestamp 1644969367
transform 1 0 4184 0 1 65290
box 0 0 1 1
use contact_14  contact_14_194
timestamp 1644969367
transform 1 0 3428 0 1 65376
box 0 0 1 1
use contact_14  contact_14_195
timestamp 1644969367
transform 1 0 4520 0 1 65462
box 0 0 1 1
use contact_14  contact_14_196
timestamp 1644969367
transform 1 0 4184 0 1 65548
box 0 0 1 1
use contact_14  contact_14_197
timestamp 1644969367
transform 1 0 3344 0 1 65634
box 0 0 1 1
use contact_14  contact_14_198
timestamp 1644969367
transform 1 0 4520 0 1 64182
box 0 0 1 1
use contact_14  contact_14_199
timestamp 1644969367
transform 1 0 4184 0 1 64096
box 0 0 1 1
use contact_14  contact_14_200
timestamp 1644969367
transform 1 0 3260 0 1 64010
box 0 0 1 1
use contact_14  contact_14_201
timestamp 1644969367
transform 1 0 4520 0 1 63924
box 0 0 1 1
use contact_14  contact_14_202
timestamp 1644969367
transform 1 0 4100 0 1 63838
box 0 0 1 1
use contact_14  contact_14_203
timestamp 1644969367
transform 1 0 3512 0 1 63752
box 0 0 1 1
use contact_14  contact_14_204
timestamp 1644969367
transform 1 0 4520 0 1 63666
box 0 0 1 1
use contact_14  contact_14_205
timestamp 1644969367
transform 1 0 4100 0 1 63580
box 0 0 1 1
use contact_14  contact_14_206
timestamp 1644969367
transform 1 0 3428 0 1 63494
box 0 0 1 1
use contact_14  contact_14_207
timestamp 1644969367
transform 1 0 4520 0 1 61870
box 0 0 1 1
use contact_14  contact_14_208
timestamp 1644969367
transform 1 0 4100 0 1 61956
box 0 0 1 1
use contact_14  contact_14_209
timestamp 1644969367
transform 1 0 3344 0 1 62042
box 0 0 1 1
use contact_14  contact_14_210
timestamp 1644969367
transform 1 0 4520 0 1 62128
box 0 0 1 1
use contact_14  contact_14_211
timestamp 1644969367
transform 1 0 4100 0 1 62214
box 0 0 1 1
use contact_14  contact_14_212
timestamp 1644969367
transform 1 0 3260 0 1 62300
box 0 0 1 1
use contact_14  contact_14_213
timestamp 1644969367
transform 1 0 4520 0 1 62386
box 0 0 1 1
use contact_14  contact_14_214
timestamp 1644969367
transform 1 0 4016 0 1 62472
box 0 0 1 1
use contact_14  contact_14_215
timestamp 1644969367
transform 1 0 3512 0 1 62558
box 0 0 1 1
use contact_14  contact_14_216
timestamp 1644969367
transform 1 0 4520 0 1 61106
box 0 0 1 1
use contact_14  contact_14_217
timestamp 1644969367
transform 1 0 4016 0 1 61020
box 0 0 1 1
use contact_14  contact_14_218
timestamp 1644969367
transform 1 0 3428 0 1 60934
box 0 0 1 1
use contact_14  contact_14_219
timestamp 1644969367
transform 1 0 4520 0 1 60848
box 0 0 1 1
use contact_14  contact_14_220
timestamp 1644969367
transform 1 0 4016 0 1 60762
box 0 0 1 1
use contact_14  contact_14_221
timestamp 1644969367
transform 1 0 3344 0 1 60676
box 0 0 1 1
use contact_14  contact_14_222
timestamp 1644969367
transform 1 0 4520 0 1 60590
box 0 0 1 1
use contact_14  contact_14_223
timestamp 1644969367
transform 1 0 4016 0 1 60504
box 0 0 1 1
use contact_14  contact_14_224
timestamp 1644969367
transform 1 0 3260 0 1 60418
box 0 0 1 1
use contact_14  contact_14_225
timestamp 1644969367
transform 1 0 4520 0 1 58794
box 0 0 1 1
use contact_14  contact_14_226
timestamp 1644969367
transform 1 0 3932 0 1 58880
box 0 0 1 1
use contact_14  contact_14_227
timestamp 1644969367
transform 1 0 3512 0 1 58966
box 0 0 1 1
use contact_14  contact_14_228
timestamp 1644969367
transform 1 0 4520 0 1 59052
box 0 0 1 1
use contact_14  contact_14_229
timestamp 1644969367
transform 1 0 3932 0 1 59138
box 0 0 1 1
use contact_14  contact_14_230
timestamp 1644969367
transform 1 0 3428 0 1 59224
box 0 0 1 1
use contact_14  contact_14_231
timestamp 1644969367
transform 1 0 4520 0 1 59310
box 0 0 1 1
use contact_14  contact_14_232
timestamp 1644969367
transform 1 0 3932 0 1 59396
box 0 0 1 1
use contact_14  contact_14_233
timestamp 1644969367
transform 1 0 3344 0 1 59482
box 0 0 1 1
use contact_14  contact_14_234
timestamp 1644969367
transform 1 0 4520 0 1 58030
box 0 0 1 1
use contact_14  contact_14_235
timestamp 1644969367
transform 1 0 3932 0 1 57944
box 0 0 1 1
use contact_14  contact_14_236
timestamp 1644969367
transform 1 0 3260 0 1 57858
box 0 0 1 1
use contact_14  contact_14_237
timestamp 1644969367
transform 1 0 4520 0 1 57772
box 0 0 1 1
use contact_14  contact_14_238
timestamp 1644969367
transform 1 0 3848 0 1 57686
box 0 0 1 1
use contact_14  contact_14_239
timestamp 1644969367
transform 1 0 3512 0 1 57600
box 0 0 1 1
use contact_14  contact_14_240
timestamp 1644969367
transform 1 0 4520 0 1 57514
box 0 0 1 1
use contact_14  contact_14_241
timestamp 1644969367
transform 1 0 3848 0 1 57428
box 0 0 1 1
use contact_14  contact_14_242
timestamp 1644969367
transform 1 0 3428 0 1 57342
box 0 0 1 1
use contact_14  contact_14_243
timestamp 1644969367
transform 1 0 4520 0 1 55718
box 0 0 1 1
use contact_14  contact_14_244
timestamp 1644969367
transform 1 0 3848 0 1 55804
box 0 0 1 1
use contact_14  contact_14_245
timestamp 1644969367
transform 1 0 3344 0 1 55890
box 0 0 1 1
use contact_14  contact_14_246
timestamp 1644969367
transform 1 0 4520 0 1 55976
box 0 0 1 1
use contact_14  contact_14_247
timestamp 1644969367
transform 1 0 3848 0 1 56062
box 0 0 1 1
use contact_14  contact_14_248
timestamp 1644969367
transform 1 0 3260 0 1 56148
box 0 0 1 1
use contact_14  contact_14_249
timestamp 1644969367
transform 1 0 4520 0 1 56234
box 0 0 1 1
use contact_14  contact_14_250
timestamp 1644969367
transform 1 0 3764 0 1 56320
box 0 0 1 1
use contact_14  contact_14_251
timestamp 1644969367
transform 1 0 3512 0 1 56406
box 0 0 1 1
use contact_14  contact_14_252
timestamp 1644969367
transform 1 0 4520 0 1 54954
box 0 0 1 1
use contact_14  contact_14_253
timestamp 1644969367
transform 1 0 3764 0 1 54868
box 0 0 1 1
use contact_14  contact_14_254
timestamp 1644969367
transform 1 0 3428 0 1 54782
box 0 0 1 1
use contact_14  contact_14_255
timestamp 1644969367
transform 1 0 4520 0 1 54696
box 0 0 1 1
use contact_14  contact_14_256
timestamp 1644969367
transform 1 0 3764 0 1 54610
box 0 0 1 1
use contact_14  contact_14_257
timestamp 1644969367
transform 1 0 3344 0 1 54524
box 0 0 1 1
use contact_14  contact_14_258
timestamp 1644969367
transform 1 0 4520 0 1 54438
box 0 0 1 1
use contact_14  contact_14_259
timestamp 1644969367
transform 1 0 3764 0 1 54352
box 0 0 1 1
use contact_14  contact_14_260
timestamp 1644969367
transform 1 0 3260 0 1 54266
box 0 0 1 1
use contact_14  contact_14_261
timestamp 1644969367
transform 1 0 4520 0 1 52642
box 0 0 1 1
use contact_14  contact_14_262
timestamp 1644969367
transform 1 0 3680 0 1 52728
box 0 0 1 1
use contact_14  contact_14_263
timestamp 1644969367
transform 1 0 3512 0 1 52814
box 0 0 1 1
use contact_14  contact_14_264
timestamp 1644969367
transform 1 0 4520 0 1 52900
box 0 0 1 1
use contact_14  contact_14_265
timestamp 1644969367
transform 1 0 3680 0 1 52986
box 0 0 1 1
use contact_14  contact_14_266
timestamp 1644969367
transform 1 0 3428 0 1 53072
box 0 0 1 1
use contact_14  contact_14_267
timestamp 1644969367
transform 1 0 4520 0 1 53158
box 0 0 1 1
use contact_14  contact_14_268
timestamp 1644969367
transform 1 0 3680 0 1 53244
box 0 0 1 1
use contact_14  contact_14_269
timestamp 1644969367
transform 1 0 3344 0 1 53330
box 0 0 1 1
use contact_14  contact_14_270
timestamp 1644969367
transform 1 0 4520 0 1 51878
box 0 0 1 1
use contact_14  contact_14_271
timestamp 1644969367
transform 1 0 3680 0 1 51792
box 0 0 1 1
use contact_14  contact_14_272
timestamp 1644969367
transform 1 0 3260 0 1 51706
box 0 0 1 1
use contact_14  contact_14_273
timestamp 1644969367
transform 1 0 4520 0 1 51620
box 0 0 1 1
use contact_14  contact_14_274
timestamp 1644969367
transform 1 0 3596 0 1 51534
box 0 0 1 1
use contact_14  contact_14_275
timestamp 1644969367
transform 1 0 3512 0 1 51448
box 0 0 1 1
use contact_14  contact_14_276
timestamp 1644969367
transform 1 0 4520 0 1 51362
box 0 0 1 1
use contact_14  contact_14_277
timestamp 1644969367
transform 1 0 3596 0 1 51276
box 0 0 1 1
use contact_14  contact_14_278
timestamp 1644969367
transform 1 0 3428 0 1 51190
box 0 0 1 1
use contact_14  contact_14_279
timestamp 1644969367
transform 1 0 4520 0 1 49566
box 0 0 1 1
use contact_14  contact_14_280
timestamp 1644969367
transform 1 0 3596 0 1 49652
box 0 0 1 1
use contact_14  contact_14_281
timestamp 1644969367
transform 1 0 3344 0 1 49738
box 0 0 1 1
use contact_14  contact_14_282
timestamp 1644969367
transform 1 0 4520 0 1 49824
box 0 0 1 1
use contact_14  contact_14_283
timestamp 1644969367
transform 1 0 3596 0 1 49910
box 0 0 1 1
use contact_14  contact_14_284
timestamp 1644969367
transform 1 0 3260 0 1 49996
box 0 0 1 1
use contact_14  contact_14_285
timestamp 1644969367
transform 1 0 4436 0 1 50082
box 0 0 1 1
use contact_14  contact_14_286
timestamp 1644969367
transform 1 0 4184 0 1 50168
box 0 0 1 1
use contact_14  contact_14_287
timestamp 1644969367
transform 1 0 3512 0 1 50254
box 0 0 1 1
use contact_14  contact_14_288
timestamp 1644969367
transform 1 0 4436 0 1 48802
box 0 0 1 1
use contact_14  contact_14_289
timestamp 1644969367
transform 1 0 4184 0 1 48716
box 0 0 1 1
use contact_14  contact_14_290
timestamp 1644969367
transform 1 0 3428 0 1 48630
box 0 0 1 1
use contact_14  contact_14_291
timestamp 1644969367
transform 1 0 4436 0 1 48544
box 0 0 1 1
use contact_14  contact_14_292
timestamp 1644969367
transform 1 0 4184 0 1 48458
box 0 0 1 1
use contact_14  contact_14_293
timestamp 1644969367
transform 1 0 3344 0 1 48372
box 0 0 1 1
use contact_14  contact_14_294
timestamp 1644969367
transform 1 0 4436 0 1 48286
box 0 0 1 1
use contact_14  contact_14_295
timestamp 1644969367
transform 1 0 4184 0 1 48200
box 0 0 1 1
use contact_14  contact_14_296
timestamp 1644969367
transform 1 0 3260 0 1 48114
box 0 0 1 1
use contact_14  contact_14_297
timestamp 1644969367
transform 1 0 4436 0 1 46490
box 0 0 1 1
use contact_14  contact_14_298
timestamp 1644969367
transform 1 0 4100 0 1 46576
box 0 0 1 1
use contact_14  contact_14_299
timestamp 1644969367
transform 1 0 3512 0 1 46662
box 0 0 1 1
use contact_14  contact_14_300
timestamp 1644969367
transform 1 0 4436 0 1 46748
box 0 0 1 1
use contact_14  contact_14_301
timestamp 1644969367
transform 1 0 4100 0 1 46834
box 0 0 1 1
use contact_14  contact_14_302
timestamp 1644969367
transform 1 0 3428 0 1 46920
box 0 0 1 1
use contact_14  contact_14_303
timestamp 1644969367
transform 1 0 4436 0 1 47006
box 0 0 1 1
use contact_14  contact_14_304
timestamp 1644969367
transform 1 0 4100 0 1 47092
box 0 0 1 1
use contact_14  contact_14_305
timestamp 1644969367
transform 1 0 3344 0 1 47178
box 0 0 1 1
use contact_14  contact_14_306
timestamp 1644969367
transform 1 0 4436 0 1 45726
box 0 0 1 1
use contact_14  contact_14_307
timestamp 1644969367
transform 1 0 4100 0 1 45640
box 0 0 1 1
use contact_14  contact_14_308
timestamp 1644969367
transform 1 0 3260 0 1 45554
box 0 0 1 1
use contact_14  contact_14_309
timestamp 1644969367
transform 1 0 4436 0 1 45468
box 0 0 1 1
use contact_14  contact_14_310
timestamp 1644969367
transform 1 0 4016 0 1 45382
box 0 0 1 1
use contact_14  contact_14_311
timestamp 1644969367
transform 1 0 3512 0 1 45296
box 0 0 1 1
use contact_14  contact_14_312
timestamp 1644969367
transform 1 0 4436 0 1 45210
box 0 0 1 1
use contact_14  contact_14_313
timestamp 1644969367
transform 1 0 4016 0 1 45124
box 0 0 1 1
use contact_14  contact_14_314
timestamp 1644969367
transform 1 0 3428 0 1 45038
box 0 0 1 1
use contact_14  contact_14_315
timestamp 1644969367
transform 1 0 4436 0 1 43414
box 0 0 1 1
use contact_14  contact_14_316
timestamp 1644969367
transform 1 0 4016 0 1 43500
box 0 0 1 1
use contact_14  contact_14_317
timestamp 1644969367
transform 1 0 3344 0 1 43586
box 0 0 1 1
use contact_14  contact_14_318
timestamp 1644969367
transform 1 0 4436 0 1 43672
box 0 0 1 1
use contact_14  contact_14_319
timestamp 1644969367
transform 1 0 4016 0 1 43758
box 0 0 1 1
use contact_14  contact_14_320
timestamp 1644969367
transform 1 0 3260 0 1 43844
box 0 0 1 1
use contact_14  contact_14_321
timestamp 1644969367
transform 1 0 4436 0 1 43930
box 0 0 1 1
use contact_14  contact_14_322
timestamp 1644969367
transform 1 0 3932 0 1 44016
box 0 0 1 1
use contact_14  contact_14_323
timestamp 1644969367
transform 1 0 3512 0 1 44102
box 0 0 1 1
use contact_14  contact_14_324
timestamp 1644969367
transform 1 0 4436 0 1 42650
box 0 0 1 1
use contact_14  contact_14_325
timestamp 1644969367
transform 1 0 3932 0 1 42564
box 0 0 1 1
use contact_14  contact_14_326
timestamp 1644969367
transform 1 0 3428 0 1 42478
box 0 0 1 1
use contact_14  contact_14_327
timestamp 1644969367
transform 1 0 4436 0 1 42392
box 0 0 1 1
use contact_14  contact_14_328
timestamp 1644969367
transform 1 0 3932 0 1 42306
box 0 0 1 1
use contact_14  contact_14_329
timestamp 1644969367
transform 1 0 3344 0 1 42220
box 0 0 1 1
use contact_14  contact_14_330
timestamp 1644969367
transform 1 0 4436 0 1 42134
box 0 0 1 1
use contact_14  contact_14_331
timestamp 1644969367
transform 1 0 3932 0 1 42048
box 0 0 1 1
use contact_14  contact_14_332
timestamp 1644969367
transform 1 0 3260 0 1 41962
box 0 0 1 1
use contact_14  contact_14_333
timestamp 1644969367
transform 1 0 4436 0 1 40338
box 0 0 1 1
use contact_14  contact_14_334
timestamp 1644969367
transform 1 0 3848 0 1 40424
box 0 0 1 1
use contact_14  contact_14_335
timestamp 1644969367
transform 1 0 3512 0 1 40510
box 0 0 1 1
use contact_14  contact_14_336
timestamp 1644969367
transform 1 0 4436 0 1 40596
box 0 0 1 1
use contact_14  contact_14_337
timestamp 1644969367
transform 1 0 3848 0 1 40682
box 0 0 1 1
use contact_14  contact_14_338
timestamp 1644969367
transform 1 0 3428 0 1 40768
box 0 0 1 1
use contact_14  contact_14_339
timestamp 1644969367
transform 1 0 4436 0 1 40854
box 0 0 1 1
use contact_14  contact_14_340
timestamp 1644969367
transform 1 0 3848 0 1 40940
box 0 0 1 1
use contact_14  contact_14_341
timestamp 1644969367
transform 1 0 3344 0 1 41026
box 0 0 1 1
use contact_14  contact_14_342
timestamp 1644969367
transform 1 0 4436 0 1 39574
box 0 0 1 1
use contact_14  contact_14_343
timestamp 1644969367
transform 1 0 3848 0 1 39488
box 0 0 1 1
use contact_14  contact_14_344
timestamp 1644969367
transform 1 0 3260 0 1 39402
box 0 0 1 1
use contact_14  contact_14_345
timestamp 1644969367
transform 1 0 4436 0 1 39316
box 0 0 1 1
use contact_14  contact_14_346
timestamp 1644969367
transform 1 0 3764 0 1 39230
box 0 0 1 1
use contact_14  contact_14_347
timestamp 1644969367
transform 1 0 3512 0 1 39144
box 0 0 1 1
use contact_14  contact_14_348
timestamp 1644969367
transform 1 0 4436 0 1 39058
box 0 0 1 1
use contact_14  contact_14_349
timestamp 1644969367
transform 1 0 3764 0 1 38972
box 0 0 1 1
use contact_14  contact_14_350
timestamp 1644969367
transform 1 0 3428 0 1 38886
box 0 0 1 1
use contact_14  contact_14_351
timestamp 1644969367
transform 1 0 4436 0 1 37262
box 0 0 1 1
use contact_14  contact_14_352
timestamp 1644969367
transform 1 0 3764 0 1 37348
box 0 0 1 1
use contact_14  contact_14_353
timestamp 1644969367
transform 1 0 3344 0 1 37434
box 0 0 1 1
use contact_14  contact_14_354
timestamp 1644969367
transform 1 0 4436 0 1 37520
box 0 0 1 1
use contact_14  contact_14_355
timestamp 1644969367
transform 1 0 3764 0 1 37606
box 0 0 1 1
use contact_14  contact_14_356
timestamp 1644969367
transform 1 0 3260 0 1 37692
box 0 0 1 1
use contact_14  contact_14_357
timestamp 1644969367
transform 1 0 4436 0 1 37778
box 0 0 1 1
use contact_14  contact_14_358
timestamp 1644969367
transform 1 0 3680 0 1 37864
box 0 0 1 1
use contact_14  contact_14_359
timestamp 1644969367
transform 1 0 3512 0 1 37950
box 0 0 1 1
use contact_14  contact_14_360
timestamp 1644969367
transform 1 0 4436 0 1 36498
box 0 0 1 1
use contact_14  contact_14_361
timestamp 1644969367
transform 1 0 3680 0 1 36412
box 0 0 1 1
use contact_14  contact_14_362
timestamp 1644969367
transform 1 0 3428 0 1 36326
box 0 0 1 1
use contact_14  contact_14_363
timestamp 1644969367
transform 1 0 4436 0 1 36240
box 0 0 1 1
use contact_14  contact_14_364
timestamp 1644969367
transform 1 0 3680 0 1 36154
box 0 0 1 1
use contact_14  contact_14_365
timestamp 1644969367
transform 1 0 3344 0 1 36068
box 0 0 1 1
use contact_14  contact_14_366
timestamp 1644969367
transform 1 0 4436 0 1 35982
box 0 0 1 1
use contact_14  contact_14_367
timestamp 1644969367
transform 1 0 3680 0 1 35896
box 0 0 1 1
use contact_14  contact_14_368
timestamp 1644969367
transform 1 0 3260 0 1 35810
box 0 0 1 1
use contact_14  contact_14_369
timestamp 1644969367
transform 1 0 4436 0 1 34186
box 0 0 1 1
use contact_14  contact_14_370
timestamp 1644969367
transform 1 0 3596 0 1 34272
box 0 0 1 1
use contact_14  contact_14_371
timestamp 1644969367
transform 1 0 3512 0 1 34358
box 0 0 1 1
use contact_14  contact_14_372
timestamp 1644969367
transform 1 0 4436 0 1 34444
box 0 0 1 1
use contact_14  contact_14_373
timestamp 1644969367
transform 1 0 3596 0 1 34530
box 0 0 1 1
use contact_14  contact_14_374
timestamp 1644969367
transform 1 0 3428 0 1 34616
box 0 0 1 1
use contact_14  contact_14_375
timestamp 1644969367
transform 1 0 4436 0 1 34702
box 0 0 1 1
use contact_14  contact_14_376
timestamp 1644969367
transform 1 0 3596 0 1 34788
box 0 0 1 1
use contact_14  contact_14_377
timestamp 1644969367
transform 1 0 3344 0 1 34874
box 0 0 1 1
use contact_14  contact_14_378
timestamp 1644969367
transform 1 0 4436 0 1 33422
box 0 0 1 1
use contact_14  contact_14_379
timestamp 1644969367
transform 1 0 3596 0 1 33336
box 0 0 1 1
use contact_14  contact_14_380
timestamp 1644969367
transform 1 0 3260 0 1 33250
box 0 0 1 1
use contact_14  contact_14_381
timestamp 1644969367
transform 1 0 4352 0 1 33164
box 0 0 1 1
use contact_14  contact_14_382
timestamp 1644969367
transform 1 0 4184 0 1 33078
box 0 0 1 1
use contact_14  contact_14_383
timestamp 1644969367
transform 1 0 3512 0 1 32992
box 0 0 1 1
use contact_14  contact_14_384
timestamp 1644969367
transform 1 0 4352 0 1 32906
box 0 0 1 1
use contact_14  contact_14_385
timestamp 1644969367
transform 1 0 4184 0 1 32820
box 0 0 1 1
use contact_14  contact_14_386
timestamp 1644969367
transform 1 0 3428 0 1 32734
box 0 0 1 1
use contact_14  contact_14_387
timestamp 1644969367
transform 1 0 4352 0 1 31110
box 0 0 1 1
use contact_14  contact_14_388
timestamp 1644969367
transform 1 0 4184 0 1 31196
box 0 0 1 1
use contact_14  contact_14_389
timestamp 1644969367
transform 1 0 3344 0 1 31282
box 0 0 1 1
use contact_14  contact_14_390
timestamp 1644969367
transform 1 0 4352 0 1 31368
box 0 0 1 1
use contact_14  contact_14_391
timestamp 1644969367
transform 1 0 4184 0 1 31454
box 0 0 1 1
use contact_14  contact_14_392
timestamp 1644969367
transform 1 0 3260 0 1 31540
box 0 0 1 1
use contact_14  contact_14_393
timestamp 1644969367
transform 1 0 4352 0 1 31626
box 0 0 1 1
use contact_14  contact_14_394
timestamp 1644969367
transform 1 0 4100 0 1 31712
box 0 0 1 1
use contact_14  contact_14_395
timestamp 1644969367
transform 1 0 3512 0 1 31798
box 0 0 1 1
use contact_14  contact_14_396
timestamp 1644969367
transform 1 0 4352 0 1 30346
box 0 0 1 1
use contact_14  contact_14_397
timestamp 1644969367
transform 1 0 4100 0 1 30260
box 0 0 1 1
use contact_14  contact_14_398
timestamp 1644969367
transform 1 0 3428 0 1 30174
box 0 0 1 1
use contact_14  contact_14_399
timestamp 1644969367
transform 1 0 4352 0 1 30088
box 0 0 1 1
use contact_14  contact_14_400
timestamp 1644969367
transform 1 0 4100 0 1 30002
box 0 0 1 1
use contact_14  contact_14_401
timestamp 1644969367
transform 1 0 3344 0 1 29916
box 0 0 1 1
use contact_14  contact_14_402
timestamp 1644969367
transform 1 0 4352 0 1 29830
box 0 0 1 1
use contact_14  contact_14_403
timestamp 1644969367
transform 1 0 4100 0 1 29744
box 0 0 1 1
use contact_14  contact_14_404
timestamp 1644969367
transform 1 0 3260 0 1 29658
box 0 0 1 1
use contact_14  contact_14_405
timestamp 1644969367
transform 1 0 4352 0 1 28034
box 0 0 1 1
use contact_14  contact_14_406
timestamp 1644969367
transform 1 0 4016 0 1 28120
box 0 0 1 1
use contact_14  contact_14_407
timestamp 1644969367
transform 1 0 3512 0 1 28206
box 0 0 1 1
use contact_14  contact_14_408
timestamp 1644969367
transform 1 0 4352 0 1 28292
box 0 0 1 1
use contact_14  contact_14_409
timestamp 1644969367
transform 1 0 4016 0 1 28378
box 0 0 1 1
use contact_14  contact_14_410
timestamp 1644969367
transform 1 0 3428 0 1 28464
box 0 0 1 1
use contact_14  contact_14_411
timestamp 1644969367
transform 1 0 4352 0 1 28550
box 0 0 1 1
use contact_14  contact_14_412
timestamp 1644969367
transform 1 0 4016 0 1 28636
box 0 0 1 1
use contact_14  contact_14_413
timestamp 1644969367
transform 1 0 3344 0 1 28722
box 0 0 1 1
use contact_14  contact_14_414
timestamp 1644969367
transform 1 0 4352 0 1 27270
box 0 0 1 1
use contact_14  contact_14_415
timestamp 1644969367
transform 1 0 4016 0 1 27184
box 0 0 1 1
use contact_14  contact_14_416
timestamp 1644969367
transform 1 0 3260 0 1 27098
box 0 0 1 1
use contact_14  contact_14_417
timestamp 1644969367
transform 1 0 4352 0 1 27012
box 0 0 1 1
use contact_14  contact_14_418
timestamp 1644969367
transform 1 0 3932 0 1 26926
box 0 0 1 1
use contact_14  contact_14_419
timestamp 1644969367
transform 1 0 3512 0 1 26840
box 0 0 1 1
use contact_14  contact_14_420
timestamp 1644969367
transform 1 0 4352 0 1 26754
box 0 0 1 1
use contact_14  contact_14_421
timestamp 1644969367
transform 1 0 3932 0 1 26668
box 0 0 1 1
use contact_14  contact_14_422
timestamp 1644969367
transform 1 0 3428 0 1 26582
box 0 0 1 1
use contact_14  contact_14_423
timestamp 1644969367
transform 1 0 4352 0 1 24958
box 0 0 1 1
use contact_14  contact_14_424
timestamp 1644969367
transform 1 0 3932 0 1 25044
box 0 0 1 1
use contact_14  contact_14_425
timestamp 1644969367
transform 1 0 3344 0 1 25130
box 0 0 1 1
use contact_14  contact_14_426
timestamp 1644969367
transform 1 0 4352 0 1 25216
box 0 0 1 1
use contact_14  contact_14_427
timestamp 1644969367
transform 1 0 3932 0 1 25302
box 0 0 1 1
use contact_14  contact_14_428
timestamp 1644969367
transform 1 0 3260 0 1 25388
box 0 0 1 1
use contact_14  contact_14_429
timestamp 1644969367
transform 1 0 4352 0 1 25474
box 0 0 1 1
use contact_14  contact_14_430
timestamp 1644969367
transform 1 0 3848 0 1 25560
box 0 0 1 1
use contact_14  contact_14_431
timestamp 1644969367
transform 1 0 3512 0 1 25646
box 0 0 1 1
use contact_14  contact_14_432
timestamp 1644969367
transform 1 0 4352 0 1 24194
box 0 0 1 1
use contact_14  contact_14_433
timestamp 1644969367
transform 1 0 3848 0 1 24108
box 0 0 1 1
use contact_14  contact_14_434
timestamp 1644969367
transform 1 0 3428 0 1 24022
box 0 0 1 1
use contact_14  contact_14_435
timestamp 1644969367
transform 1 0 4352 0 1 23936
box 0 0 1 1
use contact_14  contact_14_436
timestamp 1644969367
transform 1 0 3848 0 1 23850
box 0 0 1 1
use contact_14  contact_14_437
timestamp 1644969367
transform 1 0 3344 0 1 23764
box 0 0 1 1
use contact_14  contact_14_438
timestamp 1644969367
transform 1 0 4352 0 1 23678
box 0 0 1 1
use contact_14  contact_14_439
timestamp 1644969367
transform 1 0 3848 0 1 23592
box 0 0 1 1
use contact_14  contact_14_440
timestamp 1644969367
transform 1 0 3260 0 1 23506
box 0 0 1 1
use contact_14  contact_14_441
timestamp 1644969367
transform 1 0 4352 0 1 21882
box 0 0 1 1
use contact_14  contact_14_442
timestamp 1644969367
transform 1 0 3764 0 1 21968
box 0 0 1 1
use contact_14  contact_14_443
timestamp 1644969367
transform 1 0 3512 0 1 22054
box 0 0 1 1
use contact_14  contact_14_444
timestamp 1644969367
transform 1 0 4352 0 1 22140
box 0 0 1 1
use contact_14  contact_14_445
timestamp 1644969367
transform 1 0 3764 0 1 22226
box 0 0 1 1
use contact_14  contact_14_446
timestamp 1644969367
transform 1 0 3428 0 1 22312
box 0 0 1 1
use contact_14  contact_14_447
timestamp 1644969367
transform 1 0 4352 0 1 22398
box 0 0 1 1
use contact_14  contact_14_448
timestamp 1644969367
transform 1 0 3764 0 1 22484
box 0 0 1 1
use contact_14  contact_14_449
timestamp 1644969367
transform 1 0 3344 0 1 22570
box 0 0 1 1
use contact_14  contact_14_450
timestamp 1644969367
transform 1 0 4352 0 1 21118
box 0 0 1 1
use contact_14  contact_14_451
timestamp 1644969367
transform 1 0 3764 0 1 21032
box 0 0 1 1
use contact_14  contact_14_452
timestamp 1644969367
transform 1 0 3260 0 1 20946
box 0 0 1 1
use contact_14  contact_14_453
timestamp 1644969367
transform 1 0 4352 0 1 20860
box 0 0 1 1
use contact_14  contact_14_454
timestamp 1644969367
transform 1 0 3680 0 1 20774
box 0 0 1 1
use contact_14  contact_14_455
timestamp 1644969367
transform 1 0 3512 0 1 20688
box 0 0 1 1
use contact_14  contact_14_456
timestamp 1644969367
transform 1 0 4352 0 1 20602
box 0 0 1 1
use contact_14  contact_14_457
timestamp 1644969367
transform 1 0 3680 0 1 20516
box 0 0 1 1
use contact_14  contact_14_458
timestamp 1644969367
transform 1 0 3428 0 1 20430
box 0 0 1 1
use contact_14  contact_14_459
timestamp 1644969367
transform 1 0 4352 0 1 18806
box 0 0 1 1
use contact_14  contact_14_460
timestamp 1644969367
transform 1 0 3680 0 1 18892
box 0 0 1 1
use contact_14  contact_14_461
timestamp 1644969367
transform 1 0 3344 0 1 18978
box 0 0 1 1
use contact_14  contact_14_462
timestamp 1644969367
transform 1 0 4352 0 1 19064
box 0 0 1 1
use contact_14  contact_14_463
timestamp 1644969367
transform 1 0 3680 0 1 19150
box 0 0 1 1
use contact_14  contact_14_464
timestamp 1644969367
transform 1 0 3260 0 1 19236
box 0 0 1 1
use contact_14  contact_14_465
timestamp 1644969367
transform 1 0 4352 0 1 19322
box 0 0 1 1
use contact_14  contact_14_466
timestamp 1644969367
transform 1 0 3596 0 1 19408
box 0 0 1 1
use contact_14  contact_14_467
timestamp 1644969367
transform 1 0 3512 0 1 19494
box 0 0 1 1
use contact_14  contact_14_468
timestamp 1644969367
transform 1 0 4352 0 1 18042
box 0 0 1 1
use contact_14  contact_14_469
timestamp 1644969367
transform 1 0 3596 0 1 17956
box 0 0 1 1
use contact_14  contact_14_470
timestamp 1644969367
transform 1 0 3428 0 1 17870
box 0 0 1 1
use contact_14  contact_14_471
timestamp 1644969367
transform 1 0 4352 0 1 17784
box 0 0 1 1
use contact_14  contact_14_472
timestamp 1644969367
transform 1 0 3596 0 1 17698
box 0 0 1 1
use contact_14  contact_14_473
timestamp 1644969367
transform 1 0 3344 0 1 17612
box 0 0 1 1
use contact_14  contact_14_474
timestamp 1644969367
transform 1 0 4352 0 1 17526
box 0 0 1 1
use contact_14  contact_14_475
timestamp 1644969367
transform 1 0 3596 0 1 17440
box 0 0 1 1
use contact_14  contact_14_476
timestamp 1644969367
transform 1 0 3260 0 1 17354
box 0 0 1 1
use contact_14  contact_14_477
timestamp 1644969367
transform 1 0 4268 0 1 15730
box 0 0 1 1
use contact_14  contact_14_478
timestamp 1644969367
transform 1 0 4184 0 1 15816
box 0 0 1 1
use contact_14  contact_14_479
timestamp 1644969367
transform 1 0 3512 0 1 15902
box 0 0 1 1
use contact_14  contact_14_480
timestamp 1644969367
transform 1 0 4268 0 1 15988
box 0 0 1 1
use contact_14  contact_14_481
timestamp 1644969367
transform 1 0 4184 0 1 16074
box 0 0 1 1
use contact_14  contact_14_482
timestamp 1644969367
transform 1 0 3428 0 1 16160
box 0 0 1 1
use contact_14  contact_14_483
timestamp 1644969367
transform 1 0 4268 0 1 16246
box 0 0 1 1
use contact_14  contact_14_484
timestamp 1644969367
transform 1 0 4184 0 1 16332
box 0 0 1 1
use contact_14  contact_14_485
timestamp 1644969367
transform 1 0 3344 0 1 16418
box 0 0 1 1
use contact_14  contact_14_486
timestamp 1644969367
transform 1 0 4268 0 1 14966
box 0 0 1 1
use contact_14  contact_14_487
timestamp 1644969367
transform 1 0 4184 0 1 14880
box 0 0 1 1
use contact_14  contact_14_488
timestamp 1644969367
transform 1 0 3260 0 1 14794
box 0 0 1 1
use contact_14  contact_14_489
timestamp 1644969367
transform 1 0 4268 0 1 14708
box 0 0 1 1
use contact_14  contact_14_490
timestamp 1644969367
transform 1 0 4100 0 1 14622
box 0 0 1 1
use contact_14  contact_14_491
timestamp 1644969367
transform 1 0 3512 0 1 14536
box 0 0 1 1
use contact_14  contact_14_492
timestamp 1644969367
transform 1 0 4268 0 1 14450
box 0 0 1 1
use contact_14  contact_14_493
timestamp 1644969367
transform 1 0 4100 0 1 14364
box 0 0 1 1
use contact_14  contact_14_494
timestamp 1644969367
transform 1 0 3428 0 1 14278
box 0 0 1 1
use contact_14  contact_14_495
timestamp 1644969367
transform 1 0 4268 0 1 12654
box 0 0 1 1
use contact_14  contact_14_496
timestamp 1644969367
transform 1 0 4100 0 1 12740
box 0 0 1 1
use contact_14  contact_14_497
timestamp 1644969367
transform 1 0 3344 0 1 12826
box 0 0 1 1
use contact_14  contact_14_498
timestamp 1644969367
transform 1 0 4268 0 1 12912
box 0 0 1 1
use contact_14  contact_14_499
timestamp 1644969367
transform 1 0 4100 0 1 12998
box 0 0 1 1
use contact_14  contact_14_500
timestamp 1644969367
transform 1 0 3260 0 1 13084
box 0 0 1 1
use contact_14  contact_14_501
timestamp 1644969367
transform 1 0 4268 0 1 13170
box 0 0 1 1
use contact_14  contact_14_502
timestamp 1644969367
transform 1 0 4016 0 1 13256
box 0 0 1 1
use contact_14  contact_14_503
timestamp 1644969367
transform 1 0 3512 0 1 13342
box 0 0 1 1
use contact_14  contact_14_504
timestamp 1644969367
transform 1 0 4268 0 1 11890
box 0 0 1 1
use contact_14  contact_14_505
timestamp 1644969367
transform 1 0 4016 0 1 11804
box 0 0 1 1
use contact_14  contact_14_506
timestamp 1644969367
transform 1 0 3428 0 1 11718
box 0 0 1 1
use contact_14  contact_14_507
timestamp 1644969367
transform 1 0 4268 0 1 11632
box 0 0 1 1
use contact_14  contact_14_508
timestamp 1644969367
transform 1 0 4016 0 1 11546
box 0 0 1 1
use contact_14  contact_14_509
timestamp 1644969367
transform 1 0 3344 0 1 11460
box 0 0 1 1
use contact_14  contact_14_510
timestamp 1644969367
transform 1 0 4268 0 1 11374
box 0 0 1 1
use contact_14  contact_14_511
timestamp 1644969367
transform 1 0 4016 0 1 11288
box 0 0 1 1
use contact_14  contact_14_512
timestamp 1644969367
transform 1 0 3260 0 1 11202
box 0 0 1 1
use contact_14  contact_14_513
timestamp 1644969367
transform 1 0 4268 0 1 9578
box 0 0 1 1
use contact_14  contact_14_514
timestamp 1644969367
transform 1 0 3932 0 1 9664
box 0 0 1 1
use contact_14  contact_14_515
timestamp 1644969367
transform 1 0 3512 0 1 9750
box 0 0 1 1
use contact_14  contact_14_516
timestamp 1644969367
transform 1 0 4268 0 1 9836
box 0 0 1 1
use contact_14  contact_14_517
timestamp 1644969367
transform 1 0 3932 0 1 9922
box 0 0 1 1
use contact_14  contact_14_518
timestamp 1644969367
transform 1 0 3428 0 1 10008
box 0 0 1 1
use contact_14  contact_14_519
timestamp 1644969367
transform 1 0 4268 0 1 10094
box 0 0 1 1
use contact_14  contact_14_520
timestamp 1644969367
transform 1 0 3932 0 1 10180
box 0 0 1 1
use contact_14  contact_14_521
timestamp 1644969367
transform 1 0 3344 0 1 10266
box 0 0 1 1
use contact_14  contact_14_522
timestamp 1644969367
transform 1 0 4268 0 1 8814
box 0 0 1 1
use contact_14  contact_14_523
timestamp 1644969367
transform 1 0 3932 0 1 8728
box 0 0 1 1
use contact_14  contact_14_524
timestamp 1644969367
transform 1 0 3260 0 1 8642
box 0 0 1 1
use contact_14  contact_14_525
timestamp 1644969367
transform 1 0 4268 0 1 8556
box 0 0 1 1
use contact_14  contact_14_526
timestamp 1644969367
transform 1 0 3848 0 1 8470
box 0 0 1 1
use contact_14  contact_14_527
timestamp 1644969367
transform 1 0 3512 0 1 8384
box 0 0 1 1
use contact_14  contact_14_528
timestamp 1644969367
transform 1 0 4268 0 1 8298
box 0 0 1 1
use contact_14  contact_14_529
timestamp 1644969367
transform 1 0 3848 0 1 8212
box 0 0 1 1
use contact_14  contact_14_530
timestamp 1644969367
transform 1 0 3428 0 1 8126
box 0 0 1 1
use contact_14  contact_14_531
timestamp 1644969367
transform 1 0 4268 0 1 6502
box 0 0 1 1
use contact_14  contact_14_532
timestamp 1644969367
transform 1 0 3848 0 1 6588
box 0 0 1 1
use contact_14  contact_14_533
timestamp 1644969367
transform 1 0 3344 0 1 6674
box 0 0 1 1
use contact_14  contact_14_534
timestamp 1644969367
transform 1 0 4268 0 1 6760
box 0 0 1 1
use contact_14  contact_14_535
timestamp 1644969367
transform 1 0 3848 0 1 6846
box 0 0 1 1
use contact_14  contact_14_536
timestamp 1644969367
transform 1 0 3260 0 1 6932
box 0 0 1 1
use contact_14  contact_14_537
timestamp 1644969367
transform 1 0 4268 0 1 7018
box 0 0 1 1
use contact_14  contact_14_538
timestamp 1644969367
transform 1 0 3764 0 1 7104
box 0 0 1 1
use contact_14  contact_14_539
timestamp 1644969367
transform 1 0 3512 0 1 7190
box 0 0 1 1
use contact_14  contact_14_540
timestamp 1644969367
transform 1 0 4268 0 1 5738
box 0 0 1 1
use contact_14  contact_14_541
timestamp 1644969367
transform 1 0 3764 0 1 5652
box 0 0 1 1
use contact_14  contact_14_542
timestamp 1644969367
transform 1 0 3428 0 1 5566
box 0 0 1 1
use contact_14  contact_14_543
timestamp 1644969367
transform 1 0 4268 0 1 5480
box 0 0 1 1
use contact_14  contact_14_544
timestamp 1644969367
transform 1 0 3764 0 1 5394
box 0 0 1 1
use contact_14  contact_14_545
timestamp 1644969367
transform 1 0 3344 0 1 5308
box 0 0 1 1
use contact_14  contact_14_546
timestamp 1644969367
transform 1 0 4268 0 1 5222
box 0 0 1 1
use contact_14  contact_14_547
timestamp 1644969367
transform 1 0 3764 0 1 5136
box 0 0 1 1
use contact_14  contact_14_548
timestamp 1644969367
transform 1 0 3260 0 1 5050
box 0 0 1 1
use contact_14  contact_14_549
timestamp 1644969367
transform 1 0 4268 0 1 3426
box 0 0 1 1
use contact_14  contact_14_550
timestamp 1644969367
transform 1 0 3680 0 1 3512
box 0 0 1 1
use contact_14  contact_14_551
timestamp 1644969367
transform 1 0 3512 0 1 3598
box 0 0 1 1
use contact_14  contact_14_552
timestamp 1644969367
transform 1 0 4268 0 1 3684
box 0 0 1 1
use contact_14  contact_14_553
timestamp 1644969367
transform 1 0 3680 0 1 3770
box 0 0 1 1
use contact_14  contact_14_554
timestamp 1644969367
transform 1 0 3428 0 1 3856
box 0 0 1 1
use contact_14  contact_14_555
timestamp 1644969367
transform 1 0 4268 0 1 3942
box 0 0 1 1
use contact_14  contact_14_556
timestamp 1644969367
transform 1 0 3680 0 1 4028
box 0 0 1 1
use contact_14  contact_14_557
timestamp 1644969367
transform 1 0 3344 0 1 4114
box 0 0 1 1
use contact_14  contact_14_558
timestamp 1644969367
transform 1 0 4268 0 1 2662
box 0 0 1 1
use contact_14  contact_14_559
timestamp 1644969367
transform 1 0 3680 0 1 2576
box 0 0 1 1
use contact_14  contact_14_560
timestamp 1644969367
transform 1 0 3260 0 1 2490
box 0 0 1 1
use contact_14  contact_14_561
timestamp 1644969367
transform 1 0 4268 0 1 2404
box 0 0 1 1
use contact_14  contact_14_562
timestamp 1644969367
transform 1 0 3596 0 1 2318
box 0 0 1 1
use contact_14  contact_14_563
timestamp 1644969367
transform 1 0 3512 0 1 2232
box 0 0 1 1
use contact_14  contact_14_564
timestamp 1644969367
transform 1 0 4268 0 1 2146
box 0 0 1 1
use contact_14  contact_14_565
timestamp 1644969367
transform 1 0 3596 0 1 2060
box 0 0 1 1
use contact_14  contact_14_566
timestamp 1644969367
transform 1 0 3428 0 1 1974
box 0 0 1 1
use contact_14  contact_14_567
timestamp 1644969367
transform 1 0 4268 0 1 350
box 0 0 1 1
use contact_14  contact_14_568
timestamp 1644969367
transform 1 0 3596 0 1 436
box 0 0 1 1
use contact_14  contact_14_569
timestamp 1644969367
transform 1 0 3344 0 1 522
box 0 0 1 1
use contact_14  contact_14_570
timestamp 1644969367
transform 1 0 4268 0 1 608
box 0 0 1 1
use contact_14  contact_14_571
timestamp 1644969367
transform 1 0 3596 0 1 694
box 0 0 1 1
use contact_14  contact_14_572
timestamp 1644969367
transform 1 0 3260 0 1 780
box 0 0 1 1
use contact_14  contact_14_573
timestamp 1644969367
transform 1 0 588 0 1 28408
box 0 0 1 1
use contact_17  contact_17_148
timestamp 1644969367
transform 1 0 952 0 1 28408
box 0 0 1 1
use contact_14  contact_14_574
timestamp 1644969367
transform 1 0 504 0 1 26952
box 0 0 1 1
use contact_17  contact_17_149
timestamp 1644969367
transform 1 0 868 0 1 26952
box 0 0 1 1
use contact_14  contact_14_575
timestamp 1644969367
transform 1 0 420 0 1 25328
box 0 0 1 1
use contact_17  contact_17_150
timestamp 1644969367
transform 1 0 784 0 1 25328
box 0 0 1 1
use contact_14  contact_14_576
timestamp 1644969367
transform 1 0 336 0 1 13012
box 0 0 1 1
use contact_17  contact_17_151
timestamp 1644969367
transform 1 0 952 0 1 13012
box 0 0 1 1
use contact_14  contact_14_577
timestamp 1644969367
transform 1 0 252 0 1 11556
box 0 0 1 1
use contact_17  contact_17_152
timestamp 1644969367
transform 1 0 868 0 1 11556
box 0 0 1 1
use contact_14  contact_14_578
timestamp 1644969367
transform 1 0 168 0 1 9932
box 0 0 1 1
use contact_17  contact_17_153
timestamp 1644969367
transform 1 0 784 0 1 9932
box 0 0 1 1
use contact_14  contact_14_579
timestamp 1644969367
transform 1 0 84 0 1 2320
box 0 0 1 1
use contact_17  contact_17_154
timestamp 1644969367
transform 1 0 1300 0 1 2320
box 0 0 1 1
use contact_14  contact_14_580
timestamp 1644969367
transform 1 0 0 0 1 696
box 0 0 1 1
use contact_17  contact_17_155
timestamp 1644969367
transform 1 0 1216 0 1 696
box 0 0 1 1
use dec_cell3_2r1w  dec_cell3_2r1w_0
timestamp 1644969367
transform 1 0 4958 0 -1 98432
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_1
timestamp 1644969367
transform 1 0 4958 0 1 95356
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_2
timestamp 1644969367
transform 1 0 4958 0 -1 95356
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_3
timestamp 1644969367
transform 1 0 4958 0 1 92280
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_4
timestamp 1644969367
transform 1 0 4958 0 -1 92280
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_5
timestamp 1644969367
transform 1 0 4958 0 1 89204
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_6
timestamp 1644969367
transform 1 0 4958 0 -1 89204
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_7
timestamp 1644969367
transform 1 0 4958 0 1 86128
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_8
timestamp 1644969367
transform 1 0 4958 0 -1 86128
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_9
timestamp 1644969367
transform 1 0 4958 0 1 83052
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_10
timestamp 1644969367
transform 1 0 4958 0 -1 83052
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_11
timestamp 1644969367
transform 1 0 4958 0 1 79976
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_12
timestamp 1644969367
transform 1 0 4958 0 -1 79976
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_13
timestamp 1644969367
transform 1 0 4958 0 1 76900
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_14
timestamp 1644969367
transform 1 0 4958 0 -1 76900
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_15
timestamp 1644969367
transform 1 0 4958 0 1 73824
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_16
timestamp 1644969367
transform 1 0 4958 0 -1 73824
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_17
timestamp 1644969367
transform 1 0 4958 0 1 70748
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_18
timestamp 1644969367
transform 1 0 4958 0 -1 70748
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_19
timestamp 1644969367
transform 1 0 4958 0 1 67672
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_20
timestamp 1644969367
transform 1 0 4958 0 -1 67672
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_21
timestamp 1644969367
transform 1 0 4958 0 1 64596
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_22
timestamp 1644969367
transform 1 0 4958 0 -1 64596
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_23
timestamp 1644969367
transform 1 0 4958 0 1 61520
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_24
timestamp 1644969367
transform 1 0 4958 0 -1 61520
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_25
timestamp 1644969367
transform 1 0 4958 0 1 58444
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_26
timestamp 1644969367
transform 1 0 4958 0 -1 58444
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_27
timestamp 1644969367
transform 1 0 4958 0 1 55368
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_28
timestamp 1644969367
transform 1 0 4958 0 -1 55368
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_29
timestamp 1644969367
transform 1 0 4958 0 1 52292
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_30
timestamp 1644969367
transform 1 0 4958 0 -1 52292
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_31
timestamp 1644969367
transform 1 0 4958 0 1 49216
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_32
timestamp 1644969367
transform 1 0 4958 0 -1 49216
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_33
timestamp 1644969367
transform 1 0 4958 0 1 46140
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_34
timestamp 1644969367
transform 1 0 4958 0 -1 46140
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_35
timestamp 1644969367
transform 1 0 4958 0 1 43064
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_36
timestamp 1644969367
transform 1 0 4958 0 -1 43064
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_37
timestamp 1644969367
transform 1 0 4958 0 1 39988
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_38
timestamp 1644969367
transform 1 0 4958 0 -1 39988
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_39
timestamp 1644969367
transform 1 0 4958 0 1 36912
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_40
timestamp 1644969367
transform 1 0 4958 0 -1 36912
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_41
timestamp 1644969367
transform 1 0 4958 0 1 33836
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_42
timestamp 1644969367
transform 1 0 4958 0 -1 33836
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_43
timestamp 1644969367
transform 1 0 4958 0 1 30760
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_44
timestamp 1644969367
transform 1 0 4958 0 -1 30760
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_45
timestamp 1644969367
transform 1 0 4958 0 1 27684
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_46
timestamp 1644969367
transform 1 0 4958 0 -1 27684
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_47
timestamp 1644969367
transform 1 0 4958 0 1 24608
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_48
timestamp 1644969367
transform 1 0 4958 0 -1 24608
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_49
timestamp 1644969367
transform 1 0 4958 0 1 21532
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_50
timestamp 1644969367
transform 1 0 4958 0 -1 21532
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_51
timestamp 1644969367
transform 1 0 4958 0 1 18456
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_52
timestamp 1644969367
transform 1 0 4958 0 -1 18456
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_53
timestamp 1644969367
transform 1 0 4958 0 1 15380
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_54
timestamp 1644969367
transform 1 0 4958 0 -1 15380
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_55
timestamp 1644969367
transform 1 0 4958 0 1 12304
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_56
timestamp 1644969367
transform 1 0 4958 0 -1 12304
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_57
timestamp 1644969367
transform 1 0 4958 0 1 9228
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_58
timestamp 1644969367
transform 1 0 4958 0 -1 9228
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_59
timestamp 1644969367
transform 1 0 4958 0 1 6152
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_60
timestamp 1644969367
transform 1 0 4958 0 -1 6152
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_61
timestamp 1644969367
transform 1 0 4958 0 1 3076
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_62
timestamp 1644969367
transform 1 0 4958 0 -1 3076
box 0 -42 1494 1616
use dec_cell3_2r1w  dec_cell3_2r1w_63
timestamp 1644969367
transform 1 0 4958 0 1 0
box 0 -42 1494 1616
use hierarchical_predecode3x8  hierarchical_predecode3x8_0
timestamp 1644969367
transform 1 0 718 0 1 24632
box 0 -37 2512 12357
use hierarchical_predecode3x8  hierarchical_predecode3x8_1
timestamp 1644969367
transform 1 0 718 0 1 9236
box 0 -37 2512 12357
use hierarchical_predecode2x4  hierarchical_predecode2x4_0
timestamp 1644969367
transform 1 0 1150 0 1 0
box 0 -37 2080 6197
<< labels >>
rlabel metal2 s 18 0 46 36952 4 addr_0
rlabel metal2 s 102 0 130 36952 4 addr_1
rlabel metal2 s 186 0 214 36952 4 addr_2
rlabel metal2 s 270 0 298 36952 4 addr_3
rlabel metal2 s 354 0 382 36952 4 addr_4
rlabel metal2 s 438 0 466 36952 4 addr_5
rlabel metal2 s 522 0 550 36952 4 addr_6
rlabel metal2 s 606 0 634 36952 4 addr_7
rlabel metal1 s 6376 848 6452 876 4 decode0_0
rlabel metal1 s 6168 702 6452 730 4 decode1_0
rlabel metal1 s 6086 580 6452 608 4 decode2_0
rlabel metal1 s 6376 2200 6452 2228 4 decode0_1
rlabel metal1 s 6168 2346 6452 2374 4 decode1_1
rlabel metal1 s 6086 2468 6452 2496 4 decode2_1
rlabel metal1 s 6376 3924 6452 3952 4 decode0_2
rlabel metal1 s 6168 3778 6452 3806 4 decode1_2
rlabel metal1 s 6086 3656 6452 3684 4 decode2_2
rlabel metal1 s 6376 5276 6452 5304 4 decode0_3
rlabel metal1 s 6168 5422 6452 5450 4 decode1_3
rlabel metal1 s 6086 5544 6452 5572 4 decode2_3
rlabel metal1 s 6376 7000 6452 7028 4 decode0_4
rlabel metal1 s 6168 6854 6452 6882 4 decode1_4
rlabel metal1 s 6086 6732 6452 6760 4 decode2_4
rlabel metal1 s 6376 8352 6452 8380 4 decode0_5
rlabel metal1 s 6168 8498 6452 8526 4 decode1_5
rlabel metal1 s 6086 8620 6452 8648 4 decode2_5
rlabel metal1 s 6376 10076 6452 10104 4 decode0_6
rlabel metal1 s 6168 9930 6452 9958 4 decode1_6
rlabel metal1 s 6086 9808 6452 9836 4 decode2_6
rlabel metal1 s 6376 11428 6452 11456 4 decode0_7
rlabel metal1 s 6168 11574 6452 11602 4 decode1_7
rlabel metal1 s 6086 11696 6452 11724 4 decode2_7
rlabel metal1 s 6376 13152 6452 13180 4 decode0_8
rlabel metal1 s 6168 13006 6452 13034 4 decode1_8
rlabel metal1 s 6086 12884 6452 12912 4 decode2_8
rlabel metal1 s 6376 14504 6452 14532 4 decode0_9
rlabel metal1 s 6168 14650 6452 14678 4 decode1_9
rlabel metal1 s 6086 14772 6452 14800 4 decode2_9
rlabel metal1 s 6376 16228 6452 16256 4 decode0_10
rlabel metal1 s 6168 16082 6452 16110 4 decode1_10
rlabel metal1 s 6086 15960 6452 15988 4 decode2_10
rlabel metal1 s 6376 17580 6452 17608 4 decode0_11
rlabel metal1 s 6168 17726 6452 17754 4 decode1_11
rlabel metal1 s 6086 17848 6452 17876 4 decode2_11
rlabel metal1 s 6376 19304 6452 19332 4 decode0_12
rlabel metal1 s 6168 19158 6452 19186 4 decode1_12
rlabel metal1 s 6086 19036 6452 19064 4 decode2_12
rlabel metal1 s 6376 20656 6452 20684 4 decode0_13
rlabel metal1 s 6168 20802 6452 20830 4 decode1_13
rlabel metal1 s 6086 20924 6452 20952 4 decode2_13
rlabel metal1 s 6376 22380 6452 22408 4 decode0_14
rlabel metal1 s 6168 22234 6452 22262 4 decode1_14
rlabel metal1 s 6086 22112 6452 22140 4 decode2_14
rlabel metal1 s 6376 23732 6452 23760 4 decode0_15
rlabel metal1 s 6168 23878 6452 23906 4 decode1_15
rlabel metal1 s 6086 24000 6452 24028 4 decode2_15
rlabel metal1 s 6376 25456 6452 25484 4 decode0_16
rlabel metal1 s 6168 25310 6452 25338 4 decode1_16
rlabel metal1 s 6086 25188 6452 25216 4 decode2_16
rlabel metal1 s 6376 26808 6452 26836 4 decode0_17
rlabel metal1 s 6168 26954 6452 26982 4 decode1_17
rlabel metal1 s 6086 27076 6452 27104 4 decode2_17
rlabel metal1 s 6376 28532 6452 28560 4 decode0_18
rlabel metal1 s 6168 28386 6452 28414 4 decode1_18
rlabel metal1 s 6086 28264 6452 28292 4 decode2_18
rlabel metal1 s 6376 29884 6452 29912 4 decode0_19
rlabel metal1 s 6168 30030 6452 30058 4 decode1_19
rlabel metal1 s 6086 30152 6452 30180 4 decode2_19
rlabel metal1 s 6376 31608 6452 31636 4 decode0_20
rlabel metal1 s 6168 31462 6452 31490 4 decode1_20
rlabel metal1 s 6086 31340 6452 31368 4 decode2_20
rlabel metal1 s 6376 32960 6452 32988 4 decode0_21
rlabel metal1 s 6168 33106 6452 33134 4 decode1_21
rlabel metal1 s 6086 33228 6452 33256 4 decode2_21
rlabel metal1 s 6376 34684 6452 34712 4 decode0_22
rlabel metal1 s 6168 34538 6452 34566 4 decode1_22
rlabel metal1 s 6086 34416 6452 34444 4 decode2_22
rlabel metal1 s 6376 36036 6452 36064 4 decode0_23
rlabel metal1 s 6168 36182 6452 36210 4 decode1_23
rlabel metal1 s 6086 36304 6452 36332 4 decode2_23
rlabel metal1 s 6376 37760 6452 37788 4 decode0_24
rlabel metal1 s 6168 37614 6452 37642 4 decode1_24
rlabel metal1 s 6086 37492 6452 37520 4 decode2_24
rlabel metal1 s 6376 39112 6452 39140 4 decode0_25
rlabel metal1 s 6168 39258 6452 39286 4 decode1_25
rlabel metal1 s 6086 39380 6452 39408 4 decode2_25
rlabel metal1 s 6376 40836 6452 40864 4 decode0_26
rlabel metal1 s 6168 40690 6452 40718 4 decode1_26
rlabel metal1 s 6086 40568 6452 40596 4 decode2_26
rlabel metal1 s 6376 42188 6452 42216 4 decode0_27
rlabel metal1 s 6168 42334 6452 42362 4 decode1_27
rlabel metal1 s 6086 42456 6452 42484 4 decode2_27
rlabel metal1 s 6376 43912 6452 43940 4 decode0_28
rlabel metal1 s 6168 43766 6452 43794 4 decode1_28
rlabel metal1 s 6086 43644 6452 43672 4 decode2_28
rlabel metal1 s 6376 45264 6452 45292 4 decode0_29
rlabel metal1 s 6168 45410 6452 45438 4 decode1_29
rlabel metal1 s 6086 45532 6452 45560 4 decode2_29
rlabel metal1 s 6376 46988 6452 47016 4 decode0_30
rlabel metal1 s 6168 46842 6452 46870 4 decode1_30
rlabel metal1 s 6086 46720 6452 46748 4 decode2_30
rlabel metal1 s 6376 48340 6452 48368 4 decode0_31
rlabel metal1 s 6168 48486 6452 48514 4 decode1_31
rlabel metal1 s 6086 48608 6452 48636 4 decode2_31
rlabel metal1 s 6376 50064 6452 50092 4 decode0_32
rlabel metal1 s 6168 49918 6452 49946 4 decode1_32
rlabel metal1 s 6086 49796 6452 49824 4 decode2_32
rlabel metal1 s 6376 51416 6452 51444 4 decode0_33
rlabel metal1 s 6168 51562 6452 51590 4 decode1_33
rlabel metal1 s 6086 51684 6452 51712 4 decode2_33
rlabel metal1 s 6376 53140 6452 53168 4 decode0_34
rlabel metal1 s 6168 52994 6452 53022 4 decode1_34
rlabel metal1 s 6086 52872 6452 52900 4 decode2_34
rlabel metal1 s 6376 54492 6452 54520 4 decode0_35
rlabel metal1 s 6168 54638 6452 54666 4 decode1_35
rlabel metal1 s 6086 54760 6452 54788 4 decode2_35
rlabel metal1 s 6376 56216 6452 56244 4 decode0_36
rlabel metal1 s 6168 56070 6452 56098 4 decode1_36
rlabel metal1 s 6086 55948 6452 55976 4 decode2_36
rlabel metal1 s 6376 57568 6452 57596 4 decode0_37
rlabel metal1 s 6168 57714 6452 57742 4 decode1_37
rlabel metal1 s 6086 57836 6452 57864 4 decode2_37
rlabel metal1 s 6376 59292 6452 59320 4 decode0_38
rlabel metal1 s 6168 59146 6452 59174 4 decode1_38
rlabel metal1 s 6086 59024 6452 59052 4 decode2_38
rlabel metal1 s 6376 60644 6452 60672 4 decode0_39
rlabel metal1 s 6168 60790 6452 60818 4 decode1_39
rlabel metal1 s 6086 60912 6452 60940 4 decode2_39
rlabel metal1 s 6376 62368 6452 62396 4 decode0_40
rlabel metal1 s 6168 62222 6452 62250 4 decode1_40
rlabel metal1 s 6086 62100 6452 62128 4 decode2_40
rlabel metal1 s 6376 63720 6452 63748 4 decode0_41
rlabel metal1 s 6168 63866 6452 63894 4 decode1_41
rlabel metal1 s 6086 63988 6452 64016 4 decode2_41
rlabel metal1 s 6376 65444 6452 65472 4 decode0_42
rlabel metal1 s 6168 65298 6452 65326 4 decode1_42
rlabel metal1 s 6086 65176 6452 65204 4 decode2_42
rlabel metal1 s 6376 66796 6452 66824 4 decode0_43
rlabel metal1 s 6168 66942 6452 66970 4 decode1_43
rlabel metal1 s 6086 67064 6452 67092 4 decode2_43
rlabel metal1 s 6376 68520 6452 68548 4 decode0_44
rlabel metal1 s 6168 68374 6452 68402 4 decode1_44
rlabel metal1 s 6086 68252 6452 68280 4 decode2_44
rlabel metal1 s 6376 69872 6452 69900 4 decode0_45
rlabel metal1 s 6168 70018 6452 70046 4 decode1_45
rlabel metal1 s 6086 70140 6452 70168 4 decode2_45
rlabel metal1 s 6376 71596 6452 71624 4 decode0_46
rlabel metal1 s 6168 71450 6452 71478 4 decode1_46
rlabel metal1 s 6086 71328 6452 71356 4 decode2_46
rlabel metal1 s 6376 72948 6452 72976 4 decode0_47
rlabel metal1 s 6168 73094 6452 73122 4 decode1_47
rlabel metal1 s 6086 73216 6452 73244 4 decode2_47
rlabel metal1 s 6376 74672 6452 74700 4 decode0_48
rlabel metal1 s 6168 74526 6452 74554 4 decode1_48
rlabel metal1 s 6086 74404 6452 74432 4 decode2_48
rlabel metal1 s 6376 76024 6452 76052 4 decode0_49
rlabel metal1 s 6168 76170 6452 76198 4 decode1_49
rlabel metal1 s 6086 76292 6452 76320 4 decode2_49
rlabel metal1 s 6376 77748 6452 77776 4 decode0_50
rlabel metal1 s 6168 77602 6452 77630 4 decode1_50
rlabel metal1 s 6086 77480 6452 77508 4 decode2_50
rlabel metal1 s 6376 79100 6452 79128 4 decode0_51
rlabel metal1 s 6168 79246 6452 79274 4 decode1_51
rlabel metal1 s 6086 79368 6452 79396 4 decode2_51
rlabel metal1 s 6376 80824 6452 80852 4 decode0_52
rlabel metal1 s 6168 80678 6452 80706 4 decode1_52
rlabel metal1 s 6086 80556 6452 80584 4 decode2_52
rlabel metal1 s 6376 82176 6452 82204 4 decode0_53
rlabel metal1 s 6168 82322 6452 82350 4 decode1_53
rlabel metal1 s 6086 82444 6452 82472 4 decode2_53
rlabel metal1 s 6376 83900 6452 83928 4 decode0_54
rlabel metal1 s 6168 83754 6452 83782 4 decode1_54
rlabel metal1 s 6086 83632 6452 83660 4 decode2_54
rlabel metal1 s 6376 85252 6452 85280 4 decode0_55
rlabel metal1 s 6168 85398 6452 85426 4 decode1_55
rlabel metal1 s 6086 85520 6452 85548 4 decode2_55
rlabel metal1 s 6376 86976 6452 87004 4 decode0_56
rlabel metal1 s 6168 86830 6452 86858 4 decode1_56
rlabel metal1 s 6086 86708 6452 86736 4 decode2_56
rlabel metal1 s 6376 88328 6452 88356 4 decode0_57
rlabel metal1 s 6168 88474 6452 88502 4 decode1_57
rlabel metal1 s 6086 88596 6452 88624 4 decode2_57
rlabel metal1 s 6376 90052 6452 90080 4 decode0_58
rlabel metal1 s 6168 89906 6452 89934 4 decode1_58
rlabel metal1 s 6086 89784 6452 89812 4 decode2_58
rlabel metal1 s 6376 91404 6452 91432 4 decode0_59
rlabel metal1 s 6168 91550 6452 91578 4 decode1_59
rlabel metal1 s 6086 91672 6452 91700 4 decode2_59
rlabel metal1 s 6376 93128 6452 93156 4 decode0_60
rlabel metal1 s 6168 92982 6452 93010 4 decode1_60
rlabel metal1 s 6086 92860 6452 92888 4 decode2_60
rlabel metal1 s 6376 94480 6452 94508 4 decode0_61
rlabel metal1 s 6168 94626 6452 94654 4 decode1_61
rlabel metal1 s 6086 94748 6452 94776 4 decode2_61
rlabel metal1 s 6376 96204 6452 96232 4 decode0_62
rlabel metal1 s 6168 96058 6452 96086 4 decode1_62
rlabel metal1 s 6086 95936 6452 95964 4 decode2_62
rlabel metal1 s 6376 97556 6452 97584 4 decode0_63
rlabel metal1 s 6168 97702 6452 97730 4 decode1_63
rlabel metal1 s 6086 97824 6452 97852 4 decode2_63
rlabel metal2 s 3278 0 3306 98460 4 predecode_0
rlabel metal2 s 3362 0 3390 98460 4 predecode_1
rlabel metal2 s 3446 0 3474 98460 4 predecode_2
rlabel metal2 s 3530 0 3558 98460 4 predecode_3
rlabel metal2 s 3614 0 3642 98460 4 predecode_4
rlabel metal2 s 3698 0 3726 98460 4 predecode_5
rlabel metal2 s 3782 0 3810 98460 4 predecode_6
rlabel metal2 s 3866 0 3894 98460 4 predecode_7
rlabel metal2 s 3950 0 3978 98460 4 predecode_8
rlabel metal2 s 4034 0 4062 98460 4 predecode_9
rlabel metal2 s 4118 0 4146 98460 4 predecode_10
rlabel metal2 s 4202 0 4230 98460 4 predecode_11
rlabel metal2 s 4286 0 4314 98460 4 predecode_12
rlabel metal2 s 4370 0 4398 98460 4 predecode_13
rlabel metal2 s 4454 0 4482 98460 4 predecode_14
rlabel metal2 s 4538 0 4566 98460 4 predecode_15
rlabel metal2 s 4622 0 4650 98460 4 predecode_16
rlabel metal2 s 4706 0 4734 98460 4 predecode_17
rlabel metal2 s 4790 0 4818 98460 4 predecode_18
rlabel metal2 s 4874 0 4902 98460 4 predecode_19
rlabel metal3 s 2084 10739 2216 10813 4 vdd
rlabel metal3 s 6400 13805 6532 13879 4 vdd
rlabel metal3 s 6400 69173 6532 69247 4 vdd
rlabel metal3 s 1044 35375 1176 35449 4 vdd
rlabel metal3 s 1044 13819 1176 13893 4 vdd
rlabel metal3 s 6400 53793 6532 53867 4 vdd
rlabel metal3 s 6466 53830 6466 53830 4 vdd
rlabel metal3 s 6400 47641 6532 47715 4 vdd
rlabel metal3 s 6400 26109 6532 26183 4 vdd
rlabel metal3 s 2084 35375 2216 35449 4 vdd
rlabel metal3 s 6400 32261 6532 32335 4 vdd
rlabel metal3 s 2264 1503 2396 1577 4 vdd
rlabel metal3 s 6400 7653 6532 7727 4 vdd
rlabel metal3 s 6400 38413 6532 38487 4 vdd
rlabel metal3 s 6400 72249 6532 72323 4 vdd
rlabel metal3 s 1044 10739 1176 10813 4 vdd
rlabel metal3 s 6400 35337 6532 35411 4 vdd
rlabel metal3 s 1044 26135 1176 26209 4 vdd
rlabel metal3 s 2084 29215 2216 29289 4 vdd
rlabel metal3 s 2084 19979 2216 20053 4 vdd
rlabel metal3 s 6400 23033 6532 23107 4 vdd
rlabel metal3 s 1044 29215 1176 29289 4 vdd
rlabel metal3 s 6400 84553 6532 84627 4 vdd
rlabel metal3 s 6400 96857 6532 96931 4 vdd
rlabel metal3 s 6400 16881 6532 16955 4 vdd
rlabel metal3 s 6400 44565 6532 44639 4 vdd
rlabel metal3 s 6466 44602 6466 44602 4 vdd
rlabel metal3 s 6400 81477 6532 81551 4 vdd
rlabel metal3 s 6400 4577 6532 4651 4 vdd
rlabel metal3 s 1044 19979 1176 20053 4 vdd
rlabel metal3 s 6400 50717 6532 50791 4 vdd
rlabel metal3 s 1392 1503 1524 1577 4 vdd
rlabel metal3 s 6466 50754 6466 50754 4 vdd
rlabel metal3 s 1044 16899 1176 16973 4 vdd
rlabel metal3 s 6400 93781 6532 93855 4 vdd
rlabel metal3 s 6400 1501 6532 1575 4 vdd
rlabel metal3 s 6466 1538 6466 1538 4 vdd
rlabel metal3 s 6400 75325 6532 75399 4 vdd
rlabel metal3 s 6400 87629 6532 87703 4 vdd
rlabel metal3 s 2084 13819 2216 13893 4 vdd
rlabel metal3 s 6400 19957 6532 20031 4 vdd
rlabel metal3 s 2084 26135 2216 26209 4 vdd
rlabel metal3 s 6400 10729 6532 10803 4 vdd
rlabel metal3 s 1044 32295 1176 32369 4 vdd
rlabel metal3 s 6400 78401 6532 78475 4 vdd
rlabel metal3 s 6400 41489 6532 41563 4 vdd
rlabel metal3 s 6400 90705 6532 90779 4 vdd
rlabel metal3 s 6466 90742 6466 90742 4 vdd
rlabel metal3 s 6400 56869 6532 56943 4 vdd
rlabel metal3 s 1392 4583 1524 4657 4 vdd
rlabel metal3 s 2264 4583 2396 4657 4 vdd
rlabel metal3 s 6400 29185 6532 29259 4 vdd
rlabel metal3 s 6400 63021 6532 63095 4 vdd
rlabel metal3 s 6400 66097 6532 66171 4 vdd
rlabel metal3 s 2084 32295 2216 32369 4 vdd
rlabel metal3 s 6400 59945 6532 60019 4 vdd
rlabel metal3 s 2084 16899 2216 16973 4 vdd
rlabel metal3 s 6466 10766 6466 10766 4 vdd
rlabel metal3 s 6400 55331 6532 55405 4 gnd
rlabel metal3 s 6400 64559 6532 64633 4 gnd
rlabel metal3 s 6400 73787 6532 73861 4 gnd
rlabel metal3 s 2264 3043 2396 3117 4 gnd
rlabel metal3 s 6400 43027 6532 43101 4 gnd
rlabel metal3 s 6400 52255 6532 52329 4 gnd
rlabel metal3 s 1392 -37 1524 37 4 gnd
rlabel metal3 s 2264 -37 2396 37 4 gnd
rlabel metal3 s 6400 92243 6532 92317 4 gnd
rlabel metal3 s 6400 18419 6532 18493 4 gnd
rlabel metal3 s 2084 36915 2216 36989 4 gnd
rlabel metal3 s 2084 27675 2216 27749 4 gnd
rlabel metal3 s 6400 15343 6532 15417 4 gnd
rlabel metal3 s 6400 27647 6532 27721 4 gnd
rlabel metal3 s 1044 21519 1176 21593 4 gnd
rlabel metal3 s 6400 3039 6532 3113 4 gnd
rlabel metal3 s 6400 36875 6532 36949 4 gnd
rlabel metal3 s 6400 79939 6532 80013 4 gnd
rlabel metal3 s 2084 21519 2216 21593 4 gnd
rlabel metal3 s 1044 12279 1176 12353 4 gnd
rlabel metal3 s 1044 9199 1176 9273 4 gnd
rlabel metal3 s 1044 30755 1176 30829 4 gnd
rlabel metal3 s 6400 9191 6532 9265 4 gnd
rlabel metal3 s 6400 46103 6532 46177 4 gnd
rlabel metal3 s 2084 18439 2216 18513 4 gnd
rlabel metal3 s 6400 21495 6532 21569 4 gnd
rlabel metal3 s 2084 9199 2216 9273 4 gnd
rlabel metal3 s 6400 6115 6532 6189 4 gnd
rlabel metal3 s 6400 39951 6532 40025 4 gnd
rlabel metal3 s 6400 67635 6532 67709 4 gnd
rlabel metal3 s 2084 24595 2216 24669 4 gnd
rlabel metal3 s 1044 18439 1176 18513 4 gnd
rlabel metal3 s 2084 33835 2216 33909 4 gnd
rlabel metal3 s 6400 33799 6532 33873 4 gnd
rlabel metal3 s 6400 49179 6532 49253 4 gnd
rlabel metal3 s 2084 12279 2216 12353 4 gnd
rlabel metal3 s 6400 58407 6532 58481 4 gnd
rlabel metal3 s 6400 24571 6532 24645 4 gnd
rlabel metal3 s 6400 70711 6532 70785 4 gnd
rlabel metal3 s 6400 30723 6532 30797 4 gnd
rlabel metal3 s 6400 61483 6532 61557 4 gnd
rlabel metal3 s 6400 -37 6532 37 4 gnd
rlabel metal3 s 6400 83015 6532 83089 4 gnd
rlabel metal3 s 6400 98395 6532 98469 4 gnd
rlabel metal3 s 6400 12267 6532 12341 4 gnd
rlabel metal3 s 1044 33835 1176 33909 4 gnd
rlabel metal3 s 1044 24595 1176 24669 4 gnd
rlabel metal3 s 6400 76863 6532 76937 4 gnd
rlabel metal3 s 1044 36915 1176 36989 4 gnd
rlabel metal3 s 1044 15359 1176 15433 4 gnd
rlabel metal3 s 6400 86091 6532 86165 4 gnd
rlabel metal3 s 6400 89167 6532 89241 4 gnd
rlabel metal3 s 1044 27675 1176 27749 4 gnd
rlabel metal3 s 2084 30755 2216 30829 4 gnd
rlabel metal3 s 1392 3043 1524 3117 4 gnd
rlabel metal3 s 1392 6123 1524 6197 4 gnd
rlabel metal3 s 2084 15359 2216 15433 4 gnd
rlabel metal3 s 6400 95319 6532 95393 4 gnd
rlabel metal3 s 2264 6123 2396 6197 4 gnd
<< properties >>
string FIXED_BBOX 6400 -37 6532 0
string GDS_FILE sram_0rw2r1w_32_128_sky130A.gds
string GDS_END 3054162
string GDS_START 2861588
<< end >>
