magic
tech sky130A
magscale 1 2
timestamp 1643678851
<< checkpaint >>
rect -1296 -1277 2256 2857
<< locali >>
rect 0 1523 960 1557
rect 430 745 464 1279
rect 430 711 690 745
rect 788 711 822 745
rect 329 505 395 571
rect 196 381 262 447
rect 63 257 129 323
rect 0 -17 960 17
use pinv  pinv_0
timestamp 1643678851
transform 1 0 609 0 1 0
box -36 -17 387 1597
use pnand3  pnand3_0
timestamp 1643678851
transform 1 0 0 0 1 0
box -36 -17 645 1597
<< labels >>
rlabel locali s 805 728 805 728 4 Z
rlabel locali s 96 290 96 290 4 A
rlabel locali s 229 414 229 414 4 B
rlabel locali s 362 538 362 538 4 C
rlabel locali s 480 0 480 0 4 gnd
rlabel locali s 480 1540 480 1540 4 vdd
<< properties >>
string FIXED_BBOX 0 0 960 1540
string GDS_FILE sram_0rw2r1w_16_128_sky130A.gds
string GDS_END 1879362
string GDS_START 1878244
<< end >>
