magic
tech sky130A
magscale 1 2
timestamp 1643671299
<< checkpaint >>
rect -1260 -1228 26186 3058
<< poly >>
rect 374 221 404 318
rect 1152 279 1182 318
rect 1134 263 1200 279
rect 1134 229 1150 263
rect 1184 229 1200 263
rect 356 205 422 221
rect 1134 213 1200 229
rect 1930 221 1960 318
rect 2708 279 2738 318
rect 2690 263 2756 279
rect 2690 229 2706 263
rect 2740 229 2756 263
rect 356 171 372 205
rect 406 171 422 205
rect 356 155 422 171
rect 1912 205 1978 221
rect 2690 213 2756 229
rect 3486 221 3516 318
rect 4264 279 4294 318
rect 4246 263 4312 279
rect 4246 229 4262 263
rect 4296 229 4312 263
rect 1912 171 1928 205
rect 1962 171 1978 205
rect 1912 155 1978 171
rect 3468 205 3534 221
rect 4246 213 4312 229
rect 5042 221 5072 318
rect 5820 279 5850 318
rect 5802 263 5868 279
rect 5802 229 5818 263
rect 5852 229 5868 263
rect 3468 171 3484 205
rect 3518 171 3534 205
rect 3468 155 3534 171
rect 5024 205 5090 221
rect 5802 213 5868 229
rect 6598 221 6628 318
rect 7376 279 7406 318
rect 7358 263 7424 279
rect 7358 229 7374 263
rect 7408 229 7424 263
rect 5024 171 5040 205
rect 5074 171 5090 205
rect 5024 155 5090 171
rect 6580 205 6646 221
rect 7358 213 7424 229
rect 8154 221 8184 318
rect 8932 279 8962 318
rect 8914 263 8980 279
rect 8914 229 8930 263
rect 8964 229 8980 263
rect 6580 171 6596 205
rect 6630 171 6646 205
rect 6580 155 6646 171
rect 8136 205 8202 221
rect 8914 213 8980 229
rect 9710 221 9740 318
rect 10488 279 10518 318
rect 10470 263 10536 279
rect 10470 229 10486 263
rect 10520 229 10536 263
rect 8136 171 8152 205
rect 8186 171 8202 205
rect 8136 155 8202 171
rect 9692 205 9758 221
rect 10470 213 10536 229
rect 11266 221 11296 318
rect 12044 279 12074 318
rect 12026 263 12092 279
rect 12026 229 12042 263
rect 12076 229 12092 263
rect 9692 171 9708 205
rect 9742 171 9758 205
rect 9692 155 9758 171
rect 11248 205 11314 221
rect 12026 213 12092 229
rect 12822 221 12852 318
rect 13600 279 13630 318
rect 13582 263 13648 279
rect 13582 229 13598 263
rect 13632 229 13648 263
rect 11248 171 11264 205
rect 11298 171 11314 205
rect 11248 155 11314 171
rect 12804 205 12870 221
rect 13582 213 13648 229
rect 14378 221 14408 318
rect 15156 279 15186 318
rect 15138 263 15204 279
rect 15138 229 15154 263
rect 15188 229 15204 263
rect 12804 171 12820 205
rect 12854 171 12870 205
rect 12804 155 12870 171
rect 14360 205 14426 221
rect 15138 213 15204 229
rect 15934 221 15964 318
rect 16712 279 16742 318
rect 16694 263 16760 279
rect 16694 229 16710 263
rect 16744 229 16760 263
rect 14360 171 14376 205
rect 14410 171 14426 205
rect 14360 155 14426 171
rect 15916 205 15982 221
rect 16694 213 16760 229
rect 17490 221 17520 318
rect 18268 279 18298 318
rect 18250 263 18316 279
rect 18250 229 18266 263
rect 18300 229 18316 263
rect 15916 171 15932 205
rect 15966 171 15982 205
rect 15916 155 15982 171
rect 17472 205 17538 221
rect 18250 213 18316 229
rect 19046 221 19076 318
rect 19824 279 19854 318
rect 19806 263 19872 279
rect 19806 229 19822 263
rect 19856 229 19872 263
rect 17472 171 17488 205
rect 17522 171 17538 205
rect 17472 155 17538 171
rect 19028 205 19094 221
rect 19806 213 19872 229
rect 20602 221 20632 318
rect 21380 279 21410 318
rect 21362 263 21428 279
rect 21362 229 21378 263
rect 21412 229 21428 263
rect 19028 171 19044 205
rect 19078 171 19094 205
rect 19028 155 19094 171
rect 20584 205 20650 221
rect 21362 213 21428 229
rect 22158 221 22188 318
rect 22936 279 22966 318
rect 22918 263 22984 279
rect 22918 229 22934 263
rect 22968 229 22984 263
rect 20584 171 20600 205
rect 20634 171 20650 205
rect 20584 155 20650 171
rect 22140 205 22206 221
rect 22918 213 22984 229
rect 23714 221 23744 318
rect 24492 279 24522 318
rect 24474 263 24540 279
rect 24474 229 24490 263
rect 24524 229 24540 263
rect 22140 171 22156 205
rect 22190 171 22206 205
rect 22140 155 22206 171
rect 23696 205 23762 221
rect 24474 213 24540 229
rect 23696 171 23712 205
rect 23746 171 23762 205
rect 23696 155 23762 171
<< polycont >>
rect 1150 229 1184 263
rect 2706 229 2740 263
rect 372 171 406 205
rect 4262 229 4296 263
rect 1928 171 1962 205
rect 5818 229 5852 263
rect 3484 171 3518 205
rect 7374 229 7408 263
rect 5040 171 5074 205
rect 8930 229 8964 263
rect 6596 171 6630 205
rect 10486 229 10520 263
rect 8152 171 8186 205
rect 12042 229 12076 263
rect 9708 171 9742 205
rect 13598 229 13632 263
rect 11264 171 11298 205
rect 15154 229 15188 263
rect 12820 171 12854 205
rect 16710 229 16744 263
rect 14376 171 14410 205
rect 18266 229 18300 263
rect 15932 171 15966 205
rect 19822 229 19856 263
rect 17488 171 17522 205
rect 21378 229 21412 263
rect 19044 171 19078 205
rect 22934 229 22968 263
rect 20600 171 20634 205
rect 24490 229 24524 263
rect 22156 171 22190 205
rect 23712 171 23746 205
<< locali >>
rect 1134 263 1200 279
rect 1134 229 1150 263
rect 1184 229 1200 263
rect 356 205 422 221
rect 1134 213 1200 229
rect 2690 263 2756 279
rect 2690 229 2706 263
rect 2740 229 2756 263
rect 356 171 372 205
rect 406 171 422 205
rect 356 155 422 171
rect 1912 205 1978 221
rect 2690 213 2756 229
rect 4246 263 4312 279
rect 4246 229 4262 263
rect 4296 229 4312 263
rect 1912 171 1928 205
rect 1962 171 1978 205
rect 1912 155 1978 171
rect 3468 205 3534 221
rect 4246 213 4312 229
rect 5802 263 5868 279
rect 5802 229 5818 263
rect 5852 229 5868 263
rect 3468 171 3484 205
rect 3518 171 3534 205
rect 3468 155 3534 171
rect 5024 205 5090 221
rect 5802 213 5868 229
rect 7358 263 7424 279
rect 7358 229 7374 263
rect 7408 229 7424 263
rect 5024 171 5040 205
rect 5074 171 5090 205
rect 5024 155 5090 171
rect 6580 205 6646 221
rect 7358 213 7424 229
rect 8914 263 8980 279
rect 8914 229 8930 263
rect 8964 229 8980 263
rect 6580 171 6596 205
rect 6630 171 6646 205
rect 6580 155 6646 171
rect 8136 205 8202 221
rect 8914 213 8980 229
rect 10470 263 10536 279
rect 10470 229 10486 263
rect 10520 229 10536 263
rect 8136 171 8152 205
rect 8186 171 8202 205
rect 8136 155 8202 171
rect 9692 205 9758 221
rect 10470 213 10536 229
rect 12026 263 12092 279
rect 12026 229 12042 263
rect 12076 229 12092 263
rect 9692 171 9708 205
rect 9742 171 9758 205
rect 9692 155 9758 171
rect 11248 205 11314 221
rect 12026 213 12092 229
rect 13582 263 13648 279
rect 13582 229 13598 263
rect 13632 229 13648 263
rect 11248 171 11264 205
rect 11298 171 11314 205
rect 11248 155 11314 171
rect 12804 205 12870 221
rect 13582 213 13648 229
rect 15138 263 15204 279
rect 15138 229 15154 263
rect 15188 229 15204 263
rect 12804 171 12820 205
rect 12854 171 12870 205
rect 12804 155 12870 171
rect 14360 205 14426 221
rect 15138 213 15204 229
rect 16694 263 16760 279
rect 16694 229 16710 263
rect 16744 229 16760 263
rect 14360 171 14376 205
rect 14410 171 14426 205
rect 14360 155 14426 171
rect 15916 205 15982 221
rect 16694 213 16760 229
rect 18250 263 18316 279
rect 18250 229 18266 263
rect 18300 229 18316 263
rect 15916 171 15932 205
rect 15966 171 15982 205
rect 15916 155 15982 171
rect 17472 205 17538 221
rect 18250 213 18316 229
rect 19806 263 19872 279
rect 19806 229 19822 263
rect 19856 229 19872 263
rect 17472 171 17488 205
rect 17522 171 17538 205
rect 17472 155 17538 171
rect 19028 205 19094 221
rect 19806 213 19872 229
rect 21362 263 21428 279
rect 21362 229 21378 263
rect 21412 229 21428 263
rect 19028 171 19044 205
rect 19078 171 19094 205
rect 19028 155 19094 171
rect 20584 205 20650 221
rect 21362 213 21428 229
rect 22918 263 22984 279
rect 22918 229 22934 263
rect 22968 229 22984 263
rect 20584 171 20600 205
rect 20634 171 20650 205
rect 20584 155 20650 171
rect 22140 205 22206 221
rect 22918 213 22984 229
rect 24474 263 24540 279
rect 24474 229 24490 263
rect 24524 229 24540 263
rect 22140 171 22156 205
rect 22190 171 22206 205
rect 22140 155 22206 171
rect 23696 205 23762 221
rect 24474 213 24540 229
rect 23696 171 23712 205
rect 23746 171 23762 205
rect 23696 155 23762 171
<< viali >>
rect 1150 229 1184 263
rect 2706 229 2740 263
rect 372 171 406 205
rect 4262 229 4296 263
rect 1928 171 1962 205
rect 5818 229 5852 263
rect 3484 171 3518 205
rect 7374 229 7408 263
rect 5040 171 5074 205
rect 8930 229 8964 263
rect 6596 171 6630 205
rect 10486 229 10520 263
rect 8152 171 8186 205
rect 12042 229 12076 263
rect 9708 171 9742 205
rect 13598 229 13632 263
rect 11264 171 11298 205
rect 15154 229 15188 263
rect 12820 171 12854 205
rect 16710 229 16744 263
rect 14376 171 14410 205
rect 18266 229 18300 263
rect 15932 171 15966 205
rect 19822 229 19856 263
rect 17488 171 17522 205
rect 21378 229 21412 263
rect 19044 171 19078 205
rect 22934 229 22968 263
rect 20600 171 20634 205
rect 24490 229 24524 263
rect 22156 171 22190 205
rect 23712 171 23746 205
<< metal1 >>
rect 1138 263 1196 269
rect 1138 260 1150 263
rect 0 232 1150 260
rect 1138 229 1150 232
rect 1184 260 1196 263
rect 2694 263 2752 269
rect 2694 260 2706 263
rect 1184 232 2706 260
rect 1184 229 1196 232
rect 1138 223 1196 229
rect 2694 229 2706 232
rect 2740 260 2752 263
rect 4250 263 4308 269
rect 4250 260 4262 263
rect 2740 232 4262 260
rect 2740 229 2752 232
rect 2694 223 2752 229
rect 4250 229 4262 232
rect 4296 260 4308 263
rect 5806 263 5864 269
rect 5806 260 5818 263
rect 4296 232 5818 260
rect 4296 229 4308 232
rect 4250 223 4308 229
rect 5806 229 5818 232
rect 5852 260 5864 263
rect 7362 263 7420 269
rect 7362 260 7374 263
rect 5852 232 7374 260
rect 5852 229 5864 232
rect 5806 223 5864 229
rect 7362 229 7374 232
rect 7408 260 7420 263
rect 8918 263 8976 269
rect 8918 260 8930 263
rect 7408 232 8930 260
rect 7408 229 7420 232
rect 7362 223 7420 229
rect 8918 229 8930 232
rect 8964 260 8976 263
rect 10474 263 10532 269
rect 10474 260 10486 263
rect 8964 232 10486 260
rect 8964 229 8976 232
rect 8918 223 8976 229
rect 10474 229 10486 232
rect 10520 260 10532 263
rect 12030 263 12088 269
rect 12030 260 12042 263
rect 10520 232 12042 260
rect 10520 229 10532 232
rect 10474 223 10532 229
rect 12030 229 12042 232
rect 12076 260 12088 263
rect 13586 263 13644 269
rect 13586 260 13598 263
rect 12076 232 13598 260
rect 12076 229 12088 232
rect 12030 223 12088 229
rect 13586 229 13598 232
rect 13632 260 13644 263
rect 15142 263 15200 269
rect 15142 260 15154 263
rect 13632 232 15154 260
rect 13632 229 13644 232
rect 13586 223 13644 229
rect 15142 229 15154 232
rect 15188 260 15200 263
rect 16698 263 16756 269
rect 16698 260 16710 263
rect 15188 232 16710 260
rect 15188 229 15200 232
rect 15142 223 15200 229
rect 16698 229 16710 232
rect 16744 260 16756 263
rect 18254 263 18312 269
rect 18254 260 18266 263
rect 16744 232 18266 260
rect 16744 229 16756 232
rect 16698 223 16756 229
rect 18254 229 18266 232
rect 18300 260 18312 263
rect 19810 263 19868 269
rect 19810 260 19822 263
rect 18300 232 19822 260
rect 18300 229 18312 232
rect 18254 223 18312 229
rect 19810 229 19822 232
rect 19856 260 19868 263
rect 21366 263 21424 269
rect 21366 260 21378 263
rect 19856 232 21378 260
rect 19856 229 19868 232
rect 19810 223 19868 229
rect 21366 229 21378 232
rect 21412 260 21424 263
rect 22922 263 22980 269
rect 22922 260 22934 263
rect 21412 232 22934 260
rect 21412 229 21424 232
rect 21366 223 21424 229
rect 22922 229 22934 232
rect 22968 260 22980 263
rect 24478 263 24536 269
rect 24478 260 24490 263
rect 22968 232 24490 260
rect 22968 229 22980 232
rect 22922 223 22980 229
rect 24478 229 24490 232
rect 24524 260 24536 263
rect 24524 232 24896 260
rect 24524 229 24536 232
rect 24478 223 24536 229
rect 360 205 418 211
rect 360 202 372 205
rect 0 174 372 202
rect 360 171 372 174
rect 406 202 418 205
rect 1916 205 1974 211
rect 1916 202 1928 205
rect 406 174 1928 202
rect 406 171 418 174
rect 360 165 418 171
rect 1916 171 1928 174
rect 1962 202 1974 205
rect 3472 205 3530 211
rect 3472 202 3484 205
rect 1962 174 3484 202
rect 1962 171 1974 174
rect 1916 165 1974 171
rect 3472 171 3484 174
rect 3518 202 3530 205
rect 5028 205 5086 211
rect 5028 202 5040 205
rect 3518 174 5040 202
rect 3518 171 3530 174
rect 3472 165 3530 171
rect 5028 171 5040 174
rect 5074 202 5086 205
rect 6584 205 6642 211
rect 6584 202 6596 205
rect 5074 174 6596 202
rect 5074 171 5086 174
rect 5028 165 5086 171
rect 6584 171 6596 174
rect 6630 202 6642 205
rect 8140 205 8198 211
rect 8140 202 8152 205
rect 6630 174 8152 202
rect 6630 171 6642 174
rect 6584 165 6642 171
rect 8140 171 8152 174
rect 8186 202 8198 205
rect 9696 205 9754 211
rect 9696 202 9708 205
rect 8186 174 9708 202
rect 8186 171 8198 174
rect 8140 165 8198 171
rect 9696 171 9708 174
rect 9742 202 9754 205
rect 11252 205 11310 211
rect 11252 202 11264 205
rect 9742 174 11264 202
rect 9742 171 9754 174
rect 9696 165 9754 171
rect 11252 171 11264 174
rect 11298 202 11310 205
rect 12808 205 12866 211
rect 12808 202 12820 205
rect 11298 174 12820 202
rect 11298 171 11310 174
rect 11252 165 11310 171
rect 12808 171 12820 174
rect 12854 202 12866 205
rect 14364 205 14422 211
rect 14364 202 14376 205
rect 12854 174 14376 202
rect 12854 171 12866 174
rect 12808 165 12866 171
rect 14364 171 14376 174
rect 14410 202 14422 205
rect 15920 205 15978 211
rect 15920 202 15932 205
rect 14410 174 15932 202
rect 14410 171 14422 174
rect 14364 165 14422 171
rect 15920 171 15932 174
rect 15966 202 15978 205
rect 17476 205 17534 211
rect 17476 202 17488 205
rect 15966 174 17488 202
rect 15966 171 15978 174
rect 15920 165 15978 171
rect 17476 171 17488 174
rect 17522 202 17534 205
rect 19032 205 19090 211
rect 19032 202 19044 205
rect 17522 174 19044 202
rect 17522 171 17534 174
rect 17476 165 17534 171
rect 19032 171 19044 174
rect 19078 202 19090 205
rect 20588 205 20646 211
rect 20588 202 20600 205
rect 19078 174 20600 202
rect 19078 171 19090 174
rect 19032 165 19090 171
rect 20588 171 20600 174
rect 20634 202 20646 205
rect 22144 205 22202 211
rect 22144 202 22156 205
rect 20634 174 22156 202
rect 20634 171 20646 174
rect 20588 165 20646 171
rect 22144 171 22156 174
rect 22190 202 22202 205
rect 23700 205 23758 211
rect 23700 202 23712 205
rect 22190 174 23712 202
rect 22190 171 22202 174
rect 22144 165 22202 171
rect 23700 171 23712 174
rect 23746 202 23758 205
rect 23746 174 24896 202
rect 23746 171 23758 174
rect 23700 165 23758 171
rect 108 102 834 130
rect 1664 102 2390 130
rect 3220 102 3946 130
rect 4776 102 5502 130
rect 6332 102 7058 130
rect 7888 102 8614 130
rect 9444 102 10170 130
rect 11000 102 11726 130
rect 12556 102 13282 130
rect 14112 102 14838 130
rect 15668 102 16394 130
rect 17224 102 17950 130
rect 18780 102 19506 130
rect 20336 102 21062 130
rect 21892 102 22618 130
rect 23448 102 24174 130
rect 750 44 1476 72
rect 2306 44 3032 72
rect 3862 44 4588 72
rect 5418 44 6144 72
rect 6974 44 7700 72
rect 8530 44 9256 72
rect 10086 44 10812 72
rect 11642 44 12368 72
rect 13198 44 13924 72
rect 14754 44 15480 72
rect 16310 44 17036 72
rect 17866 44 18592 72
rect 19422 44 20148 72
rect 20978 44 21704 72
rect 22534 44 23260 72
rect 24090 44 24816 72
<< via1 >>
rect 56 90 108 142
rect 834 90 886 142
rect 1612 90 1664 142
rect 2390 90 2442 142
rect 3168 90 3220 142
rect 3946 90 3998 142
rect 4724 90 4776 142
rect 5502 90 5554 142
rect 6280 90 6332 142
rect 7058 90 7110 142
rect 7836 90 7888 142
rect 8614 90 8666 142
rect 9392 90 9444 142
rect 10170 90 10222 142
rect 10948 90 11000 142
rect 11726 90 11778 142
rect 12504 90 12556 142
rect 13282 90 13334 142
rect 14060 90 14112 142
rect 14838 90 14890 142
rect 15616 90 15668 142
rect 16394 90 16446 142
rect 17172 90 17224 142
rect 17950 90 18002 142
rect 18728 90 18780 142
rect 19506 90 19558 142
rect 20284 90 20336 142
rect 21062 90 21114 142
rect 21840 90 21892 142
rect 22618 90 22670 142
rect 23396 90 23448 142
rect 24174 90 24226 142
rect 698 32 750 84
rect 1476 32 1528 84
rect 2254 32 2306 84
rect 3032 32 3084 84
rect 3810 32 3862 84
rect 4588 32 4640 84
rect 5366 32 5418 84
rect 6144 32 6196 84
rect 6922 32 6974 84
rect 7700 32 7752 84
rect 8478 32 8530 84
rect 9256 32 9308 84
rect 10034 32 10086 84
rect 10812 32 10864 84
rect 11590 32 11642 84
rect 12368 32 12420 84
rect 13146 32 13198 84
rect 13924 32 13976 84
rect 14702 32 14754 84
rect 15480 32 15532 84
rect 16258 32 16310 84
rect 17036 32 17088 84
rect 17814 32 17866 84
rect 18592 32 18644 84
rect 19370 32 19422 84
rect 20148 32 20200 84
rect 20926 32 20978 84
rect 21704 32 21756 84
rect 22482 32 22534 84
rect 23260 32 23312 84
rect 24038 32 24090 84
rect 24816 32 24868 84
<< metal2 >>
rect 68 1742 96 1798
rect 710 1742 738 1798
rect 846 1742 874 1798
rect 1488 1742 1516 1798
rect 1624 1742 1652 1798
rect 2266 1742 2294 1798
rect 2402 1742 2430 1798
rect 3044 1742 3072 1798
rect 3180 1742 3208 1798
rect 3822 1742 3850 1798
rect 3958 1742 3986 1798
rect 4600 1742 4628 1798
rect 4736 1742 4764 1798
rect 5378 1742 5406 1798
rect 5514 1742 5542 1798
rect 6156 1742 6184 1798
rect 6292 1742 6320 1798
rect 6934 1742 6962 1798
rect 7070 1742 7098 1798
rect 7712 1742 7740 1798
rect 7848 1742 7876 1798
rect 8490 1742 8518 1798
rect 8626 1742 8654 1798
rect 9268 1742 9296 1798
rect 9404 1742 9432 1798
rect 10046 1742 10074 1798
rect 10182 1742 10210 1798
rect 10824 1742 10852 1798
rect 10960 1742 10988 1798
rect 11602 1742 11630 1798
rect 11738 1742 11766 1798
rect 12380 1742 12408 1798
rect 12516 1742 12544 1798
rect 13158 1742 13186 1798
rect 13294 1742 13322 1798
rect 13936 1742 13964 1798
rect 14072 1742 14100 1798
rect 14714 1742 14742 1798
rect 14850 1742 14878 1798
rect 15492 1742 15520 1798
rect 15628 1742 15656 1798
rect 16270 1742 16298 1798
rect 16406 1742 16434 1798
rect 17048 1742 17076 1798
rect 17184 1742 17212 1798
rect 17826 1742 17854 1798
rect 17962 1742 17990 1798
rect 18604 1742 18632 1798
rect 18740 1742 18768 1798
rect 19382 1742 19410 1798
rect 19518 1742 19546 1798
rect 20160 1742 20188 1798
rect 20296 1742 20324 1798
rect 20938 1742 20966 1798
rect 21074 1742 21102 1798
rect 21716 1742 21744 1798
rect 21852 1742 21880 1798
rect 22494 1742 22522 1798
rect 22630 1742 22658 1798
rect 23272 1742 23300 1798
rect 23408 1742 23436 1798
rect 24050 1742 24078 1798
rect 24186 1742 24214 1798
rect 24828 1742 24856 1798
rect 68 142 96 290
rect 710 84 738 290
rect 846 142 874 290
rect 1488 84 1516 290
rect 1624 142 1652 290
rect 2266 84 2294 290
rect 2402 142 2430 290
rect 3044 84 3072 290
rect 3180 142 3208 290
rect 3822 84 3850 290
rect 3958 142 3986 290
rect 4600 84 4628 290
rect 4736 142 4764 290
rect 5378 84 5406 290
rect 5514 142 5542 290
rect 6156 84 6184 290
rect 6292 142 6320 290
rect 6934 84 6962 290
rect 7070 142 7098 290
rect 7712 84 7740 290
rect 7848 142 7876 290
rect 8490 84 8518 290
rect 8626 142 8654 290
rect 9268 84 9296 290
rect 9404 142 9432 290
rect 10046 84 10074 290
rect 10182 142 10210 290
rect 10824 84 10852 290
rect 10960 142 10988 290
rect 11602 84 11630 290
rect 11738 142 11766 290
rect 12380 84 12408 290
rect 12516 142 12544 290
rect 13158 84 13186 290
rect 13294 142 13322 290
rect 13936 84 13964 290
rect 14072 142 14100 290
rect 14714 84 14742 290
rect 14850 142 14878 290
rect 15492 84 15520 290
rect 15628 142 15656 290
rect 16270 84 16298 290
rect 16406 142 16434 290
rect 17048 84 17076 290
rect 17184 142 17212 290
rect 17826 84 17854 290
rect 17962 142 17990 290
rect 18604 84 18632 290
rect 18740 142 18768 290
rect 19382 84 19410 290
rect 19518 142 19546 290
rect 20160 84 20188 290
rect 20296 142 20324 290
rect 20938 84 20966 290
rect 21074 142 21102 290
rect 21716 84 21744 290
rect 21852 142 21880 290
rect 22494 84 22522 290
rect 22630 142 22658 290
rect 23272 84 23300 290
rect 23408 142 23436 290
rect 24050 84 24078 290
rect 24186 142 24214 290
rect 24828 84 24856 290
<< metal3 >>
rect 748 1019 808 1079
rect 1526 1019 1586 1079
rect 2304 1019 2364 1079
rect 3082 1019 3142 1079
rect 3860 1019 3920 1079
rect 4638 1019 4698 1079
rect 5416 1019 5476 1079
rect 6194 1019 6254 1079
rect 6972 1019 7032 1079
rect 7750 1019 7810 1079
rect 8528 1019 8588 1079
rect 9306 1019 9366 1079
rect 10084 1019 10144 1079
rect 10862 1019 10922 1079
rect 11640 1019 11700 1079
rect 12418 1019 12478 1079
rect 13196 1019 13256 1079
rect 13974 1019 14034 1079
rect 14752 1019 14812 1079
rect 15530 1019 15590 1079
rect 16308 1019 16368 1079
rect 17086 1019 17146 1079
rect 17864 1019 17924 1079
rect 18642 1019 18702 1079
rect 19420 1019 19480 1079
rect 20198 1019 20258 1079
rect 20976 1019 21036 1079
rect 21754 1019 21814 1079
rect 22532 1019 22592 1079
rect 23310 1019 23370 1079
rect 24088 1019 24148 1079
rect 24866 1019 24926 1079
use contact_14  contact_14_0
timestamp 1643671299
transform 1 0 24827 0 1 43
box 0 0 1 1
use contact_14  contact_14_1
timestamp 1643671299
transform 1 0 24185 0 1 101
box 0 0 1 1
use contact_14  contact_14_2
timestamp 1643671299
transform 1 0 24049 0 1 43
box 0 0 1 1
use contact_14  contact_14_3
timestamp 1643671299
transform 1 0 23407 0 1 101
box 0 0 1 1
use contact_14  contact_14_4
timestamp 1643671299
transform 1 0 23271 0 1 43
box 0 0 1 1
use contact_14  contact_14_5
timestamp 1643671299
transform 1 0 22629 0 1 101
box 0 0 1 1
use contact_14  contact_14_6
timestamp 1643671299
transform 1 0 22493 0 1 43
box 0 0 1 1
use contact_14  contact_14_7
timestamp 1643671299
transform 1 0 21851 0 1 101
box 0 0 1 1
use contact_14  contact_14_8
timestamp 1643671299
transform 1 0 21715 0 1 43
box 0 0 1 1
use contact_14  contact_14_9
timestamp 1643671299
transform 1 0 21073 0 1 101
box 0 0 1 1
use contact_14  contact_14_10
timestamp 1643671299
transform 1 0 20937 0 1 43
box 0 0 1 1
use contact_14  contact_14_11
timestamp 1643671299
transform 1 0 20295 0 1 101
box 0 0 1 1
use contact_14  contact_14_12
timestamp 1643671299
transform 1 0 20159 0 1 43
box 0 0 1 1
use contact_14  contact_14_13
timestamp 1643671299
transform 1 0 19517 0 1 101
box 0 0 1 1
use contact_14  contact_14_14
timestamp 1643671299
transform 1 0 19381 0 1 43
box 0 0 1 1
use contact_14  contact_14_15
timestamp 1643671299
transform 1 0 18739 0 1 101
box 0 0 1 1
use contact_14  contact_14_16
timestamp 1643671299
transform 1 0 18603 0 1 43
box 0 0 1 1
use contact_14  contact_14_17
timestamp 1643671299
transform 1 0 17961 0 1 101
box 0 0 1 1
use contact_14  contact_14_18
timestamp 1643671299
transform 1 0 17825 0 1 43
box 0 0 1 1
use contact_14  contact_14_19
timestamp 1643671299
transform 1 0 17183 0 1 101
box 0 0 1 1
use contact_14  contact_14_20
timestamp 1643671299
transform 1 0 17047 0 1 43
box 0 0 1 1
use contact_14  contact_14_21
timestamp 1643671299
transform 1 0 16405 0 1 101
box 0 0 1 1
use contact_14  contact_14_22
timestamp 1643671299
transform 1 0 16269 0 1 43
box 0 0 1 1
use contact_14  contact_14_23
timestamp 1643671299
transform 1 0 15627 0 1 101
box 0 0 1 1
use contact_14  contact_14_24
timestamp 1643671299
transform 1 0 15491 0 1 43
box 0 0 1 1
use contact_14  contact_14_25
timestamp 1643671299
transform 1 0 14849 0 1 101
box 0 0 1 1
use contact_14  contact_14_26
timestamp 1643671299
transform 1 0 14713 0 1 43
box 0 0 1 1
use contact_14  contact_14_27
timestamp 1643671299
transform 1 0 14071 0 1 101
box 0 0 1 1
use contact_14  contact_14_28
timestamp 1643671299
transform 1 0 13935 0 1 43
box 0 0 1 1
use contact_14  contact_14_29
timestamp 1643671299
transform 1 0 13293 0 1 101
box 0 0 1 1
use contact_14  contact_14_30
timestamp 1643671299
transform 1 0 13157 0 1 43
box 0 0 1 1
use contact_14  contact_14_31
timestamp 1643671299
transform 1 0 12515 0 1 101
box 0 0 1 1
use contact_14  contact_14_32
timestamp 1643671299
transform 1 0 12379 0 1 43
box 0 0 1 1
use contact_14  contact_14_33
timestamp 1643671299
transform 1 0 11737 0 1 101
box 0 0 1 1
use contact_14  contact_14_34
timestamp 1643671299
transform 1 0 11601 0 1 43
box 0 0 1 1
use contact_14  contact_14_35
timestamp 1643671299
transform 1 0 10959 0 1 101
box 0 0 1 1
use contact_14  contact_14_36
timestamp 1643671299
transform 1 0 10823 0 1 43
box 0 0 1 1
use contact_14  contact_14_37
timestamp 1643671299
transform 1 0 10181 0 1 101
box 0 0 1 1
use contact_14  contact_14_38
timestamp 1643671299
transform 1 0 10045 0 1 43
box 0 0 1 1
use contact_14  contact_14_39
timestamp 1643671299
transform 1 0 9403 0 1 101
box 0 0 1 1
use contact_14  contact_14_40
timestamp 1643671299
transform 1 0 9267 0 1 43
box 0 0 1 1
use contact_14  contact_14_41
timestamp 1643671299
transform 1 0 8625 0 1 101
box 0 0 1 1
use contact_14  contact_14_42
timestamp 1643671299
transform 1 0 8489 0 1 43
box 0 0 1 1
use contact_14  contact_14_43
timestamp 1643671299
transform 1 0 7847 0 1 101
box 0 0 1 1
use contact_14  contact_14_44
timestamp 1643671299
transform 1 0 7711 0 1 43
box 0 0 1 1
use contact_14  contact_14_45
timestamp 1643671299
transform 1 0 7069 0 1 101
box 0 0 1 1
use contact_14  contact_14_46
timestamp 1643671299
transform 1 0 6933 0 1 43
box 0 0 1 1
use contact_14  contact_14_47
timestamp 1643671299
transform 1 0 6291 0 1 101
box 0 0 1 1
use contact_14  contact_14_48
timestamp 1643671299
transform 1 0 6155 0 1 43
box 0 0 1 1
use contact_14  contact_14_49
timestamp 1643671299
transform 1 0 5513 0 1 101
box 0 0 1 1
use contact_14  contact_14_50
timestamp 1643671299
transform 1 0 5377 0 1 43
box 0 0 1 1
use contact_14  contact_14_51
timestamp 1643671299
transform 1 0 4735 0 1 101
box 0 0 1 1
use contact_14  contact_14_52
timestamp 1643671299
transform 1 0 4599 0 1 43
box 0 0 1 1
use contact_14  contact_14_53
timestamp 1643671299
transform 1 0 3957 0 1 101
box 0 0 1 1
use contact_14  contact_14_54
timestamp 1643671299
transform 1 0 3821 0 1 43
box 0 0 1 1
use contact_14  contact_14_55
timestamp 1643671299
transform 1 0 3179 0 1 101
box 0 0 1 1
use contact_14  contact_14_56
timestamp 1643671299
transform 1 0 3043 0 1 43
box 0 0 1 1
use contact_14  contact_14_57
timestamp 1643671299
transform 1 0 2401 0 1 101
box 0 0 1 1
use contact_14  contact_14_58
timestamp 1643671299
transform 1 0 2265 0 1 43
box 0 0 1 1
use contact_14  contact_14_59
timestamp 1643671299
transform 1 0 1623 0 1 101
box 0 0 1 1
use contact_14  contact_14_60
timestamp 1643671299
transform 1 0 1487 0 1 43
box 0 0 1 1
use contact_14  contact_14_61
timestamp 1643671299
transform 1 0 845 0 1 101
box 0 0 1 1
use contact_14  contact_14_62
timestamp 1643671299
transform 1 0 709 0 1 43
box 0 0 1 1
use contact_14  contact_14_63
timestamp 1643671299
transform 1 0 67 0 1 101
box 0 0 1 1
use contact_27  contact_27_0
timestamp 1643671299
transform 1 0 24478 0 1 223
box 0 0 1 1
use contact_26  contact_26_0
timestamp 1643671299
transform 1 0 24474 0 1 213
box 0 0 1 1
use contact_27  contact_27_1
timestamp 1643671299
transform 1 0 23700 0 1 165
box 0 0 1 1
use contact_26  contact_26_1
timestamp 1643671299
transform 1 0 23696 0 1 155
box 0 0 1 1
use contact_27  contact_27_2
timestamp 1643671299
transform 1 0 22922 0 1 223
box 0 0 1 1
use contact_26  contact_26_2
timestamp 1643671299
transform 1 0 22918 0 1 213
box 0 0 1 1
use contact_27  contact_27_3
timestamp 1643671299
transform 1 0 22144 0 1 165
box 0 0 1 1
use contact_26  contact_26_3
timestamp 1643671299
transform 1 0 22140 0 1 155
box 0 0 1 1
use contact_27  contact_27_4
timestamp 1643671299
transform 1 0 21366 0 1 223
box 0 0 1 1
use contact_26  contact_26_4
timestamp 1643671299
transform 1 0 21362 0 1 213
box 0 0 1 1
use contact_27  contact_27_5
timestamp 1643671299
transform 1 0 20588 0 1 165
box 0 0 1 1
use contact_26  contact_26_5
timestamp 1643671299
transform 1 0 20584 0 1 155
box 0 0 1 1
use contact_27  contact_27_6
timestamp 1643671299
transform 1 0 19810 0 1 223
box 0 0 1 1
use contact_26  contact_26_6
timestamp 1643671299
transform 1 0 19806 0 1 213
box 0 0 1 1
use contact_27  contact_27_7
timestamp 1643671299
transform 1 0 19032 0 1 165
box 0 0 1 1
use contact_26  contact_26_7
timestamp 1643671299
transform 1 0 19028 0 1 155
box 0 0 1 1
use contact_27  contact_27_8
timestamp 1643671299
transform 1 0 18254 0 1 223
box 0 0 1 1
use contact_26  contact_26_8
timestamp 1643671299
transform 1 0 18250 0 1 213
box 0 0 1 1
use contact_27  contact_27_9
timestamp 1643671299
transform 1 0 17476 0 1 165
box 0 0 1 1
use contact_26  contact_26_9
timestamp 1643671299
transform 1 0 17472 0 1 155
box 0 0 1 1
use contact_27  contact_27_10
timestamp 1643671299
transform 1 0 16698 0 1 223
box 0 0 1 1
use contact_26  contact_26_10
timestamp 1643671299
transform 1 0 16694 0 1 213
box 0 0 1 1
use contact_27  contact_27_11
timestamp 1643671299
transform 1 0 15920 0 1 165
box 0 0 1 1
use contact_26  contact_26_11
timestamp 1643671299
transform 1 0 15916 0 1 155
box 0 0 1 1
use contact_27  contact_27_12
timestamp 1643671299
transform 1 0 15142 0 1 223
box 0 0 1 1
use contact_26  contact_26_12
timestamp 1643671299
transform 1 0 15138 0 1 213
box 0 0 1 1
use contact_27  contact_27_13
timestamp 1643671299
transform 1 0 14364 0 1 165
box 0 0 1 1
use contact_26  contact_26_13
timestamp 1643671299
transform 1 0 14360 0 1 155
box 0 0 1 1
use contact_27  contact_27_14
timestamp 1643671299
transform 1 0 13586 0 1 223
box 0 0 1 1
use contact_26  contact_26_14
timestamp 1643671299
transform 1 0 13582 0 1 213
box 0 0 1 1
use contact_27  contact_27_15
timestamp 1643671299
transform 1 0 12808 0 1 165
box 0 0 1 1
use contact_26  contact_26_15
timestamp 1643671299
transform 1 0 12804 0 1 155
box 0 0 1 1
use contact_27  contact_27_16
timestamp 1643671299
transform 1 0 12030 0 1 223
box 0 0 1 1
use contact_26  contact_26_16
timestamp 1643671299
transform 1 0 12026 0 1 213
box 0 0 1 1
use contact_27  contact_27_17
timestamp 1643671299
transform 1 0 11252 0 1 165
box 0 0 1 1
use contact_26  contact_26_17
timestamp 1643671299
transform 1 0 11248 0 1 155
box 0 0 1 1
use contact_27  contact_27_18
timestamp 1643671299
transform 1 0 10474 0 1 223
box 0 0 1 1
use contact_26  contact_26_18
timestamp 1643671299
transform 1 0 10470 0 1 213
box 0 0 1 1
use contact_27  contact_27_19
timestamp 1643671299
transform 1 0 9696 0 1 165
box 0 0 1 1
use contact_26  contact_26_19
timestamp 1643671299
transform 1 0 9692 0 1 155
box 0 0 1 1
use contact_27  contact_27_20
timestamp 1643671299
transform 1 0 8918 0 1 223
box 0 0 1 1
use contact_26  contact_26_20
timestamp 1643671299
transform 1 0 8914 0 1 213
box 0 0 1 1
use contact_27  contact_27_21
timestamp 1643671299
transform 1 0 8140 0 1 165
box 0 0 1 1
use contact_26  contact_26_21
timestamp 1643671299
transform 1 0 8136 0 1 155
box 0 0 1 1
use contact_27  contact_27_22
timestamp 1643671299
transform 1 0 7362 0 1 223
box 0 0 1 1
use contact_26  contact_26_22
timestamp 1643671299
transform 1 0 7358 0 1 213
box 0 0 1 1
use contact_27  contact_27_23
timestamp 1643671299
transform 1 0 6584 0 1 165
box 0 0 1 1
use contact_26  contact_26_23
timestamp 1643671299
transform 1 0 6580 0 1 155
box 0 0 1 1
use contact_27  contact_27_24
timestamp 1643671299
transform 1 0 5806 0 1 223
box 0 0 1 1
use contact_26  contact_26_24
timestamp 1643671299
transform 1 0 5802 0 1 213
box 0 0 1 1
use contact_27  contact_27_25
timestamp 1643671299
transform 1 0 5028 0 1 165
box 0 0 1 1
use contact_26  contact_26_25
timestamp 1643671299
transform 1 0 5024 0 1 155
box 0 0 1 1
use contact_27  contact_27_26
timestamp 1643671299
transform 1 0 4250 0 1 223
box 0 0 1 1
use contact_26  contact_26_26
timestamp 1643671299
transform 1 0 4246 0 1 213
box 0 0 1 1
use contact_27  contact_27_27
timestamp 1643671299
transform 1 0 3472 0 1 165
box 0 0 1 1
use contact_26  contact_26_27
timestamp 1643671299
transform 1 0 3468 0 1 155
box 0 0 1 1
use contact_27  contact_27_28
timestamp 1643671299
transform 1 0 2694 0 1 223
box 0 0 1 1
use contact_26  contact_26_28
timestamp 1643671299
transform 1 0 2690 0 1 213
box 0 0 1 1
use contact_27  contact_27_29
timestamp 1643671299
transform 1 0 1916 0 1 165
box 0 0 1 1
use contact_26  contact_26_29
timestamp 1643671299
transform 1 0 1912 0 1 155
box 0 0 1 1
use contact_27  contact_27_30
timestamp 1643671299
transform 1 0 1138 0 1 223
box 0 0 1 1
use contact_26  contact_26_30
timestamp 1643671299
transform 1 0 1134 0 1 213
box 0 0 1 1
use contact_27  contact_27_31
timestamp 1643671299
transform 1 0 360 0 1 165
box 0 0 1 1
use contact_26  contact_26_31
timestamp 1643671299
transform 1 0 356 0 1 155
box 0 0 1 1
use column_mux_multiport  column_mux_multiport_0
timestamp 1643671299
transform 1 0 24118 0 1 290
box 33 0 808 1508
use column_mux_multiport  column_mux_multiport_1
timestamp 1643671299
transform 1 0 23340 0 1 290
box 33 0 808 1508
use column_mux_multiport  column_mux_multiport_2
timestamp 1643671299
transform 1 0 22562 0 1 290
box 33 0 808 1508
use column_mux_multiport  column_mux_multiport_3
timestamp 1643671299
transform 1 0 21784 0 1 290
box 33 0 808 1508
use column_mux_multiport  column_mux_multiport_4
timestamp 1643671299
transform 1 0 21006 0 1 290
box 33 0 808 1508
use column_mux_multiport  column_mux_multiport_5
timestamp 1643671299
transform 1 0 20228 0 1 290
box 33 0 808 1508
use column_mux_multiport  column_mux_multiport_6
timestamp 1643671299
transform 1 0 19450 0 1 290
box 33 0 808 1508
use column_mux_multiport  column_mux_multiport_7
timestamp 1643671299
transform 1 0 18672 0 1 290
box 33 0 808 1508
use column_mux_multiport  column_mux_multiport_8
timestamp 1643671299
transform 1 0 17894 0 1 290
box 33 0 808 1508
use column_mux_multiport  column_mux_multiport_9
timestamp 1643671299
transform 1 0 17116 0 1 290
box 33 0 808 1508
use column_mux_multiport  column_mux_multiport_10
timestamp 1643671299
transform 1 0 16338 0 1 290
box 33 0 808 1508
use column_mux_multiport  column_mux_multiport_11
timestamp 1643671299
transform 1 0 15560 0 1 290
box 33 0 808 1508
use column_mux_multiport  column_mux_multiport_12
timestamp 1643671299
transform 1 0 14782 0 1 290
box 33 0 808 1508
use column_mux_multiport  column_mux_multiport_13
timestamp 1643671299
transform 1 0 14004 0 1 290
box 33 0 808 1508
use column_mux_multiport  column_mux_multiport_14
timestamp 1643671299
transform 1 0 13226 0 1 290
box 33 0 808 1508
use column_mux_multiport  column_mux_multiport_15
timestamp 1643671299
transform 1 0 12448 0 1 290
box 33 0 808 1508
use column_mux_multiport  column_mux_multiport_16
timestamp 1643671299
transform 1 0 11670 0 1 290
box 33 0 808 1508
use column_mux_multiport  column_mux_multiport_17
timestamp 1643671299
transform 1 0 10892 0 1 290
box 33 0 808 1508
use column_mux_multiport  column_mux_multiport_18
timestamp 1643671299
transform 1 0 10114 0 1 290
box 33 0 808 1508
use column_mux_multiport  column_mux_multiport_19
timestamp 1643671299
transform 1 0 9336 0 1 290
box 33 0 808 1508
use column_mux_multiport  column_mux_multiport_20
timestamp 1643671299
transform 1 0 8558 0 1 290
box 33 0 808 1508
use column_mux_multiport  column_mux_multiport_21
timestamp 1643671299
transform 1 0 7780 0 1 290
box 33 0 808 1508
use column_mux_multiport  column_mux_multiport_22
timestamp 1643671299
transform 1 0 7002 0 1 290
box 33 0 808 1508
use column_mux_multiport  column_mux_multiport_23
timestamp 1643671299
transform 1 0 6224 0 1 290
box 33 0 808 1508
use column_mux_multiport  column_mux_multiport_24
timestamp 1643671299
transform 1 0 5446 0 1 290
box 33 0 808 1508
use column_mux_multiport  column_mux_multiport_25
timestamp 1643671299
transform 1 0 4668 0 1 290
box 33 0 808 1508
use column_mux_multiport  column_mux_multiport_26
timestamp 1643671299
transform 1 0 3890 0 1 290
box 33 0 808 1508
use column_mux_multiport  column_mux_multiport_27
timestamp 1643671299
transform 1 0 3112 0 1 290
box 33 0 808 1508
use column_mux_multiport  column_mux_multiport_28
timestamp 1643671299
transform 1 0 2334 0 1 290
box 33 0 808 1508
use column_mux_multiport  column_mux_multiport_29
timestamp 1643671299
transform 1 0 1556 0 1 290
box 33 0 808 1508
use column_mux_multiport  column_mux_multiport_30
timestamp 1643671299
transform 1 0 778 0 1 290
box 33 0 808 1508
use column_mux_multiport  column_mux_multiport_31
timestamp 1643671299
transform 1 0 0 0 1 290
box 33 0 808 1508
<< labels >>
rlabel metal1 s 0 174 24896 202 4 sel_0
rlabel metal1 s 0 232 24896 260 4 sel_1
rlabel metal2 s 68 116 96 290 4 rbl0_out_0
rlabel metal2 s 710 58 738 290 4 rbl1_out_0
rlabel metal2 s 1624 116 1652 290 4 rbl0_out_1
rlabel metal2 s 2266 58 2294 290 4 rbl1_out_1
rlabel metal2 s 3180 116 3208 290 4 rbl0_out_2
rlabel metal2 s 3822 58 3850 290 4 rbl1_out_2
rlabel metal2 s 4736 116 4764 290 4 rbl0_out_3
rlabel metal2 s 5378 58 5406 290 4 rbl1_out_3
rlabel metal2 s 6292 116 6320 290 4 rbl0_out_4
rlabel metal2 s 6934 58 6962 290 4 rbl1_out_4
rlabel metal2 s 7848 116 7876 290 4 rbl0_out_5
rlabel metal2 s 8490 58 8518 290 4 rbl1_out_5
rlabel metal2 s 9404 116 9432 290 4 rbl0_out_6
rlabel metal2 s 10046 58 10074 290 4 rbl1_out_6
rlabel metal2 s 10960 116 10988 290 4 rbl0_out_7
rlabel metal2 s 11602 58 11630 290 4 rbl1_out_7
rlabel metal2 s 12516 116 12544 290 4 rbl0_out_8
rlabel metal2 s 13158 58 13186 290 4 rbl1_out_8
rlabel metal2 s 14072 116 14100 290 4 rbl0_out_9
rlabel metal2 s 14714 58 14742 290 4 rbl1_out_9
rlabel metal2 s 15628 116 15656 290 4 rbl0_out_10
rlabel metal2 s 16270 58 16298 290 4 rbl1_out_10
rlabel metal2 s 17184 116 17212 290 4 rbl0_out_11
rlabel metal2 s 17826 58 17854 290 4 rbl1_out_11
rlabel metal2 s 18740 116 18768 290 4 rbl0_out_12
rlabel metal2 s 19382 58 19410 290 4 rbl1_out_12
rlabel metal2 s 20296 116 20324 290 4 rbl0_out_13
rlabel metal2 s 20938 58 20966 290 4 rbl1_out_13
rlabel metal2 s 21852 116 21880 290 4 rbl0_out_14
rlabel metal2 s 22494 58 22522 290 4 rbl1_out_14
rlabel metal2 s 23408 116 23436 290 4 rbl0_out_15
rlabel metal2 s 24050 58 24078 290 4 rbl1_out_15
rlabel metal2 s 68 1742 96 1798 4 rbl0_0
rlabel metal2 s 710 1742 738 1798 4 rbl1_0
rlabel metal2 s 846 1742 874 1798 4 rbl0_1
rlabel metal2 s 1488 1742 1516 1798 4 rbl1_1
rlabel metal2 s 1624 1742 1652 1798 4 rbl0_2
rlabel metal2 s 2266 1742 2294 1798 4 rbl1_2
rlabel metal2 s 2402 1742 2430 1798 4 rbl0_3
rlabel metal2 s 3044 1742 3072 1798 4 rbl1_3
rlabel metal2 s 3180 1742 3208 1798 4 rbl0_4
rlabel metal2 s 3822 1742 3850 1798 4 rbl1_4
rlabel metal2 s 3958 1742 3986 1798 4 rbl0_5
rlabel metal2 s 4600 1742 4628 1798 4 rbl1_5
rlabel metal2 s 4736 1742 4764 1798 4 rbl0_6
rlabel metal2 s 5378 1742 5406 1798 4 rbl1_6
rlabel metal2 s 5514 1742 5542 1798 4 rbl0_7
rlabel metal2 s 6156 1742 6184 1798 4 rbl1_7
rlabel metal2 s 6292 1742 6320 1798 4 rbl0_8
rlabel metal2 s 6934 1742 6962 1798 4 rbl1_8
rlabel metal2 s 7070 1742 7098 1798 4 rbl0_9
rlabel metal2 s 7712 1742 7740 1798 4 rbl1_9
rlabel metal2 s 7848 1742 7876 1798 4 rbl0_10
rlabel metal2 s 8490 1742 8518 1798 4 rbl1_10
rlabel metal2 s 8626 1742 8654 1798 4 rbl0_11
rlabel metal2 s 9268 1742 9296 1798 4 rbl1_11
rlabel metal2 s 9404 1742 9432 1798 4 rbl0_12
rlabel metal2 s 10046 1742 10074 1798 4 rbl1_12
rlabel metal2 s 10182 1742 10210 1798 4 rbl0_13
rlabel metal2 s 10824 1742 10852 1798 4 rbl1_13
rlabel metal2 s 10960 1742 10988 1798 4 rbl0_14
rlabel metal2 s 11602 1742 11630 1798 4 rbl1_14
rlabel metal2 s 11738 1742 11766 1798 4 rbl0_15
rlabel metal2 s 12380 1742 12408 1798 4 rbl1_15
rlabel metal2 s 12516 1742 12544 1798 4 rbl0_16
rlabel metal2 s 13158 1742 13186 1798 4 rbl1_16
rlabel metal2 s 13294 1742 13322 1798 4 rbl0_17
rlabel metal2 s 13936 1742 13964 1798 4 rbl1_17
rlabel metal2 s 14072 1742 14100 1798 4 rbl0_18
rlabel metal2 s 14714 1742 14742 1798 4 rbl1_18
rlabel metal2 s 14850 1742 14878 1798 4 rbl0_19
rlabel metal2 s 15492 1742 15520 1798 4 rbl1_19
rlabel metal2 s 15628 1742 15656 1798 4 rbl0_20
rlabel metal2 s 16270 1742 16298 1798 4 rbl1_20
rlabel metal2 s 16406 1742 16434 1798 4 rbl0_21
rlabel metal2 s 17048 1742 17076 1798 4 rbl1_21
rlabel metal2 s 17184 1742 17212 1798 4 rbl0_22
rlabel metal2 s 17826 1742 17854 1798 4 rbl1_22
rlabel metal2 s 17962 1742 17990 1798 4 rbl0_23
rlabel metal2 s 18604 1742 18632 1798 4 rbl1_23
rlabel metal2 s 18740 1742 18768 1798 4 rbl0_24
rlabel metal2 s 19382 1742 19410 1798 4 rbl1_24
rlabel metal2 s 19518 1742 19546 1798 4 rbl0_25
rlabel metal2 s 20160 1742 20188 1798 4 rbl1_25
rlabel metal2 s 20296 1742 20324 1798 4 rbl0_26
rlabel metal2 s 20938 1742 20966 1798 4 rbl1_26
rlabel metal2 s 21074 1742 21102 1798 4 rbl0_27
rlabel metal2 s 21716 1742 21744 1798 4 rbl1_27
rlabel metal2 s 21852 1742 21880 1798 4 rbl0_28
rlabel metal2 s 22494 1742 22522 1798 4 rbl1_28
rlabel metal2 s 22630 1742 22658 1798 4 rbl0_29
rlabel metal2 s 23272 1742 23300 1798 4 rbl1_29
rlabel metal2 s 23408 1742 23436 1798 4 rbl0_30
rlabel metal2 s 24050 1742 24078 1798 4 rbl1_30
rlabel metal2 s 24186 1742 24214 1798 4 rbl0_31
rlabel metal2 s 24828 1742 24856 1798 4 rbl1_31
rlabel metal3 s 7750 1019 7810 1079 4 gnd
rlabel metal3 s 2304 1019 2364 1079 4 gnd
rlabel metal3 s 21754 1019 21814 1079 4 gnd
rlabel metal3 s 10862 1019 10922 1079 4 gnd
rlabel metal3 s 18642 1019 18702 1079 4 gnd
rlabel metal3 s 19420 1019 19480 1079 4 gnd
rlabel metal3 s 11640 1019 11700 1079 4 gnd
rlabel metal3 s 14752 1019 14812 1079 4 gnd
rlabel metal3 s 23310 1019 23370 1079 4 gnd
rlabel metal3 s 20198 1019 20258 1079 4 gnd
rlabel metal3 s 3860 1019 3920 1079 4 gnd
rlabel metal3 s 13196 1019 13256 1079 4 gnd
rlabel metal3 s 748 1019 808 1079 4 gnd
rlabel metal3 s 16308 1019 16368 1079 4 gnd
rlabel metal3 s 6194 1019 6254 1079 4 gnd
rlabel metal3 s 20976 1019 21036 1079 4 gnd
rlabel metal3 s 24088 1019 24148 1079 4 gnd
rlabel metal3 s 22532 1019 22592 1079 4 gnd
rlabel metal3 s 9306 1019 9366 1079 4 gnd
rlabel metal3 s 4638 1019 4698 1079 4 gnd
rlabel metal3 s 13974 1019 14034 1079 4 gnd
rlabel metal3 s 6972 1019 7032 1079 4 gnd
rlabel metal3 s 17864 1019 17924 1079 4 gnd
rlabel metal3 s 17086 1019 17146 1079 4 gnd
rlabel metal3 s 8528 1019 8588 1079 4 gnd
rlabel metal3 s 10084 1019 10144 1079 4 gnd
rlabel metal3 s 15530 1019 15590 1079 4 gnd
rlabel metal3 s 1526 1019 1586 1079 4 gnd
rlabel metal3 s 12418 1019 12478 1079 4 gnd
rlabel metal3 s 24866 1019 24926 1079 4 gnd
rlabel metal3 s 5416 1019 5476 1079 4 gnd
rlabel metal3 s 3082 1019 3142 1079 4 gnd
<< properties >>
string FIXED_BBOX 0 0 24896 1798
string GDS_FILE sram_0rw2r1w_16_32_sky130A.gds
string GDS_END 885624
string GDS_START 848012
<< end >>
