magic
tech sky130A
magscale 1 2
timestamp 1643671299
<< checkpaint >>
rect -1296 -1277 2835 2155
<< nwell >>
rect -36 402 1575 895
<< pwell >>
rect 1446 51 1496 133
<< psubdiff >>
rect 1446 109 1496 133
rect 1446 75 1454 109
rect 1488 75 1496 109
rect 1446 51 1496 75
<< nsubdiff >>
rect 1446 763 1496 787
rect 1446 729 1454 763
rect 1488 729 1496 763
rect 1446 705 1496 729
<< psubdiffcont >>
rect 1454 75 1488 109
<< nsubdiffcont >>
rect 1454 729 1488 763
<< poly >>
rect 114 403 144 437
rect 48 387 144 403
rect 48 353 64 387
rect 98 353 144 387
rect 48 337 144 353
rect 114 205 144 337
<< polycont >>
rect 64 353 98 387
<< locali >>
rect 0 821 1539 855
rect 62 607 96 821
rect 274 607 308 821
rect 490 607 524 821
rect 706 607 740 821
rect 922 607 956 821
rect 1138 607 1172 821
rect 1350 607 1384 821
rect 1454 763 1488 821
rect 1454 713 1488 729
rect 48 387 114 403
rect 48 353 64 387
rect 98 353 114 387
rect 48 337 114 353
rect 706 387 740 573
rect 706 353 757 387
rect 706 167 740 353
rect 1454 109 1488 125
rect 62 17 96 67
rect 274 17 308 67
rect 490 17 524 67
rect 706 17 740 67
rect 922 17 956 67
rect 1138 17 1172 67
rect 1350 17 1384 67
rect 1454 17 1488 75
rect 0 -17 1539 17
use contact_12  contact_12_0
timestamp 1643671299
transform 1 0 48 0 1 337
box 0 0 1 1
use contact_11  contact_11_0
timestamp 1643671299
transform 1 0 1446 0 1 51
box 0 0 1 1
use contact_10  contact_10_0
timestamp 1643671299
transform 1 0 1446 0 1 705
box 0 0 1 1
use nmos_m12_w0_490_sli_dli_da_p  nmos_m12_w0_490_sli_dli_da_p_0
timestamp 1643671299
transform 1 0 54 0 1 51
box 0 -26 1338 154
use pmos_m12_w1_470_sli_dli_da_p  pmos_m12_w1_470_sli_dli_da_p_0
timestamp 1643671299
transform 1 0 54 0 1 493
box -59 -56 1397 348
<< labels >>
rlabel locali s 81 370 81 370 4 A
rlabel locali s 740 370 740 370 4 Z
rlabel locali s 769 0 769 0 4 gnd
rlabel locali s 769 838 769 838 4 vdd
<< properties >>
string FIXED_BBOX 0 0 1539 662
string GDS_FILE sram_0rw2r1w_16_32_sky130A.gds
string GDS_END 1156646
string GDS_START 1154386
<< end >>
