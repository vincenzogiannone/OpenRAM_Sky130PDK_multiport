magic
tech sky130A
magscale 1 2
timestamp 1643593061
<< checkpaint >>
rect -1260 -1268 3594 2312
<< metal1 >>
rect 0 11 2334 39
<< metal2 >>
rect 70 0 98 1038
rect 532 0 560 1038
rect 848 0 876 1038
rect 1310 0 1338 1038
rect 1626 0 1654 1038
rect 2088 0 2116 1038
<< metal3 >>
rect 163 898 223 958
rect 941 898 1001 958
rect 1719 898 1779 958
use precharge_multiport_0  precharge_multiport_0_0
timestamp 1643593061
transform 1 0 1556 0 1 0
box 0 -8 778 1052
use precharge_multiport_0  precharge_multiport_0_1
timestamp 1643593061
transform 1 0 778 0 1 0
box 0 -8 778 1052
use precharge_multiport_0  precharge_multiport_0_2
timestamp 1643593061
transform 1 0 0 0 1 0
box 0 -8 778 1052
<< labels >>
rlabel metal1 s 0 10 2334 38 4 en_bar
rlabel metal3 s 1718 898 1778 958 4 vdd
rlabel metal3 s 162 898 222 958 4 vdd
rlabel metal3 s 940 898 1000 958 4 vdd
rlabel metal2 s 70 0 98 1038 4 rbl0_0
rlabel metal2 s 532 0 560 1038 4 rbl1_0
rlabel metal2 s 848 0 876 1038 4 rbl0_1
rlabel metal2 s 1310 0 1338 1038 4 rbl1_1
rlabel metal2 s 1626 0 1654 1038 4 rbl0_2
rlabel metal2 s 2088 0 2116 1038 4 rbl1_2
<< properties >>
string FIXED_BBOX 0 0 2334 1038
string GDS_FILE sram_0rw2r1w_2_16_sky130A.gds
string GDS_END 244512
string GDS_START 242158
<< end >>
