magic
tech sky130A
magscale 1 2
timestamp 1643593061
<< checkpaint >>
rect -1263 -1302 4224 2176
<< metal1 >>
rect 709 812 715 864
rect 767 812 773 864
rect 2191 812 2197 864
rect 2249 812 2255 864
rect 709 -26 715 26
rect 767 -26 773 26
rect 2191 -26 2197 26
rect 2249 -26 2255 26
<< via1 >>
rect 715 812 767 864
rect 2197 812 2249 864
rect 715 -26 767 26
rect 2197 -26 2249 26
<< metal2 >>
rect 0 328 28 838
rect 1482 328 1510 838
rect 0 0 28 272
rect 180 232 234 260
rect 1260 228 1314 256
rect 1482 0 1510 272
rect 1662 232 1716 260
rect 2742 228 2796 256
<< via2 >>
rect 713 864 769 866
rect 713 812 715 864
rect 715 812 767 864
rect 767 812 769 864
rect 2195 864 2251 866
rect 713 810 769 812
rect 2195 812 2197 864
rect 2197 812 2249 864
rect 2249 812 2251 864
rect 2195 810 2251 812
rect -1 272 55 328
rect 1481 272 1537 328
rect 713 26 769 28
rect 713 -26 715 26
rect 715 -26 767 26
rect 767 -26 769 26
rect 2195 26 2251 28
rect 713 -28 769 -26
rect 2195 -26 2197 26
rect 2197 -26 2249 26
rect 2249 -26 2251 26
rect 2195 -28 2251 -26
<< metal3 >>
rect 711 866 771 868
rect 711 810 713 866
rect 769 810 771 866
rect 711 808 771 810
rect 2193 866 2253 868
rect 2193 810 2195 866
rect 2251 810 2253 866
rect 2193 808 2253 810
rect -3 328 2964 330
rect -3 272 -1 328
rect 55 272 1481 328
rect 1537 272 2964 328
rect -3 270 2964 272
rect 711 28 771 30
rect 711 -28 713 28
rect 769 -28 771 28
rect 711 -30 771 -28
rect 2193 28 2253 30
rect 2193 -28 2195 28
rect 2251 -28 2253 28
rect 2193 -30 2253 -28
use contact_18  contact_18_0
timestamp 1643593061
transform 1 0 1479 0 1 270
box 0 0 1 1
use contact_18  contact_18_1
timestamp 1643593061
transform 1 0 -3 0 1 270
box 0 0 1 1
use contact_18  contact_18_2
timestamp 1643593061
transform 1 0 2193 0 1 -30
box 0 0 1 1
use contact_17  contact_17_0
timestamp 1643593061
transform 1 0 2191 0 1 -26
box 0 0 1 1
use contact_18  contact_18_3
timestamp 1643593061
transform 1 0 2193 0 1 808
box 0 0 1 1
use contact_17  contact_17_1
timestamp 1643593061
transform 1 0 2191 0 1 812
box 0 0 1 1
use contact_18  contact_18_4
timestamp 1643593061
transform 1 0 711 0 1 -30
box 0 0 1 1
use contact_17  contact_17_2
timestamp 1643593061
transform 1 0 709 0 1 -26
box 0 0 1 1
use contact_18  contact_18_5
timestamp 1643593061
transform 1 0 711 0 1 808
box 0 0 1 1
use contact_17  contact_17_3
timestamp 1643593061
transform 1 0 709 0 1 812
box 0 0 1 1
use dff  dff_0
timestamp 1643593061
transform 1 0 1482 0 1 0
box 0 -42 1482 916
use dff  dff_1
timestamp 1643593061
transform 1 0 0 0 1 0
box 0 -42 1482 916
<< labels >>
rlabel metal3 s 711 808 771 868 4 vdd
rlabel metal3 s 2193 808 2253 868 4 vdd
rlabel metal3 s 711 -30 771 30 4 gnd
rlabel metal3 s 2193 -30 2253 30 4 gnd
rlabel metal2 s 180 232 234 260 4 din_0
rlabel metal2 s 1260 228 1314 256 4 dout_0
rlabel metal2 s 1662 232 1716 260 4 din_1
rlabel metal2 s 2742 228 2796 256 4 dout_1
rlabel metal3 s 0 270 2964 330 4 clk
<< properties >>
string FIXED_BBOX 2193 -30 2253 -26
string GDS_FILE sram_0rw2r1w_2_16_sky130A.gds
string GDS_END 581874
string GDS_START 579208
<< end >>
