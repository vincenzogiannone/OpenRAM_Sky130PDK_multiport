magic
tech sky130A
magscale 1 2
timestamp 1643671299
<< checkpaint >>
rect -1271 -1260 60472 31678
<< locali >>
rect 3071 3327 3105 3361
<< viali >>
rect 3786 4626 3820 4660
rect 4091 4249 4125 4283
rect 3786 3788 3820 3822
rect 4091 3327 4125 3361
rect 3786 2950 3820 2984
<< metal1 >>
rect 6015 29642 6156 29670
rect 6015 29630 6043 29642
rect 5866 29602 6043 29630
rect 6015 29516 6156 29544
rect 6015 29504 6043 29516
rect 5866 29476 6043 29504
rect 6015 29290 6156 29318
rect 6015 29278 6043 29290
rect 5866 29250 6043 29278
rect 6015 28238 6156 28258
rect 5866 28230 6156 28238
rect 5866 28210 6043 28230
rect 6015 28012 6156 28032
rect 5866 28004 6156 28012
rect 5866 27984 6043 28004
rect 6015 27886 6156 27906
rect 5866 27878 6156 27886
rect 5866 27858 6043 27878
rect 6015 26562 6156 26590
rect 6015 26554 6043 26562
rect 5866 26526 6043 26554
rect 6015 26436 6156 26464
rect 6015 26428 6043 26436
rect 5866 26400 6043 26428
rect 6015 26210 6156 26238
rect 6015 26202 6043 26210
rect 5866 26174 6043 26202
rect 6015 25162 6156 25178
rect 5866 25150 6156 25162
rect 5866 25134 6043 25150
rect 6015 24936 6156 24952
rect 5866 24924 6156 24936
rect 5866 24908 6043 24924
rect 6015 24810 6156 24826
rect 5866 24798 6156 24810
rect 5866 24782 6043 24798
rect 6015 23482 6156 23510
rect 6015 23478 6043 23482
rect 5866 23450 6043 23478
rect 6015 23356 6156 23384
rect 6015 23352 6043 23356
rect 5866 23324 6043 23352
rect 6015 23130 6156 23158
rect 6015 23126 6043 23130
rect 5866 23098 6043 23126
rect 6015 22086 6156 22098
rect 5866 22070 6156 22086
rect 5866 22058 6043 22070
rect 6015 21860 6156 21872
rect 5866 21844 6156 21860
rect 5866 21832 6043 21844
rect 6015 21734 6156 21746
rect 5866 21718 6156 21734
rect 5866 21706 6043 21718
rect 6015 20402 6156 20430
rect 5866 20374 6043 20402
rect 6015 20276 6156 20304
rect 5866 20248 6043 20276
rect 6015 20050 6156 20078
rect 5866 20022 6043 20050
rect 6015 19010 6156 19018
rect 5866 18990 6156 19010
rect 5866 18982 6043 18990
rect 6015 18784 6156 18792
rect 5866 18764 6156 18784
rect 5866 18756 6043 18764
rect 6015 18658 6156 18666
rect 5866 18638 6156 18658
rect 5866 18630 6043 18638
rect 6015 17326 6156 17350
rect 5866 17322 6156 17326
rect 5866 17298 6043 17322
rect 6015 17200 6156 17224
rect 5866 17196 6156 17200
rect 5866 17172 6043 17196
rect 6015 16974 6156 16998
rect 5866 16970 6156 16974
rect 5866 16946 6043 16970
rect 6015 15934 6156 15938
rect 5866 15910 6156 15934
rect 5866 15906 6043 15910
rect 6015 15708 6156 15712
rect 5866 15684 6156 15708
rect 5866 15680 6043 15684
rect 6015 15582 6156 15586
rect 5866 15558 6156 15582
rect 5866 15554 6043 15558
rect 6015 14250 6156 14270
rect 5866 14242 6156 14250
rect 5866 14222 6043 14242
rect 6015 14124 6156 14144
rect 5866 14116 6156 14124
rect 5866 14096 6043 14116
rect 6015 13898 6156 13918
rect 5866 13890 6156 13898
rect 5866 13870 6043 13890
rect 5866 12830 6156 12858
rect 5866 12604 6156 12632
rect 5866 12478 6156 12506
rect 6015 11174 6156 11190
rect 5866 11162 6156 11174
rect 5866 11146 6043 11162
rect 6015 11048 6156 11064
rect 5866 11036 6156 11048
rect 5866 11020 6043 11036
rect 6015 10822 6156 10838
rect 5866 10810 6156 10822
rect 5866 10794 6043 10810
rect 5866 9778 6043 9782
rect 5866 9754 6156 9778
rect 6015 9750 6156 9754
rect 5866 9552 6043 9556
rect 5866 9528 6156 9552
rect 6015 9524 6156 9528
rect 5866 9426 6043 9430
rect 5866 9402 6156 9426
rect 6015 9398 6156 9402
rect 6015 8098 6156 8110
rect 5866 8082 6156 8098
rect 5866 8070 6043 8082
rect 6015 7972 6156 7984
rect 5866 7956 6156 7972
rect 5866 7944 6043 7956
rect 6015 7746 6156 7758
rect 5866 7730 6156 7746
rect 5866 7718 6043 7730
rect 5866 6698 6043 6706
rect 5866 6678 6156 6698
rect 6015 6670 6156 6678
rect 5866 6472 6043 6480
rect 5866 6452 6156 6472
rect 6015 6444 6156 6452
rect 5866 6346 6043 6354
rect 5866 6326 6156 6346
rect 6015 6318 6156 6326
rect 5836 5222 18175 5250
rect 3774 4658 3777 4666
rect 3748 4628 3777 4658
rect 3774 4620 3777 4628
rect 3829 4658 3832 4666
rect 3829 4628 3859 4658
rect 3829 4620 3832 4628
rect 4079 4283 4137 4289
rect 4079 4280 4091 4283
rect 2829 4252 4091 4280
rect 4079 4249 4091 4252
rect 4125 4249 4137 4283
rect 4079 4243 4137 4249
rect 3774 3820 3777 3828
rect 3748 3790 3777 3820
rect 3774 3782 3777 3790
rect 3829 3820 3832 3828
rect 3829 3790 3859 3820
rect 3829 3782 3832 3790
rect 4079 3361 4137 3367
rect 4079 3358 4091 3361
rect 2887 3330 4091 3358
rect 4079 3327 4091 3330
rect 4125 3327 4137 3361
rect 4079 3321 4137 3327
rect 2887 2994 6170 3022
rect 3774 2982 3777 2990
rect 3748 2964 3777 2982
rect 2829 2941 3777 2964
rect 3829 2982 3832 2990
rect 3829 2964 3859 2982
rect 3829 2941 6170 2964
rect 2829 2936 6170 2941
rect 18993 1171 31340 1199
<< via1 >>
rect 5784 5210 5836 5262
rect 3777 4660 3829 4669
rect 3777 4626 3786 4660
rect 3786 4626 3820 4660
rect 3820 4626 3829 4660
rect 3777 4617 3829 4626
rect 2777 4240 2829 4292
rect 3777 3822 3829 3831
rect 3777 3788 3786 3822
rect 3786 3788 3820 3822
rect 3820 3788 3829 3822
rect 3777 3779 3829 3788
rect 2835 3318 2887 3370
rect 2835 2982 2887 3034
rect 3777 2984 3829 2993
rect 2777 2924 2829 2976
rect 3777 2950 3786 2984
rect 3786 2950 3820 2984
rect 3820 2950 3829 2984
rect 3777 2941 3829 2950
rect 31340 1159 31392 1211
<< metal2 >>
rect 1 5674 29 30306
rect 69 5674 97 30306
rect 137 5674 165 30306
rect 205 5674 233 30306
rect 273 5674 301 30306
rect 341 5674 369 30306
rect 4662 30268 4690 30296
rect 5796 5262 5824 5606
rect 6352 5306 6406 5334
rect 7908 5306 7962 5334
rect 9464 5306 9518 5334
rect 11020 5306 11074 5334
rect 12576 5306 12630 5334
rect 14132 5306 14186 5334
rect 15688 5306 15742 5334
rect 17244 5306 17298 5334
rect 18800 5306 18854 5334
rect 20356 5306 20410 5334
rect 21912 5306 21966 5334
rect 23468 5306 23522 5334
rect 25024 5306 25078 5334
rect 26580 5306 26634 5334
rect 28136 5306 28190 5334
rect 29692 5306 29746 5334
rect 3784 4671 3824 4677
rect 3784 4609 3824 4615
rect 2789 2976 2817 4240
rect 3784 3833 3824 3839
rect 3784 3771 3824 3777
rect 2847 3034 2875 3318
rect 3784 2995 3824 3001
rect 3784 2933 3824 2939
rect 5796 0 5824 5210
rect 10906 4210 10934 4450
rect 12462 4210 12490 4450
rect 14018 4210 14046 4450
rect 15574 4210 15602 4450
rect 17130 4210 17158 4450
rect 18686 4210 18714 4450
rect 20242 4210 20270 4450
rect 21798 4210 21826 4450
rect 23354 4210 23382 4450
rect 24910 4210 24938 4450
rect 26466 4210 26494 4450
rect 28022 4210 28050 4450
rect 29578 4210 29606 4450
rect 31134 4210 31162 4450
rect 31352 1211 31380 30418
rect 32690 4210 32718 4450
rect 34246 4210 34274 4450
rect 31352 0 31380 1159
<< via2 >>
rect 3776 4669 3832 4671
rect 3776 4617 3777 4669
rect 3777 4617 3829 4669
rect 3829 4617 3832 4669
rect 3776 4615 3832 4617
rect 3776 3831 3832 3833
rect 3776 3779 3777 3831
rect 3777 3779 3829 3831
rect 3829 3779 3832 3831
rect 3776 3777 3832 3779
rect 3776 2993 3832 2995
rect 3776 2941 3777 2993
rect 3777 2941 3829 2993
rect 3829 2941 3832 2993
rect 3776 2939 3832 2941
<< metal3 >>
rect 651 30276 711 30336
rect 1410 30276 1470 30336
rect 5836 30252 5896 30312
rect 4632 29868 4692 29928
rect 651 28736 711 28796
rect 1410 28736 1470 28796
rect 5836 28714 5896 28774
rect 4632 28354 4692 28414
rect 651 27196 711 27256
rect 1410 27196 1470 27256
rect 5836 27176 5896 27236
rect 4632 26840 4692 26900
rect 651 25656 711 25716
rect 1410 25656 1470 25716
rect 5836 25638 5896 25698
rect 4632 25326 4692 25386
rect 651 24116 711 24176
rect 1410 24116 1470 24176
rect 5836 24100 5896 24160
rect 4632 23812 4692 23872
rect 5836 22562 5896 22622
rect 4632 22298 4692 22358
rect 651 21040 711 21100
rect 1410 21040 1470 21100
rect 5836 21024 5896 21084
rect 4632 20784 4692 20844
rect 651 19500 711 19560
rect 1410 19500 1470 19560
rect 5836 19486 5896 19546
rect 4632 19270 4692 19330
rect 651 17960 711 18020
rect 1410 17960 1470 18020
rect 5836 17948 5896 18008
rect 4632 17756 4692 17816
rect 651 16420 711 16480
rect 1410 16420 1470 16480
rect 5836 16410 5896 16470
rect 4632 16242 4692 16302
rect 651 14880 711 14940
rect 1410 14880 1470 14940
rect 5836 14872 5896 14932
rect 4632 14728 4692 14788
rect 5836 13334 5896 13394
rect 4632 13214 4692 13274
rect 651 11804 711 11864
rect 1410 11804 1470 11864
rect 5836 11796 5896 11856
rect 4632 11700 4692 11760
rect 651 10264 711 10324
rect 1410 10264 1470 10324
rect 5836 10258 5896 10318
rect 4632 10186 4692 10246
rect 651 8724 711 8784
rect 1410 8724 1470 8784
rect 4632 8672 4692 8732
rect 5836 8720 5896 8780
rect 651 7184 711 7244
rect 1410 7184 1470 7244
rect 4632 7158 4692 7218
rect 5836 7182 5896 7242
rect 651 5644 711 5704
rect 1410 5644 1470 5704
rect 4632 5644 4692 5704
rect 5836 5644 5896 5704
rect 6475 5534 6535 5594
rect 8031 5534 8091 5594
rect 9587 5534 9647 5594
rect 11143 5534 11203 5594
rect 12699 5534 12759 5594
rect 14255 5534 14315 5594
rect 15811 5534 15871 5594
rect 17367 5534 17427 5594
rect 18923 5534 18983 5594
rect 20479 5534 20539 5594
rect 22035 5534 22095 5594
rect 23591 5534 23651 5594
rect 25147 5534 25207 5594
rect 26703 5534 26763 5594
rect 28259 5534 28319 5594
rect 29815 5534 29875 5594
rect 6475 4702 6535 4762
rect 8031 4702 8091 4762
rect 9587 4702 9647 4762
rect 11143 4702 11203 4762
rect 12699 4702 12759 4762
rect 14255 4702 14315 4762
rect 15811 4702 15871 4762
rect 17367 4702 17427 4762
rect 18923 4702 18983 4762
rect 20479 4702 20539 4762
rect 22035 4702 22095 4762
rect 23591 4702 23651 4762
rect 25147 4702 25207 4762
rect 26703 4702 26763 4762
rect 28259 4702 28319 4762
rect 29815 4702 29875 4762
rect 3774 4671 3834 4673
rect 3774 4615 3776 4671
rect 3832 4615 3834 4671
rect 3774 4613 3834 4615
rect 10810 4386 10870 4446
rect 12366 4386 12426 4446
rect 13922 4386 13982 4446
rect 15478 4386 15538 4446
rect 17034 4386 17094 4446
rect 18590 4386 18650 4446
rect 20146 4386 20206 4446
rect 21702 4386 21762 4446
rect 23258 4386 23318 4446
rect 24814 4386 24874 4446
rect 26370 4386 26430 4446
rect 27926 4386 27986 4446
rect 29482 4386 29542 4446
rect 31038 4386 31098 4446
rect 32594 4386 32654 4446
rect 34150 4386 34210 4446
rect 35706 4386 35766 4446
rect 37262 4386 37322 4446
rect 38818 4386 38878 4446
rect 40374 4386 40434 4446
rect 41930 4386 41990 4446
rect 43486 4386 43546 4446
rect 45042 4386 45102 4446
rect 46598 4386 46658 4446
rect 48154 4386 48214 4446
rect 49710 4386 49770 4446
rect 51266 4386 51326 4446
rect 52822 4386 52882 4446
rect 54378 4386 54438 4446
rect 55934 4386 55994 4446
rect 57490 4386 57550 4446
rect 59046 4386 59106 4446
rect 3774 3833 3834 3835
rect 3774 3777 3776 3833
rect 3832 3777 3834 3833
rect 3774 3775 3834 3777
rect 10810 3440 10870 3500
rect 12366 3440 12426 3500
rect 13922 3440 13982 3500
rect 15478 3440 15538 3500
rect 17034 3440 17094 3500
rect 18590 3440 18650 3500
rect 20146 3440 20206 3500
rect 21702 3440 21762 3500
rect 23258 3440 23318 3500
rect 24814 3440 24874 3500
rect 26370 3440 26430 3500
rect 27926 3440 27986 3500
rect 29482 3440 29542 3500
rect 31038 3440 31098 3500
rect 32594 3440 32654 3500
rect 34150 3440 34210 3500
rect 35706 3440 35766 3500
rect 37262 3440 37322 3500
rect 38818 3440 38878 3500
rect 40374 3440 40434 3500
rect 41930 3440 41990 3500
rect 43486 3440 43546 3500
rect 45042 3440 45102 3500
rect 46598 3440 46658 3500
rect 48154 3440 48214 3500
rect 49710 3440 49770 3500
rect 51266 3440 51326 3500
rect 52822 3440 52882 3500
rect 54378 3440 54438 3500
rect 55934 3440 55994 3500
rect 57490 3440 57550 3500
rect 59046 3440 59106 3500
rect 3774 2995 3834 2997
rect 3774 2939 3776 2995
rect 3832 2939 3834 2995
rect 3774 2937 3834 2939
rect 6904 2117 6964 2177
rect 7682 2117 7742 2177
rect 8460 2117 8520 2177
rect 9238 2117 9298 2177
rect 10016 2117 10076 2177
rect 10794 2117 10854 2177
rect 11572 2117 11632 2177
rect 12350 2117 12410 2177
rect 13128 2117 13188 2177
rect 13906 2117 13966 2177
rect 14684 2117 14744 2177
rect 15462 2117 15522 2177
rect 16240 2117 16300 2177
rect 17018 2117 17078 2177
rect 17796 2117 17856 2177
rect 18574 2117 18634 2177
rect 19352 2117 19412 2177
rect 20130 2117 20190 2177
rect 20908 2117 20968 2177
rect 21686 2117 21746 2177
rect 22464 2117 22524 2177
rect 23242 2117 23302 2177
rect 24020 2117 24080 2177
rect 24798 2117 24858 2177
rect 25576 2117 25636 2177
rect 26354 2117 26414 2177
rect 27132 2117 27192 2177
rect 27910 2117 27970 2177
rect 28688 2117 28748 2177
rect 29466 2117 29526 2177
rect 30244 2117 30304 2177
rect 31022 2117 31082 2177
rect 6319 284 6379 344
rect 7097 284 7157 344
rect 7875 284 7935 344
rect 8653 284 8713 344
rect 9431 284 9491 344
rect 10209 284 10269 344
rect 10987 284 11047 344
rect 11765 284 11825 344
rect 12543 284 12603 344
rect 13321 284 13381 344
rect 14099 284 14159 344
rect 14877 284 14937 344
rect 15655 284 15715 344
rect 16433 284 16493 344
rect 17211 284 17271 344
rect 17989 284 18049 344
rect 18767 284 18827 344
rect 19545 284 19605 344
rect 20323 284 20383 344
rect 21101 284 21161 344
rect 21879 284 21939 344
rect 22657 284 22717 344
rect 23435 284 23495 344
rect 24213 284 24273 344
rect 24991 284 25051 344
rect 25769 284 25829 344
rect 26547 284 26607 344
rect 27325 284 27385 344
rect 28103 284 28163 344
rect 28881 284 28941 344
rect 29659 284 29719 344
rect 30437 284 30497 344
rect 31215 284 31275 344
use contact_18  contact_18_0
timestamp 1643671299
transform 1 0 3774 0 1 4613
box 0 0 1 1
use contact_17  contact_17_0
timestamp 1643671299
transform 1 0 3788 0 1 4628
box 0 0 1 1
use contact_13  contact_13_0
timestamp 1643671299
transform 1 0 3774 0 1 4620
box 0 0 1 1
use contact_18  contact_18_1
timestamp 1643671299
transform 1 0 3774 0 1 2937
box 0 0 1 1
use contact_17  contact_17_1
timestamp 1643671299
transform 1 0 3788 0 1 2952
box 0 0 1 1
use contact_13  contact_13_1
timestamp 1643671299
transform 1 0 3774 0 1 2944
box 0 0 1 1
use contact_18  contact_18_2
timestamp 1643671299
transform 1 0 3774 0 1 3775
box 0 0 1 1
use contact_17  contact_17_2
timestamp 1643671299
transform 1 0 3788 0 1 3790
box 0 0 1 1
use contact_13  contact_13_2
timestamp 1643671299
transform 1 0 3774 0 1 3782
box 0 0 1 1
use contact_17  contact_17_3
timestamp 1643671299
transform 1 0 31351 0 1 1170
box 0 0 1 1
use contact_17  contact_17_4
timestamp 1643671299
transform 1 0 5795 0 1 5221
box 0 0 1 1
use contact_17  contact_17_5
timestamp 1643671299
transform 1 0 2846 0 1 2993
box 0 0 1 1
use contact_13  contact_13_3
timestamp 1643671299
transform 1 0 4079 0 1 3321
box 0 0 1 1
use contact_17  contact_17_6
timestamp 1643671299
transform 1 0 2846 0 1 3329
box 0 0 1 1
use contact_17  contact_17_7
timestamp 1643671299
transform 1 0 2788 0 1 2935
box 0 0 1 1
use contact_13  contact_13_4
timestamp 1643671299
transform 1 0 4079 0 1 4243
box 0 0 1 1
use contact_17  contact_17_8
timestamp 1643671299
transform 1 0 2788 0 1 4251
box 0 0 1 1
use pinvbuf  pinvbuf_0
timestamp 1643671299
transform 1 0 3007 0 1 2950
box -36 0 1593 1710
use port_address  port_address_0
timestamp 1643671299
transform 1 0 0 0 1 5674
box -11 -42 5896 24666
use port_data  port_data_0
timestamp 1643671299
transform 1 0 6156 0 1 0
box 0 190 53056 5606
use replica_bitcell_array  replica_bitcell_array_0
timestamp 1643671299
transform 1 0 6156 0 1 5674
box 0 -42 24896 24682
<< labels >>
rlabel metal2 s 5796 0 5824 5606 4 w_en
rlabel metal2 s 4662 30268 4690 30296 4 wl_en
rlabel metal2 s 31352 0 31380 30418 4 p_en_bar
rlabel metal2 s 6352 5306 6406 5334 4 din0_0
rlabel metal2 s 7908 5306 7962 5334 4 din0_1
rlabel metal2 s 9464 5306 9518 5334 4 din0_2
rlabel metal2 s 11020 5306 11074 5334 4 din0_3
rlabel metal2 s 12576 5306 12630 5334 4 din0_4
rlabel metal2 s 14132 5306 14186 5334 4 din0_5
rlabel metal2 s 15688 5306 15742 5334 4 din0_6
rlabel metal2 s 17244 5306 17298 5334 4 din0_7
rlabel metal2 s 18800 5306 18854 5334 4 din0_8
rlabel metal2 s 20356 5306 20410 5334 4 din0_9
rlabel metal2 s 21912 5306 21966 5334 4 din0_10
rlabel metal2 s 23468 5306 23522 5334 4 din0_11
rlabel metal2 s 25024 5306 25078 5334 4 din0_12
rlabel metal2 s 26580 5306 26634 5334 4 din0_13
rlabel metal2 s 28136 5306 28190 5334 4 din0_14
rlabel metal2 s 29692 5306 29746 5334 4 din0_15
rlabel metal2 s 10906 4210 10934 4450 4 dout0_0
rlabel metal2 s 10920 4330 10920 4330 4 dout1_0
rlabel metal2 s 12462 4210 12490 4450 4 dout0_1
rlabel metal2 s 12476 4330 12476 4330 4 dout1_1
rlabel metal2 s 14018 4210 14046 4450 4 dout0_2
rlabel metal2 s 14032 4330 14032 4330 4 dout1_2
rlabel metal2 s 15574 4210 15602 4450 4 dout0_3
rlabel metal2 s 15588 4330 15588 4330 4 dout1_3
rlabel metal2 s 17130 4210 17158 4450 4 dout0_4
rlabel metal2 s 17144 4330 17144 4330 4 dout1_4
rlabel metal2 s 18686 4210 18714 4450 4 dout0_5
rlabel metal2 s 18700 4330 18700 4330 4 dout1_5
rlabel metal2 s 20242 4210 20270 4450 4 dout0_6
rlabel metal2 s 20256 4330 20256 4330 4 dout1_6
rlabel metal2 s 21798 4210 21826 4450 4 dout0_7
rlabel metal2 s 21812 4330 21812 4330 4 dout1_7
rlabel metal2 s 23354 4210 23382 4450 4 dout0_8
rlabel metal2 s 23368 4330 23368 4330 4 dout1_8
rlabel metal2 s 24910 4210 24938 4450 4 dout0_9
rlabel metal2 s 24924 4330 24924 4330 4 dout1_9
rlabel metal2 s 26466 4210 26494 4450 4 dout0_10
rlabel metal2 s 26480 4330 26480 4330 4 dout1_10
rlabel metal2 s 28022 4210 28050 4450 4 dout0_11
rlabel metal2 s 28036 4330 28036 4330 4 dout1_11
rlabel metal2 s 29578 4210 29606 4450 4 dout0_12
rlabel metal2 s 29592 4330 29592 4330 4 dout1_12
rlabel metal2 s 31134 4210 31162 4450 4 dout0_13
rlabel metal2 s 31148 4330 31148 4330 4 dout1_13
rlabel metal2 s 32690 4210 32718 4450 4 dout0_14
rlabel metal2 s 32704 4330 32704 4330 4 dout1_14
rlabel metal2 s 34246 4210 34274 4450 4 dout0_15
rlabel metal2 s 34260 4330 34260 4330 4 dout1_15
rlabel metal2 s 0 5674 28 30306 4 addr1
rlabel metal2 s 68 5674 96 30306 4 addr2
rlabel metal2 s 136 5674 164 30306 4 addr3
rlabel metal2 s 204 5674 232 30306 4 addr4
rlabel metal2 s 272 5674 300 30306 4 addr5
rlabel metal2 s 340 5674 368 30306 4 addr6
rlabel locali s 3088 3344 3088 3344 4 addr0
rlabel metal3 s 11764 284 11824 344 4 vdd
rlabel metal3 s 30436 284 30496 344 4 vdd
rlabel metal3 s 21878 284 21938 344 4 vdd
rlabel metal3 s 5836 16410 5896 16470 4 vdd
rlabel metal3 s 4632 7158 4692 7218 4 vdd
rlabel metal3 s 650 10264 710 10324 4 vdd
rlabel metal3 s 4632 13214 4692 13274 4 vdd
rlabel metal3 s 41930 3440 41990 3500 4 vdd
rlabel metal3 s 12366 3440 12426 3500 4 vdd
rlabel metal3 s 29658 284 29718 344 4 vdd
rlabel metal3 s 4632 28354 4692 28414 4 vdd
rlabel metal3 s 1410 28736 1470 28796 4 vdd
rlabel metal3 s 650 7184 710 7244 4 vdd
rlabel metal3 s 51266 3440 51326 3500 4 vdd
rlabel metal3 s 23258 3440 23318 3500 4 vdd
rlabel metal3 s 17988 284 18048 344 4 vdd
rlabel metal3 s 15654 284 15714 344 4 vdd
rlabel metal3 s 26546 284 26606 344 4 vdd
rlabel metal3 s 17366 4702 17426 4762 4 vdd
rlabel metal3 s 650 19500 710 19560 4 vdd
rlabel metal3 s 3774 3774 3834 3834 4 vdd
rlabel metal3 s 6318 284 6378 344 4 vdd
rlabel metal3 s 29814 4702 29874 4762 4 vdd
rlabel metal3 s 7874 284 7934 344 4 vdd
rlabel metal3 s 24212 284 24272 344 4 vdd
rlabel metal3 s 14098 284 14158 344 4 vdd
rlabel metal3 s 4632 16242 4692 16302 4 vdd
rlabel metal3 s 7096 284 7156 344 4 vdd
rlabel metal3 s 5836 7182 5896 7242 4 vdd
rlabel metal3 s 31214 284 31274 344 4 vdd
rlabel metal3 s 18922 4702 18982 4762 4 vdd
rlabel metal3 s 5836 25638 5896 25698 4 vdd
rlabel metal3 s 13320 284 13380 344 4 vdd
rlabel metal3 s 25768 284 25828 344 4 vdd
rlabel metal3 s 48154 3440 48214 3500 4 vdd
rlabel metal3 s 16432 284 16492 344 4 vdd
rlabel metal3 s 11142 4702 11202 4762 4 vdd
rlabel metal3 s 4632 19270 4692 19330 4 vdd
rlabel metal3 s 5836 10258 5896 10318 4 vdd
rlabel metal3 s 26702 4702 26762 4762 4 vdd
rlabel metal3 s 1410 7184 1470 7244 4 vdd
rlabel metal3 s 15810 4702 15870 4762 4 vdd
rlabel metal3 s 24814 3440 24874 3500 4 vdd
rlabel metal3 s 43486 3440 43546 3500 4 vdd
rlabel metal3 s 14876 284 14936 344 4 vdd
rlabel metal3 s 20322 284 20382 344 4 vdd
rlabel metal3 s 20478 4702 20538 4762 4 vdd
rlabel metal3 s 650 16420 710 16480 4 vdd
rlabel metal3 s 22034 4702 22094 4762 4 vdd
rlabel metal3 s 45042 3440 45102 3500 4 vdd
rlabel metal3 s 18766 284 18826 344 4 vdd
rlabel metal3 s 28102 284 28162 344 4 vdd
rlabel metal3 s 5836 28714 5896 28774 4 vdd
rlabel metal3 s 55934 3440 55994 3500 4 vdd
rlabel metal3 s 1410 25656 1470 25716 4 vdd
rlabel metal3 s 17210 284 17270 344 4 vdd
rlabel metal3 s 23434 284 23494 344 4 vdd
rlabel metal3 s 14254 4702 14314 4762 4 vdd
rlabel metal3 s 18590 3440 18650 3500 4 vdd
rlabel metal3 s 13922 3440 13982 3500 4 vdd
rlabel metal3 s 20146 3440 20206 3500 4 vdd
rlabel metal3 s 52822 3440 52882 3500 4 vdd
rlabel metal3 s 4632 22298 4692 22358 4 vdd
rlabel metal3 s 12698 4702 12758 4762 4 vdd
rlabel metal3 s 10810 3440 10870 3500 4 vdd
rlabel metal3 s 26370 3440 26430 3500 4 vdd
rlabel metal3 s 35706 3440 35766 3500 4 vdd
rlabel metal3 s 22656 284 22716 344 4 vdd
rlabel metal3 s 10986 284 11046 344 4 vdd
rlabel metal3 s 29482 3440 29542 3500 4 vdd
rlabel metal3 s 650 25656 710 25716 4 vdd
rlabel metal3 s 27926 3440 27986 3500 4 vdd
rlabel metal3 s 34150 3440 34210 3500 4 vdd
rlabel metal3 s 38818 3440 38878 3500 4 vdd
rlabel metal3 s 21100 284 21160 344 4 vdd
rlabel metal3 s 31038 3440 31098 3500 4 vdd
rlabel metal3 s 37262 3440 37322 3500 4 vdd
rlabel metal3 s 1410 10264 1470 10324 4 vdd
rlabel metal3 s 27324 284 27384 344 4 vdd
rlabel metal3 s 21702 3440 21762 3500 4 vdd
rlabel metal3 s 5836 19486 5896 19546 4 vdd
rlabel metal3 s 49710 3440 49770 3500 4 vdd
rlabel metal3 s 59046 3440 59106 3500 4 vdd
rlabel metal3 s 12542 284 12602 344 4 vdd
rlabel metal3 s 4632 10186 4692 10246 4 vdd
rlabel metal3 s 25146 4702 25206 4762 4 vdd
rlabel metal3 s 17034 3440 17094 3500 4 vdd
rlabel metal3 s 15478 3440 15538 3500 4 vdd
rlabel metal3 s 46598 3440 46658 3500 4 vdd
rlabel metal3 s 54378 3440 54438 3500 4 vdd
rlabel metal3 s 1410 16420 1470 16480 4 vdd
rlabel metal3 s 24990 284 25050 344 4 vdd
rlabel metal3 s 5836 22562 5896 22622 4 vdd
rlabel metal3 s 1410 19500 1470 19560 4 vdd
rlabel metal3 s 32594 3440 32654 3500 4 vdd
rlabel metal3 s 4632 25326 4692 25386 4 vdd
rlabel metal3 s 40374 3440 40434 3500 4 vdd
rlabel metal3 s 28258 4702 28318 4762 4 vdd
rlabel metal3 s 10208 284 10268 344 4 vdd
rlabel metal3 s 6474 4702 6534 4762 4 vdd
rlabel metal3 s 9586 4702 9646 4762 4 vdd
rlabel metal3 s 28880 284 28940 344 4 vdd
rlabel metal3 s 8652 284 8712 344 4 vdd
rlabel metal3 s 8030 4702 8090 4762 4 vdd
rlabel metal3 s 23590 4702 23650 4762 4 vdd
rlabel metal3 s 57490 3440 57550 3500 4 vdd
rlabel metal3 s 19544 284 19604 344 4 vdd
rlabel metal3 s 9430 284 9490 344 4 vdd
rlabel metal3 s 650 28736 710 28796 4 vdd
rlabel metal3 s 5836 13334 5896 13394 4 vdd
rlabel metal3 s 14684 2116 14744 2176 4 gnd
rlabel metal3 s 1410 24116 1470 24176 4 gnd
rlabel metal3 s 1410 14880 1470 14940 4 gnd
rlabel metal3 s 17796 2116 17856 2176 4 gnd
rlabel metal3 s 24020 2116 24080 2176 4 gnd
rlabel metal3 s 20130 2116 20190 2176 4 gnd
rlabel metal3 s 1410 21040 1470 21100 4 gnd
rlabel metal3 s 10794 2116 10854 2176 4 gnd
rlabel metal3 s 4632 8672 4692 8732 4 gnd
rlabel metal3 s 45042 4386 45102 4446 4 gnd
rlabel metal3 s 13128 2116 13188 2176 4 gnd
rlabel metal3 s 28688 2116 28748 2176 4 gnd
rlabel metal3 s 13906 2116 13966 2176 4 gnd
rlabel metal3 s 23242 2116 23302 2176 4 gnd
rlabel metal3 s 31038 4386 31098 4446 4 gnd
rlabel metal3 s 49710 4386 49770 4446 4 gnd
rlabel metal3 s 13922 4386 13982 4446 4 gnd
rlabel metal3 s 27926 4386 27986 4446 4 gnd
rlabel metal3 s 38818 4386 38878 4446 4 gnd
rlabel metal3 s 650 30276 710 30336 4 gnd
rlabel metal3 s 22464 2116 22524 2176 4 gnd
rlabel metal3 s 27910 2116 27970 2176 4 gnd
rlabel metal3 s 5836 17948 5896 18008 4 gnd
rlabel metal3 s 650 24116 710 24176 4 gnd
rlabel metal3 s 8460 2116 8520 2176 4 gnd
rlabel metal3 s 650 17960 710 18020 4 gnd
rlabel metal3 s 46598 4386 46658 4446 4 gnd
rlabel metal3 s 650 8724 710 8784 4 gnd
rlabel metal3 s 650 27196 710 27256 4 gnd
rlabel metal3 s 21686 2116 21746 2176 4 gnd
rlabel metal3 s 3774 2936 3834 2996 4 gnd
rlabel metal3 s 29482 4386 29542 4446 4 gnd
rlabel metal3 s 26354 2116 26414 2176 4 gnd
rlabel metal3 s 57490 4386 57550 4446 4 gnd
rlabel metal3 s 1410 11804 1470 11864 4 gnd
rlabel metal3 s 34150 4386 34210 4446 4 gnd
rlabel metal3 s 48154 4386 48214 4446 4 gnd
rlabel metal3 s 15462 2116 15522 2176 4 gnd
rlabel metal3 s 8030 5534 8090 5594 4 gnd
rlabel metal3 s 650 21040 710 21100 4 gnd
rlabel metal3 s 29814 5534 29874 5594 4 gnd
rlabel metal3 s 26702 5534 26762 5594 4 gnd
rlabel metal3 s 5836 11796 5896 11856 4 gnd
rlabel metal3 s 17018 2116 17078 2176 4 gnd
rlabel metal3 s 4632 14728 4692 14788 4 gnd
rlabel metal3 s 18922 5534 18982 5594 4 gnd
rlabel metal3 s 31022 2116 31082 2176 4 gnd
rlabel metal3 s 59046 4386 59106 4446 4 gnd
rlabel metal3 s 14254 5534 14314 5594 4 gnd
rlabel metal3 s 11142 5534 11202 5594 4 gnd
rlabel metal3 s 12350 2116 12410 2176 4 gnd
rlabel metal3 s 40374 4386 40434 4446 4 gnd
rlabel metal3 s 20908 2116 20968 2176 4 gnd
rlabel metal3 s 43486 4386 43546 4446 4 gnd
rlabel metal3 s 23590 5534 23650 5594 4 gnd
rlabel metal3 s 10016 2116 10076 2176 4 gnd
rlabel metal3 s 1410 27196 1470 27256 4 gnd
rlabel metal3 s 19352 2116 19412 2176 4 gnd
rlabel metal3 s 4632 20784 4692 20844 4 gnd
rlabel metal3 s 4632 29868 4692 29928 4 gnd
rlabel metal3 s 17034 4386 17094 4446 4 gnd
rlabel metal3 s 27132 2116 27192 2176 4 gnd
rlabel metal3 s 18574 2116 18634 2176 4 gnd
rlabel metal3 s 15478 4386 15538 4446 4 gnd
rlabel metal3 s 20478 5534 20538 5594 4 gnd
rlabel metal3 s 5836 14872 5896 14932 4 gnd
rlabel metal3 s 21702 4386 21762 4446 4 gnd
rlabel metal3 s 1410 17960 1470 18020 4 gnd
rlabel metal3 s 9586 5534 9646 5594 4 gnd
rlabel metal3 s 28258 5534 28318 5594 4 gnd
rlabel metal3 s 18590 4386 18650 4446 4 gnd
rlabel metal3 s 54378 4386 54438 4446 4 gnd
rlabel metal3 s 12698 5534 12758 5594 4 gnd
rlabel metal3 s 25576 2116 25636 2176 4 gnd
rlabel metal3 s 12366 4386 12426 4446 4 gnd
rlabel metal3 s 5836 5644 5896 5704 4 gnd
rlabel metal3 s 55934 4386 55994 4446 4 gnd
rlabel metal3 s 1410 5644 1470 5704 4 gnd
rlabel metal3 s 10810 4386 10870 4446 4 gnd
rlabel metal3 s 5836 8720 5896 8780 4 gnd
rlabel metal3 s 1410 8724 1470 8784 4 gnd
rlabel metal3 s 5836 21024 5896 21084 4 gnd
rlabel metal3 s 5836 24100 5896 24160 4 gnd
rlabel metal3 s 41930 4386 41990 4446 4 gnd
rlabel metal3 s 51266 4386 51326 4446 4 gnd
rlabel metal3 s 32594 4386 32654 4446 4 gnd
rlabel metal3 s 3774 4612 3834 4672 4 gnd
rlabel metal3 s 650 14880 710 14940 4 gnd
rlabel metal3 s 6904 2116 6964 2176 4 gnd
rlabel metal3 s 22034 5534 22094 5594 4 gnd
rlabel metal3 s 4632 23812 4692 23872 4 gnd
rlabel metal3 s 37262 4386 37322 4446 4 gnd
rlabel metal3 s 24814 4386 24874 4446 4 gnd
rlabel metal3 s 6474 5534 6534 5594 4 gnd
rlabel metal3 s 9238 2116 9298 2176 4 gnd
rlabel metal3 s 29466 2116 29526 2176 4 gnd
rlabel metal3 s 15810 5534 15870 5594 4 gnd
rlabel metal3 s 16240 2116 16300 2176 4 gnd
rlabel metal3 s 650 5644 710 5704 4 gnd
rlabel metal3 s 26370 4386 26430 4446 4 gnd
rlabel metal3 s 25146 5534 25206 5594 4 gnd
rlabel metal3 s 30244 2116 30304 2176 4 gnd
rlabel metal3 s 7682 2116 7742 2176 4 gnd
rlabel metal3 s 52822 4386 52882 4446 4 gnd
rlabel metal3 s 17366 5534 17426 5594 4 gnd
rlabel metal3 s 1410 30276 1470 30336 4 gnd
rlabel metal3 s 11572 2116 11632 2176 4 gnd
rlabel metal3 s 650 11804 710 11864 4 gnd
rlabel metal3 s 35706 4386 35766 4446 4 gnd
rlabel metal3 s 4632 17756 4692 17816 4 gnd
rlabel metal3 s 5836 27176 5896 27236 4 gnd
rlabel metal3 s 5836 30252 5896 30312 4 gnd
rlabel metal3 s 4632 11700 4692 11760 4 gnd
rlabel metal3 s 24798 2116 24858 2176 4 gnd
rlabel metal3 s 4632 26840 4692 26900 4 gnd
rlabel metal3 s 23258 4386 23318 4446 4 gnd
rlabel metal3 s 4632 5644 4692 5704 4 gnd
rlabel metal3 s 20146 4386 20206 4446 4 gnd
<< properties >>
string FIXED_BBOX 0 0 59296 30418
string GDS_FILE sram_0rw2r1w_16_32_sky130A.gds
string GDS_END 389026
string GDS_START 318910
<< end >>
