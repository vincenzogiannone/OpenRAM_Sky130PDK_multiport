magic
tech sky130A
timestamp 1647371806
<< nwell >>
rect 0 158 105 525
<< nmos >>
rect 45 61 60 103
<< pmos >>
rect 45 176 60 446
<< ndiff >>
rect 17 91 45 103
rect 17 74 21 91
rect 39 74 45 91
rect 17 61 45 74
rect 60 91 87 103
rect 60 74 66 91
rect 83 74 87 91
rect 60 61 87 74
<< pdiff >>
rect 18 415 45 446
rect 18 398 22 415
rect 39 398 45 415
rect 18 367 45 398
rect 18 350 22 367
rect 39 350 45 367
rect 18 319 45 350
rect 18 302 22 319
rect 39 302 45 319
rect 18 271 45 302
rect 18 254 22 271
rect 39 254 45 271
rect 18 223 45 254
rect 18 206 22 223
rect 39 206 45 223
rect 18 176 45 206
rect 60 415 87 446
rect 60 398 66 415
rect 83 398 87 415
rect 60 367 87 398
rect 60 350 66 367
rect 83 350 87 367
rect 60 319 87 350
rect 60 302 66 319
rect 83 302 87 319
rect 60 271 87 302
rect 60 254 66 271
rect 83 254 87 271
rect 60 223 87 254
rect 60 206 66 223
rect 83 206 87 223
rect 60 176 87 206
<< ndiffc >>
rect 21 74 39 91
rect 66 74 83 91
<< pdiffc >>
rect 22 398 39 415
rect 22 350 39 367
rect 22 302 39 319
rect 22 254 39 271
rect 22 206 39 223
rect 66 398 83 415
rect 66 350 83 367
rect 66 302 83 319
rect 66 254 83 271
rect 66 206 83 223
<< psubdiff >>
rect 31 26 73 34
rect 31 8 43 26
rect 61 8 73 26
rect 31 0 73 8
<< nsubdiff >>
rect 31 499 73 507
rect 31 481 43 499
rect 61 481 73 499
rect 31 473 73 481
<< psubdiffcont >>
rect 43 8 61 26
<< nsubdiffcont >>
rect 43 481 61 499
<< poly >>
rect 45 446 60 466
rect 45 153 60 176
rect 0 145 60 153
rect 0 128 5 145
rect 22 128 60 145
rect 0 120 60 128
rect 45 103 60 120
rect 45 48 60 61
<< polycont >>
rect 5 128 22 145
<< locali >>
rect 43 499 61 507
rect 25 481 43 490
rect 25 473 61 481
rect 25 446 43 473
rect 18 415 43 446
rect 18 398 22 415
rect 39 398 43 415
rect 18 367 43 398
rect 18 350 22 367
rect 39 350 43 367
rect 18 319 43 350
rect 18 302 22 319
rect 39 302 43 319
rect 18 271 43 302
rect 18 254 22 271
rect 39 254 43 271
rect 18 223 43 254
rect 18 206 22 223
rect 39 206 43 223
rect 18 176 43 206
rect 62 415 87 446
rect 62 398 66 415
rect 83 398 87 415
rect 62 367 87 398
rect 62 350 66 367
rect 83 350 87 367
rect 62 319 87 350
rect 62 302 66 319
rect 83 302 87 319
rect 62 271 87 302
rect 62 254 66 271
rect 83 254 87 271
rect 62 223 87 254
rect 62 206 66 223
rect 83 206 87 223
rect 62 176 87 206
rect 5 145 22 153
rect 5 120 22 128
rect 70 146 87 176
rect 70 103 87 129
rect 17 91 43 103
rect 17 74 21 91
rect 39 74 43 91
rect 17 61 43 74
rect 62 91 87 103
rect 62 74 66 91
rect 83 74 87 91
rect 62 61 87 74
rect 26 34 43 61
rect 26 26 61 34
rect 26 17 43 26
rect 43 0 61 8
<< viali >>
rect 43 481 61 499
rect 5 128 22 145
rect 70 129 87 146
rect 43 8 61 26
<< metal1 >>
rect 0 499 105 505
rect 0 481 43 499
rect 61 481 105 499
rect 0 475 105 481
rect 0 150 27 153
rect 0 124 1 150
rect 0 120 27 124
rect 62 151 94 154
rect 62 125 65 151
rect 91 125 94 151
rect 62 122 94 125
rect 0 26 105 32
rect 0 8 43 26
rect 61 8 105 26
rect 0 2 105 8
<< via1 >>
rect 1 145 27 150
rect 1 128 5 145
rect 5 128 22 145
rect 22 128 27 145
rect 1 124 27 128
rect 65 146 91 151
rect 65 129 70 146
rect 70 129 87 146
rect 87 129 91 146
rect 65 125 91 129
<< metal2 >>
rect 5 153 19 525
rect 74 154 88 525
rect 1 150 27 153
rect 1 120 27 124
rect 62 151 94 154
rect 62 125 65 151
rect 91 125 94 151
rect 62 122 94 125
rect 5 0 19 120
rect 74 0 88 122
<< labels >>
flabel metal2 81 49 81 49 0 FreeSans 80 0 0 0 dout
port 11 nsew
flabel metal1 18 17 18 17 0 FreeSans 80 0 0 0 gnd
port 7 nsew
flabel metal2 12 116 12 116 0 FreeSans 80 0 0 0 rbl
port 10 nsew
flabel metal1 15 491 15 491 0 FreeSans 80 0 0 0 vdd
port 6 nsew
<< properties >>
string FIXED_BBOX 0 0 105 525
<< end >>
