magic
tech sky130A
magscale 1 2
timestamp 1643671299
<< checkpaint >>
rect -1296 -1277 3240 2155
<< nwell >>
rect -36 402 1980 895
<< locali >>
rect 0 821 1944 855
rect 48 344 114 410
rect 196 360 432 394
rect 547 360 783 394
rect 902 360 1242 394
rect 1558 360 1592 394
rect 0 -17 1944 17
use pinv_8  pinv_8_0
timestamp 1643671299
transform 1 0 1161 0 1 0
box -36 -17 819 895
use pinv_7  pinv_7_0
timestamp 1643671299
transform 1 0 702 0 1 0
box -36 -17 495 895
use pinv_6  pinv_6_0
timestamp 1643671299
transform 1 0 351 0 1 0
box -36 -17 387 895
use pinv_6  pinv_6_1
timestamp 1643671299
transform 1 0 0 0 1 0
box -36 -17 387 895
<< labels >>
rlabel locali s 1575 377 1575 377 4 Z
rlabel locali s 81 377 81 377 4 A
rlabel locali s 972 0 972 0 4 gnd
rlabel locali s 972 838 972 838 4 vdd
<< properties >>
string FIXED_BBOX 0 0 1944 838
string GDS_FILE sram_0rw2r1w_16_32_sky130A.gds
string GDS_END 1195700
string GDS_START 1194556
<< end >>
