magic
tech sky130A
magscale 1 2
timestamp 1643678851
<< checkpaint >>
rect -1260 -1070 98552 7006
<< metal1 >>
rect 0 5338 47378 5366
rect 0 3110 49792 3138
rect 0 3052 49792 3080
rect 0 2994 49792 3022
rect 0 2936 49792 2964
rect 0 1171 50570 1199
<< metal2 >>
rect 196 5422 250 5450
rect 3308 5422 3362 5450
rect 6420 5422 6474 5450
rect 9532 5422 9586 5450
rect 12644 5422 12698 5450
rect 15756 5422 15810 5450
rect 18868 5422 18922 5450
rect 21980 5422 22034 5450
rect 25092 5422 25146 5450
rect 28204 5422 28258 5450
rect 31316 5422 31370 5450
rect 34428 5422 34482 5450
rect 37540 5422 37594 5450
rect 40652 5422 40706 5450
rect 43764 5422 43818 5450
rect 46876 5422 46930 5450
rect 630 4770 658 5400
rect 3742 4770 3770 5400
rect 6854 4770 6882 5400
rect 9966 4770 9994 5400
rect 750 4326 778 4566
rect 3862 4326 3890 4566
rect 6974 4326 7002 4566
rect 10086 4326 10114 4566
rect 13198 4326 13226 4566
rect 16310 4326 16338 4566
rect 19422 4326 19450 4566
rect 22534 4326 22562 4566
rect 25646 4326 25674 4566
rect 28758 4326 28786 4566
rect 31870 4326 31898 4566
rect 34982 4326 35010 4566
rect 38094 4326 38122 4566
rect 41206 4326 41234 4566
rect 44318 4326 44346 4566
rect 47430 4326 47458 4566
rect 68 1344 96 1398
rect 54 1316 96 1344
rect 54 204 82 1316
rect 710 1276 738 1398
rect 846 1344 874 1398
rect 532 1248 738 1276
rect 832 1316 874 1344
rect 532 204 560 1248
rect 832 204 860 1316
rect 1488 1276 1516 1398
rect 1624 1344 1652 1398
rect 1310 1248 1516 1276
rect 1610 1316 1652 1344
rect 1310 204 1338 1248
rect 1610 204 1638 1316
rect 2266 1276 2294 1398
rect 2402 1344 2430 1398
rect 2088 1248 2294 1276
rect 2388 1316 2430 1344
rect 2088 204 2116 1248
rect 2388 204 2416 1316
rect 3044 1276 3072 1398
rect 3180 1344 3208 1398
rect 2866 1248 3072 1276
rect 3166 1316 3208 1344
rect 2866 204 2894 1248
rect 3166 204 3194 1316
rect 3822 1276 3850 1398
rect 3958 1344 3986 1398
rect 3644 1248 3850 1276
rect 3944 1316 3986 1344
rect 3644 204 3672 1248
rect 3944 204 3972 1316
rect 4600 1276 4628 1398
rect 4736 1344 4764 1398
rect 4422 1248 4628 1276
rect 4722 1316 4764 1344
rect 4422 204 4450 1248
rect 4722 204 4750 1316
rect 5378 1276 5406 1398
rect 5514 1344 5542 1398
rect 5200 1248 5406 1276
rect 5500 1316 5542 1344
rect 5200 204 5228 1248
rect 5500 204 5528 1316
rect 6156 1276 6184 1398
rect 6292 1344 6320 1398
rect 5978 1248 6184 1276
rect 6278 1316 6320 1344
rect 5978 204 6006 1248
rect 6278 204 6306 1316
rect 6934 1276 6962 1398
rect 7070 1344 7098 1398
rect 6756 1248 6962 1276
rect 7056 1316 7098 1344
rect 6756 204 6784 1248
rect 7056 204 7084 1316
rect 7712 1276 7740 1398
rect 7848 1344 7876 1398
rect 7534 1248 7740 1276
rect 7834 1316 7876 1344
rect 7534 204 7562 1248
rect 7834 204 7862 1316
rect 8490 1276 8518 1398
rect 8626 1344 8654 1398
rect 8312 1248 8518 1276
rect 8612 1316 8654 1344
rect 8312 204 8340 1248
rect 8612 204 8640 1316
rect 9268 1276 9296 1398
rect 9404 1344 9432 1398
rect 9090 1248 9296 1276
rect 9390 1316 9432 1344
rect 9090 204 9118 1248
rect 9390 204 9418 1316
rect 10046 1276 10074 1398
rect 10182 1344 10210 1398
rect 9868 1248 10074 1276
rect 10168 1316 10210 1344
rect 9868 204 9896 1248
rect 10168 204 10196 1316
rect 10824 1276 10852 1398
rect 10960 1344 10988 1398
rect 10646 1248 10852 1276
rect 10946 1316 10988 1344
rect 10646 204 10674 1248
rect 10946 204 10974 1316
rect 11602 1276 11630 1398
rect 11738 1344 11766 1398
rect 11424 1248 11630 1276
rect 11724 1316 11766 1344
rect 11424 204 11452 1248
rect 11724 204 11752 1316
rect 12380 1276 12408 1398
rect 12516 1344 12544 1398
rect 12202 1248 12408 1276
rect 12502 1316 12544 1344
rect 12202 204 12230 1248
rect 12502 204 12530 1316
rect 13158 1276 13186 1398
rect 13294 1344 13322 1398
rect 12980 1248 13186 1276
rect 13280 1316 13322 1344
rect 12980 204 13008 1248
rect 13280 204 13308 1316
rect 13936 1276 13964 1398
rect 14072 1344 14100 1398
rect 13758 1248 13964 1276
rect 14058 1316 14100 1344
rect 13758 204 13786 1248
rect 14058 204 14086 1316
rect 14714 1276 14742 1398
rect 14850 1344 14878 1398
rect 14536 1248 14742 1276
rect 14836 1316 14878 1344
rect 14536 204 14564 1248
rect 14836 204 14864 1316
rect 15492 1276 15520 1398
rect 15628 1344 15656 1398
rect 15314 1248 15520 1276
rect 15614 1316 15656 1344
rect 15314 204 15342 1248
rect 15614 204 15642 1316
rect 16270 1276 16298 1398
rect 16406 1344 16434 1398
rect 16092 1248 16298 1276
rect 16392 1316 16434 1344
rect 16092 204 16120 1248
rect 16392 204 16420 1316
rect 17048 1276 17076 1398
rect 17184 1344 17212 1398
rect 16870 1248 17076 1276
rect 17170 1316 17212 1344
rect 16870 204 16898 1248
rect 17170 204 17198 1316
rect 17826 1276 17854 1398
rect 17962 1344 17990 1398
rect 17648 1248 17854 1276
rect 17948 1316 17990 1344
rect 17648 204 17676 1248
rect 17948 204 17976 1316
rect 18604 1276 18632 1398
rect 18740 1344 18768 1398
rect 18426 1248 18632 1276
rect 18726 1316 18768 1344
rect 18426 204 18454 1248
rect 18726 204 18754 1316
rect 19382 1276 19410 1398
rect 19518 1344 19546 1398
rect 19204 1248 19410 1276
rect 19504 1316 19546 1344
rect 19204 204 19232 1248
rect 19504 204 19532 1316
rect 20160 1276 20188 1398
rect 20296 1344 20324 1398
rect 19982 1248 20188 1276
rect 20282 1316 20324 1344
rect 19982 204 20010 1248
rect 20282 204 20310 1316
rect 20938 1276 20966 1398
rect 21074 1344 21102 1398
rect 20760 1248 20966 1276
rect 21060 1316 21102 1344
rect 20760 204 20788 1248
rect 21060 204 21088 1316
rect 21716 1276 21744 1398
rect 21852 1344 21880 1398
rect 21538 1248 21744 1276
rect 21838 1316 21880 1344
rect 21538 204 21566 1248
rect 21838 204 21866 1316
rect 22494 1276 22522 1398
rect 22630 1344 22658 1398
rect 22316 1248 22522 1276
rect 22616 1316 22658 1344
rect 22316 204 22344 1248
rect 22616 204 22644 1316
rect 23272 1276 23300 1398
rect 23408 1344 23436 1398
rect 23094 1248 23300 1276
rect 23394 1316 23436 1344
rect 23094 204 23122 1248
rect 23394 204 23422 1316
rect 24050 1276 24078 1398
rect 24186 1344 24214 1398
rect 23872 1248 24078 1276
rect 24172 1316 24214 1344
rect 23872 204 23900 1248
rect 24172 204 24200 1316
rect 24828 1276 24856 1398
rect 24964 1344 24992 1398
rect 24650 1248 24856 1276
rect 24950 1316 24992 1344
rect 24650 204 24678 1248
rect 24950 204 24978 1316
rect 25606 1276 25634 1398
rect 25742 1344 25770 1398
rect 25428 1248 25634 1276
rect 25728 1316 25770 1344
rect 25428 204 25456 1248
rect 25728 204 25756 1316
rect 26384 1276 26412 1398
rect 26520 1344 26548 1398
rect 26206 1248 26412 1276
rect 26506 1316 26548 1344
rect 26206 204 26234 1248
rect 26506 204 26534 1316
rect 27162 1276 27190 1398
rect 27298 1344 27326 1398
rect 26984 1248 27190 1276
rect 27284 1316 27326 1344
rect 26984 204 27012 1248
rect 27284 204 27312 1316
rect 27940 1276 27968 1398
rect 28076 1344 28104 1398
rect 27762 1248 27968 1276
rect 28062 1316 28104 1344
rect 27762 204 27790 1248
rect 28062 204 28090 1316
rect 28718 1276 28746 1398
rect 28854 1344 28882 1398
rect 28540 1248 28746 1276
rect 28840 1316 28882 1344
rect 28540 204 28568 1248
rect 28840 204 28868 1316
rect 29496 1276 29524 1398
rect 29632 1344 29660 1398
rect 29318 1248 29524 1276
rect 29618 1316 29660 1344
rect 29318 204 29346 1248
rect 29618 204 29646 1316
rect 30274 1276 30302 1398
rect 30410 1344 30438 1398
rect 30096 1248 30302 1276
rect 30396 1316 30438 1344
rect 30096 204 30124 1248
rect 30396 204 30424 1316
rect 31052 1276 31080 1398
rect 31188 1344 31216 1398
rect 30874 1248 31080 1276
rect 31174 1316 31216 1344
rect 30874 204 30902 1248
rect 31174 204 31202 1316
rect 31830 1276 31858 1398
rect 31966 1344 31994 1398
rect 31652 1248 31858 1276
rect 31952 1316 31994 1344
rect 31652 204 31680 1248
rect 31952 204 31980 1316
rect 32608 1276 32636 1398
rect 32744 1344 32772 1398
rect 32430 1248 32636 1276
rect 32730 1316 32772 1344
rect 32430 204 32458 1248
rect 32730 204 32758 1316
rect 33386 1276 33414 1398
rect 33522 1344 33550 1398
rect 33208 1248 33414 1276
rect 33508 1316 33550 1344
rect 33208 204 33236 1248
rect 33508 204 33536 1316
rect 34164 1276 34192 1398
rect 34300 1344 34328 1398
rect 33986 1248 34192 1276
rect 34286 1316 34328 1344
rect 33986 204 34014 1248
rect 34286 204 34314 1316
rect 34942 1276 34970 1398
rect 35078 1344 35106 1398
rect 34764 1248 34970 1276
rect 35064 1316 35106 1344
rect 34764 204 34792 1248
rect 35064 204 35092 1316
rect 35720 1276 35748 1398
rect 35856 1344 35884 1398
rect 35542 1248 35748 1276
rect 35842 1316 35884 1344
rect 35542 204 35570 1248
rect 35842 204 35870 1316
rect 36498 1276 36526 1398
rect 36634 1344 36662 1398
rect 36320 1248 36526 1276
rect 36620 1316 36662 1344
rect 36320 204 36348 1248
rect 36620 204 36648 1316
rect 37276 1276 37304 1398
rect 37412 1344 37440 1398
rect 37098 1248 37304 1276
rect 37398 1316 37440 1344
rect 37098 204 37126 1248
rect 37398 204 37426 1316
rect 38054 1276 38082 1398
rect 38190 1344 38218 1398
rect 37876 1248 38082 1276
rect 38176 1316 38218 1344
rect 37876 204 37904 1248
rect 38176 204 38204 1316
rect 38832 1276 38860 1398
rect 38968 1344 38996 1398
rect 38654 1248 38860 1276
rect 38954 1316 38996 1344
rect 38654 204 38682 1248
rect 38954 204 38982 1316
rect 39610 1276 39638 1398
rect 39746 1344 39774 1398
rect 39432 1248 39638 1276
rect 39732 1316 39774 1344
rect 39432 204 39460 1248
rect 39732 204 39760 1316
rect 40388 1276 40416 1398
rect 40524 1344 40552 1398
rect 40210 1248 40416 1276
rect 40510 1316 40552 1344
rect 40210 204 40238 1248
rect 40510 204 40538 1316
rect 41166 1276 41194 1398
rect 41302 1344 41330 1398
rect 40988 1248 41194 1276
rect 41288 1316 41330 1344
rect 40988 204 41016 1248
rect 41288 204 41316 1316
rect 41944 1276 41972 1398
rect 42080 1344 42108 1398
rect 41766 1248 41972 1276
rect 42066 1316 42108 1344
rect 41766 204 41794 1248
rect 42066 204 42094 1316
rect 42722 1276 42750 1398
rect 42858 1344 42886 1398
rect 42544 1248 42750 1276
rect 42844 1316 42886 1344
rect 42544 204 42572 1248
rect 42844 204 42872 1316
rect 43500 1276 43528 1398
rect 43636 1344 43664 1398
rect 43322 1248 43528 1276
rect 43622 1316 43664 1344
rect 43322 204 43350 1248
rect 43622 204 43650 1316
rect 44278 1276 44306 1398
rect 44414 1344 44442 1398
rect 44100 1248 44306 1276
rect 44400 1316 44442 1344
rect 44100 204 44128 1248
rect 44400 204 44428 1316
rect 45056 1276 45084 1398
rect 45192 1344 45220 1398
rect 44878 1248 45084 1276
rect 45178 1316 45220 1344
rect 44878 204 44906 1248
rect 45178 204 45206 1316
rect 45834 1276 45862 1398
rect 45970 1344 45998 1398
rect 45656 1248 45862 1276
rect 45956 1316 45998 1344
rect 45656 204 45684 1248
rect 45956 204 45984 1316
rect 46612 1276 46640 1398
rect 46748 1344 46776 1398
rect 46434 1248 46640 1276
rect 46734 1316 46776 1344
rect 46434 204 46462 1248
rect 46734 204 46762 1316
rect 47390 1276 47418 1398
rect 47526 1344 47554 1398
rect 47212 1248 47418 1276
rect 47512 1316 47554 1344
rect 47212 204 47240 1248
rect 47512 204 47540 1316
rect 48168 1276 48196 1398
rect 48304 1344 48332 1398
rect 47990 1248 48196 1276
rect 48290 1316 48332 1344
rect 47990 204 48018 1248
rect 48290 204 48318 1316
rect 48946 1276 48974 1398
rect 49082 1344 49110 1398
rect 48768 1248 48974 1276
rect 49068 1316 49110 1344
rect 48768 204 48796 1248
rect 49068 204 49096 1316
rect 49724 1276 49752 1398
rect 49546 1248 49752 1276
rect 49546 204 49574 1248
<< metal3 >>
rect 316 5614 382 5746
rect 3428 5614 3494 5746
rect 6540 5614 6606 5746
rect 9652 5614 9718 5746
rect 12764 5614 12830 5746
rect 15876 5614 15942 5746
rect 18988 5614 19054 5746
rect 22100 5614 22166 5746
rect 25212 5614 25278 5746
rect 28324 5614 28390 5746
rect 31436 5614 31502 5746
rect 34548 5614 34614 5746
rect 37660 5614 37726 5746
rect 40772 5614 40838 5746
rect 43884 5614 43950 5746
rect 46996 5614 47062 5746
rect 316 4782 382 4914
rect 3428 4782 3494 4914
rect 6540 4782 6606 4914
rect 9652 4782 9718 4914
rect 12764 4782 12830 4914
rect 15876 4782 15942 4914
rect 18988 4782 19054 4914
rect 22100 4782 22166 4914
rect 25212 4782 25278 4914
rect 28324 4782 28390 4914
rect 31436 4782 31502 4914
rect 34548 4782 34614 4914
rect 37660 4782 37726 4914
rect 40772 4782 40838 4914
rect 43884 4782 43950 4914
rect 46996 4782 47062 4914
rect 618 4499 750 4565
rect 3730 4499 3862 4565
rect 6842 4499 6974 4565
rect 9954 4499 10086 4565
rect 13066 4499 13198 4565
rect 16178 4499 16310 4565
rect 19290 4499 19422 4565
rect 22402 4499 22534 4565
rect 25514 4499 25646 4565
rect 28626 4499 28758 4565
rect 31738 4499 31870 4565
rect 34850 4499 34982 4565
rect 37962 4499 38094 4565
rect 41074 4499 41206 4565
rect 44186 4499 44318 4565
rect 47298 4499 47430 4565
rect 50410 4499 50542 4565
rect 53522 4499 53654 4565
rect 56634 4499 56766 4565
rect 59746 4499 59878 4565
rect 62858 4499 62990 4565
rect 65970 4499 66102 4565
rect 69082 4499 69214 4565
rect 72194 4499 72326 4565
rect 75306 4499 75438 4565
rect 78418 4499 78550 4565
rect 81530 4499 81662 4565
rect 84642 4499 84774 4565
rect 87754 4499 87886 4565
rect 90866 4499 90998 4565
rect 93978 4499 94110 4565
rect 97090 4499 97222 4565
rect 618 3553 750 3619
rect 3730 3553 3862 3619
rect 6842 3553 6974 3619
rect 9954 3553 10086 3619
rect 13066 3553 13198 3619
rect 16178 3553 16310 3619
rect 19290 3553 19422 3619
rect 22402 3553 22534 3619
rect 25514 3553 25646 3619
rect 28626 3553 28758 3619
rect 31738 3553 31870 3619
rect 34850 3553 34982 3619
rect 37962 3553 38094 3619
rect 41074 3553 41206 3619
rect 44186 3553 44318 3619
rect 47298 3553 47430 3619
rect 50410 3553 50542 3619
rect 53522 3553 53654 3619
rect 56634 3553 56766 3619
rect 59746 3553 59878 3619
rect 62858 3553 62990 3619
rect 65970 3553 66102 3619
rect 69082 3553 69214 3619
rect 72194 3553 72326 3619
rect 75306 3553 75438 3619
rect 78418 3553 78550 3619
rect 81530 3553 81662 3619
rect 84642 3553 84774 3619
rect 87754 3553 87886 3619
rect 90866 3553 90998 3619
rect 93978 3553 94110 3619
rect 97090 3553 97222 3619
rect 712 2114 844 2180
rect 1490 2114 1622 2180
rect 2268 2114 2400 2180
rect 3046 2114 3178 2180
rect 3824 2114 3956 2180
rect 4602 2114 4734 2180
rect 5380 2114 5512 2180
rect 6158 2114 6290 2180
rect 6936 2114 7068 2180
rect 7714 2114 7846 2180
rect 8492 2114 8624 2180
rect 9270 2114 9402 2180
rect 10048 2114 10180 2180
rect 10826 2114 10958 2180
rect 11604 2114 11736 2180
rect 12382 2114 12514 2180
rect 13160 2114 13292 2180
rect 13938 2114 14070 2180
rect 14716 2114 14848 2180
rect 15494 2114 15626 2180
rect 16272 2114 16404 2180
rect 17050 2114 17182 2180
rect 17828 2114 17960 2180
rect 18606 2114 18738 2180
rect 19384 2114 19516 2180
rect 20162 2114 20294 2180
rect 20940 2114 21072 2180
rect 21718 2114 21850 2180
rect 22496 2114 22628 2180
rect 23274 2114 23406 2180
rect 24052 2114 24184 2180
rect 24830 2114 24962 2180
rect 25608 2114 25740 2180
rect 26386 2114 26518 2180
rect 27164 2114 27296 2180
rect 27942 2114 28074 2180
rect 28720 2114 28852 2180
rect 29498 2114 29630 2180
rect 30276 2114 30408 2180
rect 31054 2114 31186 2180
rect 31832 2114 31964 2180
rect 32610 2114 32742 2180
rect 33388 2114 33520 2180
rect 34166 2114 34298 2180
rect 34944 2114 35076 2180
rect 35722 2114 35854 2180
rect 36500 2114 36632 2180
rect 37278 2114 37410 2180
rect 38056 2114 38188 2180
rect 38834 2114 38966 2180
rect 39612 2114 39744 2180
rect 40390 2114 40522 2180
rect 41168 2114 41300 2180
rect 41946 2114 42078 2180
rect 42724 2114 42856 2180
rect 43502 2114 43634 2180
rect 44280 2114 44412 2180
rect 45058 2114 45190 2180
rect 45836 2114 45968 2180
rect 46614 2114 46746 2180
rect 47392 2114 47524 2180
rect 48170 2114 48302 2180
rect 48948 2114 49080 2180
rect 49726 2114 49858 2180
rect 160 248 226 380
rect 938 248 1004 380
rect 1716 248 1782 380
rect 2494 248 2560 380
rect 3272 248 3338 380
rect 4050 248 4116 380
rect 4828 248 4894 380
rect 5606 248 5672 380
rect 6384 248 6450 380
rect 7162 248 7228 380
rect 7940 248 8006 380
rect 8718 248 8784 380
rect 9496 248 9562 380
rect 10274 248 10340 380
rect 11052 248 11118 380
rect 11830 248 11896 380
rect 12608 248 12674 380
rect 13386 248 13452 380
rect 14164 248 14230 380
rect 14942 248 15008 380
rect 15720 248 15786 380
rect 16498 248 16564 380
rect 17276 248 17342 380
rect 18054 248 18120 380
rect 18832 248 18898 380
rect 19610 248 19676 380
rect 20388 248 20454 380
rect 21166 248 21232 380
rect 21944 248 22010 380
rect 22722 248 22788 380
rect 23500 248 23566 380
rect 24278 248 24344 380
rect 25056 248 25122 380
rect 25834 248 25900 380
rect 26612 248 26678 380
rect 27390 248 27456 380
rect 28168 248 28234 380
rect 28946 248 29012 380
rect 29724 248 29790 380
rect 30502 248 30568 380
rect 31280 248 31346 380
rect 32058 248 32124 380
rect 32836 248 32902 380
rect 33614 248 33680 380
rect 34392 248 34458 380
rect 35170 248 35236 380
rect 35948 248 36014 380
rect 36726 248 36792 380
rect 37504 248 37570 380
rect 38282 248 38348 380
rect 39060 248 39126 380
rect 39838 248 39904 380
rect 40616 248 40682 380
rect 41394 248 41460 380
rect 42172 248 42238 380
rect 42950 248 43016 380
rect 43728 248 43794 380
rect 44506 248 44572 380
rect 45284 248 45350 380
rect 46062 248 46128 380
rect 46840 248 46906 380
rect 47618 248 47684 380
rect 48396 248 48462 380
rect 49174 248 49240 380
rect 49952 248 50018 380
use column_mux_array_multiport  column_mux_array_multiport_0
timestamp 1643678851
transform 1 0 0 0 -1 3312
box 0 32 49858 1914
use write_driver_array  write_driver_array_0
timestamp 1643678851
transform 1 0 0 0 -1 5722
box 0 -24 47378 952
use sense_amp_array  sense_amp_array_0
timestamp 1643678851
transform 1 0 0 0 -1 4566
box 548 0 97292 1050
use precharge_array_multiport  precharge_array_multiport_0
timestamp 1643678851
transform 1 0 0 0 -1 1194
box 0 -24 50570 1004
<< labels >>
rlabel metal2 s 196 5422 250 5450 4 din0_0
rlabel metal2 s 3308 5422 3362 5450 4 din0_1
rlabel metal2 s 6420 5422 6474 5450 4 din0_2
rlabel metal2 s 9532 5422 9586 5450 4 din0_3
rlabel metal2 s 12644 5422 12698 5450 4 din0_4
rlabel metal2 s 15756 5422 15810 5450 4 din0_5
rlabel metal2 s 18868 5422 18922 5450 4 din0_6
rlabel metal2 s 21980 5422 22034 5450 4 din0_7
rlabel metal2 s 25092 5422 25146 5450 4 din0_8
rlabel metal2 s 28204 5422 28258 5450 4 din0_9
rlabel metal2 s 31316 5422 31370 5450 4 din0_10
rlabel metal2 s 34428 5422 34482 5450 4 din0_11
rlabel metal2 s 37540 5422 37594 5450 4 din0_12
rlabel metal2 s 40652 5422 40706 5450 4 din0_13
rlabel metal2 s 43764 5422 43818 5450 4 din0_14
rlabel metal2 s 46876 5422 46930 5450 4 din0_15
rlabel metal2 s 750 4326 778 4566 4 dout0_0
rlabel metal2 s 764 4446 764 4446 4 dout1_0
rlabel metal2 s 3862 4326 3890 4566 4 dout0_1
rlabel metal2 s 3876 4446 3876 4446 4 dout1_1
rlabel metal2 s 6974 4326 7002 4566 4 dout0_2
rlabel metal2 s 6988 4446 6988 4446 4 dout1_2
rlabel metal2 s 10086 4326 10114 4566 4 dout0_3
rlabel metal2 s 10100 4446 10100 4446 4 dout1_3
rlabel metal2 s 13198 4326 13226 4566 4 dout0_4
rlabel metal2 s 13212 4446 13212 4446 4 dout1_4
rlabel metal2 s 16310 4326 16338 4566 4 dout0_5
rlabel metal2 s 16324 4446 16324 4446 4 dout1_5
rlabel metal2 s 19422 4326 19450 4566 4 dout0_6
rlabel metal2 s 19436 4446 19436 4446 4 dout1_6
rlabel metal2 s 22534 4326 22562 4566 4 dout0_7
rlabel metal2 s 22548 4446 22548 4446 4 dout1_7
rlabel metal2 s 25646 4326 25674 4566 4 dout0_8
rlabel metal2 s 25660 4446 25660 4446 4 dout1_8
rlabel metal2 s 28758 4326 28786 4566 4 dout0_9
rlabel metal2 s 28772 4446 28772 4446 4 dout1_9
rlabel metal2 s 31870 4326 31898 4566 4 dout0_10
rlabel metal2 s 31884 4446 31884 4446 4 dout1_10
rlabel metal2 s 34982 4326 35010 4566 4 dout0_11
rlabel metal2 s 34996 4446 34996 4446 4 dout1_11
rlabel metal2 s 38094 4326 38122 4566 4 dout0_12
rlabel metal2 s 38108 4446 38108 4446 4 dout1_12
rlabel metal2 s 41206 4326 41234 4566 4 dout0_13
rlabel metal2 s 41220 4446 41220 4446 4 dout1_13
rlabel metal2 s 44318 4326 44346 4566 4 dout0_14
rlabel metal2 s 44332 4446 44332 4446 4 dout1_14
rlabel metal2 s 47430 4326 47458 4566 4 dout0_15
rlabel metal2 s 47444 4446 47444 4446 4 dout1_15
rlabel metal2 s 54 204 82 1194 4 rbl0_0
rlabel metal2 s 532 204 560 1194 4 rbl1_0
rlabel metal2 s 832 204 860 1194 4 rbl0_1
rlabel metal2 s 1310 204 1338 1194 4 rbl1_1
rlabel metal2 s 1610 204 1638 1194 4 rbl0_2
rlabel metal2 s 2088 204 2116 1194 4 rbl1_2
rlabel metal2 s 2388 204 2416 1194 4 rbl0_3
rlabel metal2 s 2866 204 2894 1194 4 rbl1_3
rlabel metal2 s 3166 204 3194 1194 4 rbl0_4
rlabel metal2 s 3644 204 3672 1194 4 rbl1_4
rlabel metal2 s 3944 204 3972 1194 4 rbl0_5
rlabel metal2 s 4422 204 4450 1194 4 rbl1_5
rlabel metal2 s 4722 204 4750 1194 4 rbl0_6
rlabel metal2 s 5200 204 5228 1194 4 rbl1_6
rlabel metal2 s 5500 204 5528 1194 4 rbl0_7
rlabel metal2 s 5978 204 6006 1194 4 rbl1_7
rlabel metal2 s 6278 204 6306 1194 4 rbl0_8
rlabel metal2 s 6756 204 6784 1194 4 rbl1_8
rlabel metal2 s 7056 204 7084 1194 4 rbl0_9
rlabel metal2 s 7534 204 7562 1194 4 rbl1_9
rlabel metal2 s 7834 204 7862 1194 4 rbl0_10
rlabel metal2 s 8312 204 8340 1194 4 rbl1_10
rlabel metal2 s 8612 204 8640 1194 4 rbl0_11
rlabel metal2 s 9090 204 9118 1194 4 rbl1_11
rlabel metal2 s 9390 204 9418 1194 4 rbl0_12
rlabel metal2 s 9868 204 9896 1194 4 rbl1_12
rlabel metal2 s 10168 204 10196 1194 4 rbl0_13
rlabel metal2 s 10646 204 10674 1194 4 rbl1_13
rlabel metal2 s 10946 204 10974 1194 4 rbl0_14
rlabel metal2 s 11424 204 11452 1194 4 rbl1_14
rlabel metal2 s 11724 204 11752 1194 4 rbl0_15
rlabel metal2 s 12202 204 12230 1194 4 rbl1_15
rlabel metal2 s 12502 204 12530 1194 4 rbl0_16
rlabel metal2 s 12980 204 13008 1194 4 rbl1_16
rlabel metal2 s 13280 204 13308 1194 4 rbl0_17
rlabel metal2 s 13758 204 13786 1194 4 rbl1_17
rlabel metal2 s 14058 204 14086 1194 4 rbl0_18
rlabel metal2 s 14536 204 14564 1194 4 rbl1_18
rlabel metal2 s 14836 204 14864 1194 4 rbl0_19
rlabel metal2 s 15314 204 15342 1194 4 rbl1_19
rlabel metal2 s 15614 204 15642 1194 4 rbl0_20
rlabel metal2 s 16092 204 16120 1194 4 rbl1_20
rlabel metal2 s 16392 204 16420 1194 4 rbl0_21
rlabel metal2 s 16870 204 16898 1194 4 rbl1_21
rlabel metal2 s 17170 204 17198 1194 4 rbl0_22
rlabel metal2 s 17648 204 17676 1194 4 rbl1_22
rlabel metal2 s 17948 204 17976 1194 4 rbl0_23
rlabel metal2 s 18426 204 18454 1194 4 rbl1_23
rlabel metal2 s 18726 204 18754 1194 4 rbl0_24
rlabel metal2 s 19204 204 19232 1194 4 rbl1_24
rlabel metal2 s 19504 204 19532 1194 4 rbl0_25
rlabel metal2 s 19982 204 20010 1194 4 rbl1_25
rlabel metal2 s 20282 204 20310 1194 4 rbl0_26
rlabel metal2 s 20760 204 20788 1194 4 rbl1_26
rlabel metal2 s 21060 204 21088 1194 4 rbl0_27
rlabel metal2 s 21538 204 21566 1194 4 rbl1_27
rlabel metal2 s 21838 204 21866 1194 4 rbl0_28
rlabel metal2 s 22316 204 22344 1194 4 rbl1_28
rlabel metal2 s 22616 204 22644 1194 4 rbl0_29
rlabel metal2 s 23094 204 23122 1194 4 rbl1_29
rlabel metal2 s 23394 204 23422 1194 4 rbl0_30
rlabel metal2 s 23872 204 23900 1194 4 rbl1_30
rlabel metal2 s 24172 204 24200 1194 4 rbl0_31
rlabel metal2 s 24650 204 24678 1194 4 rbl1_31
rlabel metal2 s 24950 204 24978 1194 4 rbl0_32
rlabel metal2 s 25428 204 25456 1194 4 rbl1_32
rlabel metal2 s 25728 204 25756 1194 4 rbl0_33
rlabel metal2 s 26206 204 26234 1194 4 rbl1_33
rlabel metal2 s 26506 204 26534 1194 4 rbl0_34
rlabel metal2 s 26984 204 27012 1194 4 rbl1_34
rlabel metal2 s 27284 204 27312 1194 4 rbl0_35
rlabel metal2 s 27762 204 27790 1194 4 rbl1_35
rlabel metal2 s 28062 204 28090 1194 4 rbl0_36
rlabel metal2 s 28540 204 28568 1194 4 rbl1_36
rlabel metal2 s 28840 204 28868 1194 4 rbl0_37
rlabel metal2 s 29318 204 29346 1194 4 rbl1_37
rlabel metal2 s 29618 204 29646 1194 4 rbl0_38
rlabel metal2 s 30096 204 30124 1194 4 rbl1_38
rlabel metal2 s 30396 204 30424 1194 4 rbl0_39
rlabel metal2 s 30874 204 30902 1194 4 rbl1_39
rlabel metal2 s 31174 204 31202 1194 4 rbl0_40
rlabel metal2 s 31652 204 31680 1194 4 rbl1_40
rlabel metal2 s 31952 204 31980 1194 4 rbl0_41
rlabel metal2 s 32430 204 32458 1194 4 rbl1_41
rlabel metal2 s 32730 204 32758 1194 4 rbl0_42
rlabel metal2 s 33208 204 33236 1194 4 rbl1_42
rlabel metal2 s 33508 204 33536 1194 4 rbl0_43
rlabel metal2 s 33986 204 34014 1194 4 rbl1_43
rlabel metal2 s 34286 204 34314 1194 4 rbl0_44
rlabel metal2 s 34764 204 34792 1194 4 rbl1_44
rlabel metal2 s 35064 204 35092 1194 4 rbl0_45
rlabel metal2 s 35542 204 35570 1194 4 rbl1_45
rlabel metal2 s 35842 204 35870 1194 4 rbl0_46
rlabel metal2 s 36320 204 36348 1194 4 rbl1_46
rlabel metal2 s 36620 204 36648 1194 4 rbl0_47
rlabel metal2 s 37098 204 37126 1194 4 rbl1_47
rlabel metal2 s 37398 204 37426 1194 4 rbl0_48
rlabel metal2 s 37876 204 37904 1194 4 rbl1_48
rlabel metal2 s 38176 204 38204 1194 4 rbl0_49
rlabel metal2 s 38654 204 38682 1194 4 rbl1_49
rlabel metal2 s 38954 204 38982 1194 4 rbl0_50
rlabel metal2 s 39432 204 39460 1194 4 rbl1_50
rlabel metal2 s 39732 204 39760 1194 4 rbl0_51
rlabel metal2 s 40210 204 40238 1194 4 rbl1_51
rlabel metal2 s 40510 204 40538 1194 4 rbl0_52
rlabel metal2 s 40988 204 41016 1194 4 rbl1_52
rlabel metal2 s 41288 204 41316 1194 4 rbl0_53
rlabel metal2 s 41766 204 41794 1194 4 rbl1_53
rlabel metal2 s 42066 204 42094 1194 4 rbl0_54
rlabel metal2 s 42544 204 42572 1194 4 rbl1_54
rlabel metal2 s 42844 204 42872 1194 4 rbl0_55
rlabel metal2 s 43322 204 43350 1194 4 rbl1_55
rlabel metal2 s 43622 204 43650 1194 4 rbl0_56
rlabel metal2 s 44100 204 44128 1194 4 rbl1_56
rlabel metal2 s 44400 204 44428 1194 4 rbl0_57
rlabel metal2 s 44878 204 44906 1194 4 rbl1_57
rlabel metal2 s 45178 204 45206 1194 4 rbl0_58
rlabel metal2 s 45656 204 45684 1194 4 rbl1_58
rlabel metal2 s 45956 204 45984 1194 4 rbl0_59
rlabel metal2 s 46434 204 46462 1194 4 rbl1_59
rlabel metal2 s 46734 204 46762 1194 4 rbl0_60
rlabel metal2 s 47212 204 47240 1194 4 rbl1_60
rlabel metal2 s 47512 204 47540 1194 4 rbl0_61
rlabel metal2 s 47990 204 48018 1194 4 rbl1_61
rlabel metal2 s 48290 204 48318 1194 4 rbl0_62
rlabel metal2 s 48768 204 48796 1194 4 rbl1_62
rlabel metal2 s 49068 204 49096 1194 4 rbl0_63
rlabel metal2 s 49546 204 49574 1194 4 rbl1_63
rlabel metal2 s 630 4770 658 5400 4 wbl0_0
rlabel metal2 s 3742 4770 3770 5400 4 wbl0_1
rlabel metal2 s 6854 4770 6882 5400 4 wbl0_2
rlabel metal2 s 9966 4770 9994 5400 4 wbl0_3
rlabel metal1 s 0 1170 50570 1198 4 p_en_bar
rlabel metal1 s 0 3110 49792 3138 4 sel_0
rlabel metal1 s 0 3052 49792 3080 4 sel_1
rlabel metal1 s 0 2994 49792 3022 4 sel_2
rlabel metal1 s 0 2936 49792 2964 4 sel_3
rlabel metal1 s 0 5338 47378 5366 4 w_en
rlabel metal3 s 15720 248 15786 380 4 vdd
rlabel metal3 s 62858 3552 62990 3618 4 vdd
rlabel metal3 s 44506 248 44572 380 4 vdd
rlabel metal3 s 27390 248 27456 380 4 vdd
rlabel metal3 s 34850 3552 34982 3618 4 vdd
rlabel metal3 s 87754 3552 87886 3618 4 vdd
rlabel metal3 s 13386 248 13452 380 4 vdd
rlabel metal3 s 48396 248 48462 380 4 vdd
rlabel metal3 s 31436 4782 31502 4914 4 vdd
rlabel metal3 s 16498 248 16564 380 4 vdd
rlabel metal3 s 40772 4782 40838 4914 4 vdd
rlabel metal3 s 31280 248 31346 380 4 vdd
rlabel metal3 s 31738 3552 31870 3618 4 vdd
rlabel metal3 s 9954 3552 10086 3618 4 vdd
rlabel metal3 s 56634 3552 56766 3618 4 vdd
rlabel metal3 s 11052 248 11118 380 4 vdd
rlabel metal3 s 8718 248 8784 380 4 vdd
rlabel metal3 s 97090 3552 97222 3618 4 vdd
rlabel metal3 s 618 3552 750 3618 4 vdd
rlabel metal3 s 12764 4782 12830 4914 4 vdd
rlabel metal3 s 40616 248 40682 380 4 vdd
rlabel metal3 s 6842 3552 6974 3618 4 vdd
rlabel metal3 s 28324 4782 28390 4914 4 vdd
rlabel metal3 s 11830 248 11896 380 4 vdd
rlabel metal3 s 7940 248 8006 380 4 vdd
rlabel metal3 s 19290 3552 19422 3618 4 vdd
rlabel metal3 s 7162 248 7228 380 4 vdd
rlabel metal3 s 10274 248 10340 380 4 vdd
rlabel metal3 s 65970 3552 66102 3618 4 vdd
rlabel metal3 s 46996 4782 47062 4914 4 vdd
rlabel metal3 s 34392 248 34458 380 4 vdd
rlabel metal3 s 47298 3552 47430 3618 4 vdd
rlabel metal3 s 35948 248 36014 380 4 vdd
rlabel metal3 s 39060 248 39126 380 4 vdd
rlabel metal3 s 22100 4782 22166 4914 4 vdd
rlabel metal3 s 42172 248 42238 380 4 vdd
rlabel metal3 s 18832 248 18898 380 4 vdd
rlabel metal3 s 53522 3552 53654 3618 4 vdd
rlabel metal3 s 43728 248 43794 380 4 vdd
rlabel metal3 s 28626 3552 28758 3618 4 vdd
rlabel metal3 s 36726 248 36792 380 4 vdd
rlabel metal3 s 5606 248 5672 380 4 vdd
rlabel metal3 s 28946 248 29012 380 4 vdd
rlabel metal3 s 47618 248 47684 380 4 vdd
rlabel metal3 s 37962 3552 38094 3618 4 vdd
rlabel metal3 s 26612 248 26678 380 4 vdd
rlabel metal3 s 32836 248 32902 380 4 vdd
rlabel metal3 s 12608 248 12674 380 4 vdd
rlabel metal3 s 16178 3552 16310 3618 4 vdd
rlabel metal3 s 6384 248 6450 380 4 vdd
rlabel metal3 s 75306 3552 75438 3618 4 vdd
rlabel metal3 s 6540 4782 6606 4914 4 vdd
rlabel metal3 s 90866 3552 90998 3618 4 vdd
rlabel metal3 s 9496 248 9562 380 4 vdd
rlabel metal3 s 30502 248 30568 380 4 vdd
rlabel metal3 s 44186 3552 44318 3618 4 vdd
rlabel metal3 s 81530 3552 81662 3618 4 vdd
rlabel metal3 s 22402 3552 22534 3618 4 vdd
rlabel metal3 s 34548 4782 34614 4914 4 vdd
rlabel metal3 s 3272 248 3338 380 4 vdd
rlabel metal3 s 19610 248 19676 380 4 vdd
rlabel metal3 s 4050 248 4116 380 4 vdd
rlabel metal3 s 3428 4782 3494 4914 4 vdd
rlabel metal3 s 22722 248 22788 380 4 vdd
rlabel metal3 s 25834 248 25900 380 4 vdd
rlabel metal3 s 72194 3552 72326 3618 4 vdd
rlabel metal3 s 35170 248 35236 380 4 vdd
rlabel metal3 s 45284 248 45350 380 4 vdd
rlabel metal3 s 316 4782 382 4914 4 vdd
rlabel metal3 s 1716 248 1782 380 4 vdd
rlabel metal3 s 69082 3552 69214 3618 4 vdd
rlabel metal3 s 2494 248 2560 380 4 vdd
rlabel metal3 s 37660 4782 37726 4914 4 vdd
rlabel metal3 s 25212 4782 25278 4914 4 vdd
rlabel metal3 s 78418 3552 78550 3618 4 vdd
rlabel metal3 s 3730 3552 3862 3618 4 vdd
rlabel metal3 s 42950 248 43016 380 4 vdd
rlabel metal3 s 9652 4782 9718 4914 4 vdd
rlabel metal3 s 59746 3552 59878 3618 4 vdd
rlabel metal3 s 20388 248 20454 380 4 vdd
rlabel metal3 s 46840 248 46906 380 4 vdd
rlabel metal3 s 4828 248 4894 380 4 vdd
rlabel metal3 s 14942 248 15008 380 4 vdd
rlabel metal3 s 50410 3552 50542 3618 4 vdd
rlabel metal3 s 32058 248 32124 380 4 vdd
rlabel metal3 s 21166 248 21232 380 4 vdd
rlabel metal3 s 160 248 226 380 4 vdd
rlabel metal3 s 29724 248 29790 380 4 vdd
rlabel metal3 s 17276 248 17342 380 4 vdd
rlabel metal3 s 41394 248 41460 380 4 vdd
rlabel metal3 s 37504 248 37570 380 4 vdd
rlabel metal3 s 18054 248 18120 380 4 vdd
rlabel metal3 s 49174 248 49240 380 4 vdd
rlabel metal3 s 84642 3552 84774 3618 4 vdd
rlabel metal3 s 93978 3552 94110 3618 4 vdd
rlabel metal3 s 21944 248 22010 380 4 vdd
rlabel metal3 s 23500 248 23566 380 4 vdd
rlabel metal3 s 43884 4782 43950 4914 4 vdd
rlabel metal3 s 14164 248 14230 380 4 vdd
rlabel metal3 s 24278 248 24344 380 4 vdd
rlabel metal3 s 15876 4782 15942 4914 4 vdd
rlabel metal3 s 33614 248 33680 380 4 vdd
rlabel metal3 s 49952 248 50018 380 4 vdd
rlabel metal3 s 46062 248 46128 380 4 vdd
rlabel metal3 s 38282 248 38348 380 4 vdd
rlabel metal3 s 39838 248 39904 380 4 vdd
rlabel metal3 s 25056 248 25122 380 4 vdd
rlabel metal3 s 938 248 1004 380 4 vdd
rlabel metal3 s 28168 248 28234 380 4 vdd
rlabel metal3 s 13066 3552 13198 3618 4 vdd
rlabel metal3 s 18988 4782 19054 4914 4 vdd
rlabel metal3 s 25514 3552 25646 3618 4 vdd
rlabel metal3 s 41074 3552 41206 3618 4 vdd
rlabel metal3 s 28720 2114 28852 2180 4 gnd
rlabel metal3 s 72194 4498 72326 4564 4 gnd
rlabel metal3 s 24052 2114 24184 2180 4 gnd
rlabel metal3 s 2268 2114 2400 2180 4 gnd
rlabel metal3 s 38834 2114 38966 2180 4 gnd
rlabel metal3 s 1490 2114 1622 2180 4 gnd
rlabel metal3 s 87754 4498 87886 4564 4 gnd
rlabel metal3 s 43502 2114 43634 2180 4 gnd
rlabel metal3 s 19384 2114 19516 2180 4 gnd
rlabel metal3 s 25212 5614 25278 5746 4 gnd
rlabel metal3 s 21718 2114 21850 2180 4 gnd
rlabel metal3 s 78418 4498 78550 4564 4 gnd
rlabel metal3 s 56634 4498 56766 4564 4 gnd
rlabel metal3 s 34548 5614 34614 5746 4 gnd
rlabel metal3 s 35722 2114 35854 2180 4 gnd
rlabel metal3 s 11604 2114 11736 2180 4 gnd
rlabel metal3 s 46614 2114 46746 2180 4 gnd
rlabel metal3 s 45836 2114 45968 2180 4 gnd
rlabel metal3 s 37278 2114 37410 2180 4 gnd
rlabel metal3 s 37660 5614 37726 5746 4 gnd
rlabel metal3 s 37962 4498 38094 4564 4 gnd
rlabel metal3 s 42724 2114 42856 2180 4 gnd
rlabel metal3 s 16272 2114 16404 2180 4 gnd
rlabel metal3 s 48948 2114 49080 2180 4 gnd
rlabel metal3 s 75306 4498 75438 4564 4 gnd
rlabel metal3 s 16178 4498 16310 4564 4 gnd
rlabel metal3 s 45058 2114 45190 2180 4 gnd
rlabel metal3 s 28626 4498 28758 4564 4 gnd
rlabel metal3 s 24830 2114 24962 2180 4 gnd
rlabel metal3 s 40390 2114 40522 2180 4 gnd
rlabel metal3 s 13938 2114 14070 2180 4 gnd
rlabel metal3 s 43884 5614 43950 5746 4 gnd
rlabel metal3 s 41074 4498 41206 4564 4 gnd
rlabel metal3 s 32610 2114 32742 2180 4 gnd
rlabel metal3 s 97090 4498 97222 4564 4 gnd
rlabel metal3 s 17828 2114 17960 2180 4 gnd
rlabel metal3 s 29498 2114 29630 2180 4 gnd
rlabel metal3 s 6842 4498 6974 4564 4 gnd
rlabel metal3 s 22496 2114 22628 2180 4 gnd
rlabel metal3 s 9270 2114 9402 2180 4 gnd
rlabel metal3 s 48170 2114 48302 2180 4 gnd
rlabel metal3 s 93978 4498 94110 4564 4 gnd
rlabel metal3 s 30276 2114 30408 2180 4 gnd
rlabel metal3 s 47392 2114 47524 2180 4 gnd
rlabel metal3 s 3730 4498 3862 4564 4 gnd
rlabel metal3 s 13160 2114 13292 2180 4 gnd
rlabel metal3 s 18988 5614 19054 5746 4 gnd
rlabel metal3 s 34944 2114 35076 2180 4 gnd
rlabel metal3 s 31738 4498 31870 4564 4 gnd
rlabel metal3 s 3428 5614 3494 5746 4 gnd
rlabel metal3 s 41946 2114 42078 2180 4 gnd
rlabel metal3 s 44280 2114 44412 2180 4 gnd
rlabel metal3 s 9652 5614 9718 5746 4 gnd
rlabel metal3 s 12764 5614 12830 5746 4 gnd
rlabel metal3 s 7714 2114 7846 2180 4 gnd
rlabel metal3 s 53522 4498 53654 4564 4 gnd
rlabel metal3 s 12382 2114 12514 2180 4 gnd
rlabel metal3 s 618 4498 750 4564 4 gnd
rlabel metal3 s 10048 2114 10180 2180 4 gnd
rlabel metal3 s 22402 4498 22534 4564 4 gnd
rlabel metal3 s 26386 2114 26518 2180 4 gnd
rlabel metal3 s 84642 4498 84774 4564 4 gnd
rlabel metal3 s 50410 4498 50542 4564 4 gnd
rlabel metal3 s 25514 4498 25646 4564 4 gnd
rlabel metal3 s 40772 5614 40838 5746 4 gnd
rlabel metal3 s 17050 2114 17182 2180 4 gnd
rlabel metal3 s 6540 5614 6606 5746 4 gnd
rlabel metal3 s 9954 4498 10086 4564 4 gnd
rlabel metal3 s 6936 2114 7068 2180 4 gnd
rlabel metal3 s 34166 2114 34298 2180 4 gnd
rlabel metal3 s 39612 2114 39744 2180 4 gnd
rlabel metal3 s 62858 4498 62990 4564 4 gnd
rlabel metal3 s 31054 2114 31186 2180 4 gnd
rlabel metal3 s 19290 4498 19422 4564 4 gnd
rlabel metal3 s 14716 2114 14848 2180 4 gnd
rlabel metal3 s 47298 4498 47430 4564 4 gnd
rlabel metal3 s 49726 2114 49858 2180 4 gnd
rlabel metal3 s 31436 5614 31502 5746 4 gnd
rlabel metal3 s 46996 5614 47062 5746 4 gnd
rlabel metal3 s 44186 4498 44318 4564 4 gnd
rlabel metal3 s 712 2114 844 2180 4 gnd
rlabel metal3 s 316 5614 382 5746 4 gnd
rlabel metal3 s 10826 2114 10958 2180 4 gnd
rlabel metal3 s 65970 4498 66102 4564 4 gnd
rlabel metal3 s 28324 5614 28390 5746 4 gnd
rlabel metal3 s 22100 5614 22166 5746 4 gnd
rlabel metal3 s 5380 2114 5512 2180 4 gnd
rlabel metal3 s 31832 2114 31964 2180 4 gnd
rlabel metal3 s 34850 4498 34982 4564 4 gnd
rlabel metal3 s 27164 2114 27296 2180 4 gnd
rlabel metal3 s 3824 2114 3956 2180 4 gnd
rlabel metal3 s 4602 2114 4734 2180 4 gnd
rlabel metal3 s 20940 2114 21072 2180 4 gnd
rlabel metal3 s 36500 2114 36632 2180 4 gnd
rlabel metal3 s 33388 2114 33520 2180 4 gnd
rlabel metal3 s 27942 2114 28074 2180 4 gnd
rlabel metal3 s 15876 5614 15942 5746 4 gnd
rlabel metal3 s 38056 2114 38188 2180 4 gnd
rlabel metal3 s 69082 4498 69214 4564 4 gnd
rlabel metal3 s 59746 4498 59878 4564 4 gnd
rlabel metal3 s 90866 4498 90998 4564 4 gnd
rlabel metal3 s 6158 2114 6290 2180 4 gnd
rlabel metal3 s 13066 4498 13198 4564 4 gnd
rlabel metal3 s 18606 2114 18738 2180 4 gnd
rlabel metal3 s 25608 2114 25740 2180 4 gnd
rlabel metal3 s 8492 2114 8624 2180 4 gnd
rlabel metal3 s 20162 2114 20294 2180 4 gnd
rlabel metal3 s 81530 4498 81662 4564 4 gnd
rlabel metal3 s 15494 2114 15626 2180 4 gnd
rlabel metal3 s 41168 2114 41300 2180 4 gnd
rlabel metal3 s 23274 2114 23406 2180 4 gnd
rlabel metal3 s 3046 2114 3178 2180 4 gnd
<< properties >>
string FIXED_BBOX 0 0 97292 5722
string GDS_FILE sram_0rw2r1w_16_128_sky130A.gds
string GDS_END 1434000
string GDS_START 1315592
<< end >>
