magic
tech sky130A
magscale 1 2
timestamp 1644951705
<< checkpaint >>
rect -1296 -1277 1664 2155
<< nwell >>
rect -36 402 404 895
<< locali >>
rect 0 821 368 855
rect 48 344 114 410
rect 179 360 213 394
rect 0 -17 368 17
use pinv_0  pinv_0_0
timestamp 1644951705
transform 1 0 0 0 1 0
box -36 -17 404 895
<< labels >>
rlabel locali s 196 377 196 377 4 Z
rlabel locali s 81 377 81 377 4 A
rlabel locali s 184 0 184 0 4 gnd
rlabel locali s 184 838 184 838 4 vdd
<< properties >>
string FIXED_BBOX 0 0 368 838
string GDS_FILE sram_0rw2r1w_16_128_sky130A.gds
string GDS_END 1934632
string GDS_START 1933788
<< end >>
