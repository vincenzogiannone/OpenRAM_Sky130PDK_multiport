magic
tech sky130A
magscale 1 2
timestamp 1643593061
<< checkpaint >>
rect -1260 -1302 2742 2176
<< nwell >>
rect 0 436 1482 916
<< pwell >>
rect 140 -42 212 42
rect 422 -42 494 42
rect 704 -42 776 42
rect 986 -42 1058 42
rect 1268 -42 1340 42
<< nmos >>
rect 108 96 138 180
rect 220 96 250 180
rect 332 96 362 180
rect 444 96 474 180
rect 556 96 586 180
rect 668 96 698 180
rect 780 96 810 180
rect 892 96 922 180
rect 1004 96 1034 180
rect 1116 96 1146 180
rect 1344 96 1374 180
<< pmos >>
rect 108 472 138 742
rect 220 472 250 742
rect 332 472 362 742
rect 444 472 474 742
rect 556 472 586 742
rect 668 472 698 742
rect 780 472 810 742
rect 892 472 922 742
rect 1004 472 1034 742
rect 1116 472 1146 742
rect 1344 472 1374 742
<< ndiff >>
rect 36 154 108 180
rect 36 120 50 154
rect 84 120 108 154
rect 36 96 108 120
rect 138 154 220 180
rect 138 120 162 154
rect 196 120 220 154
rect 138 96 220 120
rect 250 154 332 180
rect 250 120 274 154
rect 308 120 332 154
rect 250 96 332 120
rect 362 154 444 180
rect 362 120 386 154
rect 420 120 444 154
rect 362 96 444 120
rect 474 96 556 180
rect 586 154 668 180
rect 586 120 610 154
rect 644 120 668 154
rect 586 96 668 120
rect 698 154 780 180
rect 698 120 722 154
rect 756 120 780 154
rect 698 96 780 120
rect 810 154 892 180
rect 810 120 834 154
rect 868 120 892 154
rect 810 96 892 120
rect 922 96 1004 180
rect 1034 154 1116 180
rect 1034 120 1058 154
rect 1092 120 1116 154
rect 1034 96 1116 120
rect 1146 154 1218 180
rect 1146 120 1170 154
rect 1204 120 1218 154
rect 1146 96 1218 120
rect 1272 154 1344 180
rect 1272 120 1286 154
rect 1320 120 1344 154
rect 1272 96 1344 120
rect 1374 154 1446 180
rect 1374 120 1398 154
rect 1432 120 1446 154
rect 1374 96 1446 120
<< pdiff >>
rect 36 700 108 742
rect 36 666 50 700
rect 84 666 108 700
rect 36 624 108 666
rect 36 590 50 624
rect 84 590 108 624
rect 36 548 108 590
rect 36 514 50 548
rect 84 514 108 548
rect 36 472 108 514
rect 138 700 220 742
rect 138 666 162 700
rect 196 666 220 700
rect 138 624 220 666
rect 138 590 162 624
rect 196 590 220 624
rect 138 548 220 590
rect 138 514 162 548
rect 196 514 220 548
rect 138 472 220 514
rect 250 700 332 742
rect 250 666 274 700
rect 308 666 332 700
rect 250 624 332 666
rect 250 590 274 624
rect 308 590 332 624
rect 250 548 332 590
rect 250 514 274 548
rect 308 514 332 548
rect 250 472 332 514
rect 362 700 444 742
rect 362 666 386 700
rect 420 666 444 700
rect 362 624 444 666
rect 362 590 386 624
rect 420 590 444 624
rect 362 548 444 590
rect 362 514 386 548
rect 420 514 444 548
rect 362 472 444 514
rect 474 472 556 742
rect 586 700 668 742
rect 586 666 610 700
rect 644 666 668 700
rect 586 624 668 666
rect 586 590 610 624
rect 644 590 668 624
rect 586 548 668 590
rect 586 514 610 548
rect 644 514 668 548
rect 586 472 668 514
rect 698 700 780 742
rect 698 666 722 700
rect 756 666 780 700
rect 698 624 780 666
rect 698 590 722 624
rect 756 590 780 624
rect 698 548 780 590
rect 698 514 722 548
rect 756 514 780 548
rect 698 472 780 514
rect 810 700 892 742
rect 810 666 834 700
rect 868 666 892 700
rect 810 624 892 666
rect 810 590 834 624
rect 868 590 892 624
rect 810 548 892 590
rect 810 514 834 548
rect 868 514 892 548
rect 810 472 892 514
rect 922 472 1004 742
rect 1034 700 1116 742
rect 1034 666 1058 700
rect 1092 666 1116 700
rect 1034 624 1116 666
rect 1034 590 1058 624
rect 1092 590 1116 624
rect 1034 548 1116 590
rect 1034 514 1058 548
rect 1092 514 1116 548
rect 1034 472 1116 514
rect 1146 700 1218 742
rect 1146 666 1170 700
rect 1204 666 1218 700
rect 1146 624 1218 666
rect 1146 590 1170 624
rect 1204 590 1218 624
rect 1146 548 1218 590
rect 1146 514 1170 548
rect 1204 514 1218 548
rect 1146 472 1218 514
rect 1272 700 1344 742
rect 1272 666 1286 700
rect 1320 666 1344 700
rect 1272 624 1344 666
rect 1272 590 1286 624
rect 1320 590 1344 624
rect 1272 548 1344 590
rect 1272 514 1286 548
rect 1320 514 1344 548
rect 1272 472 1344 514
rect 1374 700 1446 742
rect 1374 666 1398 700
rect 1432 666 1446 700
rect 1374 624 1446 666
rect 1374 590 1398 624
rect 1432 590 1446 624
rect 1374 548 1446 590
rect 1374 514 1398 548
rect 1432 514 1446 548
rect 1374 472 1446 514
<< ndiffc >>
rect 50 120 84 154
rect 162 120 196 154
rect 274 120 308 154
rect 386 120 420 154
rect 610 120 644 154
rect 722 120 756 154
rect 834 120 868 154
rect 1058 120 1092 154
rect 1170 120 1204 154
rect 1286 120 1320 154
rect 1398 120 1432 154
<< pdiffc >>
rect 50 666 84 700
rect 50 590 84 624
rect 50 514 84 548
rect 162 666 196 700
rect 162 590 196 624
rect 162 514 196 548
rect 274 666 308 700
rect 274 590 308 624
rect 274 514 308 548
rect 386 666 420 700
rect 386 590 420 624
rect 386 514 420 548
rect 610 666 644 700
rect 610 590 644 624
rect 610 514 644 548
rect 722 666 756 700
rect 722 590 756 624
rect 722 514 756 548
rect 834 666 868 700
rect 834 590 868 624
rect 834 514 868 548
rect 1058 666 1092 700
rect 1058 590 1092 624
rect 1058 514 1092 548
rect 1170 666 1204 700
rect 1170 590 1204 624
rect 1170 514 1204 548
rect 1286 666 1320 700
rect 1286 590 1320 624
rect 1286 514 1320 548
rect 1398 666 1432 700
rect 1398 590 1432 624
rect 1398 514 1432 548
<< psubdiff >>
rect 140 17 212 42
rect 140 -17 159 17
rect 193 -17 212 17
rect 140 -42 212 -17
rect 422 17 494 42
rect 422 -17 441 17
rect 475 -17 494 17
rect 422 -42 494 -17
rect 704 17 776 42
rect 704 -17 723 17
rect 757 -17 776 17
rect 704 -42 776 -17
rect 986 17 1058 42
rect 986 -17 1005 17
rect 1039 -17 1058 17
rect 986 -42 1058 -17
rect 1268 17 1340 42
rect 1268 -17 1287 17
rect 1321 -17 1340 17
rect 1268 -42 1340 -17
<< nsubdiff >>
rect 140 855 212 880
rect 140 821 159 855
rect 193 821 212 855
rect 140 796 212 821
rect 422 855 494 880
rect 422 821 441 855
rect 475 821 494 855
rect 422 796 494 821
rect 704 855 776 880
rect 704 821 723 855
rect 757 821 776 855
rect 704 796 776 821
rect 986 855 1058 880
rect 986 821 1005 855
rect 1039 821 1058 855
rect 986 796 1058 821
rect 1268 855 1340 880
rect 1268 821 1287 855
rect 1321 821 1340 855
rect 1268 796 1340 821
<< psubdiffcont >>
rect 159 -17 193 17
rect 441 -17 475 17
rect 723 -17 757 17
rect 1005 -17 1039 17
rect 1287 -17 1321 17
<< nsubdiffcont >>
rect 159 821 193 855
rect 441 821 475 855
rect 723 821 757 855
rect 1005 821 1039 855
rect 1287 821 1321 855
<< poly >>
rect 108 742 138 768
rect 220 742 250 768
rect 332 742 362 768
rect 444 742 474 768
rect 556 742 586 768
rect 668 742 698 768
rect 780 742 810 768
rect 892 742 922 768
rect 1004 742 1034 768
rect 1116 742 1146 768
rect 1344 742 1374 768
rect 108 370 138 472
rect 0 354 138 370
rect 0 320 10 354
rect 44 340 138 354
rect 44 320 54 340
rect 0 304 54 320
rect 108 180 138 340
rect 220 280 250 472
rect 332 438 362 472
rect 444 438 474 472
rect 556 438 586 472
rect 320 422 374 438
rect 320 388 330 422
rect 364 388 374 422
rect 320 372 374 388
rect 444 422 512 438
rect 444 388 468 422
rect 502 388 512 422
rect 444 372 512 388
rect 556 422 610 438
rect 556 388 566 422
rect 600 388 610 422
rect 556 372 610 388
rect 180 264 250 280
rect 180 230 190 264
rect 224 230 250 264
rect 180 214 250 230
rect 320 264 374 280
rect 320 230 330 264
rect 364 230 374 264
rect 320 214 374 230
rect 444 254 512 270
rect 444 220 468 254
rect 502 220 512 254
rect 220 180 250 214
rect 332 180 362 214
rect 444 204 512 220
rect 444 180 474 204
rect 556 180 586 372
rect 668 330 698 472
rect 780 438 810 472
rect 892 438 922 472
rect 1004 438 1034 472
rect 768 422 822 438
rect 768 388 778 422
rect 812 388 822 422
rect 768 372 822 388
rect 892 422 960 438
rect 892 388 916 422
rect 950 388 960 422
rect 892 372 960 388
rect 1004 422 1058 438
rect 1004 388 1014 422
rect 1048 388 1058 422
rect 1004 372 1058 388
rect 628 314 698 330
rect 628 280 638 314
rect 672 280 698 314
rect 628 264 698 280
rect 668 180 698 264
rect 768 264 822 280
rect 768 230 778 264
rect 812 230 822 264
rect 768 214 822 230
rect 892 254 960 270
rect 892 220 916 254
rect 950 220 960 254
rect 780 180 810 214
rect 892 204 960 220
rect 892 180 922 204
rect 1004 180 1034 372
rect 1116 330 1146 472
rect 1344 438 1374 472
rect 1320 422 1374 438
rect 1320 388 1330 422
rect 1364 388 1374 422
rect 1320 372 1374 388
rect 1076 314 1146 330
rect 1076 280 1086 314
rect 1120 280 1146 314
rect 1076 264 1146 280
rect 1116 180 1146 264
rect 1344 180 1374 372
rect 108 70 138 96
rect 220 70 250 96
rect 332 70 362 96
rect 444 70 474 96
rect 556 70 586 96
rect 668 70 698 96
rect 780 70 810 96
rect 892 70 922 96
rect 1004 70 1034 96
rect 1116 70 1146 96
rect 1344 70 1374 96
<< polycont >>
rect 10 320 44 354
rect 330 388 364 422
rect 468 388 502 422
rect 566 388 600 422
rect 190 230 224 264
rect 330 230 364 264
rect 468 220 502 254
rect 778 388 812 422
rect 916 388 950 422
rect 1014 388 1048 422
rect 638 280 672 314
rect 778 230 812 264
rect 916 220 950 254
rect 1330 388 1364 422
rect 1086 280 1120 314
<< locali >>
rect 158 855 194 872
rect 158 821 159 855
rect 193 821 194 855
rect 158 742 194 821
rect 440 855 476 872
rect 440 821 441 855
rect 475 821 476 855
rect 440 804 476 821
rect 722 855 758 872
rect 722 821 723 855
rect 757 821 758 855
rect 722 810 758 821
rect 624 776 758 810
rect 1004 855 1040 872
rect 1004 821 1005 855
rect 1039 821 1040 855
rect 1004 804 1040 821
rect 1286 855 1322 872
rect 1286 821 1287 855
rect 1321 821 1322 855
rect 624 742 658 776
rect 1004 770 1078 804
rect 1044 742 1078 770
rect 1286 742 1322 821
rect 36 700 98 742
rect 36 666 50 700
rect 84 666 98 700
rect 36 624 98 666
rect 36 590 50 624
rect 84 590 98 624
rect 36 548 98 590
rect 36 514 50 548
rect 84 514 98 548
rect 36 472 98 514
rect 148 700 210 742
rect 148 666 162 700
rect 196 666 210 700
rect 148 624 210 666
rect 148 590 162 624
rect 196 590 210 624
rect 148 548 210 590
rect 148 514 162 548
rect 196 514 210 548
rect 148 472 210 514
rect 260 700 322 742
rect 260 666 274 700
rect 308 666 322 700
rect 260 624 322 666
rect 260 590 274 624
rect 308 590 322 624
rect 260 548 322 590
rect 260 514 274 548
rect 308 514 322 548
rect 260 472 322 514
rect 372 700 434 742
rect 372 666 386 700
rect 420 666 434 700
rect 372 624 434 666
rect 372 590 386 624
rect 420 590 434 624
rect 372 548 434 590
rect 372 514 386 548
rect 420 514 434 548
rect 372 472 434 514
rect 596 700 658 742
rect 596 666 610 700
rect 644 666 658 700
rect 596 624 658 666
rect 596 590 610 624
rect 644 590 658 624
rect 596 548 658 590
rect 596 514 610 548
rect 644 514 658 548
rect 596 472 658 514
rect 708 700 770 742
rect 708 666 722 700
rect 756 666 770 700
rect 708 624 770 666
rect 708 590 722 624
rect 756 590 770 624
rect 708 548 770 590
rect 708 514 722 548
rect 756 514 770 548
rect 708 472 770 514
rect 820 700 882 742
rect 820 666 834 700
rect 868 666 882 700
rect 820 624 882 666
rect 820 590 834 624
rect 868 590 882 624
rect 820 548 882 590
rect 820 514 834 548
rect 868 514 882 548
rect 820 472 882 514
rect 1044 700 1106 742
rect 1044 666 1058 700
rect 1092 666 1106 700
rect 1044 624 1106 666
rect 1044 590 1058 624
rect 1092 590 1106 624
rect 1044 548 1106 590
rect 1044 514 1058 548
rect 1092 514 1106 548
rect 1044 472 1106 514
rect 1156 700 1218 742
rect 1156 666 1170 700
rect 1204 666 1218 700
rect 1156 624 1218 666
rect 1156 590 1170 624
rect 1204 590 1218 624
rect 1156 548 1218 590
rect 1156 514 1170 548
rect 1204 514 1218 548
rect 1156 472 1218 514
rect 1272 700 1334 742
rect 1272 666 1286 700
rect 1320 666 1334 700
rect 1272 624 1334 666
rect 1272 590 1286 624
rect 1320 590 1334 624
rect 1272 548 1334 590
rect 1272 514 1286 548
rect 1320 514 1334 548
rect 1272 472 1334 514
rect 1384 700 1446 742
rect 1384 666 1398 700
rect 1432 666 1446 700
rect 1384 624 1446 666
rect 1384 590 1398 624
rect 1432 590 1446 624
rect 1384 548 1446 590
rect 1384 514 1398 548
rect 1432 514 1446 548
rect 1384 472 1446 514
rect 64 438 98 472
rect 64 404 138 438
rect 10 354 44 370
rect 10 304 44 320
rect 104 270 138 404
rect 64 236 138 270
rect 190 264 224 280
rect 64 180 98 236
rect 190 214 224 230
rect 260 180 294 472
rect 330 422 364 438
rect 330 372 364 388
rect 400 338 434 472
rect 708 438 742 472
rect 468 422 502 438
rect 468 372 502 388
rect 566 422 742 438
rect 600 404 742 422
rect 566 372 600 388
rect 400 314 672 338
rect 400 304 638 314
rect 330 264 364 280
rect 330 214 364 230
rect 400 180 434 304
rect 468 254 502 270
rect 638 264 672 280
rect 468 204 502 220
rect 708 180 742 404
rect 778 422 812 438
rect 778 372 812 388
rect 848 338 882 472
rect 916 422 950 438
rect 916 372 950 388
rect 1014 422 1048 438
rect 1156 422 1190 472
rect 1330 422 1364 438
rect 1048 388 1330 422
rect 1014 372 1048 388
rect 848 314 1120 338
rect 848 304 1086 314
rect 778 264 812 280
rect 778 214 812 230
rect 848 180 882 304
rect 916 254 950 270
rect 1086 264 1120 280
rect 916 204 950 220
rect 1156 180 1190 388
rect 1330 372 1364 388
rect 1412 258 1446 472
rect 1304 224 1446 258
rect 1412 180 1446 224
rect 36 154 98 180
rect 36 120 50 154
rect 84 120 98 154
rect 36 96 98 120
rect 148 154 210 180
rect 148 120 162 154
rect 196 120 210 154
rect 148 96 210 120
rect 260 154 322 180
rect 260 120 274 154
rect 308 120 322 154
rect 260 96 322 120
rect 372 154 434 180
rect 372 120 386 154
rect 420 120 434 154
rect 372 96 434 120
rect 596 154 658 180
rect 596 120 610 154
rect 644 120 658 154
rect 596 96 658 120
rect 708 154 770 180
rect 708 120 722 154
rect 756 120 770 154
rect 708 96 770 120
rect 820 154 882 180
rect 820 120 834 154
rect 868 120 882 154
rect 820 96 882 120
rect 1044 154 1106 180
rect 1044 120 1058 154
rect 1092 120 1106 154
rect 1044 96 1106 120
rect 1156 154 1218 180
rect 1156 120 1170 154
rect 1204 120 1218 154
rect 1156 96 1218 120
rect 1272 154 1334 180
rect 1272 120 1286 154
rect 1320 120 1334 154
rect 1272 96 1334 120
rect 1384 154 1446 180
rect 1384 120 1398 154
rect 1432 120 1446 154
rect 1384 96 1446 120
rect 158 17 194 96
rect 624 62 658 96
rect 1044 68 1078 96
rect 158 -17 159 17
rect 193 -17 194 17
rect 158 -34 194 -17
rect 440 17 476 34
rect 624 28 758 62
rect 440 -17 441 17
rect 475 -17 476 17
rect 440 -34 476 -17
rect 722 17 758 28
rect 722 -17 723 17
rect 757 -17 758 17
rect 722 -34 758 -17
rect 1004 34 1078 68
rect 1004 17 1040 34
rect 1004 -17 1005 17
rect 1039 -17 1040 17
rect 1004 -34 1040 -17
rect 1286 17 1322 96
rect 1286 -17 1287 17
rect 1321 -17 1322 17
rect 1286 -34 1322 -17
<< viali >>
rect 159 821 193 855
rect 441 821 475 855
rect 723 821 757 855
rect 1005 821 1039 855
rect 1287 821 1321 855
rect 10 320 44 354
rect 190 230 224 264
rect 330 388 364 422
rect 468 388 502 422
rect 330 230 364 264
rect 468 220 502 254
rect 778 388 812 422
rect 916 388 950 422
rect 778 230 812 264
rect 916 220 950 254
rect 1270 224 1304 258
rect 50 120 84 154
rect 159 -17 193 17
rect 441 -17 475 17
rect 723 -17 757 17
rect 1005 -17 1039 17
rect 1287 -17 1321 17
<< metal1 >>
rect 0 855 1482 868
rect 0 821 159 855
rect 193 821 441 855
rect 475 821 723 855
rect 757 821 1005 855
rect 1039 821 1287 855
rect 1321 821 1482 855
rect 0 808 1482 821
rect 324 426 370 438
rect 906 434 958 440
rect 26 422 370 426
rect 26 398 330 422
rect 26 370 54 398
rect 324 388 330 398
rect 364 388 370 422
rect 324 372 370 388
rect 458 422 818 434
rect 458 388 468 422
rect 502 406 778 422
rect 502 388 508 406
rect 458 372 508 388
rect 772 388 778 406
rect 812 388 818 422
rect 772 376 818 388
rect 906 376 958 382
rect 0 364 54 370
rect 0 312 2 364
rect 458 338 486 372
rect 0 304 54 312
rect 342 310 486 338
rect 780 348 808 376
rect 780 320 946 348
rect 180 274 234 280
rect 342 276 370 310
rect 180 222 182 274
rect 180 214 234 222
rect 324 264 370 276
rect 324 230 330 264
rect 364 230 370 264
rect 324 218 370 230
rect 460 266 512 272
rect 772 264 818 276
rect 918 266 946 320
rect 1262 266 1314 272
rect 772 246 778 264
rect 512 230 778 246
rect 812 230 818 264
rect 332 166 360 218
rect 512 218 818 230
rect 910 254 956 266
rect 910 220 916 254
rect 950 220 956 254
rect 460 206 512 214
rect 910 208 956 220
rect 1262 208 1314 214
rect 38 154 360 166
rect 38 120 50 154
rect 84 138 360 154
rect 84 120 96 138
rect 38 108 96 120
rect 0 17 1482 30
rect 0 -17 159 17
rect 193 -17 441 17
rect 475 -17 723 17
rect 757 -17 1005 17
rect 1039 -17 1287 17
rect 1321 -17 1482 17
rect 0 -30 1482 -17
<< via1 >>
rect 906 422 958 434
rect 906 388 916 422
rect 916 388 950 422
rect 950 388 958 422
rect 906 382 958 388
rect 2 354 54 364
rect 2 320 10 354
rect 10 320 44 354
rect 44 320 54 354
rect 2 312 54 320
rect 182 264 234 274
rect 182 230 190 264
rect 190 230 224 264
rect 224 230 234 264
rect 182 222 234 230
rect 460 254 512 266
rect 460 220 468 254
rect 468 220 502 254
rect 502 220 512 254
rect 460 214 512 220
rect 1262 258 1314 266
rect 1262 224 1270 258
rect 1270 224 1304 258
rect 1304 224 1314 258
rect 1262 214 1314 224
<< metal2 >>
rect 906 434 958 440
rect 848 394 906 422
rect 2 364 54 370
rect 0 322 2 350
rect 2 304 54 312
rect 26 180 54 304
rect 182 274 234 280
rect 180 232 182 260
rect 182 216 234 222
rect 460 266 512 272
rect 460 208 512 214
rect 484 180 512 208
rect 848 180 876 394
rect 906 376 958 382
rect 1262 266 1314 272
rect 1260 228 1262 256
rect 1262 208 1314 214
rect 26 152 876 180
<< labels >>
rlabel metal1 s 68 112 68 112 4 clkb
rlabel locali s 276 332 276 332 4 net1
rlabel locali s 422 354 422 354 4 net2
rlabel mvpsubdiff s 516 564 516 564 4 net4
rlabel mvpsubdiff s 498 124 498 124 4 net5
rlabel locali s 724 352 724 352 4 net3
rlabel locali s 868 430 868 430 4 net6
rlabel locali s 1178 286 1178 286 4 net7
rlabel mvpsubdiff s 956 552 956 552 4 net8
rlabel mvpsubdiff s 960 136 960 136 4 net9
rlabel metal2 s 0 322 54 350 4 clk
port 1 nsew
rlabel metal1 s 0 808 1482 868 4 vdd
port 2 nsew
rlabel metal1 s 0 -30 1482 30 4 gnd
port 3 nsew
rlabel metal2 s 180 232 234 260 4 D
port 4 nsew
rlabel metal2 s 1260 228 1314 256 4 Q
port 5 nsew
rlabel metal2 s 207 246 207 246 4 D
rlabel metal2 s 1287 242 1287 242 4 Q
rlabel metal2 s 27 336 27 336 4 clk
rlabel metal1 s 741 838 741 838 4 vdd
rlabel metal1 s 741 0 741 0 4 gnd
<< properties >>
string FIXED_BBOX 0 0 1482 838
string GDS_FILE sram_0rw2r1w_2_16_sky130A.gds
string GDS_END 515886
string GDS_START 494506
<< end >>
