magic
tech sky130A
magscale 1 2
timestamp 1644969367
<< checkpaint >>
rect -1260 -1286 1410 1454
<< scnmos >>
rect 60 0 90 168
<< ndiff >>
rect 0 101 60 168
rect 0 67 8 101
rect 42 67 60 101
rect 0 0 60 67
rect 90 0 150 168
<< ndiffc >>
rect 8 67 42 101
<< poly >>
rect 60 168 90 194
rect 60 -26 90 0
<< locali >>
rect 8 101 42 117
rect 8 51 42 67
use contact_8  contact_8_0
timestamp 1644969367
transform 1 0 0 0 1 43
box 0 0 1 1
<< labels >>
rlabel mvvaractor s 75 84 75 84 4 G
rlabel locali s 25 84 25 84 4 S
rlabel mvpsubdiff s 125 84 125 84 4 D
<< properties >>
string FIXED_BBOX -25 -26 175 194
string GDS_FILE sram_0rw2r1w_32_128_sky130A.gds
string GDS_END 3073106
string GDS_START 3072382
<< end >>
