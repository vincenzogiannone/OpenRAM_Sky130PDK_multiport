magic
tech sky130A
magscale 1 2
timestamp 1643678851
<< checkpaint >>
rect -1260 -1294 3491 13614
<< locali >>
rect 0 12303 295 12337
rect 329 12303 1190 12337
rect 1224 12303 2195 12337
rect 2023 11575 2057 11609
rect 0 10763 295 10797
rect 329 10763 1190 10797
rect 1224 10763 2195 10797
rect 2023 9951 2057 9985
rect 0 9223 295 9257
rect 329 9223 1190 9257
rect 1224 9223 2195 9257
rect 2023 8495 2057 8529
rect 0 7683 295 7717
rect 329 7683 1190 7717
rect 1224 7683 2195 7717
rect 2023 6871 2057 6905
rect 0 6143 295 6177
rect 329 6143 1190 6177
rect 1224 6143 2195 6177
rect 2023 5415 2057 5449
rect 0 4603 295 4637
rect 329 4603 1190 4637
rect 1224 4603 2195 4637
rect 2023 3791 2057 3825
rect 0 3063 295 3097
rect 329 3063 1190 3097
rect 1224 3063 2195 3097
rect 2023 2335 2057 2369
rect 0 1523 295 1557
rect 329 1523 1190 1557
rect 1224 1523 2195 1557
rect 2023 711 2057 745
rect 0 -17 295 17
rect 329 -17 1190 17
rect 1224 -17 2195 17
<< viali >>
rect 295 12303 329 12337
rect 1190 12303 1224 12337
rect 1314 12013 1348 12047
rect 1447 11889 1481 11923
rect 1580 11765 1614 11799
rect 295 10763 329 10797
rect 1190 10763 1224 10797
rect 1580 9761 1614 9795
rect 1447 9637 1481 9671
rect 1314 9513 1348 9547
rect 295 9223 329 9257
rect 1190 9223 1224 9257
rect 1314 8933 1348 8967
rect 1447 8809 1481 8843
rect 1580 8685 1614 8719
rect 295 7683 329 7717
rect 1190 7683 1224 7717
rect 1580 6681 1614 6715
rect 1447 6557 1481 6591
rect 1314 6433 1348 6467
rect 295 6143 329 6177
rect 1190 6143 1224 6177
rect 1314 5853 1348 5887
rect 1447 5729 1481 5763
rect 1580 5605 1614 5639
rect 295 4603 329 4637
rect 1190 4603 1224 4637
rect 404 3791 438 3825
rect 536 3791 570 3825
rect 1580 3601 1614 3635
rect 1447 3477 1481 3511
rect 1314 3353 1348 3387
rect 295 3063 329 3097
rect 1190 3063 1224 3097
rect 1314 2773 1348 2807
rect 1447 2649 1481 2683
rect 1580 2525 1614 2559
rect 404 2335 438 2369
rect 536 2335 570 2369
rect 295 1523 329 1557
rect 1190 1523 1224 1557
rect 404 711 438 745
rect 536 711 570 745
rect 1580 521 1614 555
rect 1447 397 1481 431
rect 1314 273 1348 307
rect 295 -17 329 17
rect 1190 -17 1224 17
<< metal1 >>
rect 283 12335 286 12343
rect 257 12305 286 12335
rect 283 12297 286 12305
rect 338 12335 341 12343
rect 1178 12335 1181 12343
rect 338 12305 368 12335
rect 1152 12305 1181 12335
rect 338 12297 341 12305
rect 1178 12297 1181 12305
rect 1233 12335 1236 12343
rect 1233 12305 1263 12335
rect 1233 12297 1236 12305
rect 108 12016 951 12044
rect 1302 12047 1360 12053
rect 1302 12044 1314 12047
rect 1003 12016 1314 12044
rect 1302 12013 1314 12016
rect 1348 12013 1360 12047
rect 1302 12007 1360 12013
rect 176 11892 1019 11920
rect 1435 11923 1493 11929
rect 1435 11920 1447 11923
rect 1071 11892 1447 11920
rect 1435 11889 1447 11892
rect 1481 11889 1493 11923
rect 1435 11883 1493 11889
rect 244 11768 1087 11796
rect 1568 11799 1626 11805
rect 1568 11796 1580 11799
rect 1139 11768 1580 11796
rect 1568 11765 1580 11768
rect 1614 11765 1626 11799
rect 1568 11759 1626 11765
rect 283 10795 286 10803
rect 257 10765 286 10795
rect 283 10757 286 10765
rect 338 10795 341 10803
rect 1178 10795 1181 10803
rect 338 10765 368 10795
rect 1152 10765 1181 10795
rect 338 10757 341 10765
rect 1178 10757 1181 10765
rect 1233 10795 1236 10803
rect 1233 10765 1263 10795
rect 1233 10757 1236 10765
rect 1568 9795 1626 9801
rect 1568 9792 1580 9795
rect 1139 9764 1580 9792
rect 1568 9761 1580 9764
rect 1614 9761 1626 9795
rect 1568 9755 1626 9761
rect 1435 9671 1493 9677
rect 1435 9668 1447 9671
rect 1071 9640 1447 9668
rect 1435 9637 1447 9640
rect 1481 9637 1493 9671
rect 1435 9631 1493 9637
rect 1302 9547 1360 9553
rect 1302 9544 1314 9547
rect 799 9516 1314 9544
rect 1302 9513 1314 9516
rect 1348 9513 1360 9547
rect 1302 9507 1360 9513
rect 283 9255 286 9263
rect 257 9225 286 9255
rect 283 9217 286 9225
rect 338 9255 341 9263
rect 1178 9255 1181 9263
rect 338 9225 368 9255
rect 1152 9225 1181 9255
rect 338 9217 341 9225
rect 1178 9217 1181 9225
rect 1233 9255 1236 9263
rect 1233 9225 1263 9255
rect 1233 9217 1236 9225
rect 1302 8967 1360 8973
rect 1302 8964 1314 8967
rect 1003 8936 1314 8964
rect 1302 8933 1314 8936
rect 1348 8933 1360 8967
rect 1302 8927 1360 8933
rect 1435 8843 1493 8849
rect 1435 8840 1447 8843
rect 867 8812 1447 8840
rect 1435 8809 1447 8812
rect 1481 8809 1493 8843
rect 1435 8803 1493 8809
rect 1568 8719 1626 8725
rect 1568 8716 1580 8719
rect 1139 8688 1580 8716
rect 1568 8685 1580 8688
rect 1614 8685 1626 8719
rect 1568 8679 1626 8685
rect 283 7715 286 7723
rect 257 7685 286 7715
rect 283 7677 286 7685
rect 338 7715 341 7723
rect 1178 7715 1181 7723
rect 338 7685 368 7715
rect 1152 7685 1181 7715
rect 338 7677 341 7685
rect 1178 7677 1181 7685
rect 1233 7715 1236 7723
rect 1233 7685 1263 7715
rect 1233 7677 1236 7685
rect 1568 6715 1626 6721
rect 1568 6712 1580 6715
rect 1139 6684 1580 6712
rect 1568 6681 1580 6684
rect 1614 6681 1626 6715
rect 1568 6675 1626 6681
rect 1435 6591 1493 6597
rect 1435 6588 1447 6591
rect 867 6560 1447 6588
rect 1435 6557 1447 6560
rect 1481 6557 1493 6591
rect 1435 6551 1493 6557
rect 1302 6467 1360 6473
rect 1302 6464 1314 6467
rect 799 6436 1314 6464
rect 1302 6433 1314 6436
rect 1348 6433 1360 6467
rect 1302 6427 1360 6433
rect 283 6175 286 6183
rect 257 6145 286 6175
rect 283 6137 286 6145
rect 338 6175 341 6183
rect 1178 6175 1181 6183
rect 338 6145 368 6175
rect 1152 6145 1181 6175
rect 338 6137 341 6145
rect 1178 6137 1181 6145
rect 1233 6175 1236 6183
rect 1233 6145 1263 6175
rect 1233 6137 1236 6145
rect 1302 5887 1360 5893
rect 1302 5884 1314 5887
rect 1003 5856 1314 5884
rect 1302 5853 1314 5856
rect 1348 5853 1360 5887
rect 1302 5847 1360 5853
rect 1435 5763 1493 5769
rect 1435 5760 1447 5763
rect 1071 5732 1447 5760
rect 1435 5729 1447 5732
rect 1481 5729 1493 5763
rect 1435 5723 1493 5729
rect 1568 5639 1626 5645
rect 1568 5636 1580 5639
rect 935 5608 1580 5636
rect 1568 5605 1580 5608
rect 1614 5605 1626 5639
rect 1568 5599 1626 5605
rect 283 4635 286 4643
rect 257 4605 286 4635
rect 283 4597 286 4605
rect 338 4635 341 4643
rect 1178 4635 1181 4643
rect 338 4605 368 4635
rect 1152 4605 1181 4635
rect 338 4597 341 4605
rect 1178 4597 1181 4605
rect 1233 4635 1236 4643
rect 1233 4605 1263 4635
rect 1233 4597 1236 4605
rect 677 4548 883 4576
rect 392 3825 450 3831
rect 392 3822 404 3825
rect 244 3794 404 3822
rect 392 3791 404 3794
rect 438 3791 450 3825
rect 392 3785 450 3791
rect 524 3825 582 3831
rect 524 3791 536 3825
rect 570 3822 582 3825
rect 677 3822 705 4548
rect 570 3794 705 3822
rect 570 3791 582 3794
rect 524 3785 582 3791
rect 1568 3635 1626 3641
rect 1568 3632 1580 3635
rect 935 3604 1580 3632
rect 1568 3601 1580 3604
rect 1614 3601 1626 3635
rect 1568 3595 1626 3601
rect 1435 3511 1493 3517
rect 1435 3508 1447 3511
rect 1071 3480 1447 3508
rect 1435 3477 1447 3480
rect 1481 3477 1493 3511
rect 1435 3471 1493 3477
rect 1302 3387 1360 3393
rect 1302 3384 1314 3387
rect 799 3356 1314 3384
rect 1302 3353 1314 3356
rect 1348 3353 1360 3387
rect 1302 3347 1360 3353
rect 283 3095 286 3103
rect 257 3065 286 3095
rect 283 3057 286 3065
rect 338 3095 341 3103
rect 1178 3095 1181 3103
rect 338 3065 368 3095
rect 1152 3065 1181 3095
rect 338 3057 341 3065
rect 1178 3057 1181 3065
rect 1233 3095 1236 3103
rect 1233 3065 1263 3095
rect 1233 3057 1236 3065
rect 677 3008 815 3036
rect 392 2369 450 2375
rect 392 2366 404 2369
rect 176 2338 404 2366
rect 392 2335 404 2338
rect 438 2335 450 2369
rect 392 2329 450 2335
rect 524 2369 582 2375
rect 524 2335 536 2369
rect 570 2366 582 2369
rect 677 2366 705 3008
rect 1302 2807 1360 2813
rect 1302 2804 1314 2807
rect 1003 2776 1314 2804
rect 1302 2773 1314 2776
rect 1348 2773 1360 2807
rect 1302 2767 1360 2773
rect 1435 2683 1493 2689
rect 1435 2680 1447 2683
rect 867 2652 1447 2680
rect 1435 2649 1447 2652
rect 1481 2649 1493 2683
rect 1435 2643 1493 2649
rect 1568 2559 1626 2565
rect 1568 2556 1580 2559
rect 935 2528 1580 2556
rect 1568 2525 1580 2528
rect 1614 2525 1626 2559
rect 1568 2519 1626 2525
rect 570 2338 705 2366
rect 570 2335 582 2338
rect 524 2329 582 2335
rect 283 1555 286 1563
rect 257 1525 286 1555
rect 283 1517 286 1525
rect 338 1555 341 1563
rect 1178 1555 1181 1563
rect 338 1525 368 1555
rect 1152 1525 1181 1555
rect 338 1517 341 1525
rect 1178 1517 1181 1525
rect 1233 1555 1236 1563
rect 1233 1525 1263 1555
rect 1233 1517 1236 1525
rect 677 1468 747 1496
rect 392 745 450 751
rect 392 742 404 745
rect 108 714 404 742
rect 392 711 404 714
rect 438 711 450 745
rect 392 705 450 711
rect 524 745 582 751
rect 524 711 536 745
rect 570 742 582 745
rect 677 742 705 1468
rect 570 714 705 742
rect 570 711 582 714
rect 524 705 582 711
rect 1568 555 1626 561
rect 1568 552 1580 555
rect 935 524 1580 552
rect 1568 521 1580 524
rect 1614 521 1626 555
rect 1568 515 1626 521
rect 1435 431 1493 437
rect 1435 428 1447 431
rect 867 400 1447 428
rect 1435 397 1447 400
rect 1481 397 1493 431
rect 1435 391 1493 397
rect 1302 307 1360 313
rect 1302 304 1314 307
rect 799 276 1314 304
rect 1302 273 1314 276
rect 1348 273 1360 307
rect 1302 267 1360 273
rect 283 15 286 23
rect 257 -15 286 15
rect 283 -23 286 -15
rect 338 15 341 23
rect 1178 15 1181 23
rect 338 -15 368 15
rect 1152 -15 1181 15
rect 338 -23 341 -15
rect 1178 -23 1181 -15
rect 1233 15 1236 23
rect 1233 -15 1263 15
rect 1233 -23 1236 -15
<< via1 >>
rect 286 12337 338 12346
rect 286 12303 295 12337
rect 295 12303 329 12337
rect 329 12303 338 12337
rect 1181 12337 1233 12346
rect 286 12294 338 12303
rect 1181 12303 1190 12337
rect 1190 12303 1224 12337
rect 1224 12303 1233 12337
rect 1181 12294 1233 12303
rect 56 12004 108 12056
rect 951 12004 1003 12056
rect 124 11880 176 11932
rect 1019 11880 1071 11932
rect 192 11756 244 11808
rect 1087 11756 1139 11808
rect 286 10797 338 10806
rect 286 10763 295 10797
rect 295 10763 329 10797
rect 329 10763 338 10797
rect 1181 10797 1233 10806
rect 286 10754 338 10763
rect 1181 10763 1190 10797
rect 1190 10763 1224 10797
rect 1224 10763 1233 10797
rect 1181 10754 1233 10763
rect 1087 9752 1139 9804
rect 1019 9628 1071 9680
rect 747 9504 799 9556
rect 286 9257 338 9266
rect 286 9223 295 9257
rect 295 9223 329 9257
rect 329 9223 338 9257
rect 1181 9257 1233 9266
rect 286 9214 338 9223
rect 1181 9223 1190 9257
rect 1190 9223 1224 9257
rect 1224 9223 1233 9257
rect 1181 9214 1233 9223
rect 951 8924 1003 8976
rect 815 8800 867 8852
rect 1087 8676 1139 8728
rect 286 7717 338 7726
rect 286 7683 295 7717
rect 295 7683 329 7717
rect 329 7683 338 7717
rect 1181 7717 1233 7726
rect 286 7674 338 7683
rect 1181 7683 1190 7717
rect 1190 7683 1224 7717
rect 1224 7683 1233 7717
rect 1181 7674 1233 7683
rect 1087 6672 1139 6724
rect 815 6548 867 6600
rect 747 6424 799 6476
rect 286 6177 338 6186
rect 286 6143 295 6177
rect 295 6143 329 6177
rect 329 6143 338 6177
rect 1181 6177 1233 6186
rect 286 6134 338 6143
rect 1181 6143 1190 6177
rect 1190 6143 1224 6177
rect 1224 6143 1233 6177
rect 1181 6134 1233 6143
rect 951 5844 1003 5896
rect 1019 5720 1071 5772
rect 883 5596 935 5648
rect 286 4637 338 4646
rect 286 4603 295 4637
rect 295 4603 329 4637
rect 329 4603 338 4637
rect 1181 4637 1233 4646
rect 286 4594 338 4603
rect 1181 4603 1190 4637
rect 1190 4603 1224 4637
rect 1224 4603 1233 4637
rect 1181 4594 1233 4603
rect 192 3782 244 3834
rect 883 4536 935 4588
rect 883 3592 935 3644
rect 1019 3468 1071 3520
rect 747 3344 799 3396
rect 286 3097 338 3106
rect 286 3063 295 3097
rect 295 3063 329 3097
rect 329 3063 338 3097
rect 1181 3097 1233 3106
rect 286 3054 338 3063
rect 1181 3063 1190 3097
rect 1190 3063 1224 3097
rect 1224 3063 1233 3097
rect 1181 3054 1233 3063
rect 124 2326 176 2378
rect 815 2996 867 3048
rect 951 2764 1003 2816
rect 815 2640 867 2692
rect 883 2516 935 2568
rect 286 1557 338 1566
rect 286 1523 295 1557
rect 295 1523 329 1557
rect 329 1523 338 1557
rect 1181 1557 1233 1566
rect 286 1514 338 1523
rect 1181 1523 1190 1557
rect 1190 1523 1224 1557
rect 1224 1523 1233 1557
rect 1181 1514 1233 1523
rect 56 702 108 754
rect 747 1456 799 1508
rect 883 512 935 564
rect 815 388 867 440
rect 747 264 799 316
rect 286 17 338 26
rect 286 -17 295 17
rect 295 -17 329 17
rect 329 -17 338 17
rect 1181 17 1233 26
rect 286 -26 338 -17
rect 1181 -17 1190 17
rect 1190 -17 1224 17
rect 1224 -17 1233 17
rect 1181 -26 1233 -17
<< metal2 >>
rect 292 12348 332 12354
rect 1187 12348 1227 12354
rect 68 12056 96 12320
rect 68 754 96 12004
rect 136 11932 164 12320
rect 136 2378 164 11880
rect 204 11808 232 12320
rect 292 12286 332 12292
rect 204 3834 232 11756
rect 292 10808 332 10814
rect 292 10746 332 10752
rect 759 9556 787 12320
rect 292 9268 332 9274
rect 292 9206 332 9212
rect 292 7728 332 7734
rect 292 7666 332 7672
rect 759 6476 787 9504
rect 827 8852 855 12320
rect 827 6600 855 8800
rect 292 6188 332 6194
rect 292 6126 332 6132
rect 292 4648 332 4654
rect 292 4586 332 4592
rect 68 68 96 702
rect 136 68 164 2326
rect 204 68 232 3782
rect 759 3396 787 6424
rect 292 3108 332 3114
rect 292 3046 332 3052
rect 292 1568 332 1574
rect 292 1506 332 1512
rect 759 1508 787 3344
rect 827 3048 855 6548
rect 895 5648 923 12320
rect 963 12056 991 12320
rect 963 8976 991 12004
rect 1031 11932 1059 12320
rect 1031 9680 1059 11880
rect 1099 11808 1127 12320
rect 1187 12286 1227 12292
rect 1099 9804 1127 11756
rect 1187 10808 1227 10814
rect 1187 10746 1227 10752
rect 963 5896 991 8924
rect 895 4588 923 5596
rect 895 3644 923 4536
rect 827 2692 855 2996
rect 759 316 787 1456
rect 827 440 855 2640
rect 895 2568 923 3592
rect 963 2816 991 5844
rect 1031 5772 1059 9628
rect 1099 8728 1127 9752
rect 1187 9268 1227 9274
rect 1187 9206 1227 9212
rect 1099 6724 1127 8676
rect 1187 7728 1227 7734
rect 1187 7666 1227 7672
rect 1031 3520 1059 5720
rect 895 564 923 2516
rect 759 68 787 264
rect 827 68 855 388
rect 895 68 923 512
rect 963 68 991 2764
rect 1031 68 1059 3468
rect 1099 68 1127 6672
rect 1187 6188 1227 6194
rect 1187 6126 1227 6132
rect 1187 4648 1227 4654
rect 1187 4586 1227 4592
rect 1187 3108 1227 3114
rect 1187 3046 1227 3052
rect 1187 1568 1227 1574
rect 1187 1506 1227 1512
rect 292 28 332 34
rect 1187 28 1227 34
rect 292 -34 332 -28
rect 1187 -34 1227 -28
<< via2 >>
rect 284 12346 340 12348
rect 284 12294 286 12346
rect 286 12294 338 12346
rect 338 12294 340 12346
rect 1179 12346 1235 12348
rect 284 12292 340 12294
rect 284 10806 340 10808
rect 284 10754 286 10806
rect 286 10754 338 10806
rect 338 10754 340 10806
rect 284 10752 340 10754
rect 284 9266 340 9268
rect 284 9214 286 9266
rect 286 9214 338 9266
rect 338 9214 340 9266
rect 284 9212 340 9214
rect 284 7726 340 7728
rect 284 7674 286 7726
rect 286 7674 338 7726
rect 338 7674 340 7726
rect 284 7672 340 7674
rect 284 6186 340 6188
rect 284 6134 286 6186
rect 286 6134 338 6186
rect 338 6134 340 6186
rect 284 6132 340 6134
rect 284 4646 340 4648
rect 284 4594 286 4646
rect 286 4594 338 4646
rect 338 4594 340 4646
rect 284 4592 340 4594
rect 284 3106 340 3108
rect 284 3054 286 3106
rect 286 3054 338 3106
rect 338 3054 340 3106
rect 284 3052 340 3054
rect 284 1566 340 1568
rect 284 1514 286 1566
rect 286 1514 338 1566
rect 338 1514 340 1566
rect 284 1512 340 1514
rect 1179 12294 1181 12346
rect 1181 12294 1233 12346
rect 1233 12294 1235 12346
rect 1179 12292 1235 12294
rect 1179 10806 1235 10808
rect 1179 10754 1181 10806
rect 1181 10754 1233 10806
rect 1233 10754 1235 10806
rect 1179 10752 1235 10754
rect 1179 9266 1235 9268
rect 1179 9214 1181 9266
rect 1181 9214 1233 9266
rect 1233 9214 1235 9266
rect 1179 9212 1235 9214
rect 1179 7726 1235 7728
rect 1179 7674 1181 7726
rect 1181 7674 1233 7726
rect 1233 7674 1235 7726
rect 1179 7672 1235 7674
rect 1179 6186 1235 6188
rect 1179 6134 1181 6186
rect 1181 6134 1233 6186
rect 1233 6134 1235 6186
rect 1179 6132 1235 6134
rect 1179 4646 1235 4648
rect 1179 4594 1181 4646
rect 1181 4594 1233 4646
rect 1233 4594 1235 4646
rect 1179 4592 1235 4594
rect 1179 3106 1235 3108
rect 1179 3054 1181 3106
rect 1181 3054 1233 3106
rect 1233 3054 1235 3106
rect 1179 3052 1235 3054
rect 1179 1566 1235 1568
rect 1179 1514 1181 1566
rect 1181 1514 1233 1566
rect 1233 1514 1235 1566
rect 1179 1512 1235 1514
rect 284 26 340 28
rect 284 -26 286 26
rect 286 -26 338 26
rect 338 -26 340 26
rect 284 -28 340 -26
rect 1179 26 1235 28
rect 1179 -26 1181 26
rect 1181 -26 1233 26
rect 1233 -26 1235 26
rect 1179 -28 1235 -26
<< metal3 >>
rect 246 12348 378 12353
rect 246 12292 284 12348
rect 340 12292 378 12348
rect 246 12287 378 12292
rect 1141 12348 1273 12353
rect 1141 12292 1179 12348
rect 1235 12292 1273 12348
rect 1141 12287 1273 12292
rect 246 10808 378 10813
rect 246 10752 284 10808
rect 340 10752 378 10808
rect 246 10747 378 10752
rect 1141 10808 1273 10813
rect 1141 10752 1179 10808
rect 1235 10752 1273 10808
rect 1141 10747 1273 10752
rect 246 9268 378 9273
rect 246 9212 284 9268
rect 340 9212 378 9268
rect 246 9207 378 9212
rect 1141 9268 1273 9273
rect 1141 9212 1179 9268
rect 1235 9212 1273 9268
rect 1141 9207 1273 9212
rect 246 7728 378 7733
rect 246 7672 284 7728
rect 340 7672 378 7728
rect 246 7667 378 7672
rect 1141 7728 1273 7733
rect 1141 7672 1179 7728
rect 1235 7672 1273 7728
rect 1141 7667 1273 7672
rect 246 6188 378 6193
rect 246 6132 284 6188
rect 340 6132 378 6188
rect 246 6127 378 6132
rect 1141 6188 1273 6193
rect 1141 6132 1179 6188
rect 1235 6132 1273 6188
rect 1141 6127 1273 6132
rect 246 4648 378 4653
rect 246 4592 284 4648
rect 340 4592 378 4648
rect 246 4587 378 4592
rect 1141 4648 1273 4653
rect 1141 4592 1179 4648
rect 1235 4592 1273 4648
rect 1141 4587 1273 4592
rect 246 3108 378 3113
rect 246 3052 284 3108
rect 340 3052 378 3108
rect 246 3047 378 3052
rect 1141 3108 1273 3113
rect 1141 3052 1179 3108
rect 1235 3052 1273 3108
rect 1141 3047 1273 3052
rect 246 1568 378 1573
rect 246 1512 284 1568
rect 340 1512 378 1568
rect 246 1507 378 1512
rect 1141 1568 1273 1573
rect 1141 1512 1179 1568
rect 1235 1512 1273 1568
rect 1141 1507 1273 1512
rect 246 28 378 33
rect 246 -28 284 28
rect 340 -28 378 28
rect 246 -33 378 -28
rect 1141 28 1273 33
rect 1141 -28 1179 28
rect 1235 -28 1273 28
rect 1141 -33 1273 -28
use contact_18  contact_18_0
timestamp 1643678851
transform 1 0 1141 0 1 12287
box 0 0 1 1
use contact_17  contact_17_0
timestamp 1643678851
transform 1 0 1192 0 1 12305
box 0 0 1 1
use contact_13  contact_13_0
timestamp 1643678851
transform 1 0 1178 0 1 12297
box 0 0 1 1
use contact_18  contact_18_1
timestamp 1643678851
transform 1 0 246 0 1 12287
box 0 0 1 1
use contact_17  contact_17_1
timestamp 1643678851
transform 1 0 297 0 1 12305
box 0 0 1 1
use contact_13  contact_13_1
timestamp 1643678851
transform 1 0 283 0 1 12297
box 0 0 1 1
use contact_18  contact_18_2
timestamp 1643678851
transform 1 0 1141 0 1 10747
box 0 0 1 1
use contact_17  contact_17_2
timestamp 1643678851
transform 1 0 1192 0 1 10765
box 0 0 1 1
use contact_13  contact_13_2
timestamp 1643678851
transform 1 0 1178 0 1 10757
box 0 0 1 1
use contact_18  contact_18_3
timestamp 1643678851
transform 1 0 246 0 1 10747
box 0 0 1 1
use contact_17  contact_17_3
timestamp 1643678851
transform 1 0 297 0 1 10765
box 0 0 1 1
use contact_13  contact_13_3
timestamp 1643678851
transform 1 0 283 0 1 10757
box 0 0 1 1
use contact_18  contact_18_4
timestamp 1643678851
transform 1 0 1141 0 1 9207
box 0 0 1 1
use contact_17  contact_17_4
timestamp 1643678851
transform 1 0 1192 0 1 9225
box 0 0 1 1
use contact_13  contact_13_4
timestamp 1643678851
transform 1 0 1178 0 1 9217
box 0 0 1 1
use contact_18  contact_18_5
timestamp 1643678851
transform 1 0 246 0 1 9207
box 0 0 1 1
use contact_17  contact_17_5
timestamp 1643678851
transform 1 0 297 0 1 9225
box 0 0 1 1
use contact_13  contact_13_5
timestamp 1643678851
transform 1 0 283 0 1 9217
box 0 0 1 1
use contact_18  contact_18_6
timestamp 1643678851
transform 1 0 1141 0 1 10747
box 0 0 1 1
use contact_17  contact_17_6
timestamp 1643678851
transform 1 0 1192 0 1 10765
box 0 0 1 1
use contact_13  contact_13_6
timestamp 1643678851
transform 1 0 1178 0 1 10757
box 0 0 1 1
use contact_18  contact_18_7
timestamp 1643678851
transform 1 0 246 0 1 10747
box 0 0 1 1
use contact_17  contact_17_7
timestamp 1643678851
transform 1 0 297 0 1 10765
box 0 0 1 1
use contact_13  contact_13_7
timestamp 1643678851
transform 1 0 283 0 1 10757
box 0 0 1 1
use contact_18  contact_18_8
timestamp 1643678851
transform 1 0 1141 0 1 9207
box 0 0 1 1
use contact_17  contact_17_8
timestamp 1643678851
transform 1 0 1192 0 1 9225
box 0 0 1 1
use contact_13  contact_13_8
timestamp 1643678851
transform 1 0 1178 0 1 9217
box 0 0 1 1
use contact_18  contact_18_9
timestamp 1643678851
transform 1 0 246 0 1 9207
box 0 0 1 1
use contact_17  contact_17_9
timestamp 1643678851
transform 1 0 297 0 1 9225
box 0 0 1 1
use contact_13  contact_13_9
timestamp 1643678851
transform 1 0 283 0 1 9217
box 0 0 1 1
use contact_18  contact_18_10
timestamp 1643678851
transform 1 0 1141 0 1 7667
box 0 0 1 1
use contact_17  contact_17_10
timestamp 1643678851
transform 1 0 1192 0 1 7685
box 0 0 1 1
use contact_13  contact_13_10
timestamp 1643678851
transform 1 0 1178 0 1 7677
box 0 0 1 1
use contact_18  contact_18_11
timestamp 1643678851
transform 1 0 246 0 1 7667
box 0 0 1 1
use contact_17  contact_17_11
timestamp 1643678851
transform 1 0 297 0 1 7685
box 0 0 1 1
use contact_13  contact_13_11
timestamp 1643678851
transform 1 0 283 0 1 7677
box 0 0 1 1
use contact_18  contact_18_12
timestamp 1643678851
transform 1 0 1141 0 1 6127
box 0 0 1 1
use contact_17  contact_17_12
timestamp 1643678851
transform 1 0 1192 0 1 6145
box 0 0 1 1
use contact_13  contact_13_12
timestamp 1643678851
transform 1 0 1178 0 1 6137
box 0 0 1 1
use contact_18  contact_18_13
timestamp 1643678851
transform 1 0 246 0 1 6127
box 0 0 1 1
use contact_17  contact_17_13
timestamp 1643678851
transform 1 0 297 0 1 6145
box 0 0 1 1
use contact_13  contact_13_13
timestamp 1643678851
transform 1 0 283 0 1 6137
box 0 0 1 1
use contact_18  contact_18_14
timestamp 1643678851
transform 1 0 1141 0 1 7667
box 0 0 1 1
use contact_17  contact_17_14
timestamp 1643678851
transform 1 0 1192 0 1 7685
box 0 0 1 1
use contact_13  contact_13_14
timestamp 1643678851
transform 1 0 1178 0 1 7677
box 0 0 1 1
use contact_18  contact_18_15
timestamp 1643678851
transform 1 0 246 0 1 7667
box 0 0 1 1
use contact_17  contact_17_15
timestamp 1643678851
transform 1 0 297 0 1 7685
box 0 0 1 1
use contact_13  contact_13_15
timestamp 1643678851
transform 1 0 283 0 1 7677
box 0 0 1 1
use contact_18  contact_18_16
timestamp 1643678851
transform 1 0 1141 0 1 6127
box 0 0 1 1
use contact_17  contact_17_16
timestamp 1643678851
transform 1 0 1192 0 1 6145
box 0 0 1 1
use contact_13  contact_13_16
timestamp 1643678851
transform 1 0 1178 0 1 6137
box 0 0 1 1
use contact_18  contact_18_17
timestamp 1643678851
transform 1 0 246 0 1 6127
box 0 0 1 1
use contact_17  contact_17_17
timestamp 1643678851
transform 1 0 297 0 1 6145
box 0 0 1 1
use contact_13  contact_13_17
timestamp 1643678851
transform 1 0 283 0 1 6137
box 0 0 1 1
use contact_18  contact_18_18
timestamp 1643678851
transform 1 0 1141 0 1 4587
box 0 0 1 1
use contact_17  contact_17_18
timestamp 1643678851
transform 1 0 1192 0 1 4605
box 0 0 1 1
use contact_13  contact_13_18
timestamp 1643678851
transform 1 0 1178 0 1 4597
box 0 0 1 1
use contact_18  contact_18_19
timestamp 1643678851
transform 1 0 246 0 1 4587
box 0 0 1 1
use contact_17  contact_17_19
timestamp 1643678851
transform 1 0 297 0 1 4605
box 0 0 1 1
use contact_13  contact_13_19
timestamp 1643678851
transform 1 0 283 0 1 4597
box 0 0 1 1
use contact_18  contact_18_20
timestamp 1643678851
transform 1 0 1141 0 1 3047
box 0 0 1 1
use contact_17  contact_17_20
timestamp 1643678851
transform 1 0 1192 0 1 3065
box 0 0 1 1
use contact_13  contact_13_20
timestamp 1643678851
transform 1 0 1178 0 1 3057
box 0 0 1 1
use contact_18  contact_18_21
timestamp 1643678851
transform 1 0 246 0 1 3047
box 0 0 1 1
use contact_17  contact_17_21
timestamp 1643678851
transform 1 0 297 0 1 3065
box 0 0 1 1
use contact_13  contact_13_21
timestamp 1643678851
transform 1 0 283 0 1 3057
box 0 0 1 1
use contact_18  contact_18_22
timestamp 1643678851
transform 1 0 1141 0 1 4587
box 0 0 1 1
use contact_17  contact_17_22
timestamp 1643678851
transform 1 0 1192 0 1 4605
box 0 0 1 1
use contact_13  contact_13_22
timestamp 1643678851
transform 1 0 1178 0 1 4597
box 0 0 1 1
use contact_18  contact_18_23
timestamp 1643678851
transform 1 0 246 0 1 4587
box 0 0 1 1
use contact_17  contact_17_23
timestamp 1643678851
transform 1 0 297 0 1 4605
box 0 0 1 1
use contact_13  contact_13_23
timestamp 1643678851
transform 1 0 283 0 1 4597
box 0 0 1 1
use contact_18  contact_18_24
timestamp 1643678851
transform 1 0 1141 0 1 3047
box 0 0 1 1
use contact_17  contact_17_24
timestamp 1643678851
transform 1 0 1192 0 1 3065
box 0 0 1 1
use contact_13  contact_13_24
timestamp 1643678851
transform 1 0 1178 0 1 3057
box 0 0 1 1
use contact_18  contact_18_25
timestamp 1643678851
transform 1 0 246 0 1 3047
box 0 0 1 1
use contact_17  contact_17_25
timestamp 1643678851
transform 1 0 297 0 1 3065
box 0 0 1 1
use contact_13  contact_13_25
timestamp 1643678851
transform 1 0 283 0 1 3057
box 0 0 1 1
use contact_18  contact_18_26
timestamp 1643678851
transform 1 0 1141 0 1 1507
box 0 0 1 1
use contact_17  contact_17_26
timestamp 1643678851
transform 1 0 1192 0 1 1525
box 0 0 1 1
use contact_13  contact_13_26
timestamp 1643678851
transform 1 0 1178 0 1 1517
box 0 0 1 1
use contact_18  contact_18_27
timestamp 1643678851
transform 1 0 246 0 1 1507
box 0 0 1 1
use contact_17  contact_17_27
timestamp 1643678851
transform 1 0 297 0 1 1525
box 0 0 1 1
use contact_13  contact_13_27
timestamp 1643678851
transform 1 0 283 0 1 1517
box 0 0 1 1
use contact_18  contact_18_28
timestamp 1643678851
transform 1 0 1141 0 1 -33
box 0 0 1 1
use contact_17  contact_17_28
timestamp 1643678851
transform 1 0 1192 0 1 -15
box 0 0 1 1
use contact_13  contact_13_28
timestamp 1643678851
transform 1 0 1178 0 1 -23
box 0 0 1 1
use contact_18  contact_18_29
timestamp 1643678851
transform 1 0 246 0 1 -33
box 0 0 1 1
use contact_17  contact_17_29
timestamp 1643678851
transform 1 0 297 0 1 -15
box 0 0 1 1
use contact_13  contact_13_29
timestamp 1643678851
transform 1 0 283 0 1 -23
box 0 0 1 1
use contact_18  contact_18_30
timestamp 1643678851
transform 1 0 1141 0 1 1507
box 0 0 1 1
use contact_17  contact_17_30
timestamp 1643678851
transform 1 0 1192 0 1 1525
box 0 0 1 1
use contact_13  contact_13_30
timestamp 1643678851
transform 1 0 1178 0 1 1517
box 0 0 1 1
use contact_18  contact_18_31
timestamp 1643678851
transform 1 0 246 0 1 1507
box 0 0 1 1
use contact_17  contact_17_31
timestamp 1643678851
transform 1 0 297 0 1 1525
box 0 0 1 1
use contact_13  contact_13_31
timestamp 1643678851
transform 1 0 283 0 1 1517
box 0 0 1 1
use contact_17  contact_17_32
timestamp 1643678851
transform 1 0 1098 0 1 11767
box 0 0 1 1
use contact_17  contact_17_33
timestamp 1643678851
transform 1 0 203 0 1 11767
box 0 0 1 1
use contact_17  contact_17_34
timestamp 1643678851
transform 1 0 1030 0 1 11891
box 0 0 1 1
use contact_17  contact_17_35
timestamp 1643678851
transform 1 0 135 0 1 11891
box 0 0 1 1
use contact_17  contact_17_36
timestamp 1643678851
transform 1 0 962 0 1 12015
box 0 0 1 1
use contact_17  contact_17_37
timestamp 1643678851
transform 1 0 67 0 1 12015
box 0 0 1 1
use contact_14  contact_14_0
timestamp 1643678851
transform 1 0 894 0 1 4547
box 0 0 1 1
use contact_13  contact_13_32
timestamp 1643678851
transform 1 0 524 0 1 3785
box 0 0 1 1
use contact_14  contact_14_1
timestamp 1643678851
transform 1 0 826 0 1 3007
box 0 0 1 1
use contact_13  contact_13_33
timestamp 1643678851
transform 1 0 524 0 1 2329
box 0 0 1 1
use contact_14  contact_14_2
timestamp 1643678851
transform 1 0 758 0 1 1467
box 0 0 1 1
use contact_13  contact_13_34
timestamp 1643678851
transform 1 0 524 0 1 705
box 0 0 1 1
use contact_15  contact_15_0
timestamp 1643678851
transform 1 0 1568 0 1 11759
box 0 0 1 1
use contact_14  contact_14_3
timestamp 1643678851
transform 1 0 1098 0 1 11767
box 0 0 1 1
use contact_15  contact_15_1
timestamp 1643678851
transform 1 0 1435 0 1 11883
box 0 0 1 1
use contact_14  contact_14_4
timestamp 1643678851
transform 1 0 1030 0 1 11891
box 0 0 1 1
use contact_13  contact_13_35
timestamp 1643678851
transform 1 0 1302 0 1 12007
box 0 0 1 1
use contact_14  contact_14_5
timestamp 1643678851
transform 1 0 962 0 1 12015
box 0 0 1 1
use contact_15  contact_15_2
timestamp 1643678851
transform 1 0 1568 0 1 9755
box 0 0 1 1
use contact_14  contact_14_6
timestamp 1643678851
transform 1 0 1098 0 1 9763
box 0 0 1 1
use contact_15  contact_15_3
timestamp 1643678851
transform 1 0 1435 0 1 9631
box 0 0 1 1
use contact_14  contact_14_7
timestamp 1643678851
transform 1 0 1030 0 1 9639
box 0 0 1 1
use contact_13  contact_13_36
timestamp 1643678851
transform 1 0 1302 0 1 9507
box 0 0 1 1
use contact_14  contact_14_8
timestamp 1643678851
transform 1 0 758 0 1 9515
box 0 0 1 1
use contact_15  contact_15_4
timestamp 1643678851
transform 1 0 1568 0 1 8679
box 0 0 1 1
use contact_14  contact_14_9
timestamp 1643678851
transform 1 0 1098 0 1 8687
box 0 0 1 1
use contact_15  contact_15_5
timestamp 1643678851
transform 1 0 1435 0 1 8803
box 0 0 1 1
use contact_14  contact_14_10
timestamp 1643678851
transform 1 0 826 0 1 8811
box 0 0 1 1
use contact_13  contact_13_37
timestamp 1643678851
transform 1 0 1302 0 1 8927
box 0 0 1 1
use contact_14  contact_14_11
timestamp 1643678851
transform 1 0 962 0 1 8935
box 0 0 1 1
use contact_15  contact_15_6
timestamp 1643678851
transform 1 0 1568 0 1 6675
box 0 0 1 1
use contact_14  contact_14_12
timestamp 1643678851
transform 1 0 1098 0 1 6683
box 0 0 1 1
use contact_15  contact_15_7
timestamp 1643678851
transform 1 0 1435 0 1 6551
box 0 0 1 1
use contact_14  contact_14_13
timestamp 1643678851
transform 1 0 826 0 1 6559
box 0 0 1 1
use contact_13  contact_13_38
timestamp 1643678851
transform 1 0 1302 0 1 6427
box 0 0 1 1
use contact_14  contact_14_14
timestamp 1643678851
transform 1 0 758 0 1 6435
box 0 0 1 1
use contact_15  contact_15_8
timestamp 1643678851
transform 1 0 1568 0 1 5599
box 0 0 1 1
use contact_14  contact_14_15
timestamp 1643678851
transform 1 0 894 0 1 5607
box 0 0 1 1
use contact_15  contact_15_9
timestamp 1643678851
transform 1 0 1435 0 1 5723
box 0 0 1 1
use contact_14  contact_14_16
timestamp 1643678851
transform 1 0 1030 0 1 5731
box 0 0 1 1
use contact_13  contact_13_39
timestamp 1643678851
transform 1 0 1302 0 1 5847
box 0 0 1 1
use contact_14  contact_14_17
timestamp 1643678851
transform 1 0 962 0 1 5855
box 0 0 1 1
use contact_15  contact_15_10
timestamp 1643678851
transform 1 0 1568 0 1 3595
box 0 0 1 1
use contact_14  contact_14_18
timestamp 1643678851
transform 1 0 894 0 1 3603
box 0 0 1 1
use contact_15  contact_15_11
timestamp 1643678851
transform 1 0 1435 0 1 3471
box 0 0 1 1
use contact_14  contact_14_19
timestamp 1643678851
transform 1 0 1030 0 1 3479
box 0 0 1 1
use contact_13  contact_13_40
timestamp 1643678851
transform 1 0 1302 0 1 3347
box 0 0 1 1
use contact_14  contact_14_20
timestamp 1643678851
transform 1 0 758 0 1 3355
box 0 0 1 1
use contact_15  contact_15_12
timestamp 1643678851
transform 1 0 1568 0 1 2519
box 0 0 1 1
use contact_14  contact_14_21
timestamp 1643678851
transform 1 0 894 0 1 2527
box 0 0 1 1
use contact_15  contact_15_13
timestamp 1643678851
transform 1 0 1435 0 1 2643
box 0 0 1 1
use contact_14  contact_14_22
timestamp 1643678851
transform 1 0 826 0 1 2651
box 0 0 1 1
use contact_13  contact_13_41
timestamp 1643678851
transform 1 0 1302 0 1 2767
box 0 0 1 1
use contact_14  contact_14_23
timestamp 1643678851
transform 1 0 962 0 1 2775
box 0 0 1 1
use contact_15  contact_15_14
timestamp 1643678851
transform 1 0 1568 0 1 515
box 0 0 1 1
use contact_14  contact_14_24
timestamp 1643678851
transform 1 0 894 0 1 523
box 0 0 1 1
use contact_15  contact_15_15
timestamp 1643678851
transform 1 0 1435 0 1 391
box 0 0 1 1
use contact_14  contact_14_25
timestamp 1643678851
transform 1 0 826 0 1 399
box 0 0 1 1
use contact_13  contact_13_42
timestamp 1643678851
transform 1 0 1302 0 1 267
box 0 0 1 1
use contact_14  contact_14_26
timestamp 1643678851
transform 1 0 758 0 1 275
box 0 0 1 1
use contact_14  contact_14_27
timestamp 1643678851
transform 1 0 203 0 1 3793
box 0 0 1 1
use contact_13  contact_13_43
timestamp 1643678851
transform 1 0 392 0 1 3785
box 0 0 1 1
use contact_14  contact_14_28
timestamp 1643678851
transform 1 0 135 0 1 2337
box 0 0 1 1
use contact_13  contact_13_44
timestamp 1643678851
transform 1 0 392 0 1 2329
box 0 0 1 1
use contact_14  contact_14_29
timestamp 1643678851
transform 1 0 67 0 1 713
box 0 0 1 1
use contact_13  contact_13_45
timestamp 1643678851
transform 1 0 392 0 1 705
box 0 0 1 1
use and3_dec  and3_dec_0
timestamp 1643678851
transform 1 0 1235 0 -1 12320
box -36 -17 996 1597
use and3_dec  and3_dec_1
timestamp 1643678851
transform 1 0 1235 0 1 9240
box -36 -17 996 1597
use and3_dec  and3_dec_2
timestamp 1643678851
transform 1 0 1235 0 -1 9240
box -36 -17 996 1597
use and3_dec  and3_dec_3
timestamp 1643678851
transform 1 0 1235 0 1 6160
box -36 -17 996 1597
use and3_dec  and3_dec_4
timestamp 1643678851
transform 1 0 1235 0 -1 6160
box -36 -17 996 1597
use and3_dec  and3_dec_5
timestamp 1643678851
transform 1 0 1235 0 1 3080
box -36 -17 996 1597
use and3_dec  and3_dec_6
timestamp 1643678851
transform 1 0 1235 0 -1 3080
box -36 -17 996 1597
use and3_dec  and3_dec_7
timestamp 1643678851
transform 1 0 1235 0 1 0
box -36 -17 996 1597
use pinv  pinv_0
timestamp 1643678851
transform 1 0 340 0 1 3080
box -36 -17 387 1597
use pinv  pinv_1
timestamp 1643678851
transform 1 0 340 0 -1 3080
box -36 -17 387 1597
use pinv  pinv_2
timestamp 1643678851
transform 1 0 340 0 1 0
box -36 -17 387 1597
<< labels >>
rlabel metal2 s 67 713 97 743 4 in_0
rlabel metal2 s 135 2337 165 2367 4 in_1
rlabel metal2 s 203 3793 233 3823 4 in_2
rlabel locali s 2040 728 2040 728 4 out_0
rlabel locali s 2040 2352 2040 2352 4 out_1
rlabel locali s 2040 3808 2040 3808 4 out_2
rlabel locali s 2040 5432 2040 5432 4 out_3
rlabel locali s 2040 6888 2040 6888 4 out_4
rlabel locali s 2040 8512 2040 8512 4 out_5
rlabel locali s 2040 9968 2040 9968 4 out_6
rlabel locali s 2040 11592 2040 11592 4 out_7
rlabel metal3 s 246 4587 378 4653 4 vdd
rlabel metal3 s 246 7667 378 7733 4 vdd
rlabel metal3 s 246 1507 378 1573 4 vdd
rlabel metal3 s 1141 4587 1273 4653 4 vdd
rlabel metal3 s 1141 10747 1273 10813 4 vdd
rlabel metal3 s 246 10747 378 10813 4 vdd
rlabel metal3 s 312 10780 312 10780 4 vdd
rlabel metal3 s 1141 1507 1273 1573 4 vdd
rlabel metal3 s 1207 10780 1207 10780 4 vdd
rlabel metal3 s 1141 7667 1273 7733 4 vdd
rlabel metal3 s 1141 -33 1273 33 4 gnd
rlabel metal3 s 1141 3047 1273 3113 4 gnd
rlabel metal3 s 1141 9207 1273 9273 4 gnd
rlabel metal3 s 246 -33 378 33 4 gnd
rlabel metal3 s 246 12287 378 12353 4 gnd
rlabel metal3 s 246 9207 378 9273 4 gnd
rlabel metal3 s 246 3047 378 3113 4 gnd
rlabel metal3 s 1141 12287 1273 12353 4 gnd
rlabel metal3 s 1141 6127 1273 6193 4 gnd
rlabel metal3 s 246 6127 378 6193 4 gnd
<< properties >>
string FIXED_BBOX 1141 -33 1273 0
string GDS_FILE sram_0rw2r1w_16_128_sky130A.gds
string GDS_END 1878204
string GDS_START 1857340
<< end >>
