magic
tech sky130A
magscale 1 2
timestamp 1644951705
<< checkpaint >>
rect -1296 -1277 9660 2155
<< nwell >>
rect -36 402 8400 895
<< locali >>
rect 0 821 8364 855
rect 48 344 114 410
rect 196 360 449 394
rect 564 360 817 394
rect 936 360 1293 394
rect 1609 354 2093 388
rect 2843 352 3865 386
rect 6019 352 6053 386
rect 0 -17 8364 17
use pinv_10  pinv_10_0
timestamp 1644951705
transform 1 0 3784 0 1 0
box -36 -17 4616 895
use pinv_9  pinv_9_0
timestamp 1644951705
transform 1 0 2012 0 1 0
box -36 -17 1808 895
use pinv_8  pinv_8_0
timestamp 1644951705
transform 1 0 1212 0 1 0
box -36 -17 836 895
use pinv_7  pinv_7_0
timestamp 1644951705
transform 1 0 736 0 1 0
box -36 -17 512 895
use pinv_0  pinv_0_0
timestamp 1644951705
transform 1 0 368 0 1 0
box -36 -17 404 895
use pinv_0  pinv_0_1
timestamp 1644951705
transform 1 0 0 0 1 0
box -36 -17 404 895
<< labels >>
rlabel locali s 6036 369 6036 369 4 Z
rlabel locali s 81 377 81 377 4 A
rlabel locali s 4182 0 4182 0 4 gnd
rlabel locali s 4182 838 4182 838 4 vdd
<< properties >>
string FIXED_BBOX 0 0 8364 838
string GDS_FILE sram_0rw2r1w_16_128_sky130A.gds
string GDS_END 1982222
string GDS_START 1980620
<< end >>
