magic
tech sky130A
magscale 1 2
timestamp 1643593061
<< checkpaint >>
rect -1260 -1260 1261 1261
<< properties >>
string GDS_FILE sram_0rw2r1w_2_16_sky130A.gds
string GDS_END 407504
string GDS_START 407180
<< end >>
