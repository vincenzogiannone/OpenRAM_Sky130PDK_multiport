magic
tech sky130A
timestamp 1642458316
<< nwell >>
rect 0 619 389 808
<< nmos >>
rect 312 532 327 574
rect 60 422 75 506
rect 186 391 201 475
rect 312 391 327 475
rect 60 168 75 252
rect 186 168 201 252
rect 312 168 327 252
rect 60 48 75 90
rect 186 48 201 90
<< pmos >>
rect 60 637 75 721
rect 186 637 201 721
rect 312 637 327 721
<< ndiff >>
rect 270 561 312 574
rect 270 544 277 561
rect 294 544 312 561
rect 270 532 312 544
rect 327 561 369 574
rect 327 544 345 561
rect 362 544 369 561
rect 327 532 369 544
rect 18 490 60 506
rect 18 473 25 490
rect 42 473 60 490
rect 18 456 60 473
rect 18 439 25 456
rect 42 439 60 456
rect 18 422 60 439
rect 75 490 117 506
rect 75 473 93 490
rect 110 473 117 490
rect 75 456 117 473
rect 75 439 93 456
rect 110 439 117 456
rect 75 422 117 439
rect 144 459 186 475
rect 144 442 151 459
rect 168 442 186 459
rect 144 425 186 442
rect 144 408 151 425
rect 168 408 186 425
rect 144 391 186 408
rect 201 459 243 475
rect 201 442 219 459
rect 236 442 243 459
rect 201 425 243 442
rect 201 408 219 425
rect 236 408 243 425
rect 201 391 243 408
rect 270 459 312 475
rect 270 442 277 459
rect 294 442 312 459
rect 270 425 312 442
rect 270 408 277 425
rect 294 408 312 425
rect 270 391 312 408
rect 327 459 369 475
rect 327 442 345 459
rect 362 442 369 459
rect 327 425 369 442
rect 327 408 345 425
rect 362 408 369 425
rect 327 391 369 408
rect 18 236 60 252
rect 18 219 25 236
rect 42 219 60 236
rect 18 202 60 219
rect 18 185 25 202
rect 42 185 60 202
rect 18 168 60 185
rect 75 236 117 252
rect 75 219 93 236
rect 110 219 117 236
rect 75 202 117 219
rect 75 185 93 202
rect 110 185 117 202
rect 75 168 117 185
rect 144 236 186 252
rect 144 219 151 236
rect 168 219 186 236
rect 144 202 186 219
rect 144 185 151 202
rect 168 185 186 202
rect 144 168 186 185
rect 201 236 243 252
rect 201 219 219 236
rect 236 219 243 236
rect 201 202 243 219
rect 201 185 219 202
rect 236 185 243 202
rect 201 168 243 185
rect 270 236 312 252
rect 270 219 277 236
rect 294 219 312 236
rect 270 202 312 219
rect 270 185 277 202
rect 294 185 312 202
rect 270 168 312 185
rect 327 236 369 252
rect 327 219 345 236
rect 362 219 369 236
rect 327 202 369 219
rect 327 185 345 202
rect 362 185 369 202
rect 327 168 369 185
rect 18 77 60 90
rect 18 60 25 77
rect 42 60 60 77
rect 18 48 60 60
rect 75 77 117 90
rect 75 60 93 77
rect 110 60 117 77
rect 75 48 117 60
rect 144 77 186 90
rect 144 60 151 77
rect 168 60 186 77
rect 144 48 186 60
rect 201 77 243 90
rect 201 60 219 77
rect 236 60 243 77
rect 201 48 243 60
<< pdiff >>
rect 18 705 60 721
rect 18 688 25 705
rect 42 688 60 705
rect 18 671 60 688
rect 18 654 25 671
rect 42 654 60 671
rect 18 637 60 654
rect 75 705 117 721
rect 75 688 93 705
rect 110 688 117 705
rect 75 671 117 688
rect 75 654 93 671
rect 110 654 117 671
rect 75 637 117 654
rect 144 705 186 721
rect 144 688 151 705
rect 168 688 186 705
rect 144 671 186 688
rect 144 654 151 671
rect 168 654 186 671
rect 144 637 186 654
rect 201 705 243 721
rect 201 688 219 705
rect 236 688 243 705
rect 201 671 243 688
rect 201 654 219 671
rect 236 654 243 671
rect 201 637 243 654
rect 270 705 312 721
rect 270 688 277 705
rect 294 688 312 705
rect 270 671 312 688
rect 270 654 277 671
rect 294 654 312 671
rect 270 637 312 654
rect 327 705 369 721
rect 327 688 345 705
rect 362 688 369 705
rect 327 671 369 688
rect 327 654 345 671
rect 362 654 369 671
rect 327 637 369 654
<< ndiffc >>
rect 277 544 294 561
rect 345 544 362 561
rect 25 473 42 490
rect 25 439 42 456
rect 93 473 110 490
rect 93 439 110 456
rect 151 442 168 459
rect 151 408 168 425
rect 219 442 236 459
rect 219 408 236 425
rect 277 442 294 459
rect 277 408 294 425
rect 345 442 362 459
rect 345 408 362 425
rect 25 219 42 236
rect 25 185 42 202
rect 93 219 110 236
rect 93 185 110 202
rect 151 219 168 236
rect 151 185 168 202
rect 219 219 236 236
rect 219 185 236 202
rect 277 219 294 236
rect 277 185 294 202
rect 345 219 362 236
rect 345 185 362 202
rect 25 60 42 77
rect 93 60 110 77
rect 151 60 168 77
rect 219 60 236 77
<< pdiffc >>
rect 25 688 42 705
rect 25 654 42 671
rect 93 688 110 705
rect 93 654 110 671
rect 151 688 168 705
rect 151 654 168 671
rect 219 688 236 705
rect 219 654 236 671
rect 277 688 294 705
rect 277 654 294 671
rect 345 688 362 705
rect 345 654 362 671
<< psubdiff >>
rect 41 9 85 21
rect 41 -9 54 9
rect 72 -9 85 9
rect 41 -21 85 -9
rect 129 9 173 21
rect 129 -9 142 9
rect 160 -9 173 9
rect 129 -21 173 -9
rect 217 9 261 21
rect 217 -9 230 9
rect 248 -9 261 9
rect 217 -21 261 -9
rect 305 9 349 21
rect 305 -9 318 9
rect 336 -9 349 9
rect 305 -21 349 -9
<< nsubdiff >>
rect 41 779 85 790
rect 41 761 54 779
rect 72 761 85 779
rect 41 748 85 761
rect 129 779 173 790
rect 129 761 142 779
rect 160 761 173 779
rect 129 748 173 761
rect 217 779 261 790
rect 217 761 230 779
rect 248 761 261 779
rect 217 748 261 761
rect 305 779 349 790
rect 305 761 318 779
rect 336 761 349 779
rect 305 748 349 761
<< psubdiffcont >>
rect 54 -9 72 9
rect 142 -9 160 9
rect 230 -9 248 9
rect 318 -9 336 9
<< nsubdiffcont >>
rect 54 761 72 779
rect 142 761 160 779
rect 230 761 248 779
rect 318 761 336 779
<< poly >>
rect 60 721 75 734
rect 186 721 201 734
rect 312 721 327 734
rect 60 613 75 637
rect 60 604 165 613
rect 60 598 141 604
rect 133 587 141 598
rect 158 587 165 604
rect 133 579 165 587
rect 48 568 80 577
rect 48 551 56 568
rect 73 558 80 568
rect 186 558 201 637
rect 312 618 327 637
rect 301 613 335 618
rect 301 596 310 613
rect 327 596 335 613
rect 301 591 335 596
rect 312 574 327 591
rect 73 551 201 558
rect 48 543 201 551
rect 312 519 327 532
rect 60 506 75 519
rect 177 514 210 519
rect 177 497 185 514
rect 202 497 210 514
rect 177 492 210 497
rect 186 475 201 492
rect 312 475 327 488
rect 60 405 75 422
rect 52 400 85 405
rect 52 383 60 400
rect 77 383 85 400
rect 52 378 85 383
rect 186 378 201 391
rect 312 343 327 391
rect 304 338 337 343
rect 304 321 312 338
rect 329 321 337 338
rect 304 316 337 321
rect 50 291 83 296
rect 50 274 58 291
rect 75 274 83 291
rect 50 269 83 274
rect 178 291 211 296
rect 178 274 186 291
rect 203 274 211 291
rect 178 269 211 274
rect 60 252 75 269
rect 186 252 201 269
rect 312 252 327 316
rect 60 90 75 168
rect 186 155 201 168
rect 312 155 327 168
rect 176 129 209 134
rect 176 112 184 129
rect 201 112 209 129
rect 176 107 209 112
rect 186 90 201 107
rect 60 35 75 48
rect 186 35 201 48
<< polycont >>
rect 141 587 158 604
rect 56 551 73 568
rect 310 596 327 613
rect 185 497 202 514
rect 60 383 77 400
rect 312 321 329 338
rect 58 274 75 291
rect 186 274 203 291
rect 184 112 201 129
<< locali >>
rect 46 779 80 785
rect 46 778 54 779
rect 0 761 54 778
rect 72 778 80 779
rect 134 779 168 785
rect 134 778 142 779
rect 72 761 142 778
rect 160 778 168 779
rect 222 779 256 785
rect 222 778 230 779
rect 160 761 230 778
rect 248 778 256 779
rect 310 779 344 785
rect 310 778 318 779
rect 248 761 318 778
rect 336 778 344 779
rect 336 761 389 778
rect 31 754 80 761
rect 134 754 168 761
rect 222 754 256 761
rect 31 721 48 754
rect 226 721 243 754
rect 276 721 293 761
rect 310 754 344 761
rect 18 705 48 721
rect 18 688 25 705
rect 42 688 48 705
rect 18 671 48 688
rect 18 654 25 671
rect 42 654 48 671
rect 18 637 48 654
rect 87 705 117 721
rect 87 688 93 705
rect 110 688 117 705
rect 87 671 117 688
rect 87 654 93 671
rect 110 654 117 671
rect 87 637 117 654
rect 144 705 174 721
rect 144 688 151 705
rect 168 688 174 705
rect 144 671 174 688
rect 144 654 151 671
rect 168 654 174 671
rect 144 637 174 654
rect 213 705 243 721
rect 213 688 219 705
rect 236 688 243 705
rect 213 671 243 688
rect 213 654 219 671
rect 236 654 243 671
rect 213 637 243 654
rect 270 705 300 721
rect 270 688 277 705
rect 294 688 300 705
rect 270 671 300 688
rect 270 654 277 671
rect 294 654 300 671
rect 270 637 300 654
rect 339 705 369 721
rect 339 654 345 705
rect 362 654 369 705
rect 339 637 369 654
rect 87 577 104 637
rect 144 613 161 637
rect 301 613 335 618
rect 133 604 165 613
rect 133 587 141 604
rect 158 587 165 604
rect 133 579 165 587
rect 236 596 310 613
rect 327 596 335 613
rect 48 568 104 577
rect 48 551 56 568
rect 73 551 104 568
rect 48 543 104 551
rect 177 514 210 519
rect 18 490 48 506
rect 18 473 25 490
rect 42 473 48 490
rect 18 456 48 473
rect 18 439 25 456
rect 42 439 48 456
rect 18 422 48 439
rect 87 490 117 506
rect 177 497 185 514
rect 202 497 210 514
rect 177 492 210 497
rect 236 509 253 596
rect 301 591 335 596
rect 352 574 369 637
rect 270 561 300 574
rect 270 544 277 561
rect 294 544 300 561
rect 270 532 300 544
rect 339 561 369 574
rect 339 544 345 561
rect 362 544 369 561
rect 339 532 369 544
rect 236 492 356 509
rect 87 439 93 490
rect 110 439 117 490
rect 339 475 356 492
rect 87 422 117 439
rect 144 459 174 475
rect 144 442 151 459
rect 168 442 174 459
rect 144 425 174 442
rect 18 330 35 422
rect 144 408 151 425
rect 168 408 174 425
rect 52 400 85 405
rect 52 383 60 400
rect 77 383 85 400
rect 52 378 85 383
rect 144 391 174 408
rect 213 459 243 475
rect 213 408 219 459
rect 236 408 243 459
rect 213 391 243 408
rect 270 459 300 475
rect 270 442 277 459
rect 294 442 300 459
rect 270 425 300 442
rect 270 408 277 425
rect 294 408 300 425
rect 270 391 300 408
rect 339 459 369 475
rect 339 442 345 459
rect 362 442 369 459
rect 339 425 369 442
rect 339 408 345 425
rect 362 408 369 425
rect 339 391 369 408
rect 18 313 117 330
rect 50 291 83 296
rect 50 274 58 291
rect 75 274 83 291
rect 50 269 83 274
rect 100 252 117 313
rect 18 236 48 252
rect 18 219 25 236
rect 42 219 48 236
rect 18 202 48 219
rect 18 185 25 202
rect 42 185 48 202
rect 18 168 48 185
rect 87 236 117 252
rect 87 219 93 236
rect 110 219 117 236
rect 87 202 117 219
rect 87 185 93 202
rect 110 185 117 202
rect 87 168 117 185
rect 144 252 161 391
rect 270 296 287 391
rect 304 338 337 343
rect 304 321 312 338
rect 329 321 337 338
rect 304 316 337 321
rect 178 291 287 296
rect 178 274 186 291
rect 203 279 287 291
rect 203 274 211 279
rect 178 269 211 274
rect 144 236 174 252
rect 144 219 151 236
rect 168 219 174 236
rect 144 202 174 219
rect 144 185 151 202
rect 168 185 174 202
rect 144 168 174 185
rect 213 236 243 252
rect 213 185 219 236
rect 236 185 243 236
rect 213 168 243 185
rect 270 236 300 252
rect 270 219 277 236
rect 294 219 300 236
rect 270 202 300 219
rect 270 185 277 202
rect 294 185 300 202
rect 270 168 300 185
rect 339 236 369 252
rect 339 185 345 236
rect 362 185 369 236
rect 339 168 369 185
rect 18 90 35 168
rect 270 134 287 168
rect 100 129 287 134
rect 100 117 184 129
rect 100 90 117 117
rect 176 112 184 117
rect 201 117 287 129
rect 201 112 209 117
rect 176 107 209 112
rect 18 77 48 90
rect 18 60 25 77
rect 42 60 48 77
rect 18 48 48 60
rect 87 77 117 90
rect 87 60 93 77
rect 110 60 117 77
rect 87 48 117 60
rect 144 77 174 90
rect 144 60 151 77
rect 168 60 174 77
rect 144 48 174 60
rect 213 77 243 90
rect 213 60 219 77
rect 236 60 243 77
rect 213 48 243 60
rect 273 75 299 80
rect 273 58 279 75
rect 296 58 299 75
rect 273 54 299 58
rect 31 15 48 48
rect 226 15 243 48
rect 31 9 80 15
rect 31 8 54 9
rect 0 -9 54 8
rect 72 8 80 9
rect 134 9 168 15
rect 134 8 142 9
rect 72 -9 142 8
rect 160 8 168 9
rect 222 9 256 15
rect 222 8 230 9
rect 160 -9 230 8
rect 248 8 256 9
rect 276 8 293 54
rect 310 9 344 15
rect 310 8 318 9
rect 248 -9 318 8
rect 336 8 344 9
rect 336 -9 389 8
rect 47 -16 80 -9
rect 134 -16 168 -9
rect 222 -16 256 -9
rect 310 -16 344 -9
<< viali >>
rect 54 761 72 779
rect 142 761 160 779
rect 230 761 248 779
rect 318 761 336 779
rect 345 671 362 688
rect 141 587 158 604
rect 310 596 327 613
rect 56 551 73 568
rect 185 497 202 514
rect 277 544 294 561
rect 93 456 110 473
rect 60 383 77 400
rect 219 425 236 442
rect 58 274 75 291
rect 312 321 329 338
rect 186 274 203 291
rect 219 202 236 219
rect 345 202 362 219
rect 184 112 201 129
rect 151 60 168 77
rect 219 60 236 77
rect 279 58 296 75
rect 54 -9 72 9
rect 142 -9 160 9
rect 230 -9 248 9
rect 318 -9 336 9
<< metal1 >>
rect 0 779 389 785
rect 0 761 54 779
rect 72 761 142 779
rect 160 761 230 779
rect 248 761 318 779
rect 336 761 389 779
rect 0 754 389 761
rect 339 691 369 694
rect 339 665 341 691
rect 367 665 369 691
rect 339 662 369 665
rect 133 609 165 613
rect 133 583 136 609
rect 162 583 165 609
rect 301 592 306 618
rect 332 592 335 618
rect 301 591 335 592
rect 133 579 165 583
rect 49 573 79 576
rect 49 547 51 573
rect 77 547 79 573
rect 49 544 79 547
rect 270 566 299 569
rect 270 540 272 566
rect 298 540 299 566
rect 270 537 299 540
rect 177 514 210 519
rect 177 512 185 514
rect 176 498 185 512
rect 177 497 185 498
rect 202 512 210 514
rect 202 498 211 512
rect 202 497 210 498
rect 177 492 210 497
rect 87 474 117 477
rect 87 448 89 474
rect 115 448 117 474
rect 87 445 117 448
rect 213 446 243 449
rect 213 420 215 446
rect 241 420 243 446
rect 213 417 243 420
rect 52 400 85 405
rect 52 399 60 400
rect 51 385 60 399
rect 52 383 60 385
rect 77 399 85 400
rect 77 385 86 399
rect 77 383 85 385
rect 52 378 85 383
rect 304 338 337 343
rect 304 336 312 338
rect 303 322 312 336
rect 304 321 312 322
rect 329 336 337 338
rect 329 322 338 336
rect 329 321 337 322
rect 304 316 337 321
rect 50 270 53 296
rect 79 289 83 296
rect 178 291 211 296
rect 178 289 186 291
rect 79 275 186 289
rect 79 270 83 275
rect 50 269 83 270
rect 145 80 159 275
rect 178 274 186 275
rect 203 274 211 291
rect 178 269 211 274
rect 341 222 369 225
rect 213 219 242 222
rect 213 202 219 219
rect 236 202 242 219
rect 213 195 242 202
rect 367 196 369 222
rect 176 108 179 134
rect 205 108 208 134
rect 176 107 208 108
rect 222 82 236 195
rect 341 193 369 196
rect 145 77 174 80
rect 145 60 151 77
rect 168 60 174 77
rect 145 57 174 60
rect 213 77 242 82
rect 213 60 219 77
rect 236 60 242 77
rect 213 57 242 60
rect 270 80 299 83
rect 270 54 273 80
rect 270 51 299 54
rect 0 9 389 15
rect 0 -9 54 9
rect 72 -9 142 9
rect 160 -9 230 9
rect 248 -9 318 9
rect 336 -9 389 9
rect 0 -16 389 -9
<< via1 >>
rect 341 688 367 691
rect 341 671 345 688
rect 345 671 362 688
rect 362 671 367 688
rect 341 665 367 671
rect 136 604 162 609
rect 136 587 141 604
rect 141 587 158 604
rect 158 587 162 604
rect 136 583 162 587
rect 306 613 332 618
rect 306 596 310 613
rect 310 596 327 613
rect 327 596 332 613
rect 306 592 332 596
rect 51 568 77 573
rect 51 551 56 568
rect 56 551 73 568
rect 73 551 77 568
rect 51 547 77 551
rect 272 561 298 566
rect 272 544 277 561
rect 277 544 294 561
rect 294 544 298 561
rect 272 540 298 544
rect 89 473 115 474
rect 89 456 93 473
rect 93 456 110 473
rect 110 456 115 473
rect 89 448 115 456
rect 215 442 241 446
rect 215 425 219 442
rect 219 425 236 442
rect 236 425 241 442
rect 215 420 241 425
rect 53 291 79 296
rect 53 274 58 291
rect 58 274 75 291
rect 75 274 79 291
rect 53 270 79 274
rect 341 219 367 222
rect 341 202 345 219
rect 345 202 362 219
rect 362 202 367 219
rect 341 196 367 202
rect 179 129 205 134
rect 179 112 184 129
rect 184 112 201 129
rect 201 112 205 129
rect 179 108 205 112
rect 273 75 299 80
rect 273 58 279 75
rect 279 58 296 75
rect 296 58 299 75
rect 273 54 299 58
<< metal2 >>
rect 49 573 79 576
rect 49 547 51 573
rect 77 547 79 573
rect 49 544 79 547
rect 50 296 64 544
rect 96 477 110 808
rect 133 583 136 609
rect 162 583 165 609
rect 133 581 165 583
rect 87 474 117 477
rect 87 448 89 474
rect 115 448 117 474
rect 87 445 117 448
rect 50 270 53 296
rect 79 270 82 296
rect 50 269 82 270
rect 96 -21 110 445
rect 144 134 158 581
rect 222 449 236 808
rect 313 618 327 808
rect 341 691 369 694
rect 367 665 369 691
rect 341 662 369 665
rect 301 592 306 618
rect 332 592 335 618
rect 301 591 335 592
rect 270 566 299 569
rect 270 540 272 566
rect 298 540 299 566
rect 270 537 299 540
rect 213 446 243 449
rect 213 420 215 446
rect 241 420 243 446
rect 213 417 243 420
rect 144 120 179 134
rect 176 108 179 120
rect 205 108 208 134
rect 176 107 208 108
rect 222 -21 236 417
rect 270 83 284 537
rect 270 80 299 83
rect 270 54 273 80
rect 270 51 299 54
rect 313 -21 327 591
rect 355 225 369 662
rect 341 222 369 225
rect 367 196 369 222
rect 341 193 369 196
<< labels >>
flabel metal1 108 762 108 762 0 FreeSans 120 0 0 0 vdd
port 0 nsew
flabel metal1 104 -13 104 -13 0 FreeSans 120 0 0 0 gnd
port 1 nsew
flabel metal2 141 587 158 604 0 FreeSans 80 0 0 0 qbar
flabel metal2 359 494 359 494 0 FreeSans 80 0 0 0 net1
flabel locali 100 322 100 322 0 FreeSans 80 0 0 0 net2
flabel locali 159 332 159 332 0 FreeSans 80 0 0 0 net3
flabel metal2 56 551 73 568 0 FreeSans 80 0 0 0 q
flabel metal2 103 406 103 406 0 FreeSans 80 0 0 0 rbl0
port 11 nsew
flabel metal2 228 376 228 376 0 FreeSans 80 0 0 0 rbl1
port 12 nsew
flabel metal2 314 509 314 509 0 FreeSans 80 0 0 0 wbl0
port 13 nsew
flabel metal1 303 330 303 330 0 FreeSans 80 0 0 0 wwl0
port 14 nsew
flabel metal1 211 505 211 505 0 FreeSans 80 0 0 0 rwl1
port 15 nsew
flabel metal1 86 391 86 391 0 FreeSans 80 0 0 0 rwl0
port 16 nsew
<< properties >>
string FIXED_BBOX 0 0 389 770
<< end >>
