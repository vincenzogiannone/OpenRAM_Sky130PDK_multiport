magic
tech sky130A
magscale 1 2
timestamp 1644969367
<< checkpaint >>
rect -1319 -1316 7949 1611
<< nwell >>
rect -54 233 6684 351
rect -59 65 6689 233
rect -54 -54 6684 65
<< scpmos >>
rect 60 0 90 297
rect 168 0 198 297
rect 276 0 306 297
rect 384 0 414 297
rect 492 0 522 297
rect 600 0 630 297
rect 708 0 738 297
rect 816 0 846 297
rect 924 0 954 297
rect 1032 0 1062 297
rect 1140 0 1170 297
rect 1248 0 1278 297
rect 1356 0 1386 297
rect 1464 0 1494 297
rect 1572 0 1602 297
rect 1680 0 1710 297
rect 1788 0 1818 297
rect 1896 0 1926 297
rect 2004 0 2034 297
rect 2112 0 2142 297
rect 2220 0 2250 297
rect 2328 0 2358 297
rect 2436 0 2466 297
rect 2544 0 2574 297
rect 2652 0 2682 297
rect 2760 0 2790 297
rect 2868 0 2898 297
rect 2976 0 3006 297
rect 3084 0 3114 297
rect 3192 0 3222 297
rect 3300 0 3330 297
rect 3408 0 3438 297
rect 3516 0 3546 297
rect 3624 0 3654 297
rect 3732 0 3762 297
rect 3840 0 3870 297
rect 3948 0 3978 297
rect 4056 0 4086 297
rect 4164 0 4194 297
rect 4272 0 4302 297
rect 4380 0 4410 297
rect 4488 0 4518 297
rect 4596 0 4626 297
rect 4704 0 4734 297
rect 4812 0 4842 297
rect 4920 0 4950 297
rect 5028 0 5058 297
rect 5136 0 5166 297
rect 5244 0 5274 297
rect 5352 0 5382 297
rect 5460 0 5490 297
rect 5568 0 5598 297
rect 5676 0 5706 297
rect 5784 0 5814 297
rect 5892 0 5922 297
rect 6000 0 6030 297
rect 6108 0 6138 297
rect 6216 0 6246 297
rect 6324 0 6354 297
rect 6432 0 6462 297
rect 6540 0 6570 297
<< pdiff >>
rect 0 166 60 297
rect 0 132 8 166
rect 42 132 60 166
rect 0 0 60 132
rect 90 166 168 297
rect 90 132 112 166
rect 146 132 168 166
rect 90 0 168 132
rect 198 166 276 297
rect 198 132 220 166
rect 254 132 276 166
rect 198 0 276 132
rect 306 166 384 297
rect 306 132 328 166
rect 362 132 384 166
rect 306 0 384 132
rect 414 166 492 297
rect 414 132 436 166
rect 470 132 492 166
rect 414 0 492 132
rect 522 166 600 297
rect 522 132 544 166
rect 578 132 600 166
rect 522 0 600 132
rect 630 166 708 297
rect 630 132 652 166
rect 686 132 708 166
rect 630 0 708 132
rect 738 166 816 297
rect 738 132 760 166
rect 794 132 816 166
rect 738 0 816 132
rect 846 166 924 297
rect 846 132 868 166
rect 902 132 924 166
rect 846 0 924 132
rect 954 166 1032 297
rect 954 132 976 166
rect 1010 132 1032 166
rect 954 0 1032 132
rect 1062 166 1140 297
rect 1062 132 1084 166
rect 1118 132 1140 166
rect 1062 0 1140 132
rect 1170 166 1248 297
rect 1170 132 1192 166
rect 1226 132 1248 166
rect 1170 0 1248 132
rect 1278 166 1356 297
rect 1278 132 1300 166
rect 1334 132 1356 166
rect 1278 0 1356 132
rect 1386 166 1464 297
rect 1386 132 1408 166
rect 1442 132 1464 166
rect 1386 0 1464 132
rect 1494 166 1572 297
rect 1494 132 1516 166
rect 1550 132 1572 166
rect 1494 0 1572 132
rect 1602 166 1680 297
rect 1602 132 1624 166
rect 1658 132 1680 166
rect 1602 0 1680 132
rect 1710 166 1788 297
rect 1710 132 1732 166
rect 1766 132 1788 166
rect 1710 0 1788 132
rect 1818 166 1896 297
rect 1818 132 1840 166
rect 1874 132 1896 166
rect 1818 0 1896 132
rect 1926 166 2004 297
rect 1926 132 1948 166
rect 1982 132 2004 166
rect 1926 0 2004 132
rect 2034 166 2112 297
rect 2034 132 2056 166
rect 2090 132 2112 166
rect 2034 0 2112 132
rect 2142 166 2220 297
rect 2142 132 2164 166
rect 2198 132 2220 166
rect 2142 0 2220 132
rect 2250 166 2328 297
rect 2250 132 2272 166
rect 2306 132 2328 166
rect 2250 0 2328 132
rect 2358 166 2436 297
rect 2358 132 2380 166
rect 2414 132 2436 166
rect 2358 0 2436 132
rect 2466 166 2544 297
rect 2466 132 2488 166
rect 2522 132 2544 166
rect 2466 0 2544 132
rect 2574 166 2652 297
rect 2574 132 2596 166
rect 2630 132 2652 166
rect 2574 0 2652 132
rect 2682 166 2760 297
rect 2682 132 2704 166
rect 2738 132 2760 166
rect 2682 0 2760 132
rect 2790 166 2868 297
rect 2790 132 2812 166
rect 2846 132 2868 166
rect 2790 0 2868 132
rect 2898 166 2976 297
rect 2898 132 2920 166
rect 2954 132 2976 166
rect 2898 0 2976 132
rect 3006 166 3084 297
rect 3006 132 3028 166
rect 3062 132 3084 166
rect 3006 0 3084 132
rect 3114 166 3192 297
rect 3114 132 3136 166
rect 3170 132 3192 166
rect 3114 0 3192 132
rect 3222 166 3300 297
rect 3222 132 3244 166
rect 3278 132 3300 166
rect 3222 0 3300 132
rect 3330 166 3408 297
rect 3330 132 3352 166
rect 3386 132 3408 166
rect 3330 0 3408 132
rect 3438 166 3516 297
rect 3438 132 3460 166
rect 3494 132 3516 166
rect 3438 0 3516 132
rect 3546 166 3624 297
rect 3546 132 3568 166
rect 3602 132 3624 166
rect 3546 0 3624 132
rect 3654 166 3732 297
rect 3654 132 3676 166
rect 3710 132 3732 166
rect 3654 0 3732 132
rect 3762 166 3840 297
rect 3762 132 3784 166
rect 3818 132 3840 166
rect 3762 0 3840 132
rect 3870 166 3948 297
rect 3870 132 3892 166
rect 3926 132 3948 166
rect 3870 0 3948 132
rect 3978 166 4056 297
rect 3978 132 4000 166
rect 4034 132 4056 166
rect 3978 0 4056 132
rect 4086 166 4164 297
rect 4086 132 4108 166
rect 4142 132 4164 166
rect 4086 0 4164 132
rect 4194 166 4272 297
rect 4194 132 4216 166
rect 4250 132 4272 166
rect 4194 0 4272 132
rect 4302 166 4380 297
rect 4302 132 4324 166
rect 4358 132 4380 166
rect 4302 0 4380 132
rect 4410 166 4488 297
rect 4410 132 4432 166
rect 4466 132 4488 166
rect 4410 0 4488 132
rect 4518 166 4596 297
rect 4518 132 4540 166
rect 4574 132 4596 166
rect 4518 0 4596 132
rect 4626 166 4704 297
rect 4626 132 4648 166
rect 4682 132 4704 166
rect 4626 0 4704 132
rect 4734 166 4812 297
rect 4734 132 4756 166
rect 4790 132 4812 166
rect 4734 0 4812 132
rect 4842 166 4920 297
rect 4842 132 4864 166
rect 4898 132 4920 166
rect 4842 0 4920 132
rect 4950 166 5028 297
rect 4950 132 4972 166
rect 5006 132 5028 166
rect 4950 0 5028 132
rect 5058 166 5136 297
rect 5058 132 5080 166
rect 5114 132 5136 166
rect 5058 0 5136 132
rect 5166 166 5244 297
rect 5166 132 5188 166
rect 5222 132 5244 166
rect 5166 0 5244 132
rect 5274 166 5352 297
rect 5274 132 5296 166
rect 5330 132 5352 166
rect 5274 0 5352 132
rect 5382 166 5460 297
rect 5382 132 5404 166
rect 5438 132 5460 166
rect 5382 0 5460 132
rect 5490 166 5568 297
rect 5490 132 5512 166
rect 5546 132 5568 166
rect 5490 0 5568 132
rect 5598 166 5676 297
rect 5598 132 5620 166
rect 5654 132 5676 166
rect 5598 0 5676 132
rect 5706 166 5784 297
rect 5706 132 5728 166
rect 5762 132 5784 166
rect 5706 0 5784 132
rect 5814 166 5892 297
rect 5814 132 5836 166
rect 5870 132 5892 166
rect 5814 0 5892 132
rect 5922 166 6000 297
rect 5922 132 5944 166
rect 5978 132 6000 166
rect 5922 0 6000 132
rect 6030 166 6108 297
rect 6030 132 6052 166
rect 6086 132 6108 166
rect 6030 0 6108 132
rect 6138 166 6216 297
rect 6138 132 6160 166
rect 6194 132 6216 166
rect 6138 0 6216 132
rect 6246 166 6324 297
rect 6246 132 6268 166
rect 6302 132 6324 166
rect 6246 0 6324 132
rect 6354 166 6432 297
rect 6354 132 6376 166
rect 6410 132 6432 166
rect 6354 0 6432 132
rect 6462 166 6540 297
rect 6462 132 6484 166
rect 6518 132 6540 166
rect 6462 0 6540 132
rect 6570 166 6630 297
rect 6570 132 6588 166
rect 6622 132 6630 166
rect 6570 0 6630 132
<< pdiffc >>
rect 8 132 42 166
rect 112 132 146 166
rect 220 132 254 166
rect 328 132 362 166
rect 436 132 470 166
rect 544 132 578 166
rect 652 132 686 166
rect 760 132 794 166
rect 868 132 902 166
rect 976 132 1010 166
rect 1084 132 1118 166
rect 1192 132 1226 166
rect 1300 132 1334 166
rect 1408 132 1442 166
rect 1516 132 1550 166
rect 1624 132 1658 166
rect 1732 132 1766 166
rect 1840 132 1874 166
rect 1948 132 1982 166
rect 2056 132 2090 166
rect 2164 132 2198 166
rect 2272 132 2306 166
rect 2380 132 2414 166
rect 2488 132 2522 166
rect 2596 132 2630 166
rect 2704 132 2738 166
rect 2812 132 2846 166
rect 2920 132 2954 166
rect 3028 132 3062 166
rect 3136 132 3170 166
rect 3244 132 3278 166
rect 3352 132 3386 166
rect 3460 132 3494 166
rect 3568 132 3602 166
rect 3676 132 3710 166
rect 3784 132 3818 166
rect 3892 132 3926 166
rect 4000 132 4034 166
rect 4108 132 4142 166
rect 4216 132 4250 166
rect 4324 132 4358 166
rect 4432 132 4466 166
rect 4540 132 4574 166
rect 4648 132 4682 166
rect 4756 132 4790 166
rect 4864 132 4898 166
rect 4972 132 5006 166
rect 5080 132 5114 166
rect 5188 132 5222 166
rect 5296 132 5330 166
rect 5404 132 5438 166
rect 5512 132 5546 166
rect 5620 132 5654 166
rect 5728 132 5762 166
rect 5836 132 5870 166
rect 5944 132 5978 166
rect 6052 132 6086 166
rect 6160 132 6194 166
rect 6268 132 6302 166
rect 6376 132 6410 166
rect 6484 132 6518 166
rect 6588 132 6622 166
<< poly >>
rect 60 297 90 323
rect 168 297 198 323
rect 276 297 306 323
rect 384 297 414 323
rect 492 297 522 323
rect 600 297 630 323
rect 708 297 738 323
rect 816 297 846 323
rect 924 297 954 323
rect 1032 297 1062 323
rect 1140 297 1170 323
rect 1248 297 1278 323
rect 1356 297 1386 323
rect 1464 297 1494 323
rect 1572 297 1602 323
rect 1680 297 1710 323
rect 1788 297 1818 323
rect 1896 297 1926 323
rect 2004 297 2034 323
rect 2112 297 2142 323
rect 2220 297 2250 323
rect 2328 297 2358 323
rect 2436 297 2466 323
rect 2544 297 2574 323
rect 2652 297 2682 323
rect 2760 297 2790 323
rect 2868 297 2898 323
rect 2976 297 3006 323
rect 3084 297 3114 323
rect 3192 297 3222 323
rect 3300 297 3330 323
rect 3408 297 3438 323
rect 3516 297 3546 323
rect 3624 297 3654 323
rect 3732 297 3762 323
rect 3840 297 3870 323
rect 3948 297 3978 323
rect 4056 297 4086 323
rect 4164 297 4194 323
rect 4272 297 4302 323
rect 4380 297 4410 323
rect 4488 297 4518 323
rect 4596 297 4626 323
rect 4704 297 4734 323
rect 4812 297 4842 323
rect 4920 297 4950 323
rect 5028 297 5058 323
rect 5136 297 5166 323
rect 5244 297 5274 323
rect 5352 297 5382 323
rect 5460 297 5490 323
rect 5568 297 5598 323
rect 5676 297 5706 323
rect 5784 297 5814 323
rect 5892 297 5922 323
rect 6000 297 6030 323
rect 6108 297 6138 323
rect 6216 297 6246 323
rect 6324 297 6354 323
rect 6432 297 6462 323
rect 6540 297 6570 323
rect 60 -26 90 0
rect 168 -26 198 0
rect 276 -26 306 0
rect 384 -26 414 0
rect 492 -26 522 0
rect 600 -26 630 0
rect 708 -26 738 0
rect 816 -26 846 0
rect 924 -26 954 0
rect 1032 -26 1062 0
rect 1140 -26 1170 0
rect 1248 -26 1278 0
rect 1356 -26 1386 0
rect 1464 -26 1494 0
rect 1572 -26 1602 0
rect 1680 -26 1710 0
rect 1788 -26 1818 0
rect 1896 -26 1926 0
rect 2004 -26 2034 0
rect 2112 -26 2142 0
rect 2220 -26 2250 0
rect 2328 -26 2358 0
rect 2436 -26 2466 0
rect 2544 -26 2574 0
rect 2652 -26 2682 0
rect 2760 -26 2790 0
rect 2868 -26 2898 0
rect 2976 -26 3006 0
rect 3084 -26 3114 0
rect 3192 -26 3222 0
rect 3300 -26 3330 0
rect 3408 -26 3438 0
rect 3516 -26 3546 0
rect 3624 -26 3654 0
rect 3732 -26 3762 0
rect 3840 -26 3870 0
rect 3948 -26 3978 0
rect 4056 -26 4086 0
rect 4164 -26 4194 0
rect 4272 -26 4302 0
rect 4380 -26 4410 0
rect 4488 -26 4518 0
rect 4596 -26 4626 0
rect 4704 -26 4734 0
rect 4812 -26 4842 0
rect 4920 -26 4950 0
rect 5028 -26 5058 0
rect 5136 -26 5166 0
rect 5244 -26 5274 0
rect 5352 -26 5382 0
rect 5460 -26 5490 0
rect 5568 -26 5598 0
rect 5676 -26 5706 0
rect 5784 -26 5814 0
rect 5892 -26 5922 0
rect 6000 -26 6030 0
rect 6108 -26 6138 0
rect 6216 -26 6246 0
rect 6324 -26 6354 0
rect 6432 -26 6462 0
rect 6540 -26 6570 0
rect 60 -56 6570 -26
<< locali >>
rect 8 166 42 182
rect 8 116 42 132
rect 112 166 146 182
rect 112 82 146 132
rect 220 166 254 182
rect 220 116 254 132
rect 328 166 362 182
rect 328 82 362 132
rect 436 166 470 182
rect 436 116 470 132
rect 544 166 578 182
rect 544 82 578 132
rect 652 166 686 182
rect 652 116 686 132
rect 760 166 794 182
rect 760 82 794 132
rect 868 166 902 182
rect 868 116 902 132
rect 976 166 1010 182
rect 976 82 1010 132
rect 1084 166 1118 182
rect 1084 116 1118 132
rect 1192 166 1226 182
rect 1192 82 1226 132
rect 1300 166 1334 182
rect 1300 116 1334 132
rect 1408 166 1442 182
rect 1408 82 1442 132
rect 1516 166 1550 182
rect 1516 116 1550 132
rect 1624 166 1658 182
rect 1624 82 1658 132
rect 1732 166 1766 182
rect 1732 116 1766 132
rect 1840 166 1874 182
rect 1840 82 1874 132
rect 1948 166 1982 182
rect 1948 116 1982 132
rect 2056 166 2090 182
rect 2056 82 2090 132
rect 2164 166 2198 182
rect 2164 116 2198 132
rect 2272 166 2306 182
rect 2272 82 2306 132
rect 2380 166 2414 182
rect 2380 116 2414 132
rect 2488 166 2522 182
rect 2488 82 2522 132
rect 2596 166 2630 182
rect 2596 116 2630 132
rect 2704 166 2738 182
rect 2704 82 2738 132
rect 2812 166 2846 182
rect 2812 116 2846 132
rect 2920 166 2954 182
rect 2920 82 2954 132
rect 3028 166 3062 182
rect 3028 116 3062 132
rect 3136 166 3170 182
rect 3136 82 3170 132
rect 3244 166 3278 182
rect 3244 116 3278 132
rect 3352 166 3386 182
rect 3352 82 3386 132
rect 3460 166 3494 182
rect 3460 116 3494 132
rect 3568 166 3602 182
rect 3568 82 3602 132
rect 3676 166 3710 182
rect 3676 116 3710 132
rect 3784 166 3818 182
rect 3784 82 3818 132
rect 3892 166 3926 182
rect 3892 116 3926 132
rect 4000 166 4034 182
rect 4000 82 4034 132
rect 4108 166 4142 182
rect 4108 116 4142 132
rect 4216 166 4250 182
rect 4216 82 4250 132
rect 4324 166 4358 182
rect 4324 116 4358 132
rect 4432 166 4466 182
rect 4432 82 4466 132
rect 4540 166 4574 182
rect 4540 116 4574 132
rect 4648 166 4682 182
rect 4648 82 4682 132
rect 4756 166 4790 182
rect 4756 116 4790 132
rect 4864 166 4898 182
rect 4864 82 4898 132
rect 4972 166 5006 182
rect 4972 116 5006 132
rect 5080 166 5114 182
rect 5080 82 5114 132
rect 5188 166 5222 182
rect 5188 116 5222 132
rect 5296 166 5330 182
rect 5296 82 5330 132
rect 5404 166 5438 182
rect 5404 116 5438 132
rect 5512 166 5546 182
rect 5512 82 5546 132
rect 5620 166 5654 182
rect 5620 116 5654 132
rect 5728 166 5762 182
rect 5728 82 5762 132
rect 5836 166 5870 182
rect 5836 116 5870 132
rect 5944 166 5978 182
rect 5944 82 5978 132
rect 6052 166 6086 182
rect 6052 116 6086 132
rect 6160 166 6194 182
rect 6160 82 6194 132
rect 6268 166 6302 182
rect 6268 116 6302 132
rect 6376 166 6410 182
rect 6376 82 6410 132
rect 6484 166 6518 182
rect 6484 116 6518 132
rect 6588 166 6622 182
rect 6588 82 6622 132
rect 112 48 6622 82
use contact_9  contact_9_0
timestamp 1644969367
transform 1 0 6580 0 1 108
box 0 0 2 2
use contact_9  contact_9_1
timestamp 1644969367
transform 1 0 6476 0 1 108
box 0 0 2 2
use contact_9  contact_9_2
timestamp 1644969367
transform 1 0 6368 0 1 108
box 0 0 2 2
use contact_9  contact_9_3
timestamp 1644969367
transform 1 0 6260 0 1 108
box 0 0 2 2
use contact_9  contact_9_4
timestamp 1644969367
transform 1 0 6152 0 1 108
box 0 0 2 2
use contact_9  contact_9_5
timestamp 1644969367
transform 1 0 6044 0 1 108
box 0 0 2 2
use contact_9  contact_9_6
timestamp 1644969367
transform 1 0 5936 0 1 108
box 0 0 2 2
use contact_9  contact_9_7
timestamp 1644969367
transform 1 0 5828 0 1 108
box 0 0 2 2
use contact_9  contact_9_8
timestamp 1644969367
transform 1 0 5720 0 1 108
box 0 0 2 2
use contact_9  contact_9_9
timestamp 1644969367
transform 1 0 5612 0 1 108
box 0 0 2 2
use contact_9  contact_9_10
timestamp 1644969367
transform 1 0 5504 0 1 108
box 0 0 2 2
use contact_9  contact_9_11
timestamp 1644969367
transform 1 0 5396 0 1 108
box 0 0 2 2
use contact_9  contact_9_12
timestamp 1644969367
transform 1 0 5288 0 1 108
box 0 0 2 2
use contact_9  contact_9_13
timestamp 1644969367
transform 1 0 5180 0 1 108
box 0 0 2 2
use contact_9  contact_9_14
timestamp 1644969367
transform 1 0 5072 0 1 108
box 0 0 2 2
use contact_9  contact_9_15
timestamp 1644969367
transform 1 0 4964 0 1 108
box 0 0 2 2
use contact_9  contact_9_16
timestamp 1644969367
transform 1 0 4856 0 1 108
box 0 0 2 2
use contact_9  contact_9_17
timestamp 1644969367
transform 1 0 4748 0 1 108
box 0 0 2 2
use contact_9  contact_9_18
timestamp 1644969367
transform 1 0 4640 0 1 108
box 0 0 2 2
use contact_9  contact_9_19
timestamp 1644969367
transform 1 0 4532 0 1 108
box 0 0 2 2
use contact_9  contact_9_20
timestamp 1644969367
transform 1 0 4424 0 1 108
box 0 0 2 2
use contact_9  contact_9_21
timestamp 1644969367
transform 1 0 4316 0 1 108
box 0 0 2 2
use contact_9  contact_9_22
timestamp 1644969367
transform 1 0 4208 0 1 108
box 0 0 2 2
use contact_9  contact_9_23
timestamp 1644969367
transform 1 0 4100 0 1 108
box 0 0 2 2
use contact_9  contact_9_24
timestamp 1644969367
transform 1 0 3992 0 1 108
box 0 0 2 2
use contact_9  contact_9_25
timestamp 1644969367
transform 1 0 3884 0 1 108
box 0 0 2 2
use contact_9  contact_9_26
timestamp 1644969367
transform 1 0 3776 0 1 108
box 0 0 2 2
use contact_9  contact_9_27
timestamp 1644969367
transform 1 0 3668 0 1 108
box 0 0 2 2
use contact_9  contact_9_28
timestamp 1644969367
transform 1 0 3560 0 1 108
box 0 0 2 2
use contact_9  contact_9_29
timestamp 1644969367
transform 1 0 3452 0 1 108
box 0 0 2 2
use contact_9  contact_9_30
timestamp 1644969367
transform 1 0 3344 0 1 108
box 0 0 2 2
use contact_9  contact_9_31
timestamp 1644969367
transform 1 0 3236 0 1 108
box 0 0 2 2
use contact_9  contact_9_32
timestamp 1644969367
transform 1 0 3128 0 1 108
box 0 0 2 2
use contact_9  contact_9_33
timestamp 1644969367
transform 1 0 3020 0 1 108
box 0 0 2 2
use contact_9  contact_9_34
timestamp 1644969367
transform 1 0 2912 0 1 108
box 0 0 2 2
use contact_9  contact_9_35
timestamp 1644969367
transform 1 0 2804 0 1 108
box 0 0 2 2
use contact_9  contact_9_36
timestamp 1644969367
transform 1 0 2696 0 1 108
box 0 0 2 2
use contact_9  contact_9_37
timestamp 1644969367
transform 1 0 2588 0 1 108
box 0 0 2 2
use contact_9  contact_9_38
timestamp 1644969367
transform 1 0 2480 0 1 108
box 0 0 2 2
use contact_9  contact_9_39
timestamp 1644969367
transform 1 0 2372 0 1 108
box 0 0 2 2
use contact_9  contact_9_40
timestamp 1644969367
transform 1 0 2264 0 1 108
box 0 0 2 2
use contact_9  contact_9_41
timestamp 1644969367
transform 1 0 2156 0 1 108
box 0 0 2 2
use contact_9  contact_9_42
timestamp 1644969367
transform 1 0 2048 0 1 108
box 0 0 2 2
use contact_9  contact_9_43
timestamp 1644969367
transform 1 0 1940 0 1 108
box 0 0 2 2
use contact_9  contact_9_44
timestamp 1644969367
transform 1 0 1832 0 1 108
box 0 0 2 2
use contact_9  contact_9_45
timestamp 1644969367
transform 1 0 1724 0 1 108
box 0 0 2 2
use contact_9  contact_9_46
timestamp 1644969367
transform 1 0 1616 0 1 108
box 0 0 2 2
use contact_9  contact_9_47
timestamp 1644969367
transform 1 0 1508 0 1 108
box 0 0 2 2
use contact_9  contact_9_48
timestamp 1644969367
transform 1 0 1400 0 1 108
box 0 0 2 2
use contact_9  contact_9_49
timestamp 1644969367
transform 1 0 1292 0 1 108
box 0 0 2 2
use contact_9  contact_9_50
timestamp 1644969367
transform 1 0 1184 0 1 108
box 0 0 2 2
use contact_9  contact_9_51
timestamp 1644969367
transform 1 0 1076 0 1 108
box 0 0 2 2
use contact_9  contact_9_52
timestamp 1644969367
transform 1 0 968 0 1 108
box 0 0 2 2
use contact_9  contact_9_53
timestamp 1644969367
transform 1 0 860 0 1 108
box 0 0 2 2
use contact_9  contact_9_54
timestamp 1644969367
transform 1 0 752 0 1 108
box 0 0 2 2
use contact_9  contact_9_55
timestamp 1644969367
transform 1 0 644 0 1 108
box 0 0 2 2
use contact_9  contact_9_56
timestamp 1644969367
transform 1 0 536 0 1 108
box 0 0 2 2
use contact_9  contact_9_57
timestamp 1644969367
transform 1 0 428 0 1 108
box 0 0 2 2
use contact_9  contact_9_58
timestamp 1644969367
transform 1 0 320 0 1 108
box 0 0 2 2
use contact_9  contact_9_59
timestamp 1644969367
transform 1 0 212 0 1 108
box 0 0 2 2
use contact_9  contact_9_60
timestamp 1644969367
transform 1 0 104 0 1 108
box 0 0 2 2
use contact_9  contact_9_61
timestamp 1644969367
transform 1 0 0 0 1 108
box 0 0 2 2
<< labels >>
rlabel mvvaractor s 3315 -41 3315 -41 4 G
rlabel locali s 3909 149 3909 149 4 S
rlabel locali s 1101 149 1101 149 4 S
rlabel locali s 885 149 885 149 4 S
rlabel locali s 2181 149 2181 149 4 S
rlabel locali s 4341 149 4341 149 4 S
rlabel locali s 3045 149 3045 149 4 S
rlabel locali s 3693 149 3693 149 4 S
rlabel locali s 237 149 237 149 4 S
rlabel locali s 3261 149 3261 149 4 S
rlabel locali s 1533 149 1533 149 4 S
rlabel locali s 669 149 669 149 4 S
rlabel locali s 5853 149 5853 149 4 S
rlabel locali s 25 149 25 149 4 S
rlabel locali s 3477 149 3477 149 4 S
rlabel locali s 1965 149 1965 149 4 S
rlabel locali s 453 149 453 149 4 S
rlabel locali s 1317 149 1317 149 4 S
rlabel locali s 2397 149 2397 149 4 S
rlabel locali s 6501 149 6501 149 4 S
rlabel locali s 5421 149 5421 149 4 S
rlabel locali s 2613 149 2613 149 4 S
rlabel locali s 4557 149 4557 149 4 S
rlabel locali s 4773 149 4773 149 4 S
rlabel locali s 2829 149 2829 149 4 S
rlabel locali s 6285 149 6285 149 4 S
rlabel locali s 4125 149 4125 149 4 S
rlabel locali s 5637 149 5637 149 4 S
rlabel locali s 6069 149 6069 149 4 S
rlabel locali s 4989 149 4989 149 4 S
rlabel locali s 1749 149 1749 149 4 S
rlabel locali s 5205 149 5205 149 4 S
rlabel locali s 3367 65 3367 65 4 D
<< properties >>
string FIXED_BBOX -54 -56 6684 65
string GDS_FILE sram_0rw2r1w_32_128_sky130A.gds
string GDS_END 3347732
string GDS_START 3335080
<< end >>
