magic
tech sky130A
magscale 1 2
timestamp 1643678851
<< checkpaint >>
rect -1260 -1302 2530 50518
<< metal1 >>
rect 536 48606 618 48634
rect 1176 48536 1204 48564
rect 234 48486 318 48514
rect 1176 48410 1204 48438
rect 56 48340 126 48368
rect 1176 48184 1204 48212
rect 1176 47144 1204 47172
rect 56 46988 126 47016
rect 1176 46918 1204 46946
rect 234 46842 318 46870
rect 1176 46792 1204 46820
rect 536 46722 618 46750
rect 536 45530 618 45558
rect 1176 45460 1204 45488
rect 234 45410 318 45438
rect 1176 45334 1204 45362
rect 56 45264 126 45292
rect 1176 45108 1204 45136
rect 1176 44068 1204 44096
rect 56 43912 126 43940
rect 1176 43842 1204 43870
rect 234 43766 318 43794
rect 1176 43716 1204 43744
rect 536 43646 618 43674
rect 536 42454 618 42482
rect 1176 42384 1204 42412
rect 234 42334 318 42362
rect 1176 42258 1204 42286
rect 56 42188 126 42216
rect 1176 42032 1204 42060
rect 1176 40992 1204 41020
rect 56 40836 126 40864
rect 1176 40766 1204 40794
rect 234 40690 318 40718
rect 1176 40640 1204 40668
rect 536 40570 618 40598
rect 536 39378 618 39406
rect 1176 39308 1204 39336
rect 234 39258 318 39286
rect 1176 39182 1204 39210
rect 56 39112 126 39140
rect 1176 38956 1204 38984
rect 1176 37916 1204 37944
rect 56 37760 126 37788
rect 1176 37690 1204 37718
rect 234 37614 318 37642
rect 1176 37564 1204 37592
rect 536 37494 618 37522
rect 536 36302 618 36330
rect 1176 36232 1204 36260
rect 234 36182 318 36210
rect 1176 36106 1204 36134
rect 56 36036 126 36064
rect 1176 35880 1204 35908
rect 1176 34840 1204 34868
rect 56 34684 126 34712
rect 1176 34614 1204 34642
rect 234 34538 318 34566
rect 1176 34488 1204 34516
rect 536 34418 618 34446
rect 536 33226 618 33254
rect 1176 33156 1204 33184
rect 234 33106 318 33134
rect 1176 33030 1204 33058
rect 56 32960 126 32988
rect 1176 32804 1204 32832
rect 1176 31764 1204 31792
rect 56 31608 126 31636
rect 1176 31538 1204 31566
rect 234 31462 318 31490
rect 1176 31412 1204 31440
rect 536 31342 618 31370
rect 536 30150 618 30178
rect 1176 30080 1204 30108
rect 234 30030 318 30058
rect 1176 29954 1204 29982
rect 56 29884 126 29912
rect 1176 29728 1204 29756
rect 1176 28688 1204 28716
rect 56 28532 126 28560
rect 1176 28462 1204 28490
rect 234 28386 318 28414
rect 1176 28336 1204 28364
rect 536 28266 618 28294
rect 536 27074 618 27102
rect 1176 27004 1204 27032
rect 234 26954 318 26982
rect 1176 26878 1204 26906
rect 56 26808 126 26836
rect 1176 26652 1204 26680
rect 1176 25612 1204 25640
rect 56 25456 126 25484
rect 1176 25386 1204 25414
rect 234 25310 318 25338
rect 1176 25260 1204 25288
rect 536 25190 618 25218
rect 536 23998 618 24026
rect 1176 23928 1204 23956
rect 234 23878 318 23906
rect 1176 23802 1204 23830
rect 56 23732 126 23760
rect 1176 23576 1204 23604
rect 1176 22536 1204 22564
rect 56 22380 126 22408
rect 1176 22310 1204 22338
rect 234 22234 318 22262
rect 1176 22184 1204 22212
rect 536 22114 618 22142
rect 536 20922 618 20950
rect 1176 20852 1204 20880
rect 234 20802 318 20830
rect 1176 20726 1204 20754
rect 56 20656 126 20684
rect 1176 20500 1204 20528
rect 1176 19460 1204 19488
rect 56 19304 126 19332
rect 1176 19234 1204 19262
rect 234 19158 318 19186
rect 1176 19108 1204 19136
rect 536 19038 618 19066
rect 536 17846 618 17874
rect 1176 17776 1204 17804
rect 234 17726 318 17754
rect 1176 17650 1204 17678
rect 56 17580 126 17608
rect 1176 17424 1204 17452
rect 1176 16384 1204 16412
rect 56 16228 126 16256
rect 1176 16158 1204 16186
rect 234 16082 318 16110
rect 1176 16032 1204 16060
rect 536 15962 618 15990
rect 536 14770 618 14798
rect 1176 14700 1204 14728
rect 234 14650 318 14678
rect 1176 14574 1204 14602
rect 56 14504 126 14532
rect 1176 14348 1204 14376
rect 1176 13308 1204 13336
rect 56 13152 126 13180
rect 1176 13082 1204 13110
rect 234 13006 318 13034
rect 1176 12956 1204 12984
rect 536 12886 618 12914
rect 536 11694 618 11722
rect 1176 11624 1204 11652
rect 234 11574 318 11602
rect 1176 11498 1204 11526
rect 56 11428 126 11456
rect 1176 11272 1204 11300
rect 1176 10232 1204 10260
rect 56 10076 126 10104
rect 1176 10006 1204 10034
rect 234 9930 318 9958
rect 1176 9880 1204 9908
rect 536 9810 618 9838
rect 536 8618 618 8646
rect 1176 8548 1204 8576
rect 234 8498 318 8526
rect 1176 8422 1204 8450
rect 56 8352 126 8380
rect 1176 8196 1204 8224
rect 1176 7156 1204 7184
rect 56 7000 126 7028
rect 1176 6930 1204 6958
rect 234 6854 318 6882
rect 1176 6804 1204 6832
rect 536 6734 618 6762
rect 536 5542 618 5570
rect 1176 5472 1204 5500
rect 234 5422 318 5450
rect 1176 5346 1204 5374
rect 56 5276 126 5304
rect 1176 5120 1204 5148
rect 1176 4080 1204 4108
rect 56 3924 126 3952
rect 1176 3854 1204 3882
rect 234 3778 318 3806
rect 1176 3728 1204 3756
rect 536 3658 618 3686
rect 536 2466 618 2494
rect 1176 2396 1204 2424
rect 234 2346 318 2374
rect 1176 2270 1204 2298
rect 56 2200 126 2228
rect 1176 2044 1204 2072
rect 1176 1004 1204 1032
rect 56 848 126 876
rect 1176 778 1204 806
rect 234 702 318 730
rect 1176 652 1204 680
rect 536 582 618 610
<< via1 >>
rect 1178 49190 1230 49242
rect 1178 47652 1230 47704
rect 1178 46114 1230 46166
rect 1178 44576 1230 44628
rect 1178 43038 1230 43090
rect 1178 41500 1230 41552
rect 1178 39962 1230 40014
rect 1178 38424 1230 38476
rect 1178 36886 1230 36938
rect 1178 35348 1230 35400
rect 1178 33810 1230 33862
rect 1178 32272 1230 32324
rect 1178 30734 1230 30786
rect 1178 29196 1230 29248
rect 1178 27658 1230 27710
rect 1178 26120 1230 26172
rect 1178 24582 1230 24634
rect 1178 23044 1230 23096
rect 1178 21506 1230 21558
rect 1178 19968 1230 20020
rect 1178 18430 1230 18482
rect 1178 16892 1230 16944
rect 1178 15354 1230 15406
rect 1178 13816 1230 13868
rect 1178 12278 1230 12330
rect 1178 10740 1230 10792
rect 1178 9202 1230 9254
rect 1178 7664 1230 7716
rect 1178 6126 1230 6178
rect 1178 4588 1230 4640
rect 1178 3050 1230 3102
rect 1178 1512 1230 1564
rect 1178 -26 1230 26
<< metal2 >>
rect 1184 49244 1224 49250
rect 0 0 28 49216
rect 1184 49182 1224 49188
rect 192 48508 220 48536
rect 1184 47706 1224 47712
rect 1184 47644 1224 47650
rect 192 46820 220 46848
rect 1184 46168 1224 46174
rect 1184 46106 1224 46112
rect 192 45432 220 45460
rect 1184 44630 1224 44636
rect 1184 44568 1224 44574
rect 192 43744 220 43772
rect 1184 43092 1224 43098
rect 1184 43030 1224 43036
rect 192 42356 220 42384
rect 1184 41554 1224 41560
rect 1184 41492 1224 41498
rect 192 40668 220 40696
rect 1184 40016 1224 40022
rect 1184 39954 1224 39960
rect 192 39280 220 39308
rect 1184 38478 1224 38484
rect 1184 38416 1224 38422
rect 192 37592 220 37620
rect 1184 36940 1224 36946
rect 1184 36878 1224 36884
rect 192 36204 220 36232
rect 1184 35402 1224 35408
rect 1184 35340 1224 35346
rect 192 34516 220 34544
rect 1184 33864 1224 33870
rect 1184 33802 1224 33808
rect 192 33128 220 33156
rect 1184 32326 1224 32332
rect 1184 32264 1224 32270
rect 192 31440 220 31468
rect 1184 30788 1224 30794
rect 1184 30726 1224 30732
rect 192 30052 220 30080
rect 1184 29250 1224 29256
rect 1184 29188 1224 29194
rect 192 28364 220 28392
rect 1184 27712 1224 27718
rect 1184 27650 1224 27656
rect 192 26976 220 27004
rect 1184 26174 1224 26180
rect 1184 26112 1224 26118
rect 192 25288 220 25316
rect 1184 24636 1224 24642
rect 1184 24574 1224 24580
rect 192 23900 220 23928
rect 1184 23098 1224 23104
rect 1184 23036 1224 23042
rect 192 22212 220 22240
rect 1184 21560 1224 21566
rect 1184 21498 1224 21504
rect 192 20824 220 20852
rect 1184 20022 1224 20028
rect 1184 19960 1224 19966
rect 192 19136 220 19164
rect 1184 18484 1224 18490
rect 1184 18422 1224 18428
rect 192 17748 220 17776
rect 1184 16946 1224 16952
rect 1184 16884 1224 16890
rect 192 16060 220 16088
rect 1184 15408 1224 15414
rect 1184 15346 1224 15352
rect 192 14672 220 14700
rect 1184 13870 1224 13876
rect 1184 13808 1224 13814
rect 192 12984 220 13012
rect 1184 12332 1224 12338
rect 1184 12270 1224 12276
rect 192 11596 220 11624
rect 1184 10794 1224 10800
rect 1184 10732 1224 10738
rect 192 9908 220 9936
rect 1184 9256 1224 9262
rect 1184 9194 1224 9200
rect 192 8520 220 8548
rect 1184 7718 1224 7724
rect 1184 7656 1224 7662
rect 192 6832 220 6860
rect 1184 6180 1224 6186
rect 1184 6118 1224 6124
rect 192 5444 220 5472
rect 1184 4642 1224 4648
rect 1184 4580 1224 4586
rect 192 3756 220 3784
rect 1184 3104 1224 3110
rect 1184 3042 1224 3048
rect 192 2368 220 2396
rect 1184 1566 1224 1572
rect 1184 1504 1224 1510
rect 192 680 220 708
rect 1184 28 1224 34
rect 1184 -34 1224 -28
<< via2 >>
rect 1176 49242 1232 49244
rect 1176 49190 1178 49242
rect 1178 49190 1230 49242
rect 1230 49190 1232 49242
rect 1176 49188 1232 49190
rect 1176 47704 1232 47706
rect 1176 47652 1178 47704
rect 1178 47652 1230 47704
rect 1230 47652 1232 47704
rect 1176 47650 1232 47652
rect 1176 46166 1232 46168
rect 1176 46114 1178 46166
rect 1178 46114 1230 46166
rect 1230 46114 1232 46166
rect 1176 46112 1232 46114
rect 1176 44628 1232 44630
rect 1176 44576 1178 44628
rect 1178 44576 1230 44628
rect 1230 44576 1232 44628
rect 1176 44574 1232 44576
rect 1176 43090 1232 43092
rect 1176 43038 1178 43090
rect 1178 43038 1230 43090
rect 1230 43038 1232 43090
rect 1176 43036 1232 43038
rect 1176 41552 1232 41554
rect 1176 41500 1178 41552
rect 1178 41500 1230 41552
rect 1230 41500 1232 41552
rect 1176 41498 1232 41500
rect 1176 40014 1232 40016
rect 1176 39962 1178 40014
rect 1178 39962 1230 40014
rect 1230 39962 1232 40014
rect 1176 39960 1232 39962
rect 1176 38476 1232 38478
rect 1176 38424 1178 38476
rect 1178 38424 1230 38476
rect 1230 38424 1232 38476
rect 1176 38422 1232 38424
rect 1176 36938 1232 36940
rect 1176 36886 1178 36938
rect 1178 36886 1230 36938
rect 1230 36886 1232 36938
rect 1176 36884 1232 36886
rect 1176 35400 1232 35402
rect 1176 35348 1178 35400
rect 1178 35348 1230 35400
rect 1230 35348 1232 35400
rect 1176 35346 1232 35348
rect 1176 33862 1232 33864
rect 1176 33810 1178 33862
rect 1178 33810 1230 33862
rect 1230 33810 1232 33862
rect 1176 33808 1232 33810
rect 1176 32324 1232 32326
rect 1176 32272 1178 32324
rect 1178 32272 1230 32324
rect 1230 32272 1232 32324
rect 1176 32270 1232 32272
rect 1176 30786 1232 30788
rect 1176 30734 1178 30786
rect 1178 30734 1230 30786
rect 1230 30734 1232 30786
rect 1176 30732 1232 30734
rect 1176 29248 1232 29250
rect 1176 29196 1178 29248
rect 1178 29196 1230 29248
rect 1230 29196 1232 29248
rect 1176 29194 1232 29196
rect 1176 27710 1232 27712
rect 1176 27658 1178 27710
rect 1178 27658 1230 27710
rect 1230 27658 1232 27710
rect 1176 27656 1232 27658
rect 1176 26172 1232 26174
rect 1176 26120 1178 26172
rect 1178 26120 1230 26172
rect 1230 26120 1232 26172
rect 1176 26118 1232 26120
rect 1176 24634 1232 24636
rect 1176 24582 1178 24634
rect 1178 24582 1230 24634
rect 1230 24582 1232 24634
rect 1176 24580 1232 24582
rect 1176 23096 1232 23098
rect 1176 23044 1178 23096
rect 1178 23044 1230 23096
rect 1230 23044 1232 23096
rect 1176 23042 1232 23044
rect 1176 21558 1232 21560
rect 1176 21506 1178 21558
rect 1178 21506 1230 21558
rect 1230 21506 1232 21558
rect 1176 21504 1232 21506
rect 1176 20020 1232 20022
rect 1176 19968 1178 20020
rect 1178 19968 1230 20020
rect 1230 19968 1232 20020
rect 1176 19966 1232 19968
rect 1176 18482 1232 18484
rect 1176 18430 1178 18482
rect 1178 18430 1230 18482
rect 1230 18430 1232 18482
rect 1176 18428 1232 18430
rect 1176 16944 1232 16946
rect 1176 16892 1178 16944
rect 1178 16892 1230 16944
rect 1230 16892 1232 16944
rect 1176 16890 1232 16892
rect 1176 15406 1232 15408
rect 1176 15354 1178 15406
rect 1178 15354 1230 15406
rect 1230 15354 1232 15406
rect 1176 15352 1232 15354
rect 1176 13868 1232 13870
rect 1176 13816 1178 13868
rect 1178 13816 1230 13868
rect 1230 13816 1232 13868
rect 1176 13814 1232 13816
rect 1176 12330 1232 12332
rect 1176 12278 1178 12330
rect 1178 12278 1230 12330
rect 1230 12278 1232 12330
rect 1176 12276 1232 12278
rect 1176 10792 1232 10794
rect 1176 10740 1178 10792
rect 1178 10740 1230 10792
rect 1230 10740 1232 10792
rect 1176 10738 1232 10740
rect 1176 9254 1232 9256
rect 1176 9202 1178 9254
rect 1178 9202 1230 9254
rect 1230 9202 1232 9254
rect 1176 9200 1232 9202
rect 1176 7716 1232 7718
rect 1176 7664 1178 7716
rect 1178 7664 1230 7716
rect 1230 7664 1232 7716
rect 1176 7662 1232 7664
rect 1176 6178 1232 6180
rect 1176 6126 1178 6178
rect 1178 6126 1230 6178
rect 1230 6126 1232 6178
rect 1176 6124 1232 6126
rect 1176 4640 1232 4642
rect 1176 4588 1178 4640
rect 1178 4588 1230 4640
rect 1230 4588 1232 4640
rect 1176 4586 1232 4588
rect 1176 3102 1232 3104
rect 1176 3050 1178 3102
rect 1178 3050 1230 3102
rect 1230 3050 1232 3102
rect 1176 3048 1232 3050
rect 1176 1564 1232 1566
rect 1176 1512 1178 1564
rect 1178 1512 1230 1564
rect 1230 1512 1232 1564
rect 1176 1510 1232 1512
rect 1176 26 1232 28
rect 1176 -26 1178 26
rect 1178 -26 1230 26
rect 1230 -26 1232 26
rect 1176 -28 1232 -26
<< metal3 >>
rect 1138 49244 1270 49249
rect 1138 49188 1176 49244
rect 1232 49188 1270 49244
rect 1138 49183 1270 49188
rect 1138 47706 1270 47711
rect 1138 47650 1176 47706
rect 1232 47650 1270 47706
rect 1138 47645 1270 47650
rect 1138 46168 1270 46173
rect 1138 46112 1176 46168
rect 1232 46112 1270 46168
rect 1138 46107 1270 46112
rect 1138 44630 1270 44635
rect 1138 44574 1176 44630
rect 1232 44574 1270 44630
rect 1138 44569 1270 44574
rect 1138 43092 1270 43097
rect 1138 43036 1176 43092
rect 1232 43036 1270 43092
rect 1138 43031 1270 43036
rect 1138 41554 1270 41559
rect 1138 41498 1176 41554
rect 1232 41498 1270 41554
rect 1138 41493 1270 41498
rect 1138 40016 1270 40021
rect 1138 39960 1176 40016
rect 1232 39960 1270 40016
rect 1138 39955 1270 39960
rect 1138 38478 1270 38483
rect 1138 38422 1176 38478
rect 1232 38422 1270 38478
rect 1138 38417 1270 38422
rect 1138 36940 1270 36945
rect 1138 36884 1176 36940
rect 1232 36884 1270 36940
rect 1138 36879 1270 36884
rect 1138 35402 1270 35407
rect 1138 35346 1176 35402
rect 1232 35346 1270 35402
rect 1138 35341 1270 35346
rect 1138 33864 1270 33869
rect 1138 33808 1176 33864
rect 1232 33808 1270 33864
rect 1138 33803 1270 33808
rect 1138 32326 1270 32331
rect 1138 32270 1176 32326
rect 1232 32270 1270 32326
rect 1138 32265 1270 32270
rect 1138 30788 1270 30793
rect 1138 30732 1176 30788
rect 1232 30732 1270 30788
rect 1138 30727 1270 30732
rect 1138 29250 1270 29255
rect 1138 29194 1176 29250
rect 1232 29194 1270 29250
rect 1138 29189 1270 29194
rect 1138 27712 1270 27717
rect 1138 27656 1176 27712
rect 1232 27656 1270 27712
rect 1138 27651 1270 27656
rect 1138 26174 1270 26179
rect 1138 26118 1176 26174
rect 1232 26118 1270 26174
rect 1138 26113 1270 26118
rect 1138 24636 1270 24641
rect 1138 24580 1176 24636
rect 1232 24580 1270 24636
rect 1138 24575 1270 24580
rect 1138 23098 1270 23103
rect 1138 23042 1176 23098
rect 1232 23042 1270 23098
rect 1138 23037 1270 23042
rect 1138 21560 1270 21565
rect 1138 21504 1176 21560
rect 1232 21504 1270 21560
rect 1138 21499 1270 21504
rect 1138 20022 1270 20027
rect 1138 19966 1176 20022
rect 1232 19966 1270 20022
rect 1138 19961 1270 19966
rect 1138 18484 1270 18489
rect 1138 18428 1176 18484
rect 1232 18428 1270 18484
rect 1138 18423 1270 18428
rect 1138 16946 1270 16951
rect 1138 16890 1176 16946
rect 1232 16890 1270 16946
rect 1138 16885 1270 16890
rect 1138 15408 1270 15413
rect 1138 15352 1176 15408
rect 1232 15352 1270 15408
rect 1138 15347 1270 15352
rect 1138 13870 1270 13875
rect 1138 13814 1176 13870
rect 1232 13814 1270 13870
rect 1138 13809 1270 13814
rect 1138 12332 1270 12337
rect 1138 12276 1176 12332
rect 1232 12276 1270 12332
rect 1138 12271 1270 12276
rect 1138 10794 1270 10799
rect 1138 10738 1176 10794
rect 1232 10738 1270 10794
rect 1138 10733 1270 10738
rect 1138 9256 1270 9261
rect 1138 9200 1176 9256
rect 1232 9200 1270 9256
rect 1138 9195 1270 9200
rect 1138 7718 1270 7723
rect 1138 7662 1176 7718
rect 1232 7662 1270 7718
rect 1138 7657 1270 7662
rect 1138 6180 1270 6185
rect 1138 6124 1176 6180
rect 1232 6124 1270 6180
rect 1138 6119 1270 6124
rect 1138 4642 1270 4647
rect 1138 4586 1176 4642
rect 1232 4586 1270 4642
rect 1138 4581 1270 4586
rect 1138 3104 1270 3109
rect 1138 3048 1176 3104
rect 1232 3048 1270 3104
rect 1138 3043 1270 3048
rect 1138 1566 1270 1571
rect 1138 1510 1176 1566
rect 1232 1510 1270 1566
rect 1138 1505 1270 1510
rect 1138 28 1270 33
rect 1138 -28 1176 28
rect 1232 -28 1270 28
rect 1138 -33 1270 -28
use contact_18  contact_18_0
timestamp 1643678851
transform 1 0 1138 0 1 49183
box 0 0 1 1
use contact_17  contact_17_0
timestamp 1643678851
transform 1 0 1189 0 1 49201
box 0 0 1 1
use contact_18  contact_18_1
timestamp 1643678851
transform 1 0 1138 0 1 47645
box 0 0 1 1
use contact_17  contact_17_1
timestamp 1643678851
transform 1 0 1189 0 1 47663
box 0 0 1 1
use contact_18  contact_18_2
timestamp 1643678851
transform 1 0 1138 0 1 46107
box 0 0 1 1
use contact_17  contact_17_2
timestamp 1643678851
transform 1 0 1189 0 1 46125
box 0 0 1 1
use contact_18  contact_18_3
timestamp 1643678851
transform 1 0 1138 0 1 47645
box 0 0 1 1
use contact_17  contact_17_3
timestamp 1643678851
transform 1 0 1189 0 1 47663
box 0 0 1 1
use contact_18  contact_18_4
timestamp 1643678851
transform 1 0 1138 0 1 46107
box 0 0 1 1
use contact_17  contact_17_4
timestamp 1643678851
transform 1 0 1189 0 1 46125
box 0 0 1 1
use contact_18  contact_18_5
timestamp 1643678851
transform 1 0 1138 0 1 44569
box 0 0 1 1
use contact_17  contact_17_5
timestamp 1643678851
transform 1 0 1189 0 1 44587
box 0 0 1 1
use contact_18  contact_18_6
timestamp 1643678851
transform 1 0 1138 0 1 43031
box 0 0 1 1
use contact_17  contact_17_6
timestamp 1643678851
transform 1 0 1189 0 1 43049
box 0 0 1 1
use contact_18  contact_18_7
timestamp 1643678851
transform 1 0 1138 0 1 44569
box 0 0 1 1
use contact_17  contact_17_7
timestamp 1643678851
transform 1 0 1189 0 1 44587
box 0 0 1 1
use contact_18  contact_18_8
timestamp 1643678851
transform 1 0 1138 0 1 43031
box 0 0 1 1
use contact_17  contact_17_8
timestamp 1643678851
transform 1 0 1189 0 1 43049
box 0 0 1 1
use contact_18  contact_18_9
timestamp 1643678851
transform 1 0 1138 0 1 41493
box 0 0 1 1
use contact_17  contact_17_9
timestamp 1643678851
transform 1 0 1189 0 1 41511
box 0 0 1 1
use contact_18  contact_18_10
timestamp 1643678851
transform 1 0 1138 0 1 39955
box 0 0 1 1
use contact_17  contact_17_10
timestamp 1643678851
transform 1 0 1189 0 1 39973
box 0 0 1 1
use contact_18  contact_18_11
timestamp 1643678851
transform 1 0 1138 0 1 41493
box 0 0 1 1
use contact_17  contact_17_11
timestamp 1643678851
transform 1 0 1189 0 1 41511
box 0 0 1 1
use contact_18  contact_18_12
timestamp 1643678851
transform 1 0 1138 0 1 39955
box 0 0 1 1
use contact_17  contact_17_12
timestamp 1643678851
transform 1 0 1189 0 1 39973
box 0 0 1 1
use contact_18  contact_18_13
timestamp 1643678851
transform 1 0 1138 0 1 38417
box 0 0 1 1
use contact_17  contact_17_13
timestamp 1643678851
transform 1 0 1189 0 1 38435
box 0 0 1 1
use contact_18  contact_18_14
timestamp 1643678851
transform 1 0 1138 0 1 36879
box 0 0 1 1
use contact_17  contact_17_14
timestamp 1643678851
transform 1 0 1189 0 1 36897
box 0 0 1 1
use contact_18  contact_18_15
timestamp 1643678851
transform 1 0 1138 0 1 38417
box 0 0 1 1
use contact_17  contact_17_15
timestamp 1643678851
transform 1 0 1189 0 1 38435
box 0 0 1 1
use contact_18  contact_18_16
timestamp 1643678851
transform 1 0 1138 0 1 36879
box 0 0 1 1
use contact_17  contact_17_16
timestamp 1643678851
transform 1 0 1189 0 1 36897
box 0 0 1 1
use contact_18  contact_18_17
timestamp 1643678851
transform 1 0 1138 0 1 35341
box 0 0 1 1
use contact_17  contact_17_17
timestamp 1643678851
transform 1 0 1189 0 1 35359
box 0 0 1 1
use contact_18  contact_18_18
timestamp 1643678851
transform 1 0 1138 0 1 33803
box 0 0 1 1
use contact_17  contact_17_18
timestamp 1643678851
transform 1 0 1189 0 1 33821
box 0 0 1 1
use contact_18  contact_18_19
timestamp 1643678851
transform 1 0 1138 0 1 35341
box 0 0 1 1
use contact_17  contact_17_19
timestamp 1643678851
transform 1 0 1189 0 1 35359
box 0 0 1 1
use contact_18  contact_18_20
timestamp 1643678851
transform 1 0 1138 0 1 33803
box 0 0 1 1
use contact_17  contact_17_20
timestamp 1643678851
transform 1 0 1189 0 1 33821
box 0 0 1 1
use contact_18  contact_18_21
timestamp 1643678851
transform 1 0 1138 0 1 32265
box 0 0 1 1
use contact_17  contact_17_21
timestamp 1643678851
transform 1 0 1189 0 1 32283
box 0 0 1 1
use contact_18  contact_18_22
timestamp 1643678851
transform 1 0 1138 0 1 30727
box 0 0 1 1
use contact_17  contact_17_22
timestamp 1643678851
transform 1 0 1189 0 1 30745
box 0 0 1 1
use contact_18  contact_18_23
timestamp 1643678851
transform 1 0 1138 0 1 32265
box 0 0 1 1
use contact_17  contact_17_23
timestamp 1643678851
transform 1 0 1189 0 1 32283
box 0 0 1 1
use contact_18  contact_18_24
timestamp 1643678851
transform 1 0 1138 0 1 30727
box 0 0 1 1
use contact_17  contact_17_24
timestamp 1643678851
transform 1 0 1189 0 1 30745
box 0 0 1 1
use contact_18  contact_18_25
timestamp 1643678851
transform 1 0 1138 0 1 29189
box 0 0 1 1
use contact_17  contact_17_25
timestamp 1643678851
transform 1 0 1189 0 1 29207
box 0 0 1 1
use contact_18  contact_18_26
timestamp 1643678851
transform 1 0 1138 0 1 27651
box 0 0 1 1
use contact_17  contact_17_26
timestamp 1643678851
transform 1 0 1189 0 1 27669
box 0 0 1 1
use contact_18  contact_18_27
timestamp 1643678851
transform 1 0 1138 0 1 29189
box 0 0 1 1
use contact_17  contact_17_27
timestamp 1643678851
transform 1 0 1189 0 1 29207
box 0 0 1 1
use contact_18  contact_18_28
timestamp 1643678851
transform 1 0 1138 0 1 27651
box 0 0 1 1
use contact_17  contact_17_28
timestamp 1643678851
transform 1 0 1189 0 1 27669
box 0 0 1 1
use contact_18  contact_18_29
timestamp 1643678851
transform 1 0 1138 0 1 26113
box 0 0 1 1
use contact_17  contact_17_29
timestamp 1643678851
transform 1 0 1189 0 1 26131
box 0 0 1 1
use contact_18  contact_18_30
timestamp 1643678851
transform 1 0 1138 0 1 24575
box 0 0 1 1
use contact_17  contact_17_30
timestamp 1643678851
transform 1 0 1189 0 1 24593
box 0 0 1 1
use contact_18  contact_18_31
timestamp 1643678851
transform 1 0 1138 0 1 26113
box 0 0 1 1
use contact_17  contact_17_31
timestamp 1643678851
transform 1 0 1189 0 1 26131
box 0 0 1 1
use contact_18  contact_18_32
timestamp 1643678851
transform 1 0 1138 0 1 24575
box 0 0 1 1
use contact_17  contact_17_32
timestamp 1643678851
transform 1 0 1189 0 1 24593
box 0 0 1 1
use contact_18  contact_18_33
timestamp 1643678851
transform 1 0 1138 0 1 23037
box 0 0 1 1
use contact_17  contact_17_33
timestamp 1643678851
transform 1 0 1189 0 1 23055
box 0 0 1 1
use contact_18  contact_18_34
timestamp 1643678851
transform 1 0 1138 0 1 21499
box 0 0 1 1
use contact_17  contact_17_34
timestamp 1643678851
transform 1 0 1189 0 1 21517
box 0 0 1 1
use contact_18  contact_18_35
timestamp 1643678851
transform 1 0 1138 0 1 23037
box 0 0 1 1
use contact_17  contact_17_35
timestamp 1643678851
transform 1 0 1189 0 1 23055
box 0 0 1 1
use contact_18  contact_18_36
timestamp 1643678851
transform 1 0 1138 0 1 21499
box 0 0 1 1
use contact_17  contact_17_36
timestamp 1643678851
transform 1 0 1189 0 1 21517
box 0 0 1 1
use contact_18  contact_18_37
timestamp 1643678851
transform 1 0 1138 0 1 19961
box 0 0 1 1
use contact_17  contact_17_37
timestamp 1643678851
transform 1 0 1189 0 1 19979
box 0 0 1 1
use contact_18  contact_18_38
timestamp 1643678851
transform 1 0 1138 0 1 18423
box 0 0 1 1
use contact_17  contact_17_38
timestamp 1643678851
transform 1 0 1189 0 1 18441
box 0 0 1 1
use contact_18  contact_18_39
timestamp 1643678851
transform 1 0 1138 0 1 19961
box 0 0 1 1
use contact_17  contact_17_39
timestamp 1643678851
transform 1 0 1189 0 1 19979
box 0 0 1 1
use contact_18  contact_18_40
timestamp 1643678851
transform 1 0 1138 0 1 18423
box 0 0 1 1
use contact_17  contact_17_40
timestamp 1643678851
transform 1 0 1189 0 1 18441
box 0 0 1 1
use contact_18  contact_18_41
timestamp 1643678851
transform 1 0 1138 0 1 16885
box 0 0 1 1
use contact_17  contact_17_41
timestamp 1643678851
transform 1 0 1189 0 1 16903
box 0 0 1 1
use contact_18  contact_18_42
timestamp 1643678851
transform 1 0 1138 0 1 15347
box 0 0 1 1
use contact_17  contact_17_42
timestamp 1643678851
transform 1 0 1189 0 1 15365
box 0 0 1 1
use contact_18  contact_18_43
timestamp 1643678851
transform 1 0 1138 0 1 16885
box 0 0 1 1
use contact_17  contact_17_43
timestamp 1643678851
transform 1 0 1189 0 1 16903
box 0 0 1 1
use contact_18  contact_18_44
timestamp 1643678851
transform 1 0 1138 0 1 15347
box 0 0 1 1
use contact_17  contact_17_44
timestamp 1643678851
transform 1 0 1189 0 1 15365
box 0 0 1 1
use contact_18  contact_18_45
timestamp 1643678851
transform 1 0 1138 0 1 13809
box 0 0 1 1
use contact_17  contact_17_45
timestamp 1643678851
transform 1 0 1189 0 1 13827
box 0 0 1 1
use contact_18  contact_18_46
timestamp 1643678851
transform 1 0 1138 0 1 12271
box 0 0 1 1
use contact_17  contact_17_46
timestamp 1643678851
transform 1 0 1189 0 1 12289
box 0 0 1 1
use contact_18  contact_18_47
timestamp 1643678851
transform 1 0 1138 0 1 13809
box 0 0 1 1
use contact_17  contact_17_47
timestamp 1643678851
transform 1 0 1189 0 1 13827
box 0 0 1 1
use contact_18  contact_18_48
timestamp 1643678851
transform 1 0 1138 0 1 12271
box 0 0 1 1
use contact_17  contact_17_48
timestamp 1643678851
transform 1 0 1189 0 1 12289
box 0 0 1 1
use contact_18  contact_18_49
timestamp 1643678851
transform 1 0 1138 0 1 10733
box 0 0 1 1
use contact_17  contact_17_49
timestamp 1643678851
transform 1 0 1189 0 1 10751
box 0 0 1 1
use contact_18  contact_18_50
timestamp 1643678851
transform 1 0 1138 0 1 9195
box 0 0 1 1
use contact_17  contact_17_50
timestamp 1643678851
transform 1 0 1189 0 1 9213
box 0 0 1 1
use contact_18  contact_18_51
timestamp 1643678851
transform 1 0 1138 0 1 10733
box 0 0 1 1
use contact_17  contact_17_51
timestamp 1643678851
transform 1 0 1189 0 1 10751
box 0 0 1 1
use contact_18  contact_18_52
timestamp 1643678851
transform 1 0 1138 0 1 9195
box 0 0 1 1
use contact_17  contact_17_52
timestamp 1643678851
transform 1 0 1189 0 1 9213
box 0 0 1 1
use contact_18  contact_18_53
timestamp 1643678851
transform 1 0 1138 0 1 7657
box 0 0 1 1
use contact_17  contact_17_53
timestamp 1643678851
transform 1 0 1189 0 1 7675
box 0 0 1 1
use contact_18  contact_18_54
timestamp 1643678851
transform 1 0 1138 0 1 6119
box 0 0 1 1
use contact_17  contact_17_54
timestamp 1643678851
transform 1 0 1189 0 1 6137
box 0 0 1 1
use contact_18  contact_18_55
timestamp 1643678851
transform 1 0 1138 0 1 7657
box 0 0 1 1
use contact_17  contact_17_55
timestamp 1643678851
transform 1 0 1189 0 1 7675
box 0 0 1 1
use contact_18  contact_18_56
timestamp 1643678851
transform 1 0 1138 0 1 6119
box 0 0 1 1
use contact_17  contact_17_56
timestamp 1643678851
transform 1 0 1189 0 1 6137
box 0 0 1 1
use contact_18  contact_18_57
timestamp 1643678851
transform 1 0 1138 0 1 4581
box 0 0 1 1
use contact_17  contact_17_57
timestamp 1643678851
transform 1 0 1189 0 1 4599
box 0 0 1 1
use contact_18  contact_18_58
timestamp 1643678851
transform 1 0 1138 0 1 3043
box 0 0 1 1
use contact_17  contact_17_58
timestamp 1643678851
transform 1 0 1189 0 1 3061
box 0 0 1 1
use contact_18  contact_18_59
timestamp 1643678851
transform 1 0 1138 0 1 4581
box 0 0 1 1
use contact_17  contact_17_59
timestamp 1643678851
transform 1 0 1189 0 1 4599
box 0 0 1 1
use contact_18  contact_18_60
timestamp 1643678851
transform 1 0 1138 0 1 3043
box 0 0 1 1
use contact_17  contact_17_60
timestamp 1643678851
transform 1 0 1189 0 1 3061
box 0 0 1 1
use contact_18  contact_18_61
timestamp 1643678851
transform 1 0 1138 0 1 1505
box 0 0 1 1
use contact_17  contact_17_61
timestamp 1643678851
transform 1 0 1189 0 1 1523
box 0 0 1 1
use contact_18  contact_18_62
timestamp 1643678851
transform 1 0 1138 0 1 -33
box 0 0 1 1
use contact_17  contact_17_62
timestamp 1643678851
transform 1 0 1189 0 1 -15
box 0 0 1 1
use contact_18  contact_18_63
timestamp 1643678851
transform 1 0 1138 0 1 1505
box 0 0 1 1
use contact_17  contact_17_63
timestamp 1643678851
transform 1 0 1189 0 1 1523
box 0 0 1 1
use wordline_driver_cell  wordline_driver_cell_0
timestamp 1643678851
transform 1 0 0 0 -1 49216
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_1
timestamp 1643678851
transform 1 0 0 0 1 46140
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_2
timestamp 1643678851
transform 1 0 0 0 -1 46140
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_3
timestamp 1643678851
transform 1 0 0 0 1 43064
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_4
timestamp 1643678851
transform 1 0 0 0 -1 43064
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_5
timestamp 1643678851
transform 1 0 0 0 1 39988
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_6
timestamp 1643678851
transform 1 0 0 0 -1 39988
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_7
timestamp 1643678851
transform 1 0 0 0 1 36912
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_8
timestamp 1643678851
transform 1 0 0 0 -1 36912
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_9
timestamp 1643678851
transform 1 0 0 0 1 33836
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_10
timestamp 1643678851
transform 1 0 0 0 -1 33836
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_11
timestamp 1643678851
transform 1 0 0 0 1 30760
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_12
timestamp 1643678851
transform 1 0 0 0 -1 30760
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_13
timestamp 1643678851
transform 1 0 0 0 1 27684
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_14
timestamp 1643678851
transform 1 0 0 0 -1 27684
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_15
timestamp 1643678851
transform 1 0 0 0 1 24608
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_16
timestamp 1643678851
transform 1 0 0 0 -1 24608
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_17
timestamp 1643678851
transform 1 0 0 0 1 21532
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_18
timestamp 1643678851
transform 1 0 0 0 -1 21532
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_19
timestamp 1643678851
transform 1 0 0 0 1 18456
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_20
timestamp 1643678851
transform 1 0 0 0 -1 18456
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_21
timestamp 1643678851
transform 1 0 0 0 1 15380
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_22
timestamp 1643678851
transform 1 0 0 0 -1 15380
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_23
timestamp 1643678851
transform 1 0 0 0 1 12304
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_24
timestamp 1643678851
transform 1 0 0 0 -1 12304
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_25
timestamp 1643678851
transform 1 0 0 0 1 9228
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_26
timestamp 1643678851
transform 1 0 0 0 -1 9228
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_27
timestamp 1643678851
transform 1 0 0 0 1 6152
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_28
timestamp 1643678851
transform 1 0 0 0 -1 6152
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_29
timestamp 1643678851
transform 1 0 0 0 1 3076
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_30
timestamp 1643678851
transform 1 0 0 0 -1 3076
box 0 -42 1204 1616
use wordline_driver_cell  wordline_driver_cell_31
timestamp 1643678851
transform 1 0 0 0 1 0
box 0 -42 1204 1616
<< labels >>
rlabel metal2 s 0 0 28 49216 4 wl_en
rlabel metal1 s 56 848 126 876 4 in0_0
rlabel metal1 s 234 702 318 730 4 in1_0
rlabel metal1 s 536 582 618 610 4 in2_0
rlabel metal1 s 1176 778 1204 806 4 rwl0_0
rlabel metal1 s 1176 1004 1204 1032 4 rwl1_0
rlabel metal1 s 1176 652 1204 680 4 wwl0_0
rlabel metal1 s 56 2200 126 2228 4 in0_1
rlabel metal1 s 234 2346 318 2374 4 in1_1
rlabel metal1 s 536 2466 618 2494 4 in2_1
rlabel metal1 s 1176 2270 1204 2298 4 rwl0_1
rlabel metal1 s 1176 2044 1204 2072 4 rwl1_1
rlabel metal1 s 1176 2396 1204 2424 4 wwl0_1
rlabel metal1 s 56 3924 126 3952 4 in0_2
rlabel metal1 s 234 3778 318 3806 4 in1_2
rlabel metal1 s 536 3658 618 3686 4 in2_2
rlabel metal1 s 1176 3854 1204 3882 4 rwl0_2
rlabel metal1 s 1176 4080 1204 4108 4 rwl1_2
rlabel metal1 s 1176 3728 1204 3756 4 wwl0_2
rlabel metal1 s 56 5276 126 5304 4 in0_3
rlabel metal1 s 234 5422 318 5450 4 in1_3
rlabel metal1 s 536 5542 618 5570 4 in2_3
rlabel metal1 s 1176 5346 1204 5374 4 rwl0_3
rlabel metal1 s 1176 5120 1204 5148 4 rwl1_3
rlabel metal1 s 1176 5472 1204 5500 4 wwl0_3
rlabel metal1 s 56 7000 126 7028 4 in0_4
rlabel metal1 s 234 6854 318 6882 4 in1_4
rlabel metal1 s 536 6734 618 6762 4 in2_4
rlabel metal1 s 1176 6930 1204 6958 4 rwl0_4
rlabel metal1 s 1176 7156 1204 7184 4 rwl1_4
rlabel metal1 s 1176 6804 1204 6832 4 wwl0_4
rlabel metal1 s 56 8352 126 8380 4 in0_5
rlabel metal1 s 234 8498 318 8526 4 in1_5
rlabel metal1 s 536 8618 618 8646 4 in2_5
rlabel metal1 s 1176 8422 1204 8450 4 rwl0_5
rlabel metal1 s 1176 8196 1204 8224 4 rwl1_5
rlabel metal1 s 1176 8548 1204 8576 4 wwl0_5
rlabel metal1 s 56 10076 126 10104 4 in0_6
rlabel metal1 s 234 9930 318 9958 4 in1_6
rlabel metal1 s 536 9810 618 9838 4 in2_6
rlabel metal1 s 1176 10006 1204 10034 4 rwl0_6
rlabel metal1 s 1176 10232 1204 10260 4 rwl1_6
rlabel metal1 s 1176 9880 1204 9908 4 wwl0_6
rlabel metal1 s 56 11428 126 11456 4 in0_7
rlabel metal1 s 234 11574 318 11602 4 in1_7
rlabel metal1 s 536 11694 618 11722 4 in2_7
rlabel metal1 s 1176 11498 1204 11526 4 rwl0_7
rlabel metal1 s 1176 11272 1204 11300 4 rwl1_7
rlabel metal1 s 1176 11624 1204 11652 4 wwl0_7
rlabel metal1 s 56 13152 126 13180 4 in0_8
rlabel metal1 s 234 13006 318 13034 4 in1_8
rlabel metal1 s 536 12886 618 12914 4 in2_8
rlabel metal1 s 1176 13082 1204 13110 4 rwl0_8
rlabel metal1 s 1176 13308 1204 13336 4 rwl1_8
rlabel metal1 s 1176 12956 1204 12984 4 wwl0_8
rlabel metal1 s 56 14504 126 14532 4 in0_9
rlabel metal1 s 234 14650 318 14678 4 in1_9
rlabel metal1 s 536 14770 618 14798 4 in2_9
rlabel metal1 s 1176 14574 1204 14602 4 rwl0_9
rlabel metal1 s 1176 14348 1204 14376 4 rwl1_9
rlabel metal1 s 1176 14700 1204 14728 4 wwl0_9
rlabel metal1 s 56 16228 126 16256 4 in0_10
rlabel metal1 s 234 16082 318 16110 4 in1_10
rlabel metal1 s 536 15962 618 15990 4 in2_10
rlabel metal1 s 1176 16158 1204 16186 4 rwl0_10
rlabel metal1 s 1176 16384 1204 16412 4 rwl1_10
rlabel metal1 s 1176 16032 1204 16060 4 wwl0_10
rlabel metal1 s 56 17580 126 17608 4 in0_11
rlabel metal1 s 234 17726 318 17754 4 in1_11
rlabel metal1 s 536 17846 618 17874 4 in2_11
rlabel metal1 s 1176 17650 1204 17678 4 rwl0_11
rlabel metal1 s 1176 17424 1204 17452 4 rwl1_11
rlabel metal1 s 1176 17776 1204 17804 4 wwl0_11
rlabel metal1 s 56 19304 126 19332 4 in0_12
rlabel metal1 s 234 19158 318 19186 4 in1_12
rlabel metal1 s 536 19038 618 19066 4 in2_12
rlabel metal1 s 1176 19234 1204 19262 4 rwl0_12
rlabel metal1 s 1176 19460 1204 19488 4 rwl1_12
rlabel metal1 s 1176 19108 1204 19136 4 wwl0_12
rlabel metal1 s 56 20656 126 20684 4 in0_13
rlabel metal1 s 234 20802 318 20830 4 in1_13
rlabel metal1 s 536 20922 618 20950 4 in2_13
rlabel metal1 s 1176 20726 1204 20754 4 rwl0_13
rlabel metal1 s 1176 20500 1204 20528 4 rwl1_13
rlabel metal1 s 1176 20852 1204 20880 4 wwl0_13
rlabel metal1 s 56 22380 126 22408 4 in0_14
rlabel metal1 s 234 22234 318 22262 4 in1_14
rlabel metal1 s 536 22114 618 22142 4 in2_14
rlabel metal1 s 1176 22310 1204 22338 4 rwl0_14
rlabel metal1 s 1176 22536 1204 22564 4 rwl1_14
rlabel metal1 s 1176 22184 1204 22212 4 wwl0_14
rlabel metal1 s 56 23732 126 23760 4 in0_15
rlabel metal1 s 234 23878 318 23906 4 in1_15
rlabel metal1 s 536 23998 618 24026 4 in2_15
rlabel metal1 s 1176 23802 1204 23830 4 rwl0_15
rlabel metal1 s 1176 23576 1204 23604 4 rwl1_15
rlabel metal1 s 1176 23928 1204 23956 4 wwl0_15
rlabel metal1 s 56 25456 126 25484 4 in0_16
rlabel metal1 s 234 25310 318 25338 4 in1_16
rlabel metal1 s 536 25190 618 25218 4 in2_16
rlabel metal1 s 1176 25386 1204 25414 4 rwl0_16
rlabel metal1 s 1176 25612 1204 25640 4 rwl1_16
rlabel metal1 s 1176 25260 1204 25288 4 wwl0_16
rlabel metal1 s 56 26808 126 26836 4 in0_17
rlabel metal1 s 234 26954 318 26982 4 in1_17
rlabel metal1 s 536 27074 618 27102 4 in2_17
rlabel metal1 s 1176 26878 1204 26906 4 rwl0_17
rlabel metal1 s 1176 26652 1204 26680 4 rwl1_17
rlabel metal1 s 1176 27004 1204 27032 4 wwl0_17
rlabel metal1 s 56 28532 126 28560 4 in0_18
rlabel metal1 s 234 28386 318 28414 4 in1_18
rlabel metal1 s 536 28266 618 28294 4 in2_18
rlabel metal1 s 1176 28462 1204 28490 4 rwl0_18
rlabel metal1 s 1176 28688 1204 28716 4 rwl1_18
rlabel metal1 s 1176 28336 1204 28364 4 wwl0_18
rlabel metal1 s 56 29884 126 29912 4 in0_19
rlabel metal1 s 234 30030 318 30058 4 in1_19
rlabel metal1 s 536 30150 618 30178 4 in2_19
rlabel metal1 s 1176 29954 1204 29982 4 rwl0_19
rlabel metal1 s 1176 29728 1204 29756 4 rwl1_19
rlabel metal1 s 1176 30080 1204 30108 4 wwl0_19
rlabel metal1 s 56 31608 126 31636 4 in0_20
rlabel metal1 s 234 31462 318 31490 4 in1_20
rlabel metal1 s 536 31342 618 31370 4 in2_20
rlabel metal1 s 1176 31538 1204 31566 4 rwl0_20
rlabel metal1 s 1176 31764 1204 31792 4 rwl1_20
rlabel metal1 s 1176 31412 1204 31440 4 wwl0_20
rlabel metal1 s 56 32960 126 32988 4 in0_21
rlabel metal1 s 234 33106 318 33134 4 in1_21
rlabel metal1 s 536 33226 618 33254 4 in2_21
rlabel metal1 s 1176 33030 1204 33058 4 rwl0_21
rlabel metal1 s 1176 32804 1204 32832 4 rwl1_21
rlabel metal1 s 1176 33156 1204 33184 4 wwl0_21
rlabel metal1 s 56 34684 126 34712 4 in0_22
rlabel metal1 s 234 34538 318 34566 4 in1_22
rlabel metal1 s 536 34418 618 34446 4 in2_22
rlabel metal1 s 1176 34614 1204 34642 4 rwl0_22
rlabel metal1 s 1176 34840 1204 34868 4 rwl1_22
rlabel metal1 s 1176 34488 1204 34516 4 wwl0_22
rlabel metal1 s 56 36036 126 36064 4 in0_23
rlabel metal1 s 234 36182 318 36210 4 in1_23
rlabel metal1 s 536 36302 618 36330 4 in2_23
rlabel metal1 s 1176 36106 1204 36134 4 rwl0_23
rlabel metal1 s 1176 35880 1204 35908 4 rwl1_23
rlabel metal1 s 1176 36232 1204 36260 4 wwl0_23
rlabel metal1 s 56 37760 126 37788 4 in0_24
rlabel metal1 s 234 37614 318 37642 4 in1_24
rlabel metal1 s 536 37494 618 37522 4 in2_24
rlabel metal1 s 1176 37690 1204 37718 4 rwl0_24
rlabel metal1 s 1176 37916 1204 37944 4 rwl1_24
rlabel metal1 s 1176 37564 1204 37592 4 wwl0_24
rlabel metal1 s 56 39112 126 39140 4 in0_25
rlabel metal1 s 234 39258 318 39286 4 in1_25
rlabel metal1 s 536 39378 618 39406 4 in2_25
rlabel metal1 s 1176 39182 1204 39210 4 rwl0_25
rlabel metal1 s 1176 38956 1204 38984 4 rwl1_25
rlabel metal1 s 1176 39308 1204 39336 4 wwl0_25
rlabel metal1 s 56 40836 126 40864 4 in0_26
rlabel metal1 s 234 40690 318 40718 4 in1_26
rlabel metal1 s 536 40570 618 40598 4 in2_26
rlabel metal1 s 1176 40766 1204 40794 4 rwl0_26
rlabel metal1 s 1176 40992 1204 41020 4 rwl1_26
rlabel metal1 s 1176 40640 1204 40668 4 wwl0_26
rlabel metal1 s 56 42188 126 42216 4 in0_27
rlabel metal1 s 234 42334 318 42362 4 in1_27
rlabel metal1 s 536 42454 618 42482 4 in2_27
rlabel metal1 s 1176 42258 1204 42286 4 rwl0_27
rlabel metal1 s 1176 42032 1204 42060 4 rwl1_27
rlabel metal1 s 1176 42384 1204 42412 4 wwl0_27
rlabel metal1 s 56 43912 126 43940 4 in0_28
rlabel metal1 s 234 43766 318 43794 4 in1_28
rlabel metal1 s 536 43646 618 43674 4 in2_28
rlabel metal1 s 1176 43842 1204 43870 4 rwl0_28
rlabel metal1 s 1176 44068 1204 44096 4 rwl1_28
rlabel metal1 s 1176 43716 1204 43744 4 wwl0_28
rlabel metal1 s 56 45264 126 45292 4 in0_29
rlabel metal1 s 234 45410 318 45438 4 in1_29
rlabel metal1 s 536 45530 618 45558 4 in2_29
rlabel metal1 s 1176 45334 1204 45362 4 rwl0_29
rlabel metal1 s 1176 45108 1204 45136 4 rwl1_29
rlabel metal1 s 1176 45460 1204 45488 4 wwl0_29
rlabel metal1 s 56 46988 126 47016 4 in0_30
rlabel metal1 s 234 46842 318 46870 4 in1_30
rlabel metal1 s 536 46722 618 46750 4 in2_30
rlabel metal1 s 1176 46918 1204 46946 4 rwl0_30
rlabel metal1 s 1176 47144 1204 47172 4 rwl1_30
rlabel metal1 s 1176 46792 1204 46820 4 wwl0_30
rlabel metal1 s 56 48340 126 48368 4 in0_31
rlabel metal1 s 234 48486 318 48514 4 in1_31
rlabel metal1 s 536 48606 618 48634 4 in2_31
rlabel metal1 s 1176 48410 1204 48438 4 rwl0_31
rlabel metal1 s 1176 48184 1204 48212 4 rwl1_31
rlabel metal1 s 1176 48536 1204 48564 4 wwl0_31
rlabel metal3 s 1138 32265 1270 32331 4 vdd
rlabel metal3 s 1138 7657 1270 7723 4 vdd
rlabel metal3 s 1138 44569 1270 44635 4 vdd
rlabel metal3 s 1204 44602 1204 44602 4 vdd
rlabel metal3 s 1138 47645 1270 47711 4 vdd
rlabel metal3 s 1138 13809 1270 13875 4 vdd
rlabel metal3 s 1138 16885 1270 16951 4 vdd
rlabel metal3 s 1138 19961 1270 20027 4 vdd
rlabel metal3 s 1138 35341 1270 35407 4 vdd
rlabel metal3 s 1138 38417 1270 38483 4 vdd
rlabel metal3 s 1138 29189 1270 29255 4 vdd
rlabel metal3 s 1138 26113 1270 26179 4 vdd
rlabel metal3 s 1138 1505 1270 1571 4 vdd
rlabel metal3 s 1204 1538 1204 1538 4 vdd
rlabel metal3 s 1138 4581 1270 4647 4 vdd
rlabel metal3 s 1138 10733 1270 10799 4 vdd
rlabel metal3 s 1204 10766 1204 10766 4 vdd
rlabel metal3 s 1138 41493 1270 41559 4 vdd
rlabel metal3 s 1138 23037 1270 23103 4 vdd
rlabel metal3 s 1138 43031 1270 43097 4 gnd
rlabel metal3 s 1138 12271 1270 12337 4 gnd
rlabel metal3 s 1138 18423 1270 18489 4 gnd
rlabel metal3 s 1138 9195 1270 9261 4 gnd
rlabel metal3 s 1138 49183 1270 49249 4 gnd
rlabel metal3 s 1138 30727 1270 30793 4 gnd
rlabel metal3 s 1138 15347 1270 15413 4 gnd
rlabel metal3 s 1138 27651 1270 27717 4 gnd
rlabel metal3 s 1138 36879 1270 36945 4 gnd
rlabel metal3 s 1138 46107 1270 46173 4 gnd
rlabel metal3 s 1138 3043 1270 3109 4 gnd
rlabel metal3 s 1138 21499 1270 21565 4 gnd
rlabel metal3 s 1138 24575 1270 24641 4 gnd
rlabel metal3 s 1138 33803 1270 33869 4 gnd
rlabel metal3 s 1138 39955 1270 40021 4 gnd
rlabel metal3 s 1138 6119 1270 6185 4 gnd
rlabel metal3 s 1138 -33 1270 33 4 gnd
<< properties >>
string FIXED_BBOX 1138 -33 1270 0
string GDS_FILE sram_0rw2r1w_16_128_sky130A.gds
string GDS_END 1964026
string GDS_START 1907918
<< end >>
